magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1403 -1396 17394 41260
<< nwell >>
rect 10643 39191 11403 39832
rect -83 28976 1049 35795
rect -83 26133 1049 28076
rect 15910 5957 16090 7211
rect 15910 3831 16090 5069
rect 8286 0 8321 701
<< pwell >>
rect 3120 35861 15603 36067
rect -43 19217 1009 26071
rect 7911 19217 9168 19247
rect -43 19025 9168 19217
rect -43 18587 1826 19025
rect 5746 18999 9168 19025
rect 1272 17764 1826 18587
rect 312 9083 943 9169
rect 13907 2063 14356 2311
rect 13252 1940 14356 2063
rect 13106 1923 14356 1940
rect 13106 1889 13959 1923
rect 13106 1272 13446 1889
rect 1535 1054 13446 1272
rect 12197 1020 13446 1054
rect 12248 990 13446 1020
rect 12849 24 13241 226
<< psubdiff >>
rect 13925 35981 15577 36041
rect 13959 35947 13996 35981
rect 14030 35947 14067 35981
rect 14101 35947 14138 35981
rect 14172 35947 14209 35981
rect 14243 35947 14280 35981
rect 14314 35947 14351 35981
rect 14385 35947 14422 35981
rect 14456 35947 14493 35981
rect 14527 35947 14563 35981
rect 14597 35947 14633 35981
rect 14667 35947 14703 35981
rect 14737 35947 14773 35981
rect 14807 35947 14843 35981
rect 14877 35947 14913 35981
rect 14947 35947 14983 35981
rect 15017 35947 15053 35981
rect 15087 35947 15123 35981
rect 15157 35947 15193 35981
rect 15227 35947 15263 35981
rect 15297 35947 15333 35981
rect 15367 35947 15403 35981
rect 15437 35947 15473 35981
rect 15507 35947 15543 35981
rect 13925 35887 15577 35947
rect 12875 176 13215 200
rect 12909 142 12977 176
rect 13011 142 13079 176
rect 13113 142 13181 176
rect 12875 108 13215 142
rect 12909 74 12977 108
rect 13011 74 13079 108
rect 13113 74 13181 108
rect 12875 50 13215 74
<< mvpsubdiff >>
rect 3146 35981 13785 36041
rect 3180 35947 3215 35981
rect 3249 35947 3284 35981
rect 3318 35947 3353 35981
rect 3387 35947 3422 35981
rect 3456 35947 3491 35981
rect 3525 35947 3560 35981
rect 3594 35947 3629 35981
rect 3663 35947 3698 35981
rect 3732 35947 3767 35981
rect 3801 35947 3836 35981
rect 3870 35947 3905 35981
rect 3939 35947 3974 35981
rect 4008 35947 4043 35981
rect 4077 35947 4112 35981
rect 4146 35947 4181 35981
rect 4215 35947 4250 35981
rect 4284 35947 4319 35981
rect 4353 35947 4388 35981
rect 4422 35947 4457 35981
rect 4491 35947 4526 35981
rect 4560 35947 4595 35981
rect 4629 35947 4664 35981
rect 4698 35947 4733 35981
rect 4767 35947 4802 35981
rect 4836 35947 4871 35981
rect 4905 35947 4940 35981
rect 4974 35947 5009 35981
rect 5043 35947 5078 35981
rect 5112 35947 5147 35981
rect 5181 35947 5216 35981
rect 5250 35947 5285 35981
rect 5319 35947 5354 35981
rect 5388 35947 5423 35981
rect 5457 35947 5492 35981
rect 5526 35947 5561 35981
rect 5595 35947 5630 35981
rect 5664 35947 5699 35981
rect 5733 35947 5768 35981
rect 5802 35947 5837 35981
rect 5871 35947 5906 35981
rect 5940 35947 5975 35981
rect 6009 35947 6044 35981
rect 6078 35947 6113 35981
rect 6147 35947 6182 35981
rect 6216 35947 6251 35981
rect 6285 35947 6320 35981
rect 6354 35947 6389 35981
rect 6423 35947 6458 35981
rect 6492 35947 6527 35981
rect 6561 35947 6596 35981
rect 6630 35947 6665 35981
rect 6699 35947 6734 35981
rect 6768 35947 6803 35981
rect 6837 35947 6872 35981
rect 6906 35947 6941 35981
rect 6975 35947 7010 35981
rect 7044 35947 7079 35981
rect 7113 35947 7148 35981
rect 7182 35947 7217 35981
rect 7251 35947 7286 35981
rect 7320 35947 7355 35981
rect 7389 35947 7424 35981
rect 7458 35947 7493 35981
rect 7527 35947 7562 35981
rect 7596 35947 7631 35981
rect 7665 35947 7699 35981
rect 7733 35947 7767 35981
rect 7801 35947 7835 35981
rect 7869 35947 7903 35981
rect 7937 35947 7971 35981
rect 8005 35947 8039 35981
rect 8073 35947 8107 35981
rect 8141 35947 8175 35981
rect 8209 35947 8243 35981
rect 8277 35947 8311 35981
rect 8345 35947 8379 35981
rect 8413 35947 8447 35981
rect 8481 35947 8515 35981
rect 8549 35947 8583 35981
rect 8617 35947 8651 35981
rect 8685 35947 8719 35981
rect 8753 35947 8787 35981
rect 8821 35947 8855 35981
rect 8889 35947 8923 35981
rect 8957 35947 8991 35981
rect 9025 35947 9059 35981
rect 9093 35947 9127 35981
rect 9161 35947 9195 35981
rect 9229 35947 9263 35981
rect 9297 35947 9331 35981
rect 9365 35947 9399 35981
rect 9433 35947 9467 35981
rect 9501 35947 9535 35981
rect 9569 35947 9603 35981
rect 9637 35947 9671 35981
rect 9705 35947 9739 35981
rect 9773 35947 9807 35981
rect 9841 35947 9875 35981
rect 9909 35947 9943 35981
rect 9977 35947 10011 35981
rect 10045 35947 10079 35981
rect 10113 35947 10147 35981
rect 10181 35947 10215 35981
rect 10249 35947 10283 35981
rect 10317 35947 10351 35981
rect 10385 35947 10419 35981
rect 10453 35947 10487 35981
rect 10521 35947 10555 35981
rect 10589 35947 10623 35981
rect 10657 35947 10691 35981
rect 10725 35947 10759 35981
rect 10793 35947 10827 35981
rect 10861 35947 10895 35981
rect 10929 35947 10963 35981
rect 10997 35947 11031 35981
rect 11065 35947 11099 35981
rect 11133 35947 11167 35981
rect 11201 35947 11235 35981
rect 11269 35947 11303 35981
rect 11337 35947 11371 35981
rect 11405 35947 11439 35981
rect 11473 35947 11507 35981
rect 11541 35947 11575 35981
rect 11609 35947 11643 35981
rect 11677 35947 11711 35981
rect 11745 35947 11779 35981
rect 11813 35947 11847 35981
rect 11881 35947 11915 35981
rect 11949 35947 11983 35981
rect 12017 35947 12051 35981
rect 12085 35947 12119 35981
rect 12153 35947 12187 35981
rect 12221 35947 12255 35981
rect 12289 35947 12323 35981
rect 12357 35947 12391 35981
rect 12425 35947 12459 35981
rect 12493 35947 12527 35981
rect 12561 35947 12595 35981
rect 12629 35947 12663 35981
rect 12697 35947 12731 35981
rect 12765 35947 12799 35981
rect 12833 35947 12867 35981
rect 12901 35947 12935 35981
rect 12969 35947 13003 35981
rect 13037 35947 13071 35981
rect 13105 35947 13139 35981
rect 13173 35947 13207 35981
rect 13241 35947 13275 35981
rect 13309 35947 13343 35981
rect 13377 35947 13411 35981
rect 13445 35947 13479 35981
rect 13513 35947 13547 35981
rect 13581 35947 13615 35981
rect 13649 35947 13683 35981
rect 13717 35947 13751 35981
rect 3146 35887 13785 35947
rect -17 26021 843 26045
rect 17 25987 55 26021
rect 89 25987 127 26021
rect 161 25987 199 26021
rect 233 25987 271 26021
rect 305 25987 343 26021
rect 377 25987 415 26021
rect 449 25987 487 26021
rect 521 25987 559 26021
rect 593 25987 631 26021
rect 665 25987 703 26021
rect 737 25987 775 26021
rect 809 26011 843 26021
rect 877 26011 915 26045
rect 949 26011 983 26045
rect 809 25987 983 26011
rect -17 25972 983 25987
rect -17 25952 843 25972
rect 17 25918 55 25952
rect 89 25918 127 25952
rect 161 25918 199 25952
rect 233 25918 271 25952
rect 305 25918 343 25952
rect 377 25918 415 25952
rect 449 25918 487 25952
rect 521 25918 559 25952
rect 593 25918 631 25952
rect 665 25918 703 25952
rect 737 25918 775 25952
rect 809 25938 843 25952
rect 877 25938 915 25972
rect 949 25938 983 25972
rect 809 25918 983 25938
rect -17 25899 983 25918
rect -17 25883 843 25899
rect 17 25849 55 25883
rect 89 25849 127 25883
rect 161 25849 199 25883
rect 233 25849 271 25883
rect 305 25849 343 25883
rect 377 25849 415 25883
rect 449 25849 487 25883
rect 521 25849 559 25883
rect 593 25849 631 25883
rect 665 25849 703 25883
rect 737 25849 775 25883
rect 809 25865 843 25883
rect 877 25865 915 25899
rect 949 25865 983 25899
rect 809 25849 983 25865
rect -17 25826 983 25849
rect -17 25814 843 25826
rect 17 25780 55 25814
rect 89 25780 127 25814
rect 161 25780 199 25814
rect 233 25780 271 25814
rect 305 25780 343 25814
rect 377 25780 415 25814
rect 449 25780 487 25814
rect 521 25780 559 25814
rect 593 25780 631 25814
rect 665 25780 703 25814
rect 737 25780 775 25814
rect 809 25792 843 25814
rect 877 25792 915 25826
rect 949 25792 983 25826
rect 809 25780 983 25792
rect -17 25753 983 25780
rect -17 25745 843 25753
rect 17 25711 55 25745
rect 89 25711 127 25745
rect 161 25711 199 25745
rect 233 25711 271 25745
rect 305 25711 343 25745
rect 377 25711 415 25745
rect 449 25711 487 25745
rect 521 25711 559 25745
rect 593 25711 631 25745
rect 665 25711 703 25745
rect 737 25711 775 25745
rect 809 25719 843 25745
rect 877 25719 915 25753
rect 949 25719 983 25753
rect 809 25711 983 25719
rect -17 25680 983 25711
rect -17 25676 843 25680
rect 17 25642 55 25676
rect 89 25642 127 25676
rect 161 25642 199 25676
rect 233 25642 271 25676
rect 305 25642 343 25676
rect 377 25642 415 25676
rect 449 25642 487 25676
rect 521 25642 559 25676
rect 593 25642 631 25676
rect 665 25642 703 25676
rect 737 25642 775 25676
rect 809 25646 843 25676
rect 877 25646 915 25680
rect 949 25646 983 25680
rect 809 25642 983 25646
rect -17 25607 983 25642
rect 17 25573 55 25607
rect 89 25573 127 25607
rect 161 25573 199 25607
rect 233 25573 271 25607
rect 305 25573 343 25607
rect 377 25573 415 25607
rect 449 25573 487 25607
rect 521 25573 559 25607
rect 593 25573 631 25607
rect 665 25573 703 25607
rect 737 25573 775 25607
rect 809 25573 843 25607
rect 877 25573 915 25607
rect 949 25573 983 25607
rect -17 25539 983 25573
rect 17 25505 55 25539
rect 89 25505 127 25539
rect 161 25505 199 25539
rect 233 25505 271 25539
rect 305 25505 343 25539
rect 377 25505 415 25539
rect 449 25505 487 25539
rect 521 25505 559 25539
rect 593 25505 631 25539
rect 665 25505 703 25539
rect 737 25505 775 25539
rect 809 25534 983 25539
rect 809 25505 843 25534
rect -17 25500 843 25505
rect 877 25500 915 25534
rect 949 25500 983 25534
rect -17 25471 983 25500
rect 17 25437 55 25471
rect 89 25437 127 25471
rect 161 25437 199 25471
rect 233 25437 271 25471
rect 305 25437 343 25471
rect 377 25437 415 25471
rect 449 25437 487 25471
rect 521 25437 559 25471
rect 593 25437 631 25471
rect 665 25437 703 25471
rect 737 25437 775 25471
rect 809 25461 983 25471
rect 809 25437 843 25461
rect -17 25427 843 25437
rect 877 25427 915 25461
rect 949 25427 983 25461
rect -17 25403 983 25427
rect 17 25369 55 25403
rect 89 25369 127 25403
rect 161 25369 199 25403
rect 233 25369 271 25403
rect 305 25369 343 25403
rect 377 25369 415 25403
rect 449 25369 487 25403
rect 521 25369 559 25403
rect 593 25369 631 25403
rect 665 25369 703 25403
rect 737 25369 775 25403
rect 809 25388 983 25403
rect 809 25369 843 25388
rect -17 25354 843 25369
rect 877 25354 915 25388
rect 949 25354 983 25388
rect -17 25335 983 25354
rect 17 25301 55 25335
rect 89 25301 127 25335
rect 161 25301 199 25335
rect 233 25301 271 25335
rect 305 25301 343 25335
rect 377 25301 415 25335
rect 449 25301 487 25335
rect 521 25301 559 25335
rect 593 25301 631 25335
rect 665 25301 703 25335
rect 737 25301 775 25335
rect 809 25316 983 25335
rect 809 25301 843 25316
rect -17 25282 843 25301
rect 877 25282 915 25316
rect 949 25282 983 25316
rect -17 25267 983 25282
rect 17 25233 55 25267
rect 89 25233 127 25267
rect 161 25233 199 25267
rect 233 25233 271 25267
rect 305 25233 343 25267
rect 377 25233 415 25267
rect 449 25233 487 25267
rect 521 25233 559 25267
rect 593 25233 631 25267
rect 665 25233 703 25267
rect 737 25233 775 25267
rect 809 25256 983 25267
rect 809 25233 835 25256
rect -17 25199 835 25233
rect 17 25165 55 25199
rect 89 25165 127 25199
rect 161 25165 199 25199
rect 233 25165 271 25199
rect 305 25165 343 25199
rect 377 25165 415 25199
rect 449 25165 487 25199
rect 521 25165 559 25199
rect 593 25165 631 25199
rect 665 25165 703 25199
rect 737 25165 775 25199
rect 809 25165 835 25199
rect -17 25131 835 25165
rect 17 25097 55 25131
rect 89 25097 127 25131
rect 161 25097 199 25131
rect 233 25097 271 25131
rect 305 25097 343 25131
rect 377 25097 415 25131
rect 449 25097 487 25131
rect 521 25097 559 25131
rect 593 25097 631 25131
rect 665 25097 703 25131
rect 737 25097 775 25131
rect 809 25097 835 25131
rect -17 25063 835 25097
rect 17 25029 55 25063
rect 89 25029 127 25063
rect 161 25029 199 25063
rect 233 25029 271 25063
rect 305 25029 343 25063
rect 377 25029 415 25063
rect 449 25029 487 25063
rect 521 25029 559 25063
rect 593 25029 631 25063
rect 665 25029 703 25063
rect 737 25029 775 25063
rect 809 25029 835 25063
rect -17 24995 835 25029
rect 17 24961 55 24995
rect 89 24961 127 24995
rect 161 24961 199 24995
rect 233 24961 271 24995
rect 305 24961 343 24995
rect 377 24961 415 24995
rect 449 24961 487 24995
rect 521 24961 559 24995
rect 593 24961 631 24995
rect 665 24961 703 24995
rect 737 24961 775 24995
rect 809 24961 835 24995
rect -17 24927 835 24961
rect 17 24893 55 24927
rect 89 24893 127 24927
rect 161 24893 199 24927
rect 233 24893 271 24927
rect 305 24893 343 24927
rect 377 24893 415 24927
rect 449 24893 487 24927
rect 521 24893 559 24927
rect 593 24893 631 24927
rect 665 24893 703 24927
rect 737 24893 775 24927
rect 809 24893 835 24927
rect -17 24859 835 24893
rect 17 24825 55 24859
rect 89 24825 127 24859
rect 161 24825 199 24859
rect 233 24825 271 24859
rect 305 24825 343 24859
rect 377 24825 415 24859
rect 449 24825 487 24859
rect 521 24825 559 24859
rect 593 24825 631 24859
rect 665 24825 703 24859
rect 737 24825 775 24859
rect 809 24825 835 24859
rect -17 24791 835 24825
rect 17 24757 55 24791
rect 89 24757 127 24791
rect 161 24757 199 24791
rect 233 24757 271 24791
rect 305 24757 343 24791
rect 377 24757 415 24791
rect 449 24757 487 24791
rect 521 24757 559 24791
rect 593 24757 631 24791
rect 665 24757 703 24791
rect 737 24757 775 24791
rect 809 24757 835 24791
rect -17 24723 835 24757
rect 17 24689 55 24723
rect 89 24689 127 24723
rect 161 24689 199 24723
rect 233 24689 271 24723
rect 305 24689 343 24723
rect 377 24689 415 24723
rect 449 24689 487 24723
rect 521 24689 559 24723
rect 593 24689 631 24723
rect 665 24689 703 24723
rect 737 24689 775 24723
rect 809 24689 835 24723
rect -17 24655 835 24689
rect 17 24621 55 24655
rect 89 24621 127 24655
rect 161 24621 199 24655
rect 233 24621 271 24655
rect 305 24621 343 24655
rect 377 24621 415 24655
rect 449 24621 487 24655
rect 521 24621 559 24655
rect 593 24621 631 24655
rect 665 24621 703 24655
rect 737 24621 775 24655
rect 809 24621 835 24655
rect -17 24587 835 24621
rect 17 24553 55 24587
rect 89 24553 127 24587
rect 161 24553 199 24587
rect 233 24553 271 24587
rect 305 24553 343 24587
rect 377 24553 415 24587
rect 449 24553 487 24587
rect 521 24553 559 24587
rect 593 24553 631 24587
rect 665 24553 703 24587
rect 737 24553 775 24587
rect 809 24553 835 24587
rect -17 24519 835 24553
rect 17 24485 55 24519
rect 89 24485 127 24519
rect 161 24485 199 24519
rect 233 24485 271 24519
rect 305 24485 343 24519
rect 377 24485 415 24519
rect 449 24485 487 24519
rect 521 24485 559 24519
rect 593 24485 631 24519
rect 665 24485 703 24519
rect 737 24485 775 24519
rect 809 24485 835 24519
rect -17 24451 835 24485
rect 17 24417 55 24451
rect 89 24417 127 24451
rect 161 24417 199 24451
rect 233 24417 271 24451
rect 305 24417 343 24451
rect 377 24417 415 24451
rect 449 24417 487 24451
rect 521 24417 559 24451
rect 593 24417 631 24451
rect 665 24417 703 24451
rect 737 24417 775 24451
rect 809 24417 835 24451
rect -17 24383 835 24417
rect 17 24349 55 24383
rect 89 24349 127 24383
rect 161 24349 199 24383
rect 233 24349 271 24383
rect 305 24349 343 24383
rect 377 24349 415 24383
rect 449 24349 487 24383
rect 521 24349 559 24383
rect 593 24349 631 24383
rect 665 24349 703 24383
rect 737 24349 775 24383
rect 809 24349 835 24383
rect -17 24315 835 24349
rect 17 24281 55 24315
rect 89 24281 127 24315
rect 161 24281 199 24315
rect 233 24281 271 24315
rect 305 24281 343 24315
rect 377 24281 415 24315
rect 449 24281 487 24315
rect 521 24281 559 24315
rect 593 24281 631 24315
rect 665 24281 703 24315
rect 737 24281 775 24315
rect 809 24281 835 24315
rect -17 24247 835 24281
rect 17 24213 55 24247
rect 89 24213 127 24247
rect 161 24213 199 24247
rect 233 24213 271 24247
rect 305 24213 343 24247
rect 377 24213 415 24247
rect 449 24213 487 24247
rect 521 24213 559 24247
rect 593 24213 631 24247
rect 665 24213 703 24247
rect 737 24213 775 24247
rect 809 24213 835 24247
rect -17 24179 835 24213
rect 17 24145 55 24179
rect 89 24145 127 24179
rect 161 24145 199 24179
rect 233 24145 271 24179
rect 305 24145 343 24179
rect 377 24145 415 24179
rect 449 24145 487 24179
rect 521 24145 559 24179
rect 593 24145 631 24179
rect 665 24145 703 24179
rect 737 24145 775 24179
rect 809 24145 835 24179
rect -17 24111 835 24145
rect 17 24077 55 24111
rect 89 24077 127 24111
rect 161 24077 199 24111
rect 233 24077 271 24111
rect 305 24077 343 24111
rect 377 24077 415 24111
rect 449 24077 487 24111
rect 521 24077 559 24111
rect 593 24077 631 24111
rect 665 24077 703 24111
rect 737 24077 775 24111
rect 809 24077 835 24111
rect -17 24043 835 24077
rect 17 24009 55 24043
rect 89 24009 127 24043
rect 161 24009 199 24043
rect 233 24009 271 24043
rect 305 24009 343 24043
rect 377 24009 415 24043
rect 449 24009 487 24043
rect 521 24009 559 24043
rect 593 24009 631 24043
rect 665 24009 703 24043
rect 737 24009 775 24043
rect 809 24009 835 24043
rect -17 23975 835 24009
rect 17 23941 55 23975
rect 89 23941 127 23975
rect 161 23941 199 23975
rect 233 23941 271 23975
rect 305 23941 343 23975
rect 377 23941 415 23975
rect 449 23941 487 23975
rect 521 23941 559 23975
rect 593 23941 631 23975
rect 665 23941 703 23975
rect 737 23941 775 23975
rect 809 23941 835 23975
rect -17 23907 835 23941
rect 17 23873 55 23907
rect 89 23873 127 23907
rect 161 23873 199 23907
rect 233 23873 271 23907
rect 305 23873 343 23907
rect 377 23873 415 23907
rect 449 23873 487 23907
rect 521 23873 559 23907
rect 593 23873 631 23907
rect 665 23873 703 23907
rect 737 23873 775 23907
rect 809 23873 835 23907
rect -17 23839 835 23873
rect 17 23805 55 23839
rect 89 23805 127 23839
rect 161 23805 199 23839
rect 233 23805 271 23839
rect 305 23805 343 23839
rect 377 23805 415 23839
rect 449 23805 487 23839
rect 521 23805 559 23839
rect 593 23805 631 23839
rect 665 23805 703 23839
rect 737 23805 775 23839
rect 809 23805 835 23839
rect -17 23771 835 23805
rect 17 23737 55 23771
rect 89 23737 127 23771
rect 161 23737 199 23771
rect 233 23737 271 23771
rect 305 23737 343 23771
rect 377 23737 415 23771
rect 449 23737 487 23771
rect 521 23737 559 23771
rect 593 23737 631 23771
rect 665 23737 703 23771
rect 737 23737 775 23771
rect 809 23737 835 23771
rect -17 23703 835 23737
rect 17 23669 55 23703
rect 89 23669 127 23703
rect 161 23669 199 23703
rect 233 23669 271 23703
rect 305 23669 343 23703
rect 377 23669 415 23703
rect 449 23669 487 23703
rect 521 23669 559 23703
rect 593 23669 631 23703
rect 665 23669 703 23703
rect 737 23669 775 23703
rect 809 23669 835 23703
rect -17 23635 835 23669
rect 17 23601 55 23635
rect 89 23601 127 23635
rect 161 23601 199 23635
rect 233 23601 271 23635
rect 305 23601 343 23635
rect 377 23601 415 23635
rect 449 23601 487 23635
rect 521 23601 559 23635
rect 593 23601 631 23635
rect 665 23601 703 23635
rect 737 23601 775 23635
rect 809 23601 835 23635
rect -17 23567 835 23601
rect 17 23533 55 23567
rect 89 23533 127 23567
rect 161 23533 199 23567
rect 233 23533 271 23567
rect 305 23533 343 23567
rect 377 23533 415 23567
rect 449 23533 487 23567
rect 521 23533 559 23567
rect 593 23533 631 23567
rect 665 23533 703 23567
rect 737 23533 775 23567
rect 809 23533 835 23567
rect -17 23499 835 23533
rect 17 23465 55 23499
rect 89 23465 127 23499
rect 161 23465 199 23499
rect 233 23465 271 23499
rect 305 23465 343 23499
rect 377 23465 415 23499
rect 449 23465 487 23499
rect 521 23465 559 23499
rect 593 23465 631 23499
rect 665 23465 703 23499
rect 737 23465 775 23499
rect 809 23465 835 23499
rect -17 23431 835 23465
rect 17 23397 55 23431
rect 89 23397 127 23431
rect 161 23397 199 23431
rect 233 23397 271 23431
rect 305 23397 343 23431
rect 377 23397 415 23431
rect 449 23397 487 23431
rect 521 23397 559 23431
rect 593 23397 631 23431
rect 665 23397 703 23431
rect 737 23397 775 23431
rect 809 23397 835 23431
rect -17 23363 835 23397
rect 17 23329 55 23363
rect 89 23329 127 23363
rect 161 23329 199 23363
rect 233 23329 271 23363
rect 305 23329 343 23363
rect 377 23329 415 23363
rect 449 23329 487 23363
rect 521 23329 559 23363
rect 593 23329 631 23363
rect 665 23329 703 23363
rect 737 23329 775 23363
rect 809 23329 835 23363
rect -17 23295 835 23329
rect 17 23261 55 23295
rect 89 23261 127 23295
rect 161 23261 199 23295
rect 233 23261 271 23295
rect 305 23261 343 23295
rect 377 23261 415 23295
rect 449 23261 487 23295
rect 521 23261 559 23295
rect 593 23261 631 23295
rect 665 23261 703 23295
rect 737 23261 775 23295
rect 809 23261 835 23295
rect -17 23227 835 23261
rect 17 23193 55 23227
rect 89 23193 127 23227
rect 161 23193 199 23227
rect 233 23193 271 23227
rect 305 23193 343 23227
rect 377 23193 415 23227
rect 449 23193 487 23227
rect 521 23193 559 23227
rect 593 23193 631 23227
rect 665 23193 703 23227
rect 737 23193 775 23227
rect 809 23193 835 23227
rect -17 23159 835 23193
rect 17 23125 55 23159
rect 89 23125 127 23159
rect 161 23125 199 23159
rect 233 23125 271 23159
rect 305 23125 343 23159
rect 377 23125 415 23159
rect 449 23125 487 23159
rect 521 23125 559 23159
rect 593 23125 631 23159
rect 665 23125 703 23159
rect 737 23125 775 23159
rect 809 23125 835 23159
rect -17 23091 835 23125
rect 17 23057 55 23091
rect 89 23057 127 23091
rect 161 23057 199 23091
rect 233 23057 271 23091
rect 305 23057 343 23091
rect 377 23057 415 23091
rect 449 23057 487 23091
rect 521 23057 559 23091
rect 593 23057 631 23091
rect 665 23057 703 23091
rect 737 23057 775 23091
rect 809 23057 835 23091
rect -17 23023 835 23057
rect 17 22989 55 23023
rect 89 22989 127 23023
rect 161 22989 199 23023
rect 233 22989 271 23023
rect 305 22989 343 23023
rect 377 22989 415 23023
rect 449 22989 487 23023
rect 521 22989 559 23023
rect 593 22989 631 23023
rect 665 22989 703 23023
rect 737 22989 775 23023
rect 809 22989 835 23023
rect -17 22955 835 22989
rect 17 22921 55 22955
rect 89 22921 127 22955
rect 161 22921 199 22955
rect 233 22921 271 22955
rect 305 22921 343 22955
rect 377 22921 415 22955
rect 449 22921 487 22955
rect 521 22921 559 22955
rect 593 22921 631 22955
rect 665 22921 703 22955
rect 737 22921 775 22955
rect 809 22921 835 22955
rect -17 22887 835 22921
rect 17 22853 55 22887
rect 89 22853 127 22887
rect 161 22853 199 22887
rect 233 22853 271 22887
rect 305 22853 343 22887
rect 377 22853 415 22887
rect 449 22853 487 22887
rect 521 22853 559 22887
rect 593 22853 631 22887
rect 665 22853 703 22887
rect 737 22853 775 22887
rect 809 22853 835 22887
rect -17 22819 835 22853
rect 17 22785 55 22819
rect 89 22785 127 22819
rect 161 22785 199 22819
rect 233 22785 271 22819
rect 305 22785 343 22819
rect 377 22785 415 22819
rect 449 22785 487 22819
rect 521 22785 559 22819
rect 593 22785 631 22819
rect 665 22785 703 22819
rect 737 22785 775 22819
rect 809 22785 835 22819
rect -17 22751 835 22785
rect 17 22717 55 22751
rect 89 22717 127 22751
rect 161 22717 199 22751
rect 233 22717 271 22751
rect 305 22717 343 22751
rect 377 22717 415 22751
rect 449 22717 487 22751
rect 521 22717 559 22751
rect 593 22717 631 22751
rect 665 22717 703 22751
rect 737 22717 775 22751
rect 809 22717 835 22751
rect -17 22683 835 22717
rect 17 22649 55 22683
rect 89 22649 127 22683
rect 161 22649 199 22683
rect 233 22649 271 22683
rect 305 22649 343 22683
rect 377 22649 415 22683
rect 449 22649 487 22683
rect 521 22649 559 22683
rect 593 22649 631 22683
rect 665 22649 703 22683
rect 737 22649 775 22683
rect 809 22649 835 22683
rect -17 22615 835 22649
rect 17 22581 55 22615
rect 89 22581 127 22615
rect 161 22581 199 22615
rect 233 22581 271 22615
rect 305 22581 343 22615
rect 377 22581 415 22615
rect 449 22581 487 22615
rect 521 22581 559 22615
rect 593 22581 631 22615
rect 665 22581 703 22615
rect 737 22581 775 22615
rect 809 22581 835 22615
rect -17 22547 835 22581
rect 17 22513 55 22547
rect 89 22513 127 22547
rect 161 22513 199 22547
rect 233 22513 271 22547
rect 305 22513 343 22547
rect 377 22513 415 22547
rect 449 22513 487 22547
rect 521 22513 559 22547
rect 593 22513 631 22547
rect 665 22513 703 22547
rect 737 22513 775 22547
rect 809 22513 835 22547
rect -17 22479 835 22513
rect 17 22445 55 22479
rect 89 22445 127 22479
rect 161 22445 199 22479
rect 233 22445 271 22479
rect 305 22445 343 22479
rect 377 22445 415 22479
rect 449 22445 487 22479
rect 521 22445 559 22479
rect 593 22445 631 22479
rect 665 22445 703 22479
rect 737 22445 775 22479
rect 809 22445 835 22479
rect -17 22411 835 22445
rect 17 22377 55 22411
rect 89 22377 127 22411
rect 161 22377 199 22411
rect 233 22377 271 22411
rect 305 22377 343 22411
rect 377 22377 415 22411
rect 449 22377 487 22411
rect 521 22377 559 22411
rect 593 22377 631 22411
rect 665 22377 703 22411
rect 737 22377 775 22411
rect 809 22377 835 22411
rect -17 22343 835 22377
rect 17 22309 55 22343
rect 89 22309 127 22343
rect 161 22309 199 22343
rect 233 22309 271 22343
rect 305 22309 343 22343
rect 377 22309 415 22343
rect 449 22309 487 22343
rect 521 22309 559 22343
rect 593 22309 631 22343
rect 665 22309 703 22343
rect 737 22309 775 22343
rect 809 22309 835 22343
rect -17 22275 835 22309
rect 17 22241 55 22275
rect 89 22241 127 22275
rect 161 22241 199 22275
rect 233 22241 271 22275
rect 305 22241 343 22275
rect 377 22241 415 22275
rect 449 22241 487 22275
rect 521 22241 559 22275
rect 593 22241 631 22275
rect 665 22241 703 22275
rect 737 22241 775 22275
rect 809 22241 835 22275
rect -17 22207 835 22241
rect 17 22173 55 22207
rect 89 22173 127 22207
rect 161 22173 199 22207
rect 233 22173 271 22207
rect 305 22173 343 22207
rect 377 22173 415 22207
rect 449 22173 487 22207
rect 521 22173 559 22207
rect 593 22173 631 22207
rect 665 22173 703 22207
rect 737 22173 775 22207
rect 809 22173 835 22207
rect -17 22139 835 22173
rect 17 22105 55 22139
rect 89 22105 127 22139
rect 161 22105 199 22139
rect 233 22105 271 22139
rect 305 22105 343 22139
rect 377 22105 415 22139
rect 449 22105 487 22139
rect 521 22105 559 22139
rect 593 22105 631 22139
rect 665 22105 703 22139
rect 737 22105 775 22139
rect 809 22105 835 22139
rect -17 22071 835 22105
rect 17 22037 55 22071
rect 89 22037 127 22071
rect 161 22037 199 22071
rect 233 22037 271 22071
rect 305 22037 343 22071
rect 377 22037 415 22071
rect 449 22037 487 22071
rect 521 22037 559 22071
rect 593 22037 631 22071
rect 665 22037 703 22071
rect 737 22037 775 22071
rect 809 22037 835 22071
rect -17 22003 835 22037
rect 17 21969 55 22003
rect 89 21969 127 22003
rect 161 21969 199 22003
rect 233 21969 271 22003
rect 305 21969 343 22003
rect 377 21969 415 22003
rect 449 21969 487 22003
rect 521 21969 559 22003
rect 593 21969 631 22003
rect 665 21969 703 22003
rect 737 21969 775 22003
rect 809 21969 835 22003
rect -17 21935 835 21969
rect 17 21901 55 21935
rect 89 21901 127 21935
rect 161 21901 199 21935
rect 233 21901 271 21935
rect 305 21901 343 21935
rect 377 21901 415 21935
rect 449 21901 487 21935
rect 521 21901 559 21935
rect 593 21901 631 21935
rect 665 21901 703 21935
rect 737 21901 775 21935
rect 809 21901 835 21935
rect -17 21867 835 21901
rect 17 21833 55 21867
rect 89 21833 127 21867
rect 161 21833 199 21867
rect 233 21833 271 21867
rect 305 21833 343 21867
rect 377 21833 415 21867
rect 449 21833 487 21867
rect 521 21833 559 21867
rect 593 21833 631 21867
rect 665 21833 703 21867
rect 737 21833 775 21867
rect 809 21833 835 21867
rect -17 21799 835 21833
rect 17 21765 55 21799
rect 89 21765 127 21799
rect 161 21765 199 21799
rect 233 21765 271 21799
rect 305 21765 343 21799
rect 377 21765 415 21799
rect 449 21765 487 21799
rect 521 21765 559 21799
rect 593 21765 631 21799
rect 665 21765 703 21799
rect 737 21765 775 21799
rect 809 21765 835 21799
rect -17 21731 835 21765
rect 17 21697 55 21731
rect 89 21697 127 21731
rect 161 21697 199 21731
rect 233 21697 271 21731
rect 305 21697 343 21731
rect 377 21697 415 21731
rect 449 21697 487 21731
rect 521 21697 559 21731
rect 593 21697 631 21731
rect 665 21697 703 21731
rect 737 21697 775 21731
rect 809 21697 835 21731
rect -17 21663 835 21697
rect 17 21629 55 21663
rect 89 21629 127 21663
rect 161 21629 199 21663
rect 233 21629 271 21663
rect 305 21629 343 21663
rect 377 21629 415 21663
rect 449 21629 487 21663
rect 521 21629 559 21663
rect 593 21629 631 21663
rect 665 21629 703 21663
rect 737 21629 775 21663
rect 809 21629 835 21663
rect -17 21595 835 21629
rect 17 21561 55 21595
rect 89 21561 127 21595
rect 161 21561 199 21595
rect 233 21561 271 21595
rect 305 21561 343 21595
rect 377 21561 415 21595
rect 449 21561 487 21595
rect 521 21561 559 21595
rect 593 21561 631 21595
rect 665 21561 703 21595
rect 737 21561 775 21595
rect 809 21561 835 21595
rect -17 21527 835 21561
rect 17 21493 55 21527
rect 89 21493 127 21527
rect 161 21493 199 21527
rect 233 21493 271 21527
rect 305 21493 343 21527
rect 377 21493 415 21527
rect 449 21493 487 21527
rect 521 21493 559 21527
rect 593 21493 631 21527
rect 665 21493 703 21527
rect 737 21493 775 21527
rect 809 21493 835 21527
rect -17 21459 835 21493
rect 17 21425 55 21459
rect 89 21425 127 21459
rect 161 21425 199 21459
rect 233 21425 271 21459
rect 305 21425 343 21459
rect 377 21425 415 21459
rect 449 21425 487 21459
rect 521 21425 559 21459
rect 593 21425 631 21459
rect 665 21425 703 21459
rect 737 21425 775 21459
rect 809 21425 835 21459
rect -17 21391 835 21425
rect 17 21357 55 21391
rect 89 21357 127 21391
rect 161 21357 199 21391
rect 233 21357 271 21391
rect 305 21357 343 21391
rect 377 21357 415 21391
rect 449 21357 487 21391
rect 521 21357 559 21391
rect 593 21357 631 21391
rect 665 21357 703 21391
rect 737 21357 775 21391
rect 809 21357 835 21391
rect -17 21323 835 21357
rect 17 21289 55 21323
rect 89 21289 127 21323
rect 161 21289 199 21323
rect 233 21289 271 21323
rect 305 21289 343 21323
rect 377 21289 415 21323
rect 449 21289 487 21323
rect 521 21289 559 21323
rect 593 21289 631 21323
rect 665 21289 703 21323
rect 737 21289 775 21323
rect 809 21289 835 21323
rect -17 21255 835 21289
rect 17 21221 55 21255
rect 89 21221 127 21255
rect 161 21221 199 21255
rect 233 21221 271 21255
rect 305 21221 343 21255
rect 377 21221 415 21255
rect 449 21221 487 21255
rect 521 21221 559 21255
rect 593 21221 631 21255
rect 665 21221 703 21255
rect 737 21221 775 21255
rect 809 21221 835 21255
rect -17 21187 835 21221
rect 17 21153 55 21187
rect 89 21153 127 21187
rect 161 21153 199 21187
rect 233 21153 271 21187
rect 305 21153 343 21187
rect 377 21153 415 21187
rect 449 21153 487 21187
rect 521 21153 559 21187
rect 593 21153 631 21187
rect 665 21153 703 21187
rect 737 21153 775 21187
rect 809 21153 835 21187
rect -17 21119 835 21153
rect 17 21085 55 21119
rect 89 21085 127 21119
rect 161 21085 199 21119
rect 233 21085 271 21119
rect 305 21085 343 21119
rect 377 21085 415 21119
rect 449 21085 487 21119
rect 521 21085 559 21119
rect 593 21085 631 21119
rect 665 21085 703 21119
rect 737 21085 775 21119
rect 809 21085 835 21119
rect -17 21051 835 21085
rect 17 21017 55 21051
rect 89 21017 127 21051
rect 161 21017 199 21051
rect 233 21017 271 21051
rect 305 21017 343 21051
rect 377 21017 415 21051
rect 449 21017 487 21051
rect 521 21017 559 21051
rect 593 21017 631 21051
rect 665 21017 703 21051
rect 737 21017 775 21051
rect 809 21017 835 21051
rect -17 20983 835 21017
rect 17 20949 55 20983
rect 89 20949 127 20983
rect 161 20949 199 20983
rect 233 20949 271 20983
rect 305 20949 343 20983
rect 377 20949 415 20983
rect 449 20949 487 20983
rect 521 20949 559 20983
rect 593 20949 631 20983
rect 665 20949 703 20983
rect 737 20949 775 20983
rect 809 20949 835 20983
rect -17 20915 835 20949
rect 17 20881 55 20915
rect 89 20881 127 20915
rect 161 20881 199 20915
rect 233 20881 271 20915
rect 305 20881 343 20915
rect 377 20881 415 20915
rect 449 20881 487 20915
rect 521 20881 559 20915
rect 593 20881 631 20915
rect 665 20881 703 20915
rect 737 20881 775 20915
rect 809 20881 835 20915
rect -17 20847 835 20881
rect 17 20813 55 20847
rect 89 20813 127 20847
rect 161 20813 199 20847
rect 233 20813 271 20847
rect 305 20813 343 20847
rect 377 20813 415 20847
rect 449 20813 487 20847
rect 521 20813 559 20847
rect 593 20813 631 20847
rect 665 20813 703 20847
rect 737 20813 775 20847
rect 809 20813 835 20847
rect -17 20779 835 20813
rect 17 20745 55 20779
rect 89 20745 127 20779
rect 161 20745 199 20779
rect 233 20745 271 20779
rect 305 20745 343 20779
rect 377 20745 415 20779
rect 449 20745 487 20779
rect 521 20745 559 20779
rect 593 20745 631 20779
rect 665 20745 703 20779
rect 737 20745 775 20779
rect 809 20745 835 20779
rect -17 20711 835 20745
rect 17 20677 55 20711
rect 89 20677 127 20711
rect 161 20677 199 20711
rect 233 20677 271 20711
rect 305 20677 343 20711
rect 377 20677 415 20711
rect 449 20677 487 20711
rect 521 20677 559 20711
rect 593 20677 631 20711
rect 665 20677 703 20711
rect 737 20677 775 20711
rect 809 20677 835 20711
rect -17 20643 835 20677
rect 17 20609 55 20643
rect 89 20609 127 20643
rect 161 20609 199 20643
rect 233 20609 271 20643
rect 305 20609 343 20643
rect 377 20609 415 20643
rect 449 20609 487 20643
rect 521 20609 559 20643
rect 593 20609 631 20643
rect 665 20609 703 20643
rect 737 20609 775 20643
rect 809 20609 835 20643
rect -17 20575 835 20609
rect 17 20541 55 20575
rect 89 20541 127 20575
rect 161 20541 199 20575
rect 233 20541 271 20575
rect 305 20541 343 20575
rect 377 20541 415 20575
rect 449 20541 487 20575
rect 521 20541 559 20575
rect 593 20541 631 20575
rect 665 20541 703 20575
rect 737 20541 775 20575
rect 809 20541 835 20575
rect -17 20510 835 20541
rect -17 20507 983 20510
rect 17 20473 55 20507
rect 89 20473 127 20507
rect 161 20473 199 20507
rect 233 20473 271 20507
rect 305 20473 343 20507
rect 377 20473 415 20507
rect 449 20473 487 20507
rect 521 20473 559 20507
rect 593 20473 631 20507
rect 665 20473 703 20507
rect 737 20473 775 20507
rect 809 20484 983 20507
rect 809 20473 843 20484
rect -17 20450 843 20473
rect 877 20450 915 20484
rect 949 20450 983 20484
rect -17 20439 983 20450
rect 17 20405 55 20439
rect 89 20405 127 20439
rect 161 20405 199 20439
rect 233 20405 271 20439
rect 305 20405 343 20439
rect 377 20405 415 20439
rect 449 20405 487 20439
rect 521 20405 559 20439
rect 593 20405 631 20439
rect 665 20405 703 20439
rect 737 20405 775 20439
rect 809 20415 983 20439
rect -17 20371 775 20405
rect 17 20337 55 20371
rect 89 20337 127 20371
rect 161 20337 199 20371
rect 233 20337 271 20371
rect 305 20337 343 20371
rect 377 20337 415 20371
rect 449 20337 487 20371
rect 521 20337 559 20371
rect 593 20337 631 20371
rect 665 20337 703 20371
rect 737 20337 775 20371
rect -17 20303 775 20337
rect 17 20269 55 20303
rect 89 20269 127 20303
rect 161 20269 199 20303
rect 233 20269 271 20303
rect 305 20269 343 20303
rect 377 20269 415 20303
rect 449 20269 487 20303
rect 521 20269 559 20303
rect 593 20269 631 20303
rect 665 20269 703 20303
rect 737 20269 775 20303
rect -17 20235 775 20269
rect 17 20201 55 20235
rect 89 20201 127 20235
rect 161 20201 199 20235
rect 233 20201 271 20235
rect 305 20201 343 20235
rect 377 20201 415 20235
rect 449 20201 487 20235
rect 521 20201 559 20235
rect 593 20201 631 20235
rect 665 20201 703 20235
rect 737 20201 775 20235
rect -17 20167 775 20201
rect 17 20133 55 20167
rect 89 20133 127 20167
rect 161 20133 199 20167
rect 233 20133 271 20167
rect 305 20133 343 20167
rect 377 20133 415 20167
rect 449 20133 487 20167
rect 521 20133 559 20167
rect 593 20133 631 20167
rect 665 20133 703 20167
rect 737 20133 775 20167
rect -17 20099 775 20133
rect 17 20065 55 20099
rect 89 20065 127 20099
rect 161 20065 199 20099
rect 233 20065 271 20099
rect 305 20065 343 20099
rect 377 20065 415 20099
rect 449 20065 487 20099
rect 521 20065 559 20099
rect 593 20065 631 20099
rect 665 20065 703 20099
rect 737 20065 775 20099
rect -17 20031 775 20065
rect 17 19997 55 20031
rect 89 19997 127 20031
rect 161 19997 199 20031
rect 233 19997 271 20031
rect 305 19997 343 20031
rect 377 19997 415 20031
rect 449 19997 487 20031
rect 521 19997 559 20031
rect 593 19997 631 20031
rect 665 19997 703 20031
rect 737 19997 775 20031
rect -17 19963 775 19997
rect 17 19929 55 19963
rect 89 19929 127 19963
rect 161 19929 199 19963
rect 233 19929 271 19963
rect 305 19929 343 19963
rect 377 19929 415 19963
rect 449 19929 487 19963
rect 521 19929 559 19963
rect 593 19929 631 19963
rect 665 19929 703 19963
rect 737 19929 775 19963
rect -17 19895 775 19929
rect 17 19861 55 19895
rect 89 19861 127 19895
rect 161 19861 199 19895
rect 233 19861 271 19895
rect 305 19861 343 19895
rect 377 19861 415 19895
rect 449 19861 487 19895
rect 521 19861 559 19895
rect 593 19861 631 19895
rect 665 19861 703 19895
rect 737 19861 775 19895
rect -17 19827 775 19861
rect 17 19793 55 19827
rect 89 19793 127 19827
rect 161 19793 199 19827
rect 233 19793 271 19827
rect 305 19793 343 19827
rect 377 19793 415 19827
rect 449 19793 487 19827
rect 521 19793 559 19827
rect 593 19793 631 19827
rect 665 19793 703 19827
rect 737 19793 775 19827
rect -17 19759 775 19793
rect 17 19725 55 19759
rect 89 19725 127 19759
rect 161 19725 199 19759
rect 233 19725 271 19759
rect 305 19725 343 19759
rect 377 19725 415 19759
rect 449 19725 487 19759
rect 521 19725 559 19759
rect 593 19725 631 19759
rect 665 19725 703 19759
rect 737 19725 775 19759
rect -17 19691 775 19725
rect 17 19657 55 19691
rect 89 19657 127 19691
rect 161 19657 199 19691
rect 233 19657 271 19691
rect 305 19657 343 19691
rect 377 19657 415 19691
rect 449 19657 487 19691
rect 521 19657 559 19691
rect 593 19657 631 19691
rect 665 19657 703 19691
rect 737 19657 775 19691
rect -17 19623 775 19657
rect 17 19589 55 19623
rect 89 19589 127 19623
rect 161 19589 199 19623
rect 233 19589 271 19623
rect 305 19589 343 19623
rect 377 19589 415 19623
rect 449 19589 487 19623
rect 521 19589 559 19623
rect 593 19589 631 19623
rect 665 19589 703 19623
rect 737 19589 775 19623
rect -17 19555 775 19589
rect 17 19521 55 19555
rect 89 19521 127 19555
rect 161 19521 199 19555
rect 233 19521 271 19555
rect 305 19521 343 19555
rect 377 19521 415 19555
rect 449 19521 487 19555
rect 521 19521 559 19555
rect 593 19521 631 19555
rect 665 19521 703 19555
rect 737 19521 775 19555
rect -17 19487 775 19521
rect 17 19453 55 19487
rect 89 19453 127 19487
rect 161 19453 199 19487
rect 233 19453 271 19487
rect 305 19453 343 19487
rect 377 19453 415 19487
rect 449 19453 487 19487
rect 521 19453 559 19487
rect 593 19453 631 19487
rect 665 19453 703 19487
rect 737 19453 775 19487
rect -17 19419 775 19453
rect 17 19385 55 19419
rect 89 19385 127 19419
rect 161 19385 199 19419
rect 233 19385 271 19419
rect 305 19385 343 19419
rect 377 19385 415 19419
rect 449 19385 487 19419
rect 521 19385 559 19419
rect 593 19385 631 19419
rect 665 19385 703 19419
rect 737 19385 775 19419
rect -17 19351 775 19385
rect 17 19317 55 19351
rect 89 19317 127 19351
rect 161 19317 199 19351
rect 233 19317 271 19351
rect 305 19317 343 19351
rect 377 19317 415 19351
rect 449 19317 487 19351
rect 521 19317 559 19351
rect 593 19317 631 19351
rect 665 19317 703 19351
rect 737 19317 775 19351
rect -17 19283 775 19317
rect 17 19249 55 19283
rect 89 19249 127 19283
rect 161 19249 199 19283
rect 233 19249 271 19283
rect 305 19249 343 19283
rect 377 19249 415 19283
rect 449 19249 487 19283
rect 521 19249 559 19283
rect 593 19249 631 19283
rect 665 19249 703 19283
rect 737 19249 775 19283
rect -17 19215 775 19249
rect 17 19181 55 19215
rect 89 19181 127 19215
rect 161 19181 199 19215
rect 233 19181 271 19215
rect 305 19181 343 19215
rect 377 19181 415 19215
rect 449 19181 487 19215
rect 521 19181 559 19215
rect 593 19181 631 19215
rect 665 19181 703 19215
rect 737 19181 775 19215
rect -17 19147 775 19181
rect 17 19113 55 19147
rect 89 19113 127 19147
rect 161 19113 199 19147
rect 233 19113 271 19147
rect 305 19113 343 19147
rect 377 19113 415 19147
rect 449 19113 487 19147
rect 521 19113 559 19147
rect 593 19113 631 19147
rect 665 19113 703 19147
rect 737 19113 775 19147
rect -17 19079 775 19113
rect 17 19045 55 19079
rect 89 19045 127 19079
rect 161 19045 199 19079
rect 233 19045 271 19079
rect 305 19045 343 19079
rect 377 19045 415 19079
rect 449 19045 487 19079
rect 521 19045 559 19079
rect 593 19045 631 19079
rect 665 19045 703 19079
rect 737 19045 775 19079
rect -17 19011 775 19045
rect 17 18977 55 19011
rect 89 18977 127 19011
rect 161 18977 199 19011
rect 233 18977 271 19011
rect 305 18977 343 19011
rect 377 18977 415 19011
rect 449 18977 487 19011
rect 521 18977 559 19011
rect 593 18977 631 19011
rect 665 18977 703 19011
rect 737 18977 775 19011
rect -17 18943 775 18977
rect 17 18909 55 18943
rect 89 18909 127 18943
rect 161 18909 199 18943
rect 233 18909 271 18943
rect 305 18909 343 18943
rect 377 18909 415 18943
rect 449 18909 487 18943
rect 521 18909 559 18943
rect 593 18909 631 18943
rect 665 18909 703 18943
rect 737 18909 775 18943
rect -17 18875 775 18909
rect 17 18841 55 18875
rect 89 18841 127 18875
rect 161 18841 199 18875
rect 233 18841 271 18875
rect 305 18841 343 18875
rect 377 18841 415 18875
rect 449 18841 487 18875
rect 521 18841 559 18875
rect 593 18841 631 18875
rect 665 18841 703 18875
rect 737 18841 775 18875
rect -17 18807 775 18841
rect 17 18773 55 18807
rect 89 18773 127 18807
rect 161 18773 199 18807
rect 233 18773 271 18807
rect 305 18773 343 18807
rect 377 18773 415 18807
rect 449 18773 487 18807
rect 521 18773 559 18807
rect 593 18773 631 18807
rect 665 18773 703 18807
rect 737 18773 775 18807
rect -17 18739 775 18773
rect 17 18705 55 18739
rect 89 18705 127 18739
rect 161 18705 199 18739
rect 233 18705 271 18739
rect 305 18705 343 18739
rect 377 18705 415 18739
rect 449 18705 487 18739
rect 521 18705 559 18739
rect 593 18705 631 18739
rect 665 18705 703 18739
rect 737 18705 775 18739
rect -17 18671 775 18705
rect 17 18637 55 18671
rect 89 18637 127 18671
rect 161 18637 199 18671
rect 233 18637 271 18671
rect 305 18637 343 18671
rect 377 18637 415 18671
rect 449 18637 487 18671
rect 521 18637 559 18671
rect 593 18637 631 18671
rect 665 18637 703 18671
rect 737 18637 775 18671
rect 877 20381 915 20415
rect 949 20381 983 20415
rect 877 20347 983 20381
rect 877 20313 915 20347
rect 949 20313 983 20347
rect 877 20279 983 20313
rect 877 20245 915 20279
rect 949 20245 983 20279
rect 877 20211 983 20245
rect 877 20177 915 20211
rect 949 20177 983 20211
rect 877 20143 983 20177
rect 877 20109 915 20143
rect 949 20109 983 20143
rect 877 20075 983 20109
rect 877 20041 915 20075
rect 949 20041 983 20075
rect 877 20007 983 20041
rect 877 19973 915 20007
rect 949 19973 983 20007
rect 877 19939 983 19973
rect 877 19905 915 19939
rect 949 19905 983 19939
rect 877 19871 983 19905
rect 877 19837 915 19871
rect 949 19837 983 19871
rect 877 19803 983 19837
rect 877 19769 915 19803
rect 949 19769 983 19803
rect 877 19735 983 19769
rect 877 19701 915 19735
rect 949 19701 983 19735
rect 877 19667 983 19701
rect 877 19633 915 19667
rect 949 19633 983 19667
rect 877 19599 983 19633
rect 877 19565 915 19599
rect 949 19565 983 19599
rect 877 19531 983 19565
rect 877 19497 915 19531
rect 949 19497 983 19531
rect 877 19463 983 19497
rect 877 19429 915 19463
rect 949 19429 983 19463
rect 877 19395 983 19429
rect 877 19361 915 19395
rect 949 19361 983 19395
rect 877 19327 983 19361
rect 877 19293 915 19327
rect 949 19293 983 19327
rect 877 19259 983 19293
rect 877 19225 915 19259
rect 949 19225 983 19259
rect 877 19191 983 19225
rect 7937 19191 9142 19217
rect -17 18613 843 18637
rect 877 18613 915 19191
rect 949 19179 1718 19191
rect 1774 19179 9142 19191
rect 949 19157 9142 19179
rect 1017 19123 1058 19157
rect 1092 19123 1133 19157
rect 1167 19123 1208 19157
rect 1242 19123 1283 19157
rect 1317 19123 1358 19157
rect 1392 19123 1433 19157
rect 1467 19123 1508 19157
rect 1542 19123 1583 19157
rect 1617 19123 1658 19157
rect 1692 19153 9142 19157
rect 1692 19123 1729 19153
rect 1017 19119 1729 19123
rect 1763 19138 9142 19153
rect 1763 19119 1800 19138
rect 1017 19104 1800 19119
rect 1834 19104 1869 19138
rect 1903 19104 1938 19138
rect 1972 19104 2007 19138
rect 2041 19104 2076 19138
rect 2110 19104 2145 19138
rect 2179 19104 2214 19138
rect 2248 19104 2283 19138
rect 2317 19104 2352 19138
rect 2386 19104 2421 19138
rect 2455 19104 2490 19138
rect 2524 19104 2559 19138
rect 2593 19104 2628 19138
rect 2662 19104 2697 19138
rect 2731 19104 2766 19138
rect 2800 19104 2835 19138
rect 2869 19104 2904 19138
rect 2938 19104 2973 19138
rect 3007 19104 3042 19138
rect 3076 19104 3111 19138
rect 3145 19104 3180 19138
rect 3214 19104 3249 19138
rect 3283 19104 3318 19138
rect 3352 19104 3387 19138
rect 3421 19104 3456 19138
rect 3490 19104 3525 19138
rect 3559 19104 3594 19138
rect 3628 19104 3663 19138
rect 3697 19104 3732 19138
rect 3766 19104 3801 19138
rect 3835 19104 3870 19138
rect 3904 19104 3939 19138
rect 3973 19104 4008 19138
rect 4042 19104 4076 19138
rect 4110 19104 4144 19138
rect 4178 19104 4212 19138
rect 4246 19104 4280 19138
rect 4314 19104 4348 19138
rect 4382 19104 4416 19138
rect 4450 19104 4484 19138
rect 4518 19104 4552 19138
rect 4586 19104 4620 19138
rect 4654 19104 4688 19138
rect 4722 19104 4756 19138
rect 4790 19104 4824 19138
rect 4858 19104 4892 19138
rect 4926 19104 4960 19138
rect 4994 19104 5028 19138
rect 5062 19104 5096 19138
rect 5130 19104 5164 19138
rect 5198 19104 5232 19138
rect 5266 19104 5300 19138
rect 5334 19104 5368 19138
rect 5402 19104 5436 19138
rect 5470 19104 5504 19138
rect 5538 19104 5572 19138
rect 5606 19104 5640 19138
rect 5674 19104 5708 19138
rect 5742 19104 5776 19138
rect 5810 19104 5844 19138
rect 5878 19104 5912 19138
rect 5946 19104 5980 19138
rect 6014 19104 6048 19138
rect 6082 19104 6116 19138
rect 6150 19104 6184 19138
rect 6218 19104 6252 19138
rect 6286 19104 6320 19138
rect 6354 19104 6388 19138
rect 6422 19104 6456 19138
rect 6490 19104 6524 19138
rect 6558 19104 6592 19138
rect 6626 19104 6660 19138
rect 6694 19104 6728 19138
rect 6762 19104 6796 19138
rect 6830 19104 6864 19138
rect 6898 19104 6932 19138
rect 6966 19104 7000 19138
rect 7034 19104 7068 19138
rect 7102 19104 7136 19138
rect 7170 19104 7204 19138
rect 7238 19104 7272 19138
rect 7306 19104 7340 19138
rect 7374 19104 7408 19138
rect 7442 19104 7476 19138
rect 7510 19104 7544 19138
rect 7578 19104 7612 19138
rect 7646 19104 7680 19138
rect 7714 19104 7748 19138
rect 7782 19104 7816 19138
rect 7850 19104 7884 19138
rect 7918 19104 7952 19138
rect 7986 19104 8020 19138
rect 8054 19104 8088 19138
rect 8122 19104 8156 19138
rect 8190 19104 8224 19138
rect 8258 19104 8292 19138
rect 8326 19104 8360 19138
rect 8394 19104 8428 19138
rect 8462 19104 8496 19138
rect 8530 19104 8564 19138
rect 8598 19104 8632 19138
rect 8666 19104 8700 19138
rect 8734 19104 8768 19138
rect 8802 19104 8836 19138
rect 8870 19104 8904 19138
rect 8938 19104 8972 19138
rect 9006 19104 9040 19138
rect 9074 19104 9108 19138
rect 1017 19089 9142 19104
rect 1017 19055 1058 19089
rect 1092 19055 1133 19089
rect 1167 19055 1208 19089
rect 1242 19055 1283 19089
rect 1317 19055 1358 19089
rect 1392 19055 1433 19089
rect 1467 19055 1508 19089
rect 1542 19055 1583 19089
rect 1617 19055 1658 19089
rect 1692 19081 9142 19089
rect 1692 19055 1729 19081
rect 1017 19047 1729 19055
rect 1763 19051 9142 19081
rect 1763 19047 1800 19051
rect 1017 19021 1800 19047
rect 5772 19025 9142 19051
rect 1017 18987 1058 19021
rect 1092 18987 1133 19021
rect 1167 18987 1208 19021
rect 1242 18987 1283 19021
rect 1317 18987 1358 19021
rect 1392 18987 1433 19021
rect 1467 18987 1508 19021
rect 1542 18987 1583 19021
rect 1617 18987 1658 19021
rect 1692 19009 1800 19021
rect 1692 18987 1729 19009
rect 1017 18975 1729 18987
rect 1763 18975 1800 19009
rect 1017 18953 1800 18975
rect 1017 18919 1058 18953
rect 1092 18919 1133 18953
rect 1167 18919 1208 18953
rect 1242 18919 1283 18953
rect 1317 18919 1358 18953
rect 1392 18919 1433 18953
rect 1467 18919 1508 18953
rect 1542 18919 1583 18953
rect 1617 18919 1658 18953
rect 1692 18937 1800 18953
rect 1692 18919 1729 18937
rect 1017 18903 1729 18919
rect 1763 18903 1800 18937
rect 1017 18885 1800 18903
rect 1017 18851 1058 18885
rect 1092 18851 1133 18885
rect 1167 18851 1208 18885
rect 1242 18851 1283 18885
rect 1317 18851 1358 18885
rect 1392 18851 1433 18885
rect 1467 18851 1508 18885
rect 1542 18851 1583 18885
rect 1617 18851 1658 18885
rect 1692 18865 1800 18885
rect 1692 18851 1729 18865
rect 1017 18831 1729 18851
rect 1763 18831 1800 18865
rect 1017 18817 1800 18831
rect 1017 18783 1058 18817
rect 1092 18783 1133 18817
rect 1167 18783 1208 18817
rect 1242 18783 1283 18817
rect 1317 18783 1358 18817
rect 1392 18783 1433 18817
rect 1467 18783 1508 18817
rect 1542 18783 1583 18817
rect 1617 18783 1658 18817
rect 1692 18793 1800 18817
rect 1692 18783 1729 18793
rect 1017 18759 1729 18783
rect 1763 18759 1800 18793
rect 1017 18749 1800 18759
rect 1017 18715 1058 18749
rect 1092 18715 1133 18749
rect 1167 18715 1208 18749
rect 1242 18715 1283 18749
rect 1317 18715 1358 18749
rect 1392 18715 1433 18749
rect 1467 18715 1508 18749
rect 1542 18715 1583 18749
rect 1617 18715 1658 18749
rect 1692 18720 1800 18749
rect 1692 18715 1729 18720
rect 1017 18686 1729 18715
rect 1763 18686 1800 18720
rect 1017 18681 1800 18686
rect 1017 18647 1058 18681
rect 1092 18647 1133 18681
rect 1167 18647 1208 18681
rect 1242 18647 1283 18681
rect 1317 18647 1358 18681
rect 1392 18647 1433 18681
rect 1467 18647 1508 18681
rect 1542 18647 1583 18681
rect 1617 18647 1658 18681
rect 1692 18647 1800 18681
rect 949 18613 1729 18647
rect 1763 18613 1800 18647
rect 1298 18577 1800 18613
rect 1298 18543 1332 18577
rect 1366 18543 1412 18577
rect 1446 18543 1492 18577
rect 1526 18543 1572 18577
rect 1606 18543 1652 18577
rect 1686 18543 1732 18577
rect 1766 18543 1800 18577
rect 1298 18509 1800 18543
rect 1298 18475 1332 18509
rect 1366 18475 1412 18509
rect 1446 18475 1492 18509
rect 1526 18475 1572 18509
rect 1606 18475 1652 18509
rect 1686 18475 1732 18509
rect 1766 18475 1800 18509
rect 1298 18441 1800 18475
rect 1298 18407 1332 18441
rect 1366 18407 1412 18441
rect 1446 18407 1492 18441
rect 1526 18407 1572 18441
rect 1606 18407 1652 18441
rect 1686 18407 1732 18441
rect 1766 18407 1800 18441
rect 1298 18373 1800 18407
rect 1298 18339 1332 18373
rect 1366 18339 1412 18373
rect 1446 18339 1492 18373
rect 1526 18339 1572 18373
rect 1606 18339 1652 18373
rect 1686 18339 1732 18373
rect 1766 18339 1800 18373
rect 1298 18305 1800 18339
rect 1298 18271 1332 18305
rect 1366 18271 1412 18305
rect 1446 18271 1492 18305
rect 1526 18271 1572 18305
rect 1606 18271 1652 18305
rect 1686 18271 1732 18305
rect 1766 18271 1800 18305
rect 1298 18237 1800 18271
rect 1298 18203 1332 18237
rect 1366 18203 1412 18237
rect 1446 18203 1492 18237
rect 1526 18203 1572 18237
rect 1606 18203 1652 18237
rect 1686 18203 1732 18237
rect 1766 18203 1800 18237
rect 1298 18169 1800 18203
rect 1298 18135 1332 18169
rect 1366 18135 1412 18169
rect 1446 18135 1492 18169
rect 1526 18135 1572 18169
rect 1606 18135 1652 18169
rect 1686 18135 1732 18169
rect 1766 18135 1800 18169
rect 1298 18100 1800 18135
rect 1298 18066 1332 18100
rect 1366 18066 1412 18100
rect 1446 18066 1492 18100
rect 1526 18066 1572 18100
rect 1606 18066 1652 18100
rect 1686 18066 1732 18100
rect 1766 18066 1800 18100
rect 1298 18031 1800 18066
rect 1298 17997 1332 18031
rect 1366 17997 1412 18031
rect 1446 17997 1492 18031
rect 1526 17997 1572 18031
rect 1606 17997 1652 18031
rect 1686 17997 1732 18031
rect 1766 17997 1800 18031
rect 1298 17962 1800 17997
rect 1298 17928 1332 17962
rect 1366 17928 1412 17962
rect 1446 17928 1492 17962
rect 1526 17928 1572 17962
rect 1606 17928 1652 17962
rect 1686 17928 1732 17962
rect 1766 17928 1800 17962
rect 1298 17893 1800 17928
rect 1298 17859 1332 17893
rect 1366 17859 1412 17893
rect 1446 17859 1492 17893
rect 1526 17859 1572 17893
rect 1606 17859 1652 17893
rect 1686 17859 1732 17893
rect 1766 17859 1800 17893
rect 1298 17824 1800 17859
rect 1298 17790 1332 17824
rect 1366 17790 1412 17824
rect 1446 17790 1492 17824
rect 1526 17790 1572 17824
rect 1606 17790 1652 17824
rect 1686 17790 1732 17824
rect 1766 17790 1800 17824
rect 338 9109 362 9143
rect 396 9109 433 9143
rect 467 9109 504 9143
rect 538 9109 575 9143
rect 609 9109 646 9143
rect 680 9109 717 9143
rect 751 9109 788 9143
rect 822 9109 859 9143
rect 893 9109 917 9143
rect 13933 2251 14330 2285
rect 13967 2217 14006 2251
rect 14040 2217 14079 2251
rect 14113 2217 14152 2251
rect 14186 2217 14224 2251
rect 14258 2217 14296 2251
rect 13933 2173 14330 2217
rect 13967 2139 14006 2173
rect 14040 2139 14079 2173
rect 14113 2139 14152 2173
rect 14186 2139 14224 2173
rect 14258 2139 14296 2173
rect 13933 2095 14330 2139
rect 13967 2061 14006 2095
rect 14040 2061 14079 2095
rect 14113 2061 14152 2095
rect 14186 2061 14224 2095
rect 14258 2061 14296 2095
rect 13933 2037 14330 2061
rect 13278 2003 13312 2037
rect 13346 2003 13382 2037
rect 13416 2003 13451 2037
rect 13485 2003 13520 2037
rect 13554 2003 13589 2037
rect 13623 2003 13658 2037
rect 13692 2003 13727 2037
rect 13761 2003 13796 2037
rect 13830 2003 13865 2037
rect 13899 2017 14330 2037
rect 13899 2003 13933 2017
rect 13278 1983 13933 2003
rect 13967 1983 14006 2017
rect 14040 1983 14079 2017
rect 14113 1983 14152 2017
rect 14186 1983 14224 2017
rect 14258 1983 14296 2017
rect 13278 1949 14330 1983
rect 13278 1915 13312 1949
rect 13346 1915 13382 1949
rect 13416 1915 13451 1949
rect 13485 1915 13520 1949
rect 13554 1915 13589 1949
rect 13623 1915 13658 1949
rect 13692 1915 13727 1949
rect 13761 1915 13796 1949
rect 13830 1915 13865 1949
rect 13899 1915 13933 1949
rect 13278 1914 13420 1915
rect 13132 1880 13420 1914
rect 13132 1846 13133 1880
rect 13167 1846 13217 1880
rect 13251 1846 13301 1880
rect 13335 1846 13385 1880
rect 13419 1846 13420 1880
rect 13132 1810 13420 1846
rect 13132 1776 13133 1810
rect 13167 1776 13217 1810
rect 13251 1776 13301 1810
rect 13335 1776 13385 1810
rect 13419 1776 13420 1810
rect 13132 1740 13420 1776
rect 13132 1706 13133 1740
rect 13167 1706 13217 1740
rect 13251 1706 13301 1740
rect 13335 1706 13385 1740
rect 13419 1706 13420 1740
rect 13132 1669 13420 1706
rect 13132 1635 13133 1669
rect 13167 1635 13217 1669
rect 13251 1635 13301 1669
rect 13335 1635 13385 1669
rect 13419 1635 13420 1669
rect 13132 1598 13420 1635
rect 13132 1564 13133 1598
rect 13167 1564 13217 1598
rect 13251 1564 13301 1598
rect 13335 1564 13385 1598
rect 13419 1564 13420 1598
rect 13132 1527 13420 1564
rect 13132 1493 13133 1527
rect 13167 1493 13217 1527
rect 13251 1493 13301 1527
rect 13335 1493 13385 1527
rect 13419 1493 13420 1527
rect 13132 1456 13420 1493
rect 13132 1422 13133 1456
rect 13167 1422 13217 1456
rect 13251 1422 13301 1456
rect 13335 1422 13385 1456
rect 13419 1422 13420 1456
rect 13132 1385 13420 1422
rect 13132 1351 13133 1385
rect 13167 1351 13217 1385
rect 13251 1351 13301 1385
rect 13335 1351 13385 1385
rect 13419 1351 13420 1385
rect 13132 1314 13420 1351
rect 13132 1280 13133 1314
rect 13167 1280 13217 1314
rect 13251 1280 13301 1314
rect 13335 1280 13385 1314
rect 13419 1280 13420 1314
rect 13132 1246 13420 1280
rect 1561 1212 12298 1246
rect 12332 1212 12369 1246
rect 12403 1212 12440 1246
rect 12474 1212 12511 1246
rect 12545 1212 12582 1246
rect 12616 1212 12653 1246
rect 12687 1212 12724 1246
rect 12758 1212 12795 1246
rect 12829 1212 12866 1246
rect 12900 1212 12937 1246
rect 12971 1212 13008 1246
rect 13042 1212 13079 1246
rect 13113 1212 13150 1246
rect 13184 1212 13221 1246
rect 13255 1212 13292 1246
rect 13326 1212 13362 1246
rect 13396 1212 13420 1246
rect 1561 1180 13420 1212
rect 1595 1146 1630 1180
rect 1664 1146 1699 1180
rect 1733 1146 1768 1180
rect 1802 1146 1837 1180
rect 1871 1146 1906 1180
rect 1940 1146 1975 1180
rect 2009 1146 2044 1180
rect 2078 1146 2113 1180
rect 2147 1146 2182 1180
rect 2216 1146 2251 1180
rect 2285 1146 2320 1180
rect 2354 1146 2389 1180
rect 2423 1146 2458 1180
rect 2492 1146 2527 1180
rect 2561 1146 2596 1180
rect 2630 1146 2665 1180
rect 2699 1146 2734 1180
rect 2768 1146 2803 1180
rect 2837 1146 2872 1180
rect 2906 1146 2941 1180
rect 2975 1146 3009 1180
rect 3043 1146 3077 1180
rect 3111 1146 3145 1180
rect 3179 1146 3213 1180
rect 3247 1146 3281 1180
rect 3315 1146 3349 1180
rect 3383 1146 3417 1180
rect 3451 1146 3485 1180
rect 3519 1146 3553 1180
rect 3587 1146 3621 1180
rect 3655 1146 3689 1180
rect 3723 1146 3757 1180
rect 3791 1146 3825 1180
rect 3859 1146 3893 1180
rect 3927 1146 3961 1180
rect 3995 1146 4029 1180
rect 4063 1146 4097 1180
rect 4131 1146 4165 1180
rect 4199 1146 4233 1180
rect 4267 1146 4301 1180
rect 4335 1146 4369 1180
rect 4403 1146 4437 1180
rect 4471 1146 4505 1180
rect 4539 1146 4573 1180
rect 4607 1146 4641 1180
rect 4675 1146 4709 1180
rect 4743 1146 4777 1180
rect 4811 1146 4845 1180
rect 4879 1146 4913 1180
rect 4947 1146 4981 1180
rect 5015 1146 5049 1180
rect 5083 1146 5117 1180
rect 5151 1146 5185 1180
rect 5219 1146 5253 1180
rect 5287 1146 5321 1180
rect 5355 1146 5389 1180
rect 5423 1146 5457 1180
rect 5491 1146 5525 1180
rect 5559 1146 5593 1180
rect 5627 1146 5661 1180
rect 5695 1146 5729 1180
rect 5763 1146 5797 1180
rect 5831 1146 5865 1180
rect 5899 1146 5933 1180
rect 5967 1146 6001 1180
rect 6035 1146 6069 1180
rect 6103 1146 6137 1180
rect 6171 1146 6205 1180
rect 6239 1146 6273 1180
rect 6307 1146 6341 1180
rect 6375 1146 6409 1180
rect 6443 1146 6477 1180
rect 6511 1146 6545 1180
rect 6579 1146 6613 1180
rect 6647 1146 6681 1180
rect 6715 1146 6749 1180
rect 6783 1146 6817 1180
rect 6851 1146 6885 1180
rect 6919 1146 6953 1180
rect 6987 1146 7021 1180
rect 7055 1146 7089 1180
rect 7123 1146 7157 1180
rect 7191 1146 7225 1180
rect 7259 1146 7293 1180
rect 7327 1146 7361 1180
rect 7395 1146 7429 1180
rect 7463 1146 7497 1180
rect 7531 1146 7565 1180
rect 7599 1146 7633 1180
rect 7667 1146 7701 1180
rect 7735 1146 7769 1180
rect 7803 1146 7837 1180
rect 7871 1146 7905 1180
rect 7939 1146 7973 1180
rect 8007 1146 8041 1180
rect 8075 1146 8109 1180
rect 8143 1146 8177 1180
rect 8211 1146 8245 1180
rect 8279 1146 8313 1180
rect 8347 1146 8381 1180
rect 8415 1146 8449 1180
rect 8483 1146 8517 1180
rect 8551 1146 8585 1180
rect 8619 1146 8653 1180
rect 8687 1146 8721 1180
rect 8755 1146 8789 1180
rect 8823 1146 8857 1180
rect 8891 1146 8925 1180
rect 8959 1146 8993 1180
rect 9027 1146 9061 1180
rect 9095 1146 9129 1180
rect 9163 1146 9197 1180
rect 9231 1146 9265 1180
rect 9299 1146 9333 1180
rect 9367 1146 9401 1180
rect 9435 1146 9469 1180
rect 9503 1146 9537 1180
rect 9571 1146 9605 1180
rect 9639 1146 9673 1180
rect 9707 1146 9741 1180
rect 9775 1146 9809 1180
rect 9843 1146 9877 1180
rect 9911 1146 9945 1180
rect 9979 1146 10013 1180
rect 10047 1146 10081 1180
rect 10115 1146 10149 1180
rect 10183 1146 10217 1180
rect 10251 1146 10285 1180
rect 10319 1146 10353 1180
rect 10387 1146 10421 1180
rect 10455 1146 10489 1180
rect 10523 1146 10557 1180
rect 10591 1146 10625 1180
rect 10659 1146 10693 1180
rect 10727 1146 10761 1180
rect 10795 1146 10829 1180
rect 10863 1146 10897 1180
rect 10931 1146 10965 1180
rect 10999 1146 11033 1180
rect 11067 1146 11101 1180
rect 11135 1146 11169 1180
rect 11203 1146 11237 1180
rect 11271 1146 11305 1180
rect 11339 1146 11373 1180
rect 11407 1146 11441 1180
rect 11475 1146 11509 1180
rect 11543 1146 11577 1180
rect 11611 1146 11645 1180
rect 11679 1146 11713 1180
rect 11747 1146 11781 1180
rect 11815 1146 11849 1180
rect 11883 1146 11917 1180
rect 11951 1146 11985 1180
rect 12019 1146 12053 1180
rect 12087 1146 12121 1180
rect 12155 1146 12189 1180
rect 12223 1148 13420 1180
rect 12223 1146 12298 1148
rect 1561 1114 12298 1146
rect 12332 1114 12369 1148
rect 12403 1114 12440 1148
rect 12474 1114 12511 1148
rect 12545 1114 12582 1148
rect 12616 1114 12653 1148
rect 12687 1114 12724 1148
rect 12758 1114 12795 1148
rect 12829 1114 12866 1148
rect 12900 1114 12937 1148
rect 12971 1114 13008 1148
rect 13042 1114 13079 1148
rect 13113 1114 13150 1148
rect 13184 1114 13221 1148
rect 13255 1114 13292 1148
rect 13326 1114 13362 1148
rect 13396 1114 13420 1148
rect 1561 1080 13420 1114
rect 12223 1054 13420 1080
rect 12248 1050 13420 1054
rect 12248 1046 12298 1050
rect 12274 1016 12298 1046
rect 12332 1016 12369 1050
rect 12403 1016 12440 1050
rect 12474 1016 12511 1050
rect 12545 1016 12582 1050
rect 12616 1016 12653 1050
rect 12687 1016 12724 1050
rect 12758 1016 12795 1050
rect 12829 1016 12866 1050
rect 12900 1016 12937 1050
rect 12971 1016 13008 1050
rect 13042 1016 13079 1050
rect 13113 1016 13150 1050
rect 13184 1016 13221 1050
rect 13255 1016 13292 1050
rect 13326 1016 13362 1050
rect 13396 1016 13420 1050
<< mvnsubdiff >>
rect -17 35705 843 35729
rect 17 35671 55 35705
rect 89 35671 127 35705
rect 161 35671 199 35705
rect 233 35671 271 35705
rect 305 35671 343 35705
rect 377 35671 415 35705
rect 449 35671 487 35705
rect 521 35671 559 35705
rect 593 35671 631 35705
rect 665 35671 703 35705
rect 737 35671 775 35705
rect 809 35695 843 35705
rect 877 35695 915 35729
rect 949 35695 983 35729
rect 809 35671 983 35695
rect -17 35645 983 35671
rect -17 35637 843 35645
rect 17 35603 55 35637
rect 89 35603 127 35637
rect 161 35603 199 35637
rect 233 35603 271 35637
rect 305 35603 343 35637
rect 377 35603 415 35637
rect 449 35603 487 35637
rect 521 35603 559 35637
rect 593 35603 631 35637
rect 665 35603 703 35637
rect 737 35603 775 35637
rect 809 35611 843 35637
rect 877 35611 915 35645
rect 949 35611 983 35645
rect 809 35603 983 35611
rect -17 35569 983 35603
rect 17 35535 55 35569
rect 89 35535 127 35569
rect 161 35535 199 35569
rect 233 35535 271 35569
rect 305 35535 343 35569
rect 377 35535 415 35569
rect 449 35535 487 35569
rect 521 35535 559 35569
rect 593 35535 631 35569
rect 665 35535 703 35569
rect 737 35535 775 35569
rect 809 35561 983 35569
rect 809 35535 843 35561
rect -17 35527 843 35535
rect 877 35527 915 35561
rect 949 35527 983 35561
rect -17 35501 983 35527
rect 17 35467 55 35501
rect 89 35467 127 35501
rect 161 35467 199 35501
rect 233 35467 271 35501
rect 305 35467 343 35501
rect 377 35467 415 35501
rect 449 35467 487 35501
rect 521 35467 559 35501
rect 593 35467 631 35501
rect 665 35467 703 35501
rect 737 35467 775 35501
rect 809 35477 983 35501
rect 809 35467 843 35477
rect -17 35443 843 35467
rect 877 35443 915 35477
rect 949 35443 983 35477
rect -17 35433 983 35443
rect 17 35399 55 35433
rect 89 35399 127 35433
rect 161 35399 199 35433
rect 233 35399 271 35433
rect 305 35399 343 35433
rect 377 35399 415 35433
rect 449 35399 487 35433
rect 521 35399 559 35433
rect 593 35399 631 35433
rect 665 35399 703 35433
rect 737 35399 775 35433
rect 809 35399 983 35433
rect -17 35393 983 35399
rect -17 35365 843 35393
rect 17 35331 55 35365
rect 89 35331 127 35365
rect 161 35331 199 35365
rect 233 35331 271 35365
rect 305 35331 343 35365
rect 377 35331 415 35365
rect 449 35331 487 35365
rect 521 35331 559 35365
rect 593 35331 631 35365
rect 665 35331 703 35365
rect 737 35331 775 35365
rect 809 35359 843 35365
rect 877 35359 915 35393
rect 949 35359 983 35393
rect 809 35331 983 35359
rect -17 35309 983 35331
rect -17 35297 843 35309
rect 17 35263 55 35297
rect 89 35263 127 35297
rect 161 35263 199 35297
rect 233 35263 271 35297
rect 305 35263 343 35297
rect 377 35263 415 35297
rect 449 35263 487 35297
rect 521 35263 559 35297
rect 593 35263 631 35297
rect 665 35263 703 35297
rect 737 35263 775 35297
rect 809 35275 843 35297
rect 877 35275 915 35309
rect 949 35275 983 35309
rect 809 35263 983 35275
rect -17 35229 983 35263
rect 17 35195 55 35229
rect 89 35195 127 35229
rect 161 35195 199 35229
rect 233 35195 271 35229
rect 305 35195 343 35229
rect 377 35195 415 35229
rect 449 35195 487 35229
rect 521 35195 559 35229
rect 593 35195 631 35229
rect 665 35195 703 35229
rect 737 35195 775 35229
rect 809 35225 983 35229
rect 809 35195 843 35225
rect -17 35191 843 35195
rect 877 35191 915 35225
rect 949 35191 983 35225
rect -17 35161 983 35191
rect 17 35127 55 35161
rect 89 35127 127 35161
rect 161 35127 199 35161
rect 233 35127 271 35161
rect 305 35127 343 35161
rect 377 35127 415 35161
rect 449 35127 487 35161
rect 521 35127 559 35161
rect 593 35127 631 35161
rect 665 35127 703 35161
rect 737 35127 775 35161
rect 809 35141 983 35161
rect 809 35127 843 35141
rect -17 35107 843 35127
rect 877 35107 915 35141
rect 949 35107 983 35141
rect -17 35093 983 35107
rect 17 35059 55 35093
rect 89 35059 127 35093
rect 161 35059 199 35093
rect 233 35059 271 35093
rect 305 35059 343 35093
rect 377 35059 415 35093
rect 449 35059 487 35093
rect 521 35059 559 35093
rect 593 35059 631 35093
rect 665 35059 703 35093
rect 737 35059 775 35093
rect 809 35059 983 35093
rect -17 35057 983 35059
rect -17 35025 843 35057
rect 17 34991 55 35025
rect 89 34991 127 35025
rect 161 34991 199 35025
rect 233 34991 271 35025
rect 305 34991 343 35025
rect 377 34991 415 35025
rect 449 34991 487 35025
rect 521 34991 559 35025
rect 593 34991 631 35025
rect 665 34991 703 35025
rect 737 34991 775 35025
rect 809 35023 843 35025
rect 877 35023 915 35057
rect 949 35023 983 35057
rect 809 34991 983 35023
rect -17 34973 983 34991
rect -17 34957 843 34973
rect 17 34923 55 34957
rect 89 34923 127 34957
rect 161 34923 199 34957
rect 233 34923 271 34957
rect 305 34923 343 34957
rect 377 34923 415 34957
rect 449 34923 487 34957
rect 521 34923 559 34957
rect 593 34923 631 34957
rect 665 34923 703 34957
rect 737 34923 775 34957
rect 809 34939 843 34957
rect 877 34939 915 34973
rect 949 34939 983 34973
rect 809 34923 983 34939
rect -17 34889 983 34923
rect 17 34855 55 34889
rect 89 34855 127 34889
rect 161 34855 199 34889
rect 233 34855 271 34889
rect 305 34855 343 34889
rect 377 34855 415 34889
rect 449 34855 487 34889
rect 521 34855 559 34889
rect 593 34855 631 34889
rect 665 34855 703 34889
rect 737 34855 775 34889
rect 809 34855 843 34889
rect 877 34855 915 34889
rect 949 34855 983 34889
rect -17 34821 983 34855
rect 17 34787 55 34821
rect 89 34787 127 34821
rect 161 34787 199 34821
rect 233 34787 271 34821
rect 305 34787 343 34821
rect 377 34787 415 34821
rect 449 34787 487 34821
rect 521 34787 559 34821
rect 593 34787 631 34821
rect 665 34787 703 34821
rect 737 34787 775 34821
rect 809 34805 983 34821
rect 809 34787 843 34805
rect -17 34771 843 34787
rect 877 34771 915 34805
rect 949 34771 983 34805
rect -17 34753 983 34771
rect 17 34719 55 34753
rect 89 34719 127 34753
rect 161 34719 199 34753
rect 233 34719 271 34753
rect 305 34719 343 34753
rect 377 34719 415 34753
rect 449 34719 487 34753
rect 521 34719 559 34753
rect 593 34719 631 34753
rect 665 34719 703 34753
rect 737 34719 775 34753
rect 809 34721 983 34753
rect 809 34719 843 34721
rect -17 34687 843 34719
rect 877 34687 915 34721
rect 949 34687 983 34721
rect -17 34685 983 34687
rect 17 34651 55 34685
rect 89 34651 127 34685
rect 161 34651 199 34685
rect 233 34651 271 34685
rect 305 34651 343 34685
rect 377 34651 415 34685
rect 449 34651 487 34685
rect 521 34651 559 34685
rect 593 34651 631 34685
rect 665 34651 703 34685
rect 737 34651 775 34685
rect 809 34651 983 34685
rect -17 34637 983 34651
rect -17 34617 843 34637
rect 17 34583 55 34617
rect 89 34583 127 34617
rect 161 34583 199 34617
rect 233 34583 271 34617
rect 305 34583 343 34617
rect 377 34583 415 34617
rect 449 34583 487 34617
rect 521 34583 559 34617
rect 593 34583 631 34617
rect 665 34583 703 34617
rect 737 34583 775 34617
rect 809 34603 843 34617
rect 877 34603 915 34637
rect 949 34603 983 34637
rect 809 34583 983 34603
rect -17 34553 983 34583
rect -17 34549 843 34553
rect 17 34515 55 34549
rect 89 34515 127 34549
rect 161 34515 199 34549
rect 233 34515 271 34549
rect 305 34515 343 34549
rect 377 34515 415 34549
rect 449 34515 487 34549
rect 521 34515 559 34549
rect 593 34515 631 34549
rect 665 34515 703 34549
rect 737 34515 775 34549
rect 809 34519 843 34549
rect 877 34519 915 34553
rect 949 34519 983 34553
rect 809 34515 983 34519
rect -17 34481 983 34515
rect 17 34447 55 34481
rect 89 34447 127 34481
rect 161 34447 199 34481
rect 233 34447 271 34481
rect 305 34447 343 34481
rect 377 34447 415 34481
rect 449 34447 487 34481
rect 521 34447 559 34481
rect 593 34447 631 34481
rect 665 34447 703 34481
rect 737 34447 775 34481
rect 809 34469 983 34481
rect 809 34447 843 34469
rect -17 34435 843 34447
rect 877 34435 915 34469
rect 949 34435 983 34469
rect -17 34413 983 34435
rect 17 34379 55 34413
rect 89 34379 127 34413
rect 161 34379 199 34413
rect 233 34379 271 34413
rect 305 34379 343 34413
rect 377 34379 415 34413
rect 449 34379 487 34413
rect 521 34379 559 34413
rect 593 34379 631 34413
rect 665 34379 703 34413
rect 737 34379 775 34413
rect 809 34385 983 34413
rect 809 34379 843 34385
rect -17 34351 843 34379
rect 877 34351 915 34385
rect 949 34351 983 34385
rect -17 34345 983 34351
rect 17 34311 55 34345
rect 89 34311 127 34345
rect 161 34311 199 34345
rect 233 34311 271 34345
rect 305 34311 343 34345
rect 377 34311 415 34345
rect 449 34311 487 34345
rect 521 34311 559 34345
rect 593 34311 631 34345
rect 665 34311 703 34345
rect 737 34311 775 34345
rect 809 34311 983 34345
rect -17 34301 983 34311
rect -17 34277 843 34301
rect 17 34243 55 34277
rect 89 34243 127 34277
rect 161 34243 199 34277
rect 233 34243 271 34277
rect 305 34243 343 34277
rect 377 34243 415 34277
rect 449 34243 487 34277
rect 521 34243 559 34277
rect 593 34243 631 34277
rect 665 34243 703 34277
rect 737 34243 775 34277
rect 809 34267 843 34277
rect 877 34267 915 34301
rect 949 34267 983 34301
rect 809 34243 983 34267
rect -17 34217 983 34243
rect -17 34209 843 34217
rect 17 34175 55 34209
rect 89 34175 127 34209
rect 161 34175 199 34209
rect 233 34175 271 34209
rect 305 34175 343 34209
rect 377 34175 415 34209
rect 449 34175 487 34209
rect 521 34175 559 34209
rect 593 34175 631 34209
rect 665 34175 703 34209
rect 737 34175 775 34209
rect 809 34183 843 34209
rect 877 34183 915 34217
rect 949 34183 983 34217
rect 809 34175 983 34183
rect -17 34141 983 34175
rect 17 34107 55 34141
rect 89 34107 127 34141
rect 161 34107 199 34141
rect 233 34107 271 34141
rect 305 34107 343 34141
rect 377 34107 415 34141
rect 449 34107 487 34141
rect 521 34107 559 34141
rect 593 34107 631 34141
rect 665 34107 703 34141
rect 737 34107 775 34141
rect 809 34133 983 34141
rect 809 34107 843 34133
rect -17 34099 843 34107
rect 877 34099 915 34133
rect 949 34099 983 34133
rect -17 34073 983 34099
rect 17 34039 55 34073
rect 89 34039 127 34073
rect 161 34039 199 34073
rect 233 34039 271 34073
rect 305 34039 343 34073
rect 377 34039 415 34073
rect 449 34039 487 34073
rect 521 34039 559 34073
rect 593 34039 631 34073
rect 665 34039 703 34073
rect 737 34039 775 34073
rect 809 34049 983 34073
rect 809 34039 843 34049
rect -17 34015 843 34039
rect 877 34015 915 34049
rect 949 34015 983 34049
rect -17 34005 983 34015
rect 17 33971 55 34005
rect 89 33971 127 34005
rect 161 33971 199 34005
rect 233 33971 271 34005
rect 305 33971 343 34005
rect 377 33971 415 34005
rect 449 33971 487 34005
rect 521 33971 559 34005
rect 593 33971 631 34005
rect 665 33971 703 34005
rect 737 33971 775 34005
rect 809 33971 983 34005
rect -17 33965 983 33971
rect -17 33937 843 33965
rect 17 33903 55 33937
rect 89 33903 127 33937
rect 161 33903 199 33937
rect 233 33903 271 33937
rect 305 33903 343 33937
rect 377 33903 415 33937
rect 449 33903 487 33937
rect 521 33903 559 33937
rect 593 33903 631 33937
rect 665 33903 703 33937
rect 737 33903 775 33937
rect 809 33931 843 33937
rect 877 33931 915 33965
rect 949 33931 983 33965
rect 809 33903 983 33931
rect -17 33881 983 33903
rect -17 33869 843 33881
rect 17 33835 55 33869
rect 89 33835 127 33869
rect 161 33835 199 33869
rect 233 33835 271 33869
rect 305 33835 343 33869
rect 377 33835 415 33869
rect 449 33835 487 33869
rect 521 33835 559 33869
rect 593 33835 631 33869
rect 665 33835 703 33869
rect 737 33835 775 33869
rect 809 33847 843 33869
rect 877 33847 915 33881
rect 949 33847 983 33881
rect 809 33835 983 33847
rect -17 33801 983 33835
rect 17 33767 55 33801
rect 89 33767 127 33801
rect 161 33767 199 33801
rect 233 33767 271 33801
rect 305 33767 343 33801
rect 377 33767 415 33801
rect 449 33767 487 33801
rect 521 33767 559 33801
rect 593 33767 631 33801
rect 665 33767 703 33801
rect 737 33767 775 33801
rect 809 33797 983 33801
rect 809 33767 843 33797
rect -17 33763 843 33767
rect 877 33763 915 33797
rect 949 33763 983 33797
rect -17 33733 983 33763
rect 17 33699 55 33733
rect 89 33699 127 33733
rect 161 33699 199 33733
rect 233 33699 271 33733
rect 305 33699 343 33733
rect 377 33699 415 33733
rect 449 33699 487 33733
rect 521 33699 559 33733
rect 593 33699 631 33733
rect 665 33699 703 33733
rect 737 33699 775 33733
rect 809 33713 983 33733
rect 809 33699 843 33713
rect -17 33679 843 33699
rect 877 33679 915 33713
rect 949 33679 983 33713
rect -17 33665 983 33679
rect 17 33631 55 33665
rect 89 33631 127 33665
rect 161 33631 199 33665
rect 233 33631 271 33665
rect 305 33631 343 33665
rect 377 33631 415 33665
rect 449 33631 487 33665
rect 521 33631 559 33665
rect 593 33631 631 33665
rect 665 33631 703 33665
rect 737 33631 775 33665
rect 809 33631 983 33665
rect -17 33629 983 33631
rect -17 33597 843 33629
rect 17 33563 55 33597
rect 89 33563 127 33597
rect 161 33563 199 33597
rect 233 33563 271 33597
rect 305 33563 343 33597
rect 377 33563 415 33597
rect 449 33563 487 33597
rect 521 33563 559 33597
rect 593 33563 631 33597
rect 665 33563 703 33597
rect 737 33563 775 33597
rect 809 33595 843 33597
rect 877 33595 915 33629
rect 949 33595 983 33629
rect 809 33563 983 33595
rect -17 33545 983 33563
rect -17 33529 843 33545
rect 17 33495 55 33529
rect 89 33495 127 33529
rect 161 33495 199 33529
rect 233 33495 271 33529
rect 305 33495 343 33529
rect 377 33495 415 33529
rect 449 33495 487 33529
rect 521 33495 559 33529
rect 593 33495 631 33529
rect 665 33495 703 33529
rect 737 33495 775 33529
rect 809 33511 843 33529
rect 877 33511 915 33545
rect 949 33511 983 33545
rect 809 33495 983 33511
rect -17 33461 983 33495
rect 17 33427 55 33461
rect 89 33427 127 33461
rect 161 33427 199 33461
rect 233 33427 271 33461
rect 305 33427 343 33461
rect 377 33427 415 33461
rect 449 33427 487 33461
rect 521 33427 559 33461
rect 593 33427 631 33461
rect 665 33427 703 33461
rect 737 33427 775 33461
rect 809 33427 843 33461
rect 877 33427 915 33461
rect 949 33427 983 33461
rect -17 33393 983 33427
rect 17 33359 55 33393
rect 89 33359 127 33393
rect 161 33359 199 33393
rect 233 33359 271 33393
rect 305 33359 343 33393
rect 377 33359 415 33393
rect 449 33359 487 33393
rect 521 33359 559 33393
rect 593 33359 631 33393
rect 665 33359 703 33393
rect 737 33359 775 33393
rect 809 33377 983 33393
rect 809 33359 843 33377
rect -17 33343 843 33359
rect 877 33343 915 33377
rect 949 33343 983 33377
rect -17 33325 983 33343
rect 17 33291 55 33325
rect 89 33291 127 33325
rect 161 33291 199 33325
rect 233 33291 271 33325
rect 305 33291 343 33325
rect 377 33291 415 33325
rect 449 33291 487 33325
rect 521 33291 559 33325
rect 593 33291 631 33325
rect 665 33291 703 33325
rect 737 33291 775 33325
rect 809 33293 983 33325
rect 809 33291 843 33293
rect -17 33259 843 33291
rect 877 33259 915 33293
rect 949 33259 983 33293
rect -17 33257 983 33259
rect 17 33223 55 33257
rect 89 33223 127 33257
rect 161 33223 199 33257
rect 233 33223 271 33257
rect 305 33223 343 33257
rect 377 33223 415 33257
rect 449 33223 487 33257
rect 521 33223 559 33257
rect 593 33223 631 33257
rect 665 33223 703 33257
rect 737 33223 775 33257
rect 809 33223 983 33257
rect -17 33209 983 33223
rect -17 33189 843 33209
rect 17 33155 55 33189
rect 89 33155 127 33189
rect 161 33155 199 33189
rect 233 33155 271 33189
rect 305 33155 343 33189
rect 377 33155 415 33189
rect 449 33155 487 33189
rect 521 33155 559 33189
rect 593 33155 631 33189
rect 665 33155 703 33189
rect 737 33155 775 33189
rect 809 33175 843 33189
rect 877 33175 915 33209
rect 949 33175 983 33209
rect 809 33155 983 33175
rect -17 33125 983 33155
rect -17 33121 843 33125
rect 17 33087 55 33121
rect 89 33087 127 33121
rect 161 33087 199 33121
rect 233 33087 271 33121
rect 305 33087 343 33121
rect 377 33087 415 33121
rect 449 33087 487 33121
rect 521 33087 559 33121
rect 593 33087 631 33121
rect 665 33087 703 33121
rect 737 33087 775 33121
rect 809 33091 843 33121
rect 877 33091 915 33125
rect 949 33091 983 33125
rect 809 33087 983 33091
rect -17 33053 983 33087
rect 17 33019 55 33053
rect 89 33019 127 33053
rect 161 33019 199 33053
rect 233 33019 271 33053
rect 305 33019 343 33053
rect 377 33019 415 33053
rect 449 33019 487 33053
rect 521 33019 559 33053
rect 593 33019 631 33053
rect 665 33019 703 33053
rect 737 33019 775 33053
rect 809 33041 983 33053
rect 809 33019 843 33041
rect -17 33007 843 33019
rect 877 33007 915 33041
rect 949 33007 983 33041
rect -17 32985 983 33007
rect 17 32951 55 32985
rect 89 32951 127 32985
rect 161 32951 199 32985
rect 233 32951 271 32985
rect 305 32951 343 32985
rect 377 32951 415 32985
rect 449 32951 487 32985
rect 521 32951 559 32985
rect 593 32951 631 32985
rect 665 32951 703 32985
rect 737 32951 775 32985
rect 809 32957 983 32985
rect 809 32951 843 32957
rect -17 32923 843 32951
rect 877 32923 915 32957
rect 949 32923 983 32957
rect -17 32917 983 32923
rect 17 32883 55 32917
rect 89 32883 127 32917
rect 161 32883 199 32917
rect 233 32883 271 32917
rect 305 32883 343 32917
rect 377 32883 415 32917
rect 449 32883 487 32917
rect 521 32883 559 32917
rect 593 32883 631 32917
rect 665 32883 703 32917
rect 737 32883 775 32917
rect 809 32883 983 32917
rect -17 32873 983 32883
rect -17 32849 843 32873
rect 17 32815 55 32849
rect 89 32815 127 32849
rect 161 32815 199 32849
rect 233 32815 271 32849
rect 305 32815 343 32849
rect 377 32815 415 32849
rect 449 32815 487 32849
rect 521 32815 559 32849
rect 593 32815 631 32849
rect 665 32815 703 32849
rect 737 32815 775 32849
rect 809 32839 843 32849
rect 877 32839 915 32873
rect 949 32839 983 32873
rect 809 32815 983 32839
rect -17 32789 983 32815
rect -17 32781 843 32789
rect 17 32747 55 32781
rect 89 32747 127 32781
rect 161 32747 199 32781
rect 233 32747 271 32781
rect 305 32747 343 32781
rect 377 32747 415 32781
rect 449 32747 487 32781
rect 521 32747 559 32781
rect 593 32747 631 32781
rect 665 32747 703 32781
rect 737 32747 775 32781
rect 809 32755 843 32781
rect 877 32755 915 32789
rect 949 32755 983 32789
rect 809 32747 983 32755
rect -17 32713 983 32747
rect 17 32679 55 32713
rect 89 32679 127 32713
rect 161 32679 199 32713
rect 233 32679 271 32713
rect 305 32679 343 32713
rect 377 32679 415 32713
rect 449 32679 487 32713
rect 521 32679 559 32713
rect 593 32679 631 32713
rect 665 32679 703 32713
rect 737 32679 775 32713
rect 809 32705 983 32713
rect 809 32679 843 32705
rect -17 32671 843 32679
rect 877 32671 915 32705
rect 949 32671 983 32705
rect -17 32645 983 32671
rect 17 32611 55 32645
rect 89 32611 127 32645
rect 161 32611 199 32645
rect 233 32611 271 32645
rect 305 32611 343 32645
rect 377 32611 415 32645
rect 449 32611 487 32645
rect 521 32611 559 32645
rect 593 32611 631 32645
rect 665 32611 703 32645
rect 737 32611 775 32645
rect 809 32621 983 32645
rect 809 32611 843 32621
rect -17 32587 843 32611
rect 877 32587 915 32621
rect 949 32587 983 32621
rect -17 32577 983 32587
rect 17 32543 55 32577
rect 89 32543 127 32577
rect 161 32543 199 32577
rect 233 32543 271 32577
rect 305 32543 343 32577
rect 377 32543 415 32577
rect 449 32543 487 32577
rect 521 32543 559 32577
rect 593 32543 631 32577
rect 665 32543 703 32577
rect 737 32543 775 32577
rect 809 32543 983 32577
rect -17 32537 983 32543
rect -17 32509 843 32537
rect 17 32475 55 32509
rect 89 32475 127 32509
rect 161 32475 199 32509
rect 233 32475 271 32509
rect 305 32475 343 32509
rect 377 32475 415 32509
rect 449 32475 487 32509
rect 521 32475 559 32509
rect 593 32475 631 32509
rect 665 32475 703 32509
rect 737 32475 775 32509
rect 809 32503 843 32509
rect 877 32503 915 32537
rect 949 32503 983 32537
rect 809 32475 983 32503
rect -17 32453 983 32475
rect -17 32441 843 32453
rect 17 32407 55 32441
rect 89 32407 127 32441
rect 161 32407 199 32441
rect 233 32407 271 32441
rect 305 32407 343 32441
rect 377 32407 415 32441
rect 449 32407 487 32441
rect 521 32407 559 32441
rect 593 32407 631 32441
rect 665 32407 703 32441
rect 737 32407 775 32441
rect 809 32419 843 32441
rect 877 32419 915 32453
rect 949 32419 983 32453
rect 809 32407 983 32419
rect -17 32373 983 32407
rect 17 32339 55 32373
rect 89 32339 127 32373
rect 161 32339 199 32373
rect 233 32339 271 32373
rect 305 32339 343 32373
rect 377 32339 415 32373
rect 449 32339 487 32373
rect 521 32339 559 32373
rect 593 32339 631 32373
rect 665 32339 703 32373
rect 737 32339 775 32373
rect 809 32369 983 32373
rect 809 32339 843 32369
rect -17 32335 843 32339
rect 877 32335 915 32369
rect 949 32335 983 32369
rect -17 32305 983 32335
rect 17 32271 55 32305
rect 89 32271 127 32305
rect 161 32271 199 32305
rect 233 32271 271 32305
rect 305 32271 343 32305
rect 377 32271 415 32305
rect 449 32271 487 32305
rect 521 32271 559 32305
rect 593 32271 631 32305
rect 665 32271 703 32305
rect 737 32271 775 32305
rect 809 32285 983 32305
rect 809 32271 843 32285
rect -17 32251 843 32271
rect 877 32251 915 32285
rect 949 32251 983 32285
rect -17 32237 983 32251
rect 17 32203 55 32237
rect 89 32203 127 32237
rect 161 32203 199 32237
rect 233 32203 271 32237
rect 305 32203 343 32237
rect 377 32203 415 32237
rect 449 32203 487 32237
rect 521 32203 559 32237
rect 593 32203 631 32237
rect 665 32203 703 32237
rect 737 32203 775 32237
rect 809 32203 983 32237
rect -17 32201 983 32203
rect -17 32169 843 32201
rect 17 32135 55 32169
rect 89 32135 127 32169
rect 161 32135 199 32169
rect 233 32135 271 32169
rect 305 32135 343 32169
rect 377 32135 415 32169
rect 449 32135 487 32169
rect 521 32135 559 32169
rect 593 32135 631 32169
rect 665 32135 703 32169
rect 737 32135 775 32169
rect 809 32167 843 32169
rect 877 32167 915 32201
rect 949 32167 983 32201
rect 809 32135 983 32167
rect -17 32117 983 32135
rect -17 32101 843 32117
rect 17 32067 55 32101
rect 89 32067 127 32101
rect 161 32067 199 32101
rect 233 32067 271 32101
rect 305 32067 343 32101
rect 377 32067 415 32101
rect 449 32067 487 32101
rect 521 32067 559 32101
rect 593 32067 631 32101
rect 665 32067 703 32101
rect 737 32067 775 32101
rect 809 32083 843 32101
rect 877 32083 915 32117
rect 949 32083 983 32117
rect 809 32067 983 32083
rect -17 32033 983 32067
rect 17 31999 55 32033
rect 89 31999 127 32033
rect 161 31999 199 32033
rect 233 31999 271 32033
rect 305 31999 343 32033
rect 377 31999 415 32033
rect 449 31999 487 32033
rect 521 31999 559 32033
rect 593 31999 631 32033
rect 665 31999 703 32033
rect 737 31999 775 32033
rect 809 31999 843 32033
rect 877 31999 915 32033
rect 949 31999 983 32033
rect -17 31965 983 31999
rect 17 31931 55 31965
rect 89 31931 127 31965
rect 161 31931 199 31965
rect 233 31931 271 31965
rect 305 31931 343 31965
rect 377 31931 415 31965
rect 449 31931 487 31965
rect 521 31931 559 31965
rect 593 31931 631 31965
rect 665 31931 703 31965
rect 737 31931 775 31965
rect 809 31949 983 31965
rect 809 31931 843 31949
rect -17 31915 843 31931
rect 877 31915 915 31949
rect 949 31915 983 31949
rect -17 31897 983 31915
rect 17 31863 55 31897
rect 89 31863 127 31897
rect 161 31863 199 31897
rect 233 31863 271 31897
rect 305 31863 343 31897
rect 377 31863 415 31897
rect 449 31863 487 31897
rect 521 31863 559 31897
rect 593 31863 631 31897
rect 665 31863 703 31897
rect 737 31863 775 31897
rect 809 31865 983 31897
rect 809 31863 843 31865
rect -17 31831 843 31863
rect 877 31831 915 31865
rect 949 31831 983 31865
rect -17 31829 983 31831
rect 17 31795 55 31829
rect 89 31795 127 31829
rect 161 31795 199 31829
rect 233 31795 271 31829
rect 305 31795 343 31829
rect 377 31795 415 31829
rect 449 31795 487 31829
rect 521 31795 559 31829
rect 593 31795 631 31829
rect 665 31795 703 31829
rect 737 31795 775 31829
rect 809 31795 983 31829
rect -17 31781 983 31795
rect -17 31761 843 31781
rect 17 31727 55 31761
rect 89 31727 127 31761
rect 161 31727 199 31761
rect 233 31727 271 31761
rect 305 31727 343 31761
rect 377 31727 415 31761
rect 449 31727 487 31761
rect 521 31727 559 31761
rect 593 31727 631 31761
rect 665 31727 703 31761
rect 737 31727 775 31761
rect 809 31747 843 31761
rect 877 31747 915 31781
rect 949 31747 983 31781
rect 809 31727 983 31747
rect -17 31697 983 31727
rect -17 31693 843 31697
rect 17 31659 55 31693
rect 89 31659 127 31693
rect 161 31659 199 31693
rect 233 31659 271 31693
rect 305 31659 343 31693
rect 377 31659 415 31693
rect 449 31659 487 31693
rect 521 31659 559 31693
rect 593 31659 631 31693
rect 665 31659 703 31693
rect 737 31659 775 31693
rect 809 31663 843 31693
rect 877 31663 915 31697
rect 949 31663 983 31697
rect 809 31659 983 31663
rect -17 31625 983 31659
rect 17 31591 55 31625
rect 89 31591 127 31625
rect 161 31591 199 31625
rect 233 31591 271 31625
rect 305 31591 343 31625
rect 377 31591 415 31625
rect 449 31591 487 31625
rect 521 31591 559 31625
rect 593 31591 631 31625
rect 665 31591 703 31625
rect 737 31591 775 31625
rect 809 31613 983 31625
rect 809 31591 843 31613
rect -17 31579 843 31591
rect 877 31579 915 31613
rect 949 31579 983 31613
rect -17 31557 983 31579
rect 17 31523 55 31557
rect 89 31523 127 31557
rect 161 31523 199 31557
rect 233 31523 271 31557
rect 305 31523 343 31557
rect 377 31523 415 31557
rect 449 31523 487 31557
rect 521 31523 559 31557
rect 593 31523 631 31557
rect 665 31523 703 31557
rect 737 31523 775 31557
rect 809 31529 983 31557
rect 809 31523 843 31529
rect -17 31495 843 31523
rect 877 31495 915 31529
rect 949 31495 983 31529
rect -17 31489 983 31495
rect 17 31455 55 31489
rect 89 31455 127 31489
rect 161 31455 199 31489
rect 233 31455 271 31489
rect 305 31455 343 31489
rect 377 31455 415 31489
rect 449 31455 487 31489
rect 521 31455 559 31489
rect 593 31455 631 31489
rect 665 31455 703 31489
rect 737 31455 775 31489
rect 809 31455 983 31489
rect -17 31445 983 31455
rect -17 31421 843 31445
rect 17 31387 55 31421
rect 89 31387 127 31421
rect 161 31387 199 31421
rect 233 31387 271 31421
rect 305 31387 343 31421
rect 377 31387 415 31421
rect 449 31387 487 31421
rect 521 31387 559 31421
rect 593 31387 631 31421
rect 665 31387 703 31421
rect 737 31387 775 31421
rect 809 31411 843 31421
rect 877 31411 915 31445
rect 949 31411 983 31445
rect 809 31387 983 31411
rect -17 31361 983 31387
rect -17 31353 843 31361
rect 17 31319 55 31353
rect 89 31319 127 31353
rect 161 31319 199 31353
rect 233 31319 271 31353
rect 305 31319 343 31353
rect 377 31319 415 31353
rect 449 31319 487 31353
rect 521 31319 559 31353
rect 593 31319 631 31353
rect 665 31319 703 31353
rect 737 31319 775 31353
rect 809 31327 843 31353
rect 877 31327 915 31361
rect 949 31327 983 31361
rect 809 31319 983 31327
rect -17 31285 983 31319
rect 17 31251 55 31285
rect 89 31251 127 31285
rect 161 31251 199 31285
rect 233 31251 271 31285
rect 305 31251 343 31285
rect 377 31251 415 31285
rect 449 31251 487 31285
rect 521 31251 559 31285
rect 593 31251 631 31285
rect 665 31251 703 31285
rect 737 31251 775 31285
rect 809 31277 983 31285
rect 809 31251 843 31277
rect -17 31243 843 31251
rect 877 31243 915 31277
rect 949 31243 983 31277
rect -17 31217 983 31243
rect 17 31183 55 31217
rect 89 31183 127 31217
rect 161 31183 199 31217
rect 233 31183 271 31217
rect 305 31183 343 31217
rect 377 31183 415 31217
rect 449 31183 487 31217
rect 521 31183 559 31217
rect 593 31183 631 31217
rect 665 31183 703 31217
rect 737 31183 775 31217
rect 809 31193 983 31217
rect 809 31183 843 31193
rect -17 31159 843 31183
rect 877 31159 915 31193
rect 949 31159 983 31193
rect -17 31149 983 31159
rect 17 31115 55 31149
rect 89 31115 127 31149
rect 161 31115 199 31149
rect 233 31115 271 31149
rect 305 31115 343 31149
rect 377 31115 415 31149
rect 449 31115 487 31149
rect 521 31115 559 31149
rect 593 31115 631 31149
rect 665 31115 703 31149
rect 737 31115 775 31149
rect 809 31115 983 31149
rect -17 31109 983 31115
rect -17 31081 843 31109
rect 17 31047 55 31081
rect 89 31047 127 31081
rect 161 31047 199 31081
rect 233 31047 271 31081
rect 305 31047 343 31081
rect 377 31047 415 31081
rect 449 31047 487 31081
rect 521 31047 559 31081
rect 593 31047 631 31081
rect 665 31047 703 31081
rect 737 31047 775 31081
rect 809 31075 843 31081
rect 877 31075 915 31109
rect 949 31075 983 31109
rect 809 31047 983 31075
rect -17 31025 983 31047
rect -17 31013 843 31025
rect 17 30979 55 31013
rect 89 30979 127 31013
rect 161 30979 199 31013
rect 233 30979 271 31013
rect 305 30979 343 31013
rect 377 30979 415 31013
rect 449 30979 487 31013
rect 521 30979 559 31013
rect 593 30979 631 31013
rect 665 30979 703 31013
rect 737 30979 775 31013
rect 809 30991 843 31013
rect 877 30991 915 31025
rect 949 30991 983 31025
rect 809 30979 983 30991
rect -17 30945 983 30979
rect 17 30911 55 30945
rect 89 30911 127 30945
rect 161 30911 199 30945
rect 233 30911 271 30945
rect 305 30911 343 30945
rect 377 30911 415 30945
rect 449 30911 487 30945
rect 521 30911 559 30945
rect 593 30911 631 30945
rect 665 30911 703 30945
rect 737 30911 775 30945
rect 809 30941 983 30945
rect 809 30911 843 30941
rect -17 30907 843 30911
rect 877 30907 915 30941
rect 949 30907 983 30941
rect -17 30877 983 30907
rect 17 30843 55 30877
rect 89 30843 127 30877
rect 161 30843 199 30877
rect 233 30843 271 30877
rect 305 30843 343 30877
rect 377 30843 415 30877
rect 449 30843 487 30877
rect 521 30843 559 30877
rect 593 30843 631 30877
rect 665 30843 703 30877
rect 737 30843 775 30877
rect 809 30857 983 30877
rect 809 30843 843 30857
rect -17 30823 843 30843
rect 877 30823 915 30857
rect 949 30823 983 30857
rect -17 30809 983 30823
rect 17 30775 55 30809
rect 89 30775 127 30809
rect 161 30775 199 30809
rect 233 30775 271 30809
rect 305 30775 343 30809
rect 377 30775 415 30809
rect 449 30775 487 30809
rect 521 30775 559 30809
rect 593 30775 631 30809
rect 665 30775 703 30809
rect 737 30775 775 30809
rect 809 30775 983 30809
rect -17 30773 983 30775
rect -17 30741 843 30773
rect 17 30707 55 30741
rect 89 30707 127 30741
rect 161 30707 199 30741
rect 233 30707 271 30741
rect 305 30707 343 30741
rect 377 30707 415 30741
rect 449 30707 487 30741
rect 521 30707 559 30741
rect 593 30707 631 30741
rect 665 30707 703 30741
rect 737 30707 775 30741
rect 809 30739 843 30741
rect 877 30739 915 30773
rect 949 30739 983 30773
rect 809 30707 983 30739
rect -17 30689 983 30707
rect -17 30673 843 30689
rect 17 30639 55 30673
rect 89 30639 127 30673
rect 161 30639 199 30673
rect 233 30639 271 30673
rect 305 30639 343 30673
rect 377 30639 415 30673
rect 449 30639 487 30673
rect 521 30639 559 30673
rect 593 30639 631 30673
rect 665 30639 703 30673
rect 737 30639 775 30673
rect 809 30655 843 30673
rect 877 30655 915 30689
rect 949 30655 983 30689
rect 809 30639 983 30655
rect -17 30605 983 30639
rect 17 30571 55 30605
rect 89 30571 127 30605
rect 161 30571 199 30605
rect 233 30571 271 30605
rect 305 30571 343 30605
rect 377 30571 415 30605
rect 449 30571 487 30605
rect 521 30571 559 30605
rect 593 30571 631 30605
rect 665 30571 703 30605
rect 737 30571 775 30605
rect 809 30571 843 30605
rect 877 30571 915 30605
rect 949 30571 983 30605
rect -17 30537 983 30571
rect 17 30503 55 30537
rect 89 30503 127 30537
rect 161 30503 199 30537
rect 233 30503 271 30537
rect 305 30503 343 30537
rect 377 30503 415 30537
rect 449 30503 487 30537
rect 521 30503 559 30537
rect 593 30503 631 30537
rect 665 30503 703 30537
rect 737 30503 775 30537
rect 809 30521 983 30537
rect 809 30503 843 30521
rect -17 30487 843 30503
rect 877 30487 915 30521
rect 949 30487 983 30521
rect -17 30469 983 30487
rect 17 30435 55 30469
rect 89 30435 127 30469
rect 161 30435 199 30469
rect 233 30435 271 30469
rect 305 30435 343 30469
rect 377 30435 415 30469
rect 449 30435 487 30469
rect 521 30435 559 30469
rect 593 30435 631 30469
rect 665 30435 703 30469
rect 737 30435 775 30469
rect 809 30436 983 30469
rect 809 30435 843 30436
rect -17 30402 843 30435
rect 877 30402 915 30436
rect 949 30402 983 30436
rect -17 30401 983 30402
rect 17 30367 55 30401
rect 89 30367 127 30401
rect 161 30367 199 30401
rect 233 30367 271 30401
rect 305 30367 343 30401
rect 377 30367 415 30401
rect 449 30367 487 30401
rect 521 30367 559 30401
rect 593 30367 631 30401
rect 665 30367 703 30401
rect 737 30367 775 30401
rect 809 30367 983 30401
rect -17 30351 983 30367
rect -17 30333 843 30351
rect 17 30299 55 30333
rect 89 30299 127 30333
rect 161 30299 199 30333
rect 233 30299 271 30333
rect 305 30299 343 30333
rect 377 30299 415 30333
rect 449 30299 487 30333
rect 521 30299 559 30333
rect 593 30299 631 30333
rect 665 30299 703 30333
rect 737 30299 775 30333
rect 809 30317 843 30333
rect 877 30317 915 30351
rect 949 30317 983 30351
rect 809 30299 983 30317
rect -17 30266 983 30299
rect -17 30265 843 30266
rect 17 30231 55 30265
rect 89 30231 127 30265
rect 161 30231 199 30265
rect 233 30231 271 30265
rect 305 30231 343 30265
rect 377 30231 415 30265
rect 449 30231 487 30265
rect 521 30231 559 30265
rect 593 30231 631 30265
rect 665 30231 703 30265
rect 737 30231 775 30265
rect 809 30232 843 30265
rect 877 30232 915 30266
rect 949 30232 983 30266
rect 809 30231 983 30232
rect -17 30197 983 30231
rect 17 30163 55 30197
rect 89 30163 127 30197
rect 161 30163 199 30197
rect 233 30163 271 30197
rect 305 30163 343 30197
rect 377 30163 415 30197
rect 449 30163 487 30197
rect 521 30163 559 30197
rect 593 30163 631 30197
rect 665 30163 703 30197
rect 737 30163 775 30197
rect 809 30181 983 30197
rect 809 30163 843 30181
rect -17 30147 843 30163
rect 877 30147 915 30181
rect 949 30147 983 30181
rect -17 30129 983 30147
rect 17 30095 55 30129
rect 89 30095 127 30129
rect 161 30095 199 30129
rect 233 30095 271 30129
rect 305 30095 343 30129
rect 377 30095 415 30129
rect 449 30095 487 30129
rect 521 30095 559 30129
rect 593 30095 631 30129
rect 665 30095 703 30129
rect 737 30095 775 30129
rect 809 30096 983 30129
rect 809 30095 843 30096
rect -17 30062 843 30095
rect 877 30062 915 30096
rect 949 30062 983 30096
rect -17 30061 983 30062
rect 17 30027 55 30061
rect 89 30027 127 30061
rect 161 30027 199 30061
rect 233 30027 271 30061
rect 305 30027 343 30061
rect 377 30027 415 30061
rect 449 30027 487 30061
rect 521 30027 559 30061
rect 593 30027 631 30061
rect 665 30027 703 30061
rect 737 30027 775 30061
rect 809 30027 983 30061
rect -17 30011 983 30027
rect -17 29993 843 30011
rect 17 29959 55 29993
rect 89 29959 127 29993
rect 161 29959 199 29993
rect 233 29959 271 29993
rect 305 29959 343 29993
rect 377 29959 415 29993
rect 449 29959 487 29993
rect 521 29959 559 29993
rect 593 29959 631 29993
rect 665 29959 703 29993
rect 737 29959 775 29993
rect 809 29977 843 29993
rect 877 29977 915 30011
rect 949 29977 983 30011
rect 809 29959 983 29977
rect -17 29926 983 29959
rect -17 29925 843 29926
rect 17 29891 55 29925
rect 89 29891 127 29925
rect 161 29891 199 29925
rect 233 29891 271 29925
rect 305 29891 343 29925
rect 377 29891 415 29925
rect 449 29891 487 29925
rect 521 29891 559 29925
rect 593 29891 631 29925
rect 665 29891 703 29925
rect 737 29891 775 29925
rect 809 29892 843 29925
rect 877 29892 915 29926
rect 949 29892 983 29926
rect 809 29891 983 29892
rect -17 29857 983 29891
rect 17 29823 55 29857
rect 89 29823 127 29857
rect 161 29823 199 29857
rect 233 29823 271 29857
rect 305 29823 343 29857
rect 377 29823 415 29857
rect 449 29823 487 29857
rect 521 29823 559 29857
rect 593 29823 631 29857
rect 665 29823 703 29857
rect 737 29823 775 29857
rect 809 29841 983 29857
rect 809 29823 843 29841
rect -17 29807 843 29823
rect 877 29807 915 29841
rect 949 29807 983 29841
rect -17 29789 983 29807
rect 17 29755 55 29789
rect 89 29755 127 29789
rect 161 29755 199 29789
rect 233 29755 271 29789
rect 305 29755 343 29789
rect 377 29755 415 29789
rect 449 29755 487 29789
rect 521 29755 559 29789
rect 593 29755 631 29789
rect 665 29755 703 29789
rect 737 29755 775 29789
rect 809 29756 983 29789
rect 809 29755 843 29756
rect -17 29722 843 29755
rect 877 29722 915 29756
rect 949 29722 983 29756
rect -17 29721 983 29722
rect 17 29687 55 29721
rect 89 29687 127 29721
rect 161 29687 199 29721
rect 233 29687 271 29721
rect 305 29687 343 29721
rect 377 29687 415 29721
rect 449 29687 487 29721
rect 521 29687 559 29721
rect 593 29687 631 29721
rect 665 29687 703 29721
rect 737 29687 775 29721
rect 809 29687 983 29721
rect -17 29671 983 29687
rect -17 29652 843 29671
rect 17 29618 55 29652
rect 89 29618 127 29652
rect 161 29618 199 29652
rect 233 29618 271 29652
rect 305 29618 343 29652
rect 377 29618 415 29652
rect 449 29618 487 29652
rect 521 29618 559 29652
rect 593 29618 631 29652
rect 665 29618 703 29652
rect 737 29618 775 29652
rect 809 29637 843 29652
rect 877 29637 915 29671
rect 949 29637 983 29671
rect 809 29618 983 29637
rect -17 29586 983 29618
rect -17 29583 843 29586
rect 17 29549 55 29583
rect 89 29549 127 29583
rect 161 29549 199 29583
rect 233 29549 271 29583
rect 305 29549 343 29583
rect 377 29549 415 29583
rect 449 29549 487 29583
rect 521 29549 559 29583
rect 593 29549 631 29583
rect 665 29549 703 29583
rect 737 29549 775 29583
rect 809 29552 843 29583
rect 877 29552 915 29586
rect 949 29552 983 29586
rect 809 29549 983 29552
rect -17 29514 983 29549
rect 17 29480 55 29514
rect 89 29480 127 29514
rect 161 29480 199 29514
rect 233 29480 271 29514
rect 305 29480 343 29514
rect 377 29480 415 29514
rect 449 29480 487 29514
rect 521 29480 559 29514
rect 593 29480 631 29514
rect 665 29480 703 29514
rect 737 29480 775 29514
rect 809 29501 983 29514
rect 809 29480 843 29501
rect -17 29467 843 29480
rect 877 29467 915 29501
rect 949 29467 983 29501
rect -17 29445 983 29467
rect 17 29411 55 29445
rect 89 29411 127 29445
rect 161 29411 199 29445
rect 233 29411 271 29445
rect 305 29411 343 29445
rect 377 29411 415 29445
rect 449 29411 487 29445
rect 521 29411 559 29445
rect 593 29411 631 29445
rect 665 29411 703 29445
rect 737 29411 775 29445
rect 809 29416 983 29445
rect 809 29411 843 29416
rect -17 29382 843 29411
rect 877 29382 915 29416
rect 949 29382 983 29416
rect -17 29376 983 29382
rect 17 29342 55 29376
rect 89 29342 127 29376
rect 161 29342 199 29376
rect 233 29342 271 29376
rect 305 29342 343 29376
rect 377 29342 415 29376
rect 449 29342 487 29376
rect 521 29342 559 29376
rect 593 29342 631 29376
rect 665 29342 703 29376
rect 737 29342 775 29376
rect 809 29342 983 29376
rect -17 29331 983 29342
rect -17 29307 843 29331
rect 17 29273 55 29307
rect 89 29273 127 29307
rect 161 29273 199 29307
rect 233 29273 271 29307
rect 305 29273 343 29307
rect 377 29273 415 29307
rect 449 29273 487 29307
rect 521 29273 559 29307
rect 593 29273 631 29307
rect 665 29273 703 29307
rect 737 29273 775 29307
rect 809 29297 843 29307
rect 877 29297 915 29331
rect 949 29297 983 29331
rect 809 29273 983 29297
rect -17 29246 983 29273
rect -17 29238 843 29246
rect 17 29204 55 29238
rect 89 29204 127 29238
rect 161 29204 199 29238
rect 233 29204 271 29238
rect 305 29204 343 29238
rect 377 29204 415 29238
rect 449 29204 487 29238
rect 521 29204 559 29238
rect 593 29204 631 29238
rect 665 29204 703 29238
rect 737 29204 775 29238
rect 809 29212 843 29238
rect 877 29212 915 29246
rect 949 29212 983 29246
rect 809 29204 983 29212
rect -17 29169 983 29204
rect 17 29135 55 29169
rect 89 29135 127 29169
rect 161 29135 199 29169
rect 233 29135 271 29169
rect 305 29135 343 29169
rect 377 29135 415 29169
rect 449 29135 487 29169
rect 521 29135 559 29169
rect 593 29135 631 29169
rect 665 29135 703 29169
rect 737 29135 775 29169
rect 809 29161 983 29169
rect 809 29135 843 29161
rect -17 29127 843 29135
rect 877 29127 915 29161
rect 949 29127 983 29161
rect -17 29100 983 29127
rect 17 29066 55 29100
rect 89 29066 127 29100
rect 161 29066 199 29100
rect 233 29066 271 29100
rect 305 29066 343 29100
rect 377 29066 415 29100
rect 449 29066 487 29100
rect 521 29066 559 29100
rect 593 29066 631 29100
rect 665 29066 703 29100
rect 737 29066 775 29100
rect 809 29076 983 29100
rect 809 29066 843 29076
rect -17 29042 843 29066
rect 877 29042 915 29076
rect 949 29042 983 29076
rect -17 27986 843 28010
rect 17 27952 55 27986
rect 89 27952 127 27986
rect 161 27952 199 27986
rect 233 27952 271 27986
rect 305 27952 343 27986
rect 377 27952 415 27986
rect 449 27952 487 27986
rect 521 27952 559 27986
rect 593 27952 631 27986
rect 665 27952 703 27986
rect 737 27952 775 27986
rect 809 27976 843 27986
rect 877 27976 915 28010
rect 949 27976 983 28010
rect 809 27952 983 27976
rect -17 27942 983 27952
rect -17 27917 843 27942
rect 17 27883 55 27917
rect 89 27883 127 27917
rect 161 27883 199 27917
rect 233 27883 271 27917
rect 305 27883 343 27917
rect 377 27883 415 27917
rect 449 27883 487 27917
rect 521 27883 559 27917
rect 593 27883 631 27917
rect 665 27883 703 27917
rect 737 27883 775 27917
rect 809 27908 843 27917
rect 877 27908 915 27942
rect 949 27908 983 27942
rect 809 27883 983 27908
rect -17 27874 983 27883
rect -17 27848 843 27874
rect 17 27814 55 27848
rect 89 27814 127 27848
rect 161 27814 199 27848
rect 233 27814 271 27848
rect 305 27814 343 27848
rect 377 27814 415 27848
rect 449 27814 487 27848
rect 521 27814 559 27848
rect 593 27814 631 27848
rect 665 27814 703 27848
rect 737 27814 775 27848
rect 809 27840 843 27848
rect 877 27840 915 27874
rect 949 27840 983 27874
rect 809 27814 983 27840
rect -17 27806 983 27814
rect -17 27779 843 27806
rect 17 27745 55 27779
rect 89 27745 127 27779
rect 161 27745 199 27779
rect 233 27745 271 27779
rect 305 27745 343 27779
rect 377 27745 415 27779
rect 449 27745 487 27779
rect 521 27745 559 27779
rect 593 27745 631 27779
rect 665 27745 703 27779
rect 737 27745 775 27779
rect 809 27772 843 27779
rect 877 27772 915 27806
rect 949 27772 983 27806
rect 809 27745 983 27772
rect -17 27738 983 27745
rect -17 27710 843 27738
rect 17 27676 55 27710
rect 89 27676 127 27710
rect 161 27676 199 27710
rect 233 27676 271 27710
rect 305 27676 343 27710
rect 377 27676 415 27710
rect 449 27676 487 27710
rect 521 27676 559 27710
rect 593 27676 631 27710
rect 665 27676 703 27710
rect 737 27676 775 27710
rect 809 27704 843 27710
rect 877 27704 915 27738
rect 949 27704 983 27738
rect 809 27676 983 27704
rect -17 27670 983 27676
rect -17 27641 843 27670
rect 17 27607 55 27641
rect 89 27607 127 27641
rect 161 27607 199 27641
rect 233 27607 271 27641
rect 305 27607 343 27641
rect 377 27607 415 27641
rect 449 27607 487 27641
rect 521 27607 559 27641
rect 593 27607 631 27641
rect 665 27607 703 27641
rect 737 27607 775 27641
rect 809 27636 843 27641
rect 877 27636 915 27670
rect 949 27636 983 27670
rect 809 27607 983 27636
rect -17 27602 983 27607
rect -17 27572 843 27602
rect 17 27538 55 27572
rect 89 27538 127 27572
rect 161 27538 199 27572
rect 233 27538 271 27572
rect 305 27538 343 27572
rect 377 27538 415 27572
rect 449 27538 487 27572
rect 521 27538 559 27572
rect 593 27538 631 27572
rect 665 27538 703 27572
rect 737 27538 775 27572
rect 809 27568 843 27572
rect 877 27568 915 27602
rect 949 27568 983 27602
rect 809 27538 983 27568
rect -17 27534 983 27538
rect -17 27503 843 27534
rect 17 27469 55 27503
rect 89 27469 127 27503
rect 161 27469 199 27503
rect 233 27469 271 27503
rect 305 27469 343 27503
rect 377 27469 415 27503
rect 449 27469 487 27503
rect 521 27469 559 27503
rect 593 27469 631 27503
rect 665 27469 703 27503
rect 737 27469 775 27503
rect 809 27500 843 27503
rect 877 27500 915 27534
rect 949 27500 983 27534
rect 809 27469 983 27500
rect -17 27466 983 27469
rect -17 27434 843 27466
rect 17 27400 55 27434
rect 89 27400 127 27434
rect 161 27400 199 27434
rect 233 27400 271 27434
rect 305 27400 343 27434
rect 377 27400 415 27434
rect 449 27400 487 27434
rect 521 27400 559 27434
rect 593 27400 631 27434
rect 665 27400 703 27434
rect 737 27400 775 27434
rect 809 27432 843 27434
rect 877 27432 915 27466
rect 949 27432 983 27466
rect 809 27400 983 27432
rect -17 27398 983 27400
rect -17 27365 843 27398
rect 17 27331 55 27365
rect 89 27331 127 27365
rect 161 27331 199 27365
rect 233 27331 271 27365
rect 305 27331 343 27365
rect 377 27331 415 27365
rect 449 27331 487 27365
rect 521 27331 559 27365
rect 593 27331 631 27365
rect 665 27331 703 27365
rect 737 27331 775 27365
rect 809 27364 843 27365
rect 877 27364 915 27398
rect 949 27364 983 27398
rect 809 27331 983 27364
rect -17 27330 983 27331
rect -17 27296 843 27330
rect 877 27296 915 27330
rect 949 27296 983 27330
rect 17 27262 55 27296
rect 89 27262 127 27296
rect 161 27262 199 27296
rect 233 27262 271 27296
rect 305 27262 343 27296
rect 377 27262 415 27296
rect 449 27262 487 27296
rect 521 27262 559 27296
rect 593 27262 631 27296
rect 665 27262 703 27296
rect 737 27262 775 27296
rect 809 27262 983 27296
rect -17 27228 843 27262
rect 877 27228 915 27262
rect 949 27228 983 27262
rect -17 27227 983 27228
rect 17 27193 55 27227
rect 89 27193 127 27227
rect 161 27193 199 27227
rect 233 27193 271 27227
rect 305 27193 343 27227
rect 377 27193 415 27227
rect 449 27193 487 27227
rect 521 27193 559 27227
rect 593 27193 631 27227
rect 665 27193 703 27227
rect 737 27193 775 27227
rect 809 27194 983 27227
rect 809 27193 843 27194
rect -17 27160 843 27193
rect 877 27160 915 27194
rect 949 27160 983 27194
rect -17 27158 983 27160
rect 17 27124 55 27158
rect 89 27124 127 27158
rect 161 27124 199 27158
rect 233 27124 271 27158
rect 305 27124 343 27158
rect 377 27124 415 27158
rect 449 27124 487 27158
rect 521 27124 559 27158
rect 593 27124 631 27158
rect 665 27124 703 27158
rect 737 27124 775 27158
rect 809 27126 983 27158
rect 809 27124 843 27126
rect -17 27092 843 27124
rect 877 27092 915 27126
rect 949 27092 983 27126
rect -17 27089 983 27092
rect 17 27055 55 27089
rect 89 27055 127 27089
rect 161 27055 199 27089
rect 233 27055 271 27089
rect 305 27055 343 27089
rect 377 27055 415 27089
rect 449 27055 487 27089
rect 521 27055 559 27089
rect 593 27055 631 27089
rect 665 27055 703 27089
rect 737 27055 775 27089
rect 809 27058 983 27089
rect 809 27055 843 27058
rect -17 27024 843 27055
rect 877 27024 915 27058
rect 949 27024 983 27058
rect -17 27020 983 27024
rect 17 26986 55 27020
rect 89 26986 127 27020
rect 161 26986 199 27020
rect 233 26986 271 27020
rect 305 26986 343 27020
rect 377 26986 415 27020
rect 449 26986 487 27020
rect 521 26986 559 27020
rect 593 26986 631 27020
rect 665 26986 703 27020
rect 737 26986 775 27020
rect 809 26990 983 27020
rect 809 26986 843 26990
rect -17 26956 843 26986
rect 877 26956 915 26990
rect 949 26956 983 26990
rect -17 26951 983 26956
rect 17 26917 55 26951
rect 89 26917 127 26951
rect 161 26917 199 26951
rect 233 26917 271 26951
rect 305 26917 343 26951
rect 377 26917 415 26951
rect 449 26917 487 26951
rect 521 26917 559 26951
rect 593 26917 631 26951
rect 665 26917 703 26951
rect 737 26917 775 26951
rect 809 26922 983 26951
rect 809 26917 843 26922
rect -17 26888 843 26917
rect 877 26888 915 26922
rect 949 26888 983 26922
rect -17 26882 983 26888
rect 17 26848 55 26882
rect 89 26848 127 26882
rect 161 26848 199 26882
rect 233 26848 271 26882
rect 305 26848 343 26882
rect 377 26848 415 26882
rect 449 26848 487 26882
rect 521 26848 559 26882
rect 593 26848 631 26882
rect 665 26848 703 26882
rect 737 26848 775 26882
rect 809 26854 983 26882
rect 809 26848 843 26854
rect -17 26820 843 26848
rect 877 26820 915 26854
rect 949 26820 983 26854
rect -17 26813 983 26820
rect 17 26779 55 26813
rect 89 26779 127 26813
rect 161 26779 199 26813
rect 233 26779 271 26813
rect 305 26779 343 26813
rect 377 26779 415 26813
rect 449 26779 487 26813
rect 521 26779 559 26813
rect 593 26779 631 26813
rect 665 26779 703 26813
rect 737 26779 775 26813
rect 809 26785 983 26813
rect 809 26779 843 26785
rect -17 26751 843 26779
rect 877 26751 915 26785
rect 949 26751 983 26785
rect -17 26744 983 26751
rect 17 26710 55 26744
rect 89 26710 127 26744
rect 161 26710 199 26744
rect 233 26710 271 26744
rect 305 26710 343 26744
rect 377 26710 415 26744
rect 449 26710 487 26744
rect 521 26710 559 26744
rect 593 26710 631 26744
rect 665 26710 703 26744
rect 737 26710 775 26744
rect 809 26716 983 26744
rect 809 26710 843 26716
rect -17 26682 843 26710
rect 877 26682 915 26716
rect 949 26682 983 26716
rect -17 26675 983 26682
rect 17 26641 55 26675
rect 89 26641 127 26675
rect 161 26641 199 26675
rect 233 26641 271 26675
rect 305 26641 343 26675
rect 377 26641 415 26675
rect 449 26641 487 26675
rect 521 26641 559 26675
rect 593 26641 631 26675
rect 665 26641 703 26675
rect 737 26641 775 26675
rect 809 26647 983 26675
rect 809 26641 843 26647
rect -17 26613 843 26641
rect 877 26613 915 26647
rect 949 26613 983 26647
rect -17 26606 983 26613
rect 17 26572 55 26606
rect 89 26572 127 26606
rect 161 26572 199 26606
rect 233 26572 271 26606
rect 305 26572 343 26606
rect 377 26572 415 26606
rect 449 26572 487 26606
rect 521 26572 559 26606
rect 593 26572 631 26606
rect 665 26572 703 26606
rect 737 26572 775 26606
rect 809 26578 983 26606
rect 809 26572 843 26578
rect -17 26544 843 26572
rect 877 26544 915 26578
rect 949 26544 983 26578
rect -17 26537 983 26544
rect 17 26503 55 26537
rect 89 26503 127 26537
rect 161 26503 199 26537
rect 233 26503 271 26537
rect 305 26503 343 26537
rect 377 26503 415 26537
rect 449 26503 487 26537
rect 521 26503 559 26537
rect 593 26503 631 26537
rect 665 26503 703 26537
rect 737 26503 775 26537
rect 809 26509 983 26537
rect 809 26503 843 26509
rect -17 26475 843 26503
rect 877 26475 915 26509
rect 949 26475 983 26509
rect -17 26467 983 26475
rect 17 26433 55 26467
rect 89 26433 127 26467
rect 161 26433 199 26467
rect 233 26433 271 26467
rect 305 26433 343 26467
rect 377 26433 415 26467
rect 449 26433 487 26467
rect 521 26433 559 26467
rect 593 26433 631 26467
rect 665 26433 703 26467
rect 737 26433 775 26467
rect 809 26440 983 26467
rect 809 26433 843 26440
rect -17 26406 843 26433
rect 877 26406 915 26440
rect 949 26406 983 26440
rect -17 26397 983 26406
rect 17 26363 55 26397
rect 89 26363 127 26397
rect 161 26363 199 26397
rect 233 26363 271 26397
rect 305 26363 343 26397
rect 377 26363 415 26397
rect 449 26363 487 26397
rect 521 26363 559 26397
rect 593 26363 631 26397
rect 665 26363 703 26397
rect 737 26363 775 26397
rect 809 26371 983 26397
rect 809 26363 843 26371
rect -17 26337 843 26363
rect 877 26337 915 26371
rect 949 26337 983 26371
rect -17 26327 983 26337
rect 17 26293 55 26327
rect 89 26293 127 26327
rect 161 26293 199 26327
rect 233 26293 271 26327
rect 305 26293 343 26327
rect 377 26293 415 26327
rect 449 26293 487 26327
rect 521 26293 559 26327
rect 593 26293 631 26327
rect 665 26293 703 26327
rect 737 26293 775 26327
rect 809 26302 983 26327
rect 809 26293 843 26302
rect -17 26268 843 26293
rect 877 26268 915 26302
rect 949 26268 983 26302
rect -17 26257 983 26268
rect 17 26223 55 26257
rect 89 26223 127 26257
rect 161 26223 199 26257
rect 233 26223 271 26257
rect 305 26223 343 26257
rect 377 26223 415 26257
rect 449 26223 487 26257
rect 521 26223 559 26257
rect 593 26223 631 26257
rect 665 26223 703 26257
rect 737 26223 775 26257
rect 809 26233 983 26257
rect 809 26223 843 26233
rect -17 26199 843 26223
rect 877 26199 915 26233
rect 949 26199 983 26233
rect 15976 7121 16024 7145
rect 15976 7087 15983 7121
rect 16017 7087 16024 7121
rect 15976 7052 16024 7087
rect 15976 7018 15983 7052
rect 16017 7018 16024 7052
rect 15976 6983 16024 7018
rect 15976 6949 15983 6983
rect 16017 6949 16024 6983
rect 15976 6914 16024 6949
rect 15976 6880 15983 6914
rect 16017 6880 16024 6914
rect 15976 6845 16024 6880
rect 15976 6811 15983 6845
rect 16017 6811 16024 6845
rect 15976 6776 16024 6811
rect 15976 6742 15983 6776
rect 16017 6742 16024 6776
rect 15976 6707 16024 6742
rect 15976 6673 15983 6707
rect 16017 6673 16024 6707
rect 15976 6638 16024 6673
rect 15976 6604 15983 6638
rect 16017 6604 16024 6638
rect 15976 6569 16024 6604
rect 15976 6535 15983 6569
rect 16017 6535 16024 6569
rect 15976 6500 16024 6535
rect 15976 6466 15983 6500
rect 16017 6466 16024 6500
rect 15976 6431 16024 6466
rect 15976 6397 15983 6431
rect 16017 6397 16024 6431
rect 15976 6361 16024 6397
rect 15976 6327 15983 6361
rect 16017 6327 16024 6361
rect 15976 6291 16024 6327
rect 15976 6257 15983 6291
rect 16017 6257 16024 6291
rect 15976 6221 16024 6257
rect 15976 6187 15983 6221
rect 16017 6187 16024 6221
rect 15976 6151 16024 6187
rect 15976 6117 15983 6151
rect 16017 6117 16024 6151
rect 15976 6081 16024 6117
rect 15976 6047 15983 6081
rect 16017 6047 16024 6081
rect 15976 6023 16024 6047
rect 15976 4979 16024 5003
rect 15976 4945 15983 4979
rect 16017 4945 16024 4979
rect 15976 4911 16024 4945
rect 15976 4877 15983 4911
rect 16017 4877 16024 4911
rect 15976 4843 16024 4877
rect 15976 4809 15983 4843
rect 16017 4809 16024 4843
rect 15976 4775 16024 4809
rect 15976 4741 15983 4775
rect 16017 4741 16024 4775
rect 15976 4707 16024 4741
rect 15976 4673 15983 4707
rect 16017 4673 16024 4707
rect 15976 4639 16024 4673
rect 15976 4605 15983 4639
rect 16017 4605 16024 4639
rect 15976 4571 16024 4605
rect 15976 4537 15983 4571
rect 16017 4537 16024 4571
rect 15976 4503 16024 4537
rect 15976 4469 15983 4503
rect 16017 4469 16024 4503
rect 15976 4435 16024 4469
rect 15976 4401 15983 4435
rect 16017 4401 16024 4435
rect 15976 4367 16024 4401
rect 15976 4333 15983 4367
rect 16017 4333 16024 4367
rect 15976 4299 16024 4333
rect 15976 4265 15983 4299
rect 16017 4265 16024 4299
rect 15976 4231 16024 4265
rect 15976 4197 15983 4231
rect 16017 4197 16024 4231
rect 15976 4162 16024 4197
rect 15976 4128 15983 4162
rect 16017 4128 16024 4162
rect 15976 4093 16024 4128
rect 15976 4059 15983 4093
rect 16017 4059 16024 4093
rect 15976 4024 16024 4059
rect 15976 3990 15983 4024
rect 16017 3990 16024 4024
rect 15976 3955 16024 3990
rect 15976 3921 15983 3955
rect 16017 3921 16024 3955
rect 15976 3897 16024 3921
<< psubdiffcont >>
rect 13925 35947 13959 35981
rect 13996 35947 14030 35981
rect 14067 35947 14101 35981
rect 14138 35947 14172 35981
rect 14209 35947 14243 35981
rect 14280 35947 14314 35981
rect 14351 35947 14385 35981
rect 14422 35947 14456 35981
rect 14493 35947 14527 35981
rect 14563 35947 14597 35981
rect 14633 35947 14667 35981
rect 14703 35947 14737 35981
rect 14773 35947 14807 35981
rect 14843 35947 14877 35981
rect 14913 35947 14947 35981
rect 14983 35947 15017 35981
rect 15053 35947 15087 35981
rect 15123 35947 15157 35981
rect 15193 35947 15227 35981
rect 15263 35947 15297 35981
rect 15333 35947 15367 35981
rect 15403 35947 15437 35981
rect 15473 35947 15507 35981
rect 15543 35947 15577 35981
rect 12875 142 12909 176
rect 12977 142 13011 176
rect 13079 142 13113 176
rect 13181 142 13215 176
rect 12875 74 12909 108
rect 12977 74 13011 108
rect 13079 74 13113 108
rect 13181 74 13215 108
<< mvpsubdiffcont >>
rect 3146 35947 3180 35981
rect 3215 35947 3249 35981
rect 3284 35947 3318 35981
rect 3353 35947 3387 35981
rect 3422 35947 3456 35981
rect 3491 35947 3525 35981
rect 3560 35947 3594 35981
rect 3629 35947 3663 35981
rect 3698 35947 3732 35981
rect 3767 35947 3801 35981
rect 3836 35947 3870 35981
rect 3905 35947 3939 35981
rect 3974 35947 4008 35981
rect 4043 35947 4077 35981
rect 4112 35947 4146 35981
rect 4181 35947 4215 35981
rect 4250 35947 4284 35981
rect 4319 35947 4353 35981
rect 4388 35947 4422 35981
rect 4457 35947 4491 35981
rect 4526 35947 4560 35981
rect 4595 35947 4629 35981
rect 4664 35947 4698 35981
rect 4733 35947 4767 35981
rect 4802 35947 4836 35981
rect 4871 35947 4905 35981
rect 4940 35947 4974 35981
rect 5009 35947 5043 35981
rect 5078 35947 5112 35981
rect 5147 35947 5181 35981
rect 5216 35947 5250 35981
rect 5285 35947 5319 35981
rect 5354 35947 5388 35981
rect 5423 35947 5457 35981
rect 5492 35947 5526 35981
rect 5561 35947 5595 35981
rect 5630 35947 5664 35981
rect 5699 35947 5733 35981
rect 5768 35947 5802 35981
rect 5837 35947 5871 35981
rect 5906 35947 5940 35981
rect 5975 35947 6009 35981
rect 6044 35947 6078 35981
rect 6113 35947 6147 35981
rect 6182 35947 6216 35981
rect 6251 35947 6285 35981
rect 6320 35947 6354 35981
rect 6389 35947 6423 35981
rect 6458 35947 6492 35981
rect 6527 35947 6561 35981
rect 6596 35947 6630 35981
rect 6665 35947 6699 35981
rect 6734 35947 6768 35981
rect 6803 35947 6837 35981
rect 6872 35947 6906 35981
rect 6941 35947 6975 35981
rect 7010 35947 7044 35981
rect 7079 35947 7113 35981
rect 7148 35947 7182 35981
rect 7217 35947 7251 35981
rect 7286 35947 7320 35981
rect 7355 35947 7389 35981
rect 7424 35947 7458 35981
rect 7493 35947 7527 35981
rect 7562 35947 7596 35981
rect 7631 35947 7665 35981
rect 7699 35947 7733 35981
rect 7767 35947 7801 35981
rect 7835 35947 7869 35981
rect 7903 35947 7937 35981
rect 7971 35947 8005 35981
rect 8039 35947 8073 35981
rect 8107 35947 8141 35981
rect 8175 35947 8209 35981
rect 8243 35947 8277 35981
rect 8311 35947 8345 35981
rect 8379 35947 8413 35981
rect 8447 35947 8481 35981
rect 8515 35947 8549 35981
rect 8583 35947 8617 35981
rect 8651 35947 8685 35981
rect 8719 35947 8753 35981
rect 8787 35947 8821 35981
rect 8855 35947 8889 35981
rect 8923 35947 8957 35981
rect 8991 35947 9025 35981
rect 9059 35947 9093 35981
rect 9127 35947 9161 35981
rect 9195 35947 9229 35981
rect 9263 35947 9297 35981
rect 9331 35947 9365 35981
rect 9399 35947 9433 35981
rect 9467 35947 9501 35981
rect 9535 35947 9569 35981
rect 9603 35947 9637 35981
rect 9671 35947 9705 35981
rect 9739 35947 9773 35981
rect 9807 35947 9841 35981
rect 9875 35947 9909 35981
rect 9943 35947 9977 35981
rect 10011 35947 10045 35981
rect 10079 35947 10113 35981
rect 10147 35947 10181 35981
rect 10215 35947 10249 35981
rect 10283 35947 10317 35981
rect 10351 35947 10385 35981
rect 10419 35947 10453 35981
rect 10487 35947 10521 35981
rect 10555 35947 10589 35981
rect 10623 35947 10657 35981
rect 10691 35947 10725 35981
rect 10759 35947 10793 35981
rect 10827 35947 10861 35981
rect 10895 35947 10929 35981
rect 10963 35947 10997 35981
rect 11031 35947 11065 35981
rect 11099 35947 11133 35981
rect 11167 35947 11201 35981
rect 11235 35947 11269 35981
rect 11303 35947 11337 35981
rect 11371 35947 11405 35981
rect 11439 35947 11473 35981
rect 11507 35947 11541 35981
rect 11575 35947 11609 35981
rect 11643 35947 11677 35981
rect 11711 35947 11745 35981
rect 11779 35947 11813 35981
rect 11847 35947 11881 35981
rect 11915 35947 11949 35981
rect 11983 35947 12017 35981
rect 12051 35947 12085 35981
rect 12119 35947 12153 35981
rect 12187 35947 12221 35981
rect 12255 35947 12289 35981
rect 12323 35947 12357 35981
rect 12391 35947 12425 35981
rect 12459 35947 12493 35981
rect 12527 35947 12561 35981
rect 12595 35947 12629 35981
rect 12663 35947 12697 35981
rect 12731 35947 12765 35981
rect 12799 35947 12833 35981
rect 12867 35947 12901 35981
rect 12935 35947 12969 35981
rect 13003 35947 13037 35981
rect 13071 35947 13105 35981
rect 13139 35947 13173 35981
rect 13207 35947 13241 35981
rect 13275 35947 13309 35981
rect 13343 35947 13377 35981
rect 13411 35947 13445 35981
rect 13479 35947 13513 35981
rect 13547 35947 13581 35981
rect 13615 35947 13649 35981
rect 13683 35947 13717 35981
rect 13751 35947 13785 35981
rect -17 25987 17 26021
rect 55 25987 89 26021
rect 127 25987 161 26021
rect 199 25987 233 26021
rect 271 25987 305 26021
rect 343 25987 377 26021
rect 415 25987 449 26021
rect 487 25987 521 26021
rect 559 25987 593 26021
rect 631 25987 665 26021
rect 703 25987 737 26021
rect 775 25987 809 26021
rect 843 26011 877 26045
rect 915 26011 949 26045
rect -17 25918 17 25952
rect 55 25918 89 25952
rect 127 25918 161 25952
rect 199 25918 233 25952
rect 271 25918 305 25952
rect 343 25918 377 25952
rect 415 25918 449 25952
rect 487 25918 521 25952
rect 559 25918 593 25952
rect 631 25918 665 25952
rect 703 25918 737 25952
rect 775 25918 809 25952
rect 843 25938 877 25972
rect 915 25938 949 25972
rect -17 25849 17 25883
rect 55 25849 89 25883
rect 127 25849 161 25883
rect 199 25849 233 25883
rect 271 25849 305 25883
rect 343 25849 377 25883
rect 415 25849 449 25883
rect 487 25849 521 25883
rect 559 25849 593 25883
rect 631 25849 665 25883
rect 703 25849 737 25883
rect 775 25849 809 25883
rect 843 25865 877 25899
rect 915 25865 949 25899
rect -17 25780 17 25814
rect 55 25780 89 25814
rect 127 25780 161 25814
rect 199 25780 233 25814
rect 271 25780 305 25814
rect 343 25780 377 25814
rect 415 25780 449 25814
rect 487 25780 521 25814
rect 559 25780 593 25814
rect 631 25780 665 25814
rect 703 25780 737 25814
rect 775 25780 809 25814
rect 843 25792 877 25826
rect 915 25792 949 25826
rect -17 25711 17 25745
rect 55 25711 89 25745
rect 127 25711 161 25745
rect 199 25711 233 25745
rect 271 25711 305 25745
rect 343 25711 377 25745
rect 415 25711 449 25745
rect 487 25711 521 25745
rect 559 25711 593 25745
rect 631 25711 665 25745
rect 703 25711 737 25745
rect 775 25711 809 25745
rect 843 25719 877 25753
rect 915 25719 949 25753
rect -17 25642 17 25676
rect 55 25642 89 25676
rect 127 25642 161 25676
rect 199 25642 233 25676
rect 271 25642 305 25676
rect 343 25642 377 25676
rect 415 25642 449 25676
rect 487 25642 521 25676
rect 559 25642 593 25676
rect 631 25642 665 25676
rect 703 25642 737 25676
rect 775 25642 809 25676
rect 843 25646 877 25680
rect 915 25646 949 25680
rect -17 25573 17 25607
rect 55 25573 89 25607
rect 127 25573 161 25607
rect 199 25573 233 25607
rect 271 25573 305 25607
rect 343 25573 377 25607
rect 415 25573 449 25607
rect 487 25573 521 25607
rect 559 25573 593 25607
rect 631 25573 665 25607
rect 703 25573 737 25607
rect 775 25573 809 25607
rect 843 25573 877 25607
rect 915 25573 949 25607
rect -17 25505 17 25539
rect 55 25505 89 25539
rect 127 25505 161 25539
rect 199 25505 233 25539
rect 271 25505 305 25539
rect 343 25505 377 25539
rect 415 25505 449 25539
rect 487 25505 521 25539
rect 559 25505 593 25539
rect 631 25505 665 25539
rect 703 25505 737 25539
rect 775 25505 809 25539
rect 843 25500 877 25534
rect 915 25500 949 25534
rect -17 25437 17 25471
rect 55 25437 89 25471
rect 127 25437 161 25471
rect 199 25437 233 25471
rect 271 25437 305 25471
rect 343 25437 377 25471
rect 415 25437 449 25471
rect 487 25437 521 25471
rect 559 25437 593 25471
rect 631 25437 665 25471
rect 703 25437 737 25471
rect 775 25437 809 25471
rect 843 25427 877 25461
rect 915 25427 949 25461
rect -17 25369 17 25403
rect 55 25369 89 25403
rect 127 25369 161 25403
rect 199 25369 233 25403
rect 271 25369 305 25403
rect 343 25369 377 25403
rect 415 25369 449 25403
rect 487 25369 521 25403
rect 559 25369 593 25403
rect 631 25369 665 25403
rect 703 25369 737 25403
rect 775 25369 809 25403
rect 843 25354 877 25388
rect 915 25354 949 25388
rect -17 25301 17 25335
rect 55 25301 89 25335
rect 127 25301 161 25335
rect 199 25301 233 25335
rect 271 25301 305 25335
rect 343 25301 377 25335
rect 415 25301 449 25335
rect 487 25301 521 25335
rect 559 25301 593 25335
rect 631 25301 665 25335
rect 703 25301 737 25335
rect 775 25301 809 25335
rect 843 25282 877 25316
rect 915 25282 949 25316
rect -17 25233 17 25267
rect 55 25233 89 25267
rect 127 25233 161 25267
rect 199 25233 233 25267
rect 271 25233 305 25267
rect 343 25233 377 25267
rect 415 25233 449 25267
rect 487 25233 521 25267
rect 559 25233 593 25267
rect 631 25233 665 25267
rect 703 25233 737 25267
rect 775 25233 809 25267
rect -17 25165 17 25199
rect 55 25165 89 25199
rect 127 25165 161 25199
rect 199 25165 233 25199
rect 271 25165 305 25199
rect 343 25165 377 25199
rect 415 25165 449 25199
rect 487 25165 521 25199
rect 559 25165 593 25199
rect 631 25165 665 25199
rect 703 25165 737 25199
rect 775 25165 809 25199
rect -17 25097 17 25131
rect 55 25097 89 25131
rect 127 25097 161 25131
rect 199 25097 233 25131
rect 271 25097 305 25131
rect 343 25097 377 25131
rect 415 25097 449 25131
rect 487 25097 521 25131
rect 559 25097 593 25131
rect 631 25097 665 25131
rect 703 25097 737 25131
rect 775 25097 809 25131
rect -17 25029 17 25063
rect 55 25029 89 25063
rect 127 25029 161 25063
rect 199 25029 233 25063
rect 271 25029 305 25063
rect 343 25029 377 25063
rect 415 25029 449 25063
rect 487 25029 521 25063
rect 559 25029 593 25063
rect 631 25029 665 25063
rect 703 25029 737 25063
rect 775 25029 809 25063
rect -17 24961 17 24995
rect 55 24961 89 24995
rect 127 24961 161 24995
rect 199 24961 233 24995
rect 271 24961 305 24995
rect 343 24961 377 24995
rect 415 24961 449 24995
rect 487 24961 521 24995
rect 559 24961 593 24995
rect 631 24961 665 24995
rect 703 24961 737 24995
rect 775 24961 809 24995
rect -17 24893 17 24927
rect 55 24893 89 24927
rect 127 24893 161 24927
rect 199 24893 233 24927
rect 271 24893 305 24927
rect 343 24893 377 24927
rect 415 24893 449 24927
rect 487 24893 521 24927
rect 559 24893 593 24927
rect 631 24893 665 24927
rect 703 24893 737 24927
rect 775 24893 809 24927
rect -17 24825 17 24859
rect 55 24825 89 24859
rect 127 24825 161 24859
rect 199 24825 233 24859
rect 271 24825 305 24859
rect 343 24825 377 24859
rect 415 24825 449 24859
rect 487 24825 521 24859
rect 559 24825 593 24859
rect 631 24825 665 24859
rect 703 24825 737 24859
rect 775 24825 809 24859
rect -17 24757 17 24791
rect 55 24757 89 24791
rect 127 24757 161 24791
rect 199 24757 233 24791
rect 271 24757 305 24791
rect 343 24757 377 24791
rect 415 24757 449 24791
rect 487 24757 521 24791
rect 559 24757 593 24791
rect 631 24757 665 24791
rect 703 24757 737 24791
rect 775 24757 809 24791
rect -17 24689 17 24723
rect 55 24689 89 24723
rect 127 24689 161 24723
rect 199 24689 233 24723
rect 271 24689 305 24723
rect 343 24689 377 24723
rect 415 24689 449 24723
rect 487 24689 521 24723
rect 559 24689 593 24723
rect 631 24689 665 24723
rect 703 24689 737 24723
rect 775 24689 809 24723
rect -17 24621 17 24655
rect 55 24621 89 24655
rect 127 24621 161 24655
rect 199 24621 233 24655
rect 271 24621 305 24655
rect 343 24621 377 24655
rect 415 24621 449 24655
rect 487 24621 521 24655
rect 559 24621 593 24655
rect 631 24621 665 24655
rect 703 24621 737 24655
rect 775 24621 809 24655
rect -17 24553 17 24587
rect 55 24553 89 24587
rect 127 24553 161 24587
rect 199 24553 233 24587
rect 271 24553 305 24587
rect 343 24553 377 24587
rect 415 24553 449 24587
rect 487 24553 521 24587
rect 559 24553 593 24587
rect 631 24553 665 24587
rect 703 24553 737 24587
rect 775 24553 809 24587
rect -17 24485 17 24519
rect 55 24485 89 24519
rect 127 24485 161 24519
rect 199 24485 233 24519
rect 271 24485 305 24519
rect 343 24485 377 24519
rect 415 24485 449 24519
rect 487 24485 521 24519
rect 559 24485 593 24519
rect 631 24485 665 24519
rect 703 24485 737 24519
rect 775 24485 809 24519
rect -17 24417 17 24451
rect 55 24417 89 24451
rect 127 24417 161 24451
rect 199 24417 233 24451
rect 271 24417 305 24451
rect 343 24417 377 24451
rect 415 24417 449 24451
rect 487 24417 521 24451
rect 559 24417 593 24451
rect 631 24417 665 24451
rect 703 24417 737 24451
rect 775 24417 809 24451
rect -17 24349 17 24383
rect 55 24349 89 24383
rect 127 24349 161 24383
rect 199 24349 233 24383
rect 271 24349 305 24383
rect 343 24349 377 24383
rect 415 24349 449 24383
rect 487 24349 521 24383
rect 559 24349 593 24383
rect 631 24349 665 24383
rect 703 24349 737 24383
rect 775 24349 809 24383
rect -17 24281 17 24315
rect 55 24281 89 24315
rect 127 24281 161 24315
rect 199 24281 233 24315
rect 271 24281 305 24315
rect 343 24281 377 24315
rect 415 24281 449 24315
rect 487 24281 521 24315
rect 559 24281 593 24315
rect 631 24281 665 24315
rect 703 24281 737 24315
rect 775 24281 809 24315
rect -17 24213 17 24247
rect 55 24213 89 24247
rect 127 24213 161 24247
rect 199 24213 233 24247
rect 271 24213 305 24247
rect 343 24213 377 24247
rect 415 24213 449 24247
rect 487 24213 521 24247
rect 559 24213 593 24247
rect 631 24213 665 24247
rect 703 24213 737 24247
rect 775 24213 809 24247
rect -17 24145 17 24179
rect 55 24145 89 24179
rect 127 24145 161 24179
rect 199 24145 233 24179
rect 271 24145 305 24179
rect 343 24145 377 24179
rect 415 24145 449 24179
rect 487 24145 521 24179
rect 559 24145 593 24179
rect 631 24145 665 24179
rect 703 24145 737 24179
rect 775 24145 809 24179
rect -17 24077 17 24111
rect 55 24077 89 24111
rect 127 24077 161 24111
rect 199 24077 233 24111
rect 271 24077 305 24111
rect 343 24077 377 24111
rect 415 24077 449 24111
rect 487 24077 521 24111
rect 559 24077 593 24111
rect 631 24077 665 24111
rect 703 24077 737 24111
rect 775 24077 809 24111
rect -17 24009 17 24043
rect 55 24009 89 24043
rect 127 24009 161 24043
rect 199 24009 233 24043
rect 271 24009 305 24043
rect 343 24009 377 24043
rect 415 24009 449 24043
rect 487 24009 521 24043
rect 559 24009 593 24043
rect 631 24009 665 24043
rect 703 24009 737 24043
rect 775 24009 809 24043
rect -17 23941 17 23975
rect 55 23941 89 23975
rect 127 23941 161 23975
rect 199 23941 233 23975
rect 271 23941 305 23975
rect 343 23941 377 23975
rect 415 23941 449 23975
rect 487 23941 521 23975
rect 559 23941 593 23975
rect 631 23941 665 23975
rect 703 23941 737 23975
rect 775 23941 809 23975
rect -17 23873 17 23907
rect 55 23873 89 23907
rect 127 23873 161 23907
rect 199 23873 233 23907
rect 271 23873 305 23907
rect 343 23873 377 23907
rect 415 23873 449 23907
rect 487 23873 521 23907
rect 559 23873 593 23907
rect 631 23873 665 23907
rect 703 23873 737 23907
rect 775 23873 809 23907
rect -17 23805 17 23839
rect 55 23805 89 23839
rect 127 23805 161 23839
rect 199 23805 233 23839
rect 271 23805 305 23839
rect 343 23805 377 23839
rect 415 23805 449 23839
rect 487 23805 521 23839
rect 559 23805 593 23839
rect 631 23805 665 23839
rect 703 23805 737 23839
rect 775 23805 809 23839
rect -17 23737 17 23771
rect 55 23737 89 23771
rect 127 23737 161 23771
rect 199 23737 233 23771
rect 271 23737 305 23771
rect 343 23737 377 23771
rect 415 23737 449 23771
rect 487 23737 521 23771
rect 559 23737 593 23771
rect 631 23737 665 23771
rect 703 23737 737 23771
rect 775 23737 809 23771
rect -17 23669 17 23703
rect 55 23669 89 23703
rect 127 23669 161 23703
rect 199 23669 233 23703
rect 271 23669 305 23703
rect 343 23669 377 23703
rect 415 23669 449 23703
rect 487 23669 521 23703
rect 559 23669 593 23703
rect 631 23669 665 23703
rect 703 23669 737 23703
rect 775 23669 809 23703
rect -17 23601 17 23635
rect 55 23601 89 23635
rect 127 23601 161 23635
rect 199 23601 233 23635
rect 271 23601 305 23635
rect 343 23601 377 23635
rect 415 23601 449 23635
rect 487 23601 521 23635
rect 559 23601 593 23635
rect 631 23601 665 23635
rect 703 23601 737 23635
rect 775 23601 809 23635
rect -17 23533 17 23567
rect 55 23533 89 23567
rect 127 23533 161 23567
rect 199 23533 233 23567
rect 271 23533 305 23567
rect 343 23533 377 23567
rect 415 23533 449 23567
rect 487 23533 521 23567
rect 559 23533 593 23567
rect 631 23533 665 23567
rect 703 23533 737 23567
rect 775 23533 809 23567
rect -17 23465 17 23499
rect 55 23465 89 23499
rect 127 23465 161 23499
rect 199 23465 233 23499
rect 271 23465 305 23499
rect 343 23465 377 23499
rect 415 23465 449 23499
rect 487 23465 521 23499
rect 559 23465 593 23499
rect 631 23465 665 23499
rect 703 23465 737 23499
rect 775 23465 809 23499
rect -17 23397 17 23431
rect 55 23397 89 23431
rect 127 23397 161 23431
rect 199 23397 233 23431
rect 271 23397 305 23431
rect 343 23397 377 23431
rect 415 23397 449 23431
rect 487 23397 521 23431
rect 559 23397 593 23431
rect 631 23397 665 23431
rect 703 23397 737 23431
rect 775 23397 809 23431
rect -17 23329 17 23363
rect 55 23329 89 23363
rect 127 23329 161 23363
rect 199 23329 233 23363
rect 271 23329 305 23363
rect 343 23329 377 23363
rect 415 23329 449 23363
rect 487 23329 521 23363
rect 559 23329 593 23363
rect 631 23329 665 23363
rect 703 23329 737 23363
rect 775 23329 809 23363
rect -17 23261 17 23295
rect 55 23261 89 23295
rect 127 23261 161 23295
rect 199 23261 233 23295
rect 271 23261 305 23295
rect 343 23261 377 23295
rect 415 23261 449 23295
rect 487 23261 521 23295
rect 559 23261 593 23295
rect 631 23261 665 23295
rect 703 23261 737 23295
rect 775 23261 809 23295
rect -17 23193 17 23227
rect 55 23193 89 23227
rect 127 23193 161 23227
rect 199 23193 233 23227
rect 271 23193 305 23227
rect 343 23193 377 23227
rect 415 23193 449 23227
rect 487 23193 521 23227
rect 559 23193 593 23227
rect 631 23193 665 23227
rect 703 23193 737 23227
rect 775 23193 809 23227
rect -17 23125 17 23159
rect 55 23125 89 23159
rect 127 23125 161 23159
rect 199 23125 233 23159
rect 271 23125 305 23159
rect 343 23125 377 23159
rect 415 23125 449 23159
rect 487 23125 521 23159
rect 559 23125 593 23159
rect 631 23125 665 23159
rect 703 23125 737 23159
rect 775 23125 809 23159
rect -17 23057 17 23091
rect 55 23057 89 23091
rect 127 23057 161 23091
rect 199 23057 233 23091
rect 271 23057 305 23091
rect 343 23057 377 23091
rect 415 23057 449 23091
rect 487 23057 521 23091
rect 559 23057 593 23091
rect 631 23057 665 23091
rect 703 23057 737 23091
rect 775 23057 809 23091
rect -17 22989 17 23023
rect 55 22989 89 23023
rect 127 22989 161 23023
rect 199 22989 233 23023
rect 271 22989 305 23023
rect 343 22989 377 23023
rect 415 22989 449 23023
rect 487 22989 521 23023
rect 559 22989 593 23023
rect 631 22989 665 23023
rect 703 22989 737 23023
rect 775 22989 809 23023
rect -17 22921 17 22955
rect 55 22921 89 22955
rect 127 22921 161 22955
rect 199 22921 233 22955
rect 271 22921 305 22955
rect 343 22921 377 22955
rect 415 22921 449 22955
rect 487 22921 521 22955
rect 559 22921 593 22955
rect 631 22921 665 22955
rect 703 22921 737 22955
rect 775 22921 809 22955
rect -17 22853 17 22887
rect 55 22853 89 22887
rect 127 22853 161 22887
rect 199 22853 233 22887
rect 271 22853 305 22887
rect 343 22853 377 22887
rect 415 22853 449 22887
rect 487 22853 521 22887
rect 559 22853 593 22887
rect 631 22853 665 22887
rect 703 22853 737 22887
rect 775 22853 809 22887
rect -17 22785 17 22819
rect 55 22785 89 22819
rect 127 22785 161 22819
rect 199 22785 233 22819
rect 271 22785 305 22819
rect 343 22785 377 22819
rect 415 22785 449 22819
rect 487 22785 521 22819
rect 559 22785 593 22819
rect 631 22785 665 22819
rect 703 22785 737 22819
rect 775 22785 809 22819
rect -17 22717 17 22751
rect 55 22717 89 22751
rect 127 22717 161 22751
rect 199 22717 233 22751
rect 271 22717 305 22751
rect 343 22717 377 22751
rect 415 22717 449 22751
rect 487 22717 521 22751
rect 559 22717 593 22751
rect 631 22717 665 22751
rect 703 22717 737 22751
rect 775 22717 809 22751
rect -17 22649 17 22683
rect 55 22649 89 22683
rect 127 22649 161 22683
rect 199 22649 233 22683
rect 271 22649 305 22683
rect 343 22649 377 22683
rect 415 22649 449 22683
rect 487 22649 521 22683
rect 559 22649 593 22683
rect 631 22649 665 22683
rect 703 22649 737 22683
rect 775 22649 809 22683
rect -17 22581 17 22615
rect 55 22581 89 22615
rect 127 22581 161 22615
rect 199 22581 233 22615
rect 271 22581 305 22615
rect 343 22581 377 22615
rect 415 22581 449 22615
rect 487 22581 521 22615
rect 559 22581 593 22615
rect 631 22581 665 22615
rect 703 22581 737 22615
rect 775 22581 809 22615
rect -17 22513 17 22547
rect 55 22513 89 22547
rect 127 22513 161 22547
rect 199 22513 233 22547
rect 271 22513 305 22547
rect 343 22513 377 22547
rect 415 22513 449 22547
rect 487 22513 521 22547
rect 559 22513 593 22547
rect 631 22513 665 22547
rect 703 22513 737 22547
rect 775 22513 809 22547
rect -17 22445 17 22479
rect 55 22445 89 22479
rect 127 22445 161 22479
rect 199 22445 233 22479
rect 271 22445 305 22479
rect 343 22445 377 22479
rect 415 22445 449 22479
rect 487 22445 521 22479
rect 559 22445 593 22479
rect 631 22445 665 22479
rect 703 22445 737 22479
rect 775 22445 809 22479
rect -17 22377 17 22411
rect 55 22377 89 22411
rect 127 22377 161 22411
rect 199 22377 233 22411
rect 271 22377 305 22411
rect 343 22377 377 22411
rect 415 22377 449 22411
rect 487 22377 521 22411
rect 559 22377 593 22411
rect 631 22377 665 22411
rect 703 22377 737 22411
rect 775 22377 809 22411
rect -17 22309 17 22343
rect 55 22309 89 22343
rect 127 22309 161 22343
rect 199 22309 233 22343
rect 271 22309 305 22343
rect 343 22309 377 22343
rect 415 22309 449 22343
rect 487 22309 521 22343
rect 559 22309 593 22343
rect 631 22309 665 22343
rect 703 22309 737 22343
rect 775 22309 809 22343
rect -17 22241 17 22275
rect 55 22241 89 22275
rect 127 22241 161 22275
rect 199 22241 233 22275
rect 271 22241 305 22275
rect 343 22241 377 22275
rect 415 22241 449 22275
rect 487 22241 521 22275
rect 559 22241 593 22275
rect 631 22241 665 22275
rect 703 22241 737 22275
rect 775 22241 809 22275
rect -17 22173 17 22207
rect 55 22173 89 22207
rect 127 22173 161 22207
rect 199 22173 233 22207
rect 271 22173 305 22207
rect 343 22173 377 22207
rect 415 22173 449 22207
rect 487 22173 521 22207
rect 559 22173 593 22207
rect 631 22173 665 22207
rect 703 22173 737 22207
rect 775 22173 809 22207
rect -17 22105 17 22139
rect 55 22105 89 22139
rect 127 22105 161 22139
rect 199 22105 233 22139
rect 271 22105 305 22139
rect 343 22105 377 22139
rect 415 22105 449 22139
rect 487 22105 521 22139
rect 559 22105 593 22139
rect 631 22105 665 22139
rect 703 22105 737 22139
rect 775 22105 809 22139
rect -17 22037 17 22071
rect 55 22037 89 22071
rect 127 22037 161 22071
rect 199 22037 233 22071
rect 271 22037 305 22071
rect 343 22037 377 22071
rect 415 22037 449 22071
rect 487 22037 521 22071
rect 559 22037 593 22071
rect 631 22037 665 22071
rect 703 22037 737 22071
rect 775 22037 809 22071
rect -17 21969 17 22003
rect 55 21969 89 22003
rect 127 21969 161 22003
rect 199 21969 233 22003
rect 271 21969 305 22003
rect 343 21969 377 22003
rect 415 21969 449 22003
rect 487 21969 521 22003
rect 559 21969 593 22003
rect 631 21969 665 22003
rect 703 21969 737 22003
rect 775 21969 809 22003
rect -17 21901 17 21935
rect 55 21901 89 21935
rect 127 21901 161 21935
rect 199 21901 233 21935
rect 271 21901 305 21935
rect 343 21901 377 21935
rect 415 21901 449 21935
rect 487 21901 521 21935
rect 559 21901 593 21935
rect 631 21901 665 21935
rect 703 21901 737 21935
rect 775 21901 809 21935
rect -17 21833 17 21867
rect 55 21833 89 21867
rect 127 21833 161 21867
rect 199 21833 233 21867
rect 271 21833 305 21867
rect 343 21833 377 21867
rect 415 21833 449 21867
rect 487 21833 521 21867
rect 559 21833 593 21867
rect 631 21833 665 21867
rect 703 21833 737 21867
rect 775 21833 809 21867
rect -17 21765 17 21799
rect 55 21765 89 21799
rect 127 21765 161 21799
rect 199 21765 233 21799
rect 271 21765 305 21799
rect 343 21765 377 21799
rect 415 21765 449 21799
rect 487 21765 521 21799
rect 559 21765 593 21799
rect 631 21765 665 21799
rect 703 21765 737 21799
rect 775 21765 809 21799
rect -17 21697 17 21731
rect 55 21697 89 21731
rect 127 21697 161 21731
rect 199 21697 233 21731
rect 271 21697 305 21731
rect 343 21697 377 21731
rect 415 21697 449 21731
rect 487 21697 521 21731
rect 559 21697 593 21731
rect 631 21697 665 21731
rect 703 21697 737 21731
rect 775 21697 809 21731
rect -17 21629 17 21663
rect 55 21629 89 21663
rect 127 21629 161 21663
rect 199 21629 233 21663
rect 271 21629 305 21663
rect 343 21629 377 21663
rect 415 21629 449 21663
rect 487 21629 521 21663
rect 559 21629 593 21663
rect 631 21629 665 21663
rect 703 21629 737 21663
rect 775 21629 809 21663
rect -17 21561 17 21595
rect 55 21561 89 21595
rect 127 21561 161 21595
rect 199 21561 233 21595
rect 271 21561 305 21595
rect 343 21561 377 21595
rect 415 21561 449 21595
rect 487 21561 521 21595
rect 559 21561 593 21595
rect 631 21561 665 21595
rect 703 21561 737 21595
rect 775 21561 809 21595
rect -17 21493 17 21527
rect 55 21493 89 21527
rect 127 21493 161 21527
rect 199 21493 233 21527
rect 271 21493 305 21527
rect 343 21493 377 21527
rect 415 21493 449 21527
rect 487 21493 521 21527
rect 559 21493 593 21527
rect 631 21493 665 21527
rect 703 21493 737 21527
rect 775 21493 809 21527
rect -17 21425 17 21459
rect 55 21425 89 21459
rect 127 21425 161 21459
rect 199 21425 233 21459
rect 271 21425 305 21459
rect 343 21425 377 21459
rect 415 21425 449 21459
rect 487 21425 521 21459
rect 559 21425 593 21459
rect 631 21425 665 21459
rect 703 21425 737 21459
rect 775 21425 809 21459
rect -17 21357 17 21391
rect 55 21357 89 21391
rect 127 21357 161 21391
rect 199 21357 233 21391
rect 271 21357 305 21391
rect 343 21357 377 21391
rect 415 21357 449 21391
rect 487 21357 521 21391
rect 559 21357 593 21391
rect 631 21357 665 21391
rect 703 21357 737 21391
rect 775 21357 809 21391
rect -17 21289 17 21323
rect 55 21289 89 21323
rect 127 21289 161 21323
rect 199 21289 233 21323
rect 271 21289 305 21323
rect 343 21289 377 21323
rect 415 21289 449 21323
rect 487 21289 521 21323
rect 559 21289 593 21323
rect 631 21289 665 21323
rect 703 21289 737 21323
rect 775 21289 809 21323
rect -17 21221 17 21255
rect 55 21221 89 21255
rect 127 21221 161 21255
rect 199 21221 233 21255
rect 271 21221 305 21255
rect 343 21221 377 21255
rect 415 21221 449 21255
rect 487 21221 521 21255
rect 559 21221 593 21255
rect 631 21221 665 21255
rect 703 21221 737 21255
rect 775 21221 809 21255
rect -17 21153 17 21187
rect 55 21153 89 21187
rect 127 21153 161 21187
rect 199 21153 233 21187
rect 271 21153 305 21187
rect 343 21153 377 21187
rect 415 21153 449 21187
rect 487 21153 521 21187
rect 559 21153 593 21187
rect 631 21153 665 21187
rect 703 21153 737 21187
rect 775 21153 809 21187
rect -17 21085 17 21119
rect 55 21085 89 21119
rect 127 21085 161 21119
rect 199 21085 233 21119
rect 271 21085 305 21119
rect 343 21085 377 21119
rect 415 21085 449 21119
rect 487 21085 521 21119
rect 559 21085 593 21119
rect 631 21085 665 21119
rect 703 21085 737 21119
rect 775 21085 809 21119
rect -17 21017 17 21051
rect 55 21017 89 21051
rect 127 21017 161 21051
rect 199 21017 233 21051
rect 271 21017 305 21051
rect 343 21017 377 21051
rect 415 21017 449 21051
rect 487 21017 521 21051
rect 559 21017 593 21051
rect 631 21017 665 21051
rect 703 21017 737 21051
rect 775 21017 809 21051
rect -17 20949 17 20983
rect 55 20949 89 20983
rect 127 20949 161 20983
rect 199 20949 233 20983
rect 271 20949 305 20983
rect 343 20949 377 20983
rect 415 20949 449 20983
rect 487 20949 521 20983
rect 559 20949 593 20983
rect 631 20949 665 20983
rect 703 20949 737 20983
rect 775 20949 809 20983
rect -17 20881 17 20915
rect 55 20881 89 20915
rect 127 20881 161 20915
rect 199 20881 233 20915
rect 271 20881 305 20915
rect 343 20881 377 20915
rect 415 20881 449 20915
rect 487 20881 521 20915
rect 559 20881 593 20915
rect 631 20881 665 20915
rect 703 20881 737 20915
rect 775 20881 809 20915
rect -17 20813 17 20847
rect 55 20813 89 20847
rect 127 20813 161 20847
rect 199 20813 233 20847
rect 271 20813 305 20847
rect 343 20813 377 20847
rect 415 20813 449 20847
rect 487 20813 521 20847
rect 559 20813 593 20847
rect 631 20813 665 20847
rect 703 20813 737 20847
rect 775 20813 809 20847
rect -17 20745 17 20779
rect 55 20745 89 20779
rect 127 20745 161 20779
rect 199 20745 233 20779
rect 271 20745 305 20779
rect 343 20745 377 20779
rect 415 20745 449 20779
rect 487 20745 521 20779
rect 559 20745 593 20779
rect 631 20745 665 20779
rect 703 20745 737 20779
rect 775 20745 809 20779
rect -17 20677 17 20711
rect 55 20677 89 20711
rect 127 20677 161 20711
rect 199 20677 233 20711
rect 271 20677 305 20711
rect 343 20677 377 20711
rect 415 20677 449 20711
rect 487 20677 521 20711
rect 559 20677 593 20711
rect 631 20677 665 20711
rect 703 20677 737 20711
rect 775 20677 809 20711
rect -17 20609 17 20643
rect 55 20609 89 20643
rect 127 20609 161 20643
rect 199 20609 233 20643
rect 271 20609 305 20643
rect 343 20609 377 20643
rect 415 20609 449 20643
rect 487 20609 521 20643
rect 559 20609 593 20643
rect 631 20609 665 20643
rect 703 20609 737 20643
rect 775 20609 809 20643
rect -17 20541 17 20575
rect 55 20541 89 20575
rect 127 20541 161 20575
rect 199 20541 233 20575
rect 271 20541 305 20575
rect 343 20541 377 20575
rect 415 20541 449 20575
rect 487 20541 521 20575
rect 559 20541 593 20575
rect 631 20541 665 20575
rect 703 20541 737 20575
rect 775 20541 809 20575
rect -17 20473 17 20507
rect 55 20473 89 20507
rect 127 20473 161 20507
rect 199 20473 233 20507
rect 271 20473 305 20507
rect 343 20473 377 20507
rect 415 20473 449 20507
rect 487 20473 521 20507
rect 559 20473 593 20507
rect 631 20473 665 20507
rect 703 20473 737 20507
rect 775 20473 809 20507
rect 843 20450 877 20484
rect 915 20450 949 20484
rect -17 20405 17 20439
rect 55 20405 89 20439
rect 127 20405 161 20439
rect 199 20405 233 20439
rect 271 20405 305 20439
rect 343 20405 377 20439
rect 415 20405 449 20439
rect 487 20405 521 20439
rect 559 20405 593 20439
rect 631 20405 665 20439
rect 703 20405 737 20439
rect 775 20415 809 20439
rect -17 20337 17 20371
rect 55 20337 89 20371
rect 127 20337 161 20371
rect 199 20337 233 20371
rect 271 20337 305 20371
rect 343 20337 377 20371
rect 415 20337 449 20371
rect 487 20337 521 20371
rect 559 20337 593 20371
rect 631 20337 665 20371
rect 703 20337 737 20371
rect -17 20269 17 20303
rect 55 20269 89 20303
rect 127 20269 161 20303
rect 199 20269 233 20303
rect 271 20269 305 20303
rect 343 20269 377 20303
rect 415 20269 449 20303
rect 487 20269 521 20303
rect 559 20269 593 20303
rect 631 20269 665 20303
rect 703 20269 737 20303
rect -17 20201 17 20235
rect 55 20201 89 20235
rect 127 20201 161 20235
rect 199 20201 233 20235
rect 271 20201 305 20235
rect 343 20201 377 20235
rect 415 20201 449 20235
rect 487 20201 521 20235
rect 559 20201 593 20235
rect 631 20201 665 20235
rect 703 20201 737 20235
rect -17 20133 17 20167
rect 55 20133 89 20167
rect 127 20133 161 20167
rect 199 20133 233 20167
rect 271 20133 305 20167
rect 343 20133 377 20167
rect 415 20133 449 20167
rect 487 20133 521 20167
rect 559 20133 593 20167
rect 631 20133 665 20167
rect 703 20133 737 20167
rect -17 20065 17 20099
rect 55 20065 89 20099
rect 127 20065 161 20099
rect 199 20065 233 20099
rect 271 20065 305 20099
rect 343 20065 377 20099
rect 415 20065 449 20099
rect 487 20065 521 20099
rect 559 20065 593 20099
rect 631 20065 665 20099
rect 703 20065 737 20099
rect -17 19997 17 20031
rect 55 19997 89 20031
rect 127 19997 161 20031
rect 199 19997 233 20031
rect 271 19997 305 20031
rect 343 19997 377 20031
rect 415 19997 449 20031
rect 487 19997 521 20031
rect 559 19997 593 20031
rect 631 19997 665 20031
rect 703 19997 737 20031
rect -17 19929 17 19963
rect 55 19929 89 19963
rect 127 19929 161 19963
rect 199 19929 233 19963
rect 271 19929 305 19963
rect 343 19929 377 19963
rect 415 19929 449 19963
rect 487 19929 521 19963
rect 559 19929 593 19963
rect 631 19929 665 19963
rect 703 19929 737 19963
rect -17 19861 17 19895
rect 55 19861 89 19895
rect 127 19861 161 19895
rect 199 19861 233 19895
rect 271 19861 305 19895
rect 343 19861 377 19895
rect 415 19861 449 19895
rect 487 19861 521 19895
rect 559 19861 593 19895
rect 631 19861 665 19895
rect 703 19861 737 19895
rect -17 19793 17 19827
rect 55 19793 89 19827
rect 127 19793 161 19827
rect 199 19793 233 19827
rect 271 19793 305 19827
rect 343 19793 377 19827
rect 415 19793 449 19827
rect 487 19793 521 19827
rect 559 19793 593 19827
rect 631 19793 665 19827
rect 703 19793 737 19827
rect -17 19725 17 19759
rect 55 19725 89 19759
rect 127 19725 161 19759
rect 199 19725 233 19759
rect 271 19725 305 19759
rect 343 19725 377 19759
rect 415 19725 449 19759
rect 487 19725 521 19759
rect 559 19725 593 19759
rect 631 19725 665 19759
rect 703 19725 737 19759
rect -17 19657 17 19691
rect 55 19657 89 19691
rect 127 19657 161 19691
rect 199 19657 233 19691
rect 271 19657 305 19691
rect 343 19657 377 19691
rect 415 19657 449 19691
rect 487 19657 521 19691
rect 559 19657 593 19691
rect 631 19657 665 19691
rect 703 19657 737 19691
rect -17 19589 17 19623
rect 55 19589 89 19623
rect 127 19589 161 19623
rect 199 19589 233 19623
rect 271 19589 305 19623
rect 343 19589 377 19623
rect 415 19589 449 19623
rect 487 19589 521 19623
rect 559 19589 593 19623
rect 631 19589 665 19623
rect 703 19589 737 19623
rect -17 19521 17 19555
rect 55 19521 89 19555
rect 127 19521 161 19555
rect 199 19521 233 19555
rect 271 19521 305 19555
rect 343 19521 377 19555
rect 415 19521 449 19555
rect 487 19521 521 19555
rect 559 19521 593 19555
rect 631 19521 665 19555
rect 703 19521 737 19555
rect -17 19453 17 19487
rect 55 19453 89 19487
rect 127 19453 161 19487
rect 199 19453 233 19487
rect 271 19453 305 19487
rect 343 19453 377 19487
rect 415 19453 449 19487
rect 487 19453 521 19487
rect 559 19453 593 19487
rect 631 19453 665 19487
rect 703 19453 737 19487
rect -17 19385 17 19419
rect 55 19385 89 19419
rect 127 19385 161 19419
rect 199 19385 233 19419
rect 271 19385 305 19419
rect 343 19385 377 19419
rect 415 19385 449 19419
rect 487 19385 521 19419
rect 559 19385 593 19419
rect 631 19385 665 19419
rect 703 19385 737 19419
rect -17 19317 17 19351
rect 55 19317 89 19351
rect 127 19317 161 19351
rect 199 19317 233 19351
rect 271 19317 305 19351
rect 343 19317 377 19351
rect 415 19317 449 19351
rect 487 19317 521 19351
rect 559 19317 593 19351
rect 631 19317 665 19351
rect 703 19317 737 19351
rect -17 19249 17 19283
rect 55 19249 89 19283
rect 127 19249 161 19283
rect 199 19249 233 19283
rect 271 19249 305 19283
rect 343 19249 377 19283
rect 415 19249 449 19283
rect 487 19249 521 19283
rect 559 19249 593 19283
rect 631 19249 665 19283
rect 703 19249 737 19283
rect -17 19181 17 19215
rect 55 19181 89 19215
rect 127 19181 161 19215
rect 199 19181 233 19215
rect 271 19181 305 19215
rect 343 19181 377 19215
rect 415 19181 449 19215
rect 487 19181 521 19215
rect 559 19181 593 19215
rect 631 19181 665 19215
rect 703 19181 737 19215
rect -17 19113 17 19147
rect 55 19113 89 19147
rect 127 19113 161 19147
rect 199 19113 233 19147
rect 271 19113 305 19147
rect 343 19113 377 19147
rect 415 19113 449 19147
rect 487 19113 521 19147
rect 559 19113 593 19147
rect 631 19113 665 19147
rect 703 19113 737 19147
rect -17 19045 17 19079
rect 55 19045 89 19079
rect 127 19045 161 19079
rect 199 19045 233 19079
rect 271 19045 305 19079
rect 343 19045 377 19079
rect 415 19045 449 19079
rect 487 19045 521 19079
rect 559 19045 593 19079
rect 631 19045 665 19079
rect 703 19045 737 19079
rect -17 18977 17 19011
rect 55 18977 89 19011
rect 127 18977 161 19011
rect 199 18977 233 19011
rect 271 18977 305 19011
rect 343 18977 377 19011
rect 415 18977 449 19011
rect 487 18977 521 19011
rect 559 18977 593 19011
rect 631 18977 665 19011
rect 703 18977 737 19011
rect -17 18909 17 18943
rect 55 18909 89 18943
rect 127 18909 161 18943
rect 199 18909 233 18943
rect 271 18909 305 18943
rect 343 18909 377 18943
rect 415 18909 449 18943
rect 487 18909 521 18943
rect 559 18909 593 18943
rect 631 18909 665 18943
rect 703 18909 737 18943
rect -17 18841 17 18875
rect 55 18841 89 18875
rect 127 18841 161 18875
rect 199 18841 233 18875
rect 271 18841 305 18875
rect 343 18841 377 18875
rect 415 18841 449 18875
rect 487 18841 521 18875
rect 559 18841 593 18875
rect 631 18841 665 18875
rect 703 18841 737 18875
rect -17 18773 17 18807
rect 55 18773 89 18807
rect 127 18773 161 18807
rect 199 18773 233 18807
rect 271 18773 305 18807
rect 343 18773 377 18807
rect 415 18773 449 18807
rect 487 18773 521 18807
rect 559 18773 593 18807
rect 631 18773 665 18807
rect 703 18773 737 18807
rect -17 18705 17 18739
rect 55 18705 89 18739
rect 127 18705 161 18739
rect 199 18705 233 18739
rect 271 18705 305 18739
rect 343 18705 377 18739
rect 415 18705 449 18739
rect 487 18705 521 18739
rect 559 18705 593 18739
rect 631 18705 665 18739
rect 703 18705 737 18739
rect -17 18637 17 18671
rect 55 18637 89 18671
rect 127 18637 161 18671
rect 199 18637 233 18671
rect 271 18637 305 18671
rect 343 18637 377 18671
rect 415 18637 449 18671
rect 487 18637 521 18671
rect 559 18637 593 18671
rect 631 18637 665 18671
rect 703 18637 737 18671
rect 775 18637 877 20415
rect 915 20381 949 20415
rect 915 20313 949 20347
rect 915 20245 949 20279
rect 915 20177 949 20211
rect 915 20109 949 20143
rect 915 20041 949 20075
rect 915 19973 949 20007
rect 915 19905 949 19939
rect 915 19837 949 19871
rect 915 19769 949 19803
rect 915 19701 949 19735
rect 915 19633 949 19667
rect 915 19565 949 19599
rect 915 19497 949 19531
rect 915 19429 949 19463
rect 915 19361 949 19395
rect 915 19293 949 19327
rect 915 19225 949 19259
rect 843 18613 877 18637
rect 915 19157 949 19191
rect 915 18647 1017 19157
rect 1058 19123 1092 19157
rect 1133 19123 1167 19157
rect 1208 19123 1242 19157
rect 1283 19123 1317 19157
rect 1358 19123 1392 19157
rect 1433 19123 1467 19157
rect 1508 19123 1542 19157
rect 1583 19123 1617 19157
rect 1658 19123 1692 19157
rect 1729 19119 1763 19153
rect 1800 19104 1834 19138
rect 1869 19104 1903 19138
rect 1938 19104 1972 19138
rect 2007 19104 2041 19138
rect 2076 19104 2110 19138
rect 2145 19104 2179 19138
rect 2214 19104 2248 19138
rect 2283 19104 2317 19138
rect 2352 19104 2386 19138
rect 2421 19104 2455 19138
rect 2490 19104 2524 19138
rect 2559 19104 2593 19138
rect 2628 19104 2662 19138
rect 2697 19104 2731 19138
rect 2766 19104 2800 19138
rect 2835 19104 2869 19138
rect 2904 19104 2938 19138
rect 2973 19104 3007 19138
rect 3042 19104 3076 19138
rect 3111 19104 3145 19138
rect 3180 19104 3214 19138
rect 3249 19104 3283 19138
rect 3318 19104 3352 19138
rect 3387 19104 3421 19138
rect 3456 19104 3490 19138
rect 3525 19104 3559 19138
rect 3594 19104 3628 19138
rect 3663 19104 3697 19138
rect 3732 19104 3766 19138
rect 3801 19104 3835 19138
rect 3870 19104 3904 19138
rect 3939 19104 3973 19138
rect 4008 19104 4042 19138
rect 4076 19104 4110 19138
rect 4144 19104 4178 19138
rect 4212 19104 4246 19138
rect 4280 19104 4314 19138
rect 4348 19104 4382 19138
rect 4416 19104 4450 19138
rect 4484 19104 4518 19138
rect 4552 19104 4586 19138
rect 4620 19104 4654 19138
rect 4688 19104 4722 19138
rect 4756 19104 4790 19138
rect 4824 19104 4858 19138
rect 4892 19104 4926 19138
rect 4960 19104 4994 19138
rect 5028 19104 5062 19138
rect 5096 19104 5130 19138
rect 5164 19104 5198 19138
rect 5232 19104 5266 19138
rect 5300 19104 5334 19138
rect 5368 19104 5402 19138
rect 5436 19104 5470 19138
rect 5504 19104 5538 19138
rect 5572 19104 5606 19138
rect 5640 19104 5674 19138
rect 5708 19104 5742 19138
rect 5776 19104 5810 19138
rect 5844 19104 5878 19138
rect 5912 19104 5946 19138
rect 5980 19104 6014 19138
rect 6048 19104 6082 19138
rect 6116 19104 6150 19138
rect 6184 19104 6218 19138
rect 6252 19104 6286 19138
rect 6320 19104 6354 19138
rect 6388 19104 6422 19138
rect 6456 19104 6490 19138
rect 6524 19104 6558 19138
rect 6592 19104 6626 19138
rect 6660 19104 6694 19138
rect 6728 19104 6762 19138
rect 6796 19104 6830 19138
rect 6864 19104 6898 19138
rect 6932 19104 6966 19138
rect 7000 19104 7034 19138
rect 7068 19104 7102 19138
rect 7136 19104 7170 19138
rect 7204 19104 7238 19138
rect 7272 19104 7306 19138
rect 7340 19104 7374 19138
rect 7408 19104 7442 19138
rect 7476 19104 7510 19138
rect 7544 19104 7578 19138
rect 7612 19104 7646 19138
rect 7680 19104 7714 19138
rect 7748 19104 7782 19138
rect 7816 19104 7850 19138
rect 7884 19104 7918 19138
rect 7952 19104 7986 19138
rect 8020 19104 8054 19138
rect 8088 19104 8122 19138
rect 8156 19104 8190 19138
rect 8224 19104 8258 19138
rect 8292 19104 8326 19138
rect 8360 19104 8394 19138
rect 8428 19104 8462 19138
rect 8496 19104 8530 19138
rect 8564 19104 8598 19138
rect 8632 19104 8666 19138
rect 8700 19104 8734 19138
rect 8768 19104 8802 19138
rect 8836 19104 8870 19138
rect 8904 19104 8938 19138
rect 8972 19104 9006 19138
rect 9040 19104 9074 19138
rect 9108 19104 9142 19138
rect 1058 19055 1092 19089
rect 1133 19055 1167 19089
rect 1208 19055 1242 19089
rect 1283 19055 1317 19089
rect 1358 19055 1392 19089
rect 1433 19055 1467 19089
rect 1508 19055 1542 19089
rect 1583 19055 1617 19089
rect 1658 19055 1692 19089
rect 1729 19047 1763 19081
rect 1058 18987 1092 19021
rect 1133 18987 1167 19021
rect 1208 18987 1242 19021
rect 1283 18987 1317 19021
rect 1358 18987 1392 19021
rect 1433 18987 1467 19021
rect 1508 18987 1542 19021
rect 1583 18987 1617 19021
rect 1658 18987 1692 19021
rect 1729 18975 1763 19009
rect 1058 18919 1092 18953
rect 1133 18919 1167 18953
rect 1208 18919 1242 18953
rect 1283 18919 1317 18953
rect 1358 18919 1392 18953
rect 1433 18919 1467 18953
rect 1508 18919 1542 18953
rect 1583 18919 1617 18953
rect 1658 18919 1692 18953
rect 1729 18903 1763 18937
rect 1058 18851 1092 18885
rect 1133 18851 1167 18885
rect 1208 18851 1242 18885
rect 1283 18851 1317 18885
rect 1358 18851 1392 18885
rect 1433 18851 1467 18885
rect 1508 18851 1542 18885
rect 1583 18851 1617 18885
rect 1658 18851 1692 18885
rect 1729 18831 1763 18865
rect 1058 18783 1092 18817
rect 1133 18783 1167 18817
rect 1208 18783 1242 18817
rect 1283 18783 1317 18817
rect 1358 18783 1392 18817
rect 1433 18783 1467 18817
rect 1508 18783 1542 18817
rect 1583 18783 1617 18817
rect 1658 18783 1692 18817
rect 1729 18759 1763 18793
rect 1058 18715 1092 18749
rect 1133 18715 1167 18749
rect 1208 18715 1242 18749
rect 1283 18715 1317 18749
rect 1358 18715 1392 18749
rect 1433 18715 1467 18749
rect 1508 18715 1542 18749
rect 1583 18715 1617 18749
rect 1658 18715 1692 18749
rect 1729 18686 1763 18720
rect 1058 18647 1092 18681
rect 1133 18647 1167 18681
rect 1208 18647 1242 18681
rect 1283 18647 1317 18681
rect 1358 18647 1392 18681
rect 1433 18647 1467 18681
rect 1508 18647 1542 18681
rect 1583 18647 1617 18681
rect 1658 18647 1692 18681
rect 915 18613 949 18647
rect 1729 18613 1763 18647
rect 1332 18543 1366 18577
rect 1412 18543 1446 18577
rect 1492 18543 1526 18577
rect 1572 18543 1606 18577
rect 1652 18543 1686 18577
rect 1732 18543 1766 18577
rect 1332 18475 1366 18509
rect 1412 18475 1446 18509
rect 1492 18475 1526 18509
rect 1572 18475 1606 18509
rect 1652 18475 1686 18509
rect 1732 18475 1766 18509
rect 1332 18407 1366 18441
rect 1412 18407 1446 18441
rect 1492 18407 1526 18441
rect 1572 18407 1606 18441
rect 1652 18407 1686 18441
rect 1732 18407 1766 18441
rect 1332 18339 1366 18373
rect 1412 18339 1446 18373
rect 1492 18339 1526 18373
rect 1572 18339 1606 18373
rect 1652 18339 1686 18373
rect 1732 18339 1766 18373
rect 1332 18271 1366 18305
rect 1412 18271 1446 18305
rect 1492 18271 1526 18305
rect 1572 18271 1606 18305
rect 1652 18271 1686 18305
rect 1732 18271 1766 18305
rect 1332 18203 1366 18237
rect 1412 18203 1446 18237
rect 1492 18203 1526 18237
rect 1572 18203 1606 18237
rect 1652 18203 1686 18237
rect 1732 18203 1766 18237
rect 1332 18135 1366 18169
rect 1412 18135 1446 18169
rect 1492 18135 1526 18169
rect 1572 18135 1606 18169
rect 1652 18135 1686 18169
rect 1732 18135 1766 18169
rect 1332 18066 1366 18100
rect 1412 18066 1446 18100
rect 1492 18066 1526 18100
rect 1572 18066 1606 18100
rect 1652 18066 1686 18100
rect 1732 18066 1766 18100
rect 1332 17997 1366 18031
rect 1412 17997 1446 18031
rect 1492 17997 1526 18031
rect 1572 17997 1606 18031
rect 1652 17997 1686 18031
rect 1732 17997 1766 18031
rect 1332 17928 1366 17962
rect 1412 17928 1446 17962
rect 1492 17928 1526 17962
rect 1572 17928 1606 17962
rect 1652 17928 1686 17962
rect 1732 17928 1766 17962
rect 1332 17859 1366 17893
rect 1412 17859 1446 17893
rect 1492 17859 1526 17893
rect 1572 17859 1606 17893
rect 1652 17859 1686 17893
rect 1732 17859 1766 17893
rect 1332 17790 1366 17824
rect 1412 17790 1446 17824
rect 1492 17790 1526 17824
rect 1572 17790 1606 17824
rect 1652 17790 1686 17824
rect 1732 17790 1766 17824
rect 362 9109 396 9143
rect 433 9109 467 9143
rect 504 9109 538 9143
rect 575 9109 609 9143
rect 646 9109 680 9143
rect 717 9109 751 9143
rect 788 9109 822 9143
rect 859 9109 893 9143
rect 13933 2217 13967 2251
rect 14006 2217 14040 2251
rect 14079 2217 14113 2251
rect 14152 2217 14186 2251
rect 14224 2217 14258 2251
rect 14296 2217 14330 2251
rect 13933 2139 13967 2173
rect 14006 2139 14040 2173
rect 14079 2139 14113 2173
rect 14152 2139 14186 2173
rect 14224 2139 14258 2173
rect 14296 2139 14330 2173
rect 13933 2061 13967 2095
rect 14006 2061 14040 2095
rect 14079 2061 14113 2095
rect 14152 2061 14186 2095
rect 14224 2061 14258 2095
rect 14296 2061 14330 2095
rect 13312 2003 13346 2037
rect 13382 2003 13416 2037
rect 13451 2003 13485 2037
rect 13520 2003 13554 2037
rect 13589 2003 13623 2037
rect 13658 2003 13692 2037
rect 13727 2003 13761 2037
rect 13796 2003 13830 2037
rect 13865 2003 13899 2037
rect 13933 1983 13967 2017
rect 14006 1983 14040 2017
rect 14079 1983 14113 2017
rect 14152 1983 14186 2017
rect 14224 1983 14258 2017
rect 14296 1983 14330 2017
rect 13312 1915 13346 1949
rect 13382 1915 13416 1949
rect 13451 1915 13485 1949
rect 13520 1915 13554 1949
rect 13589 1915 13623 1949
rect 13658 1915 13692 1949
rect 13727 1915 13761 1949
rect 13796 1915 13830 1949
rect 13865 1915 13899 1949
rect 13133 1846 13167 1880
rect 13217 1846 13251 1880
rect 13301 1846 13335 1880
rect 13385 1846 13419 1880
rect 13133 1776 13167 1810
rect 13217 1776 13251 1810
rect 13301 1776 13335 1810
rect 13385 1776 13419 1810
rect 13133 1706 13167 1740
rect 13217 1706 13251 1740
rect 13301 1706 13335 1740
rect 13385 1706 13419 1740
rect 13133 1635 13167 1669
rect 13217 1635 13251 1669
rect 13301 1635 13335 1669
rect 13385 1635 13419 1669
rect 13133 1564 13167 1598
rect 13217 1564 13251 1598
rect 13301 1564 13335 1598
rect 13385 1564 13419 1598
rect 13133 1493 13167 1527
rect 13217 1493 13251 1527
rect 13301 1493 13335 1527
rect 13385 1493 13419 1527
rect 13133 1422 13167 1456
rect 13217 1422 13251 1456
rect 13301 1422 13335 1456
rect 13385 1422 13419 1456
rect 13133 1351 13167 1385
rect 13217 1351 13251 1385
rect 13301 1351 13335 1385
rect 13385 1351 13419 1385
rect 13133 1280 13167 1314
rect 13217 1280 13251 1314
rect 13301 1280 13335 1314
rect 13385 1280 13419 1314
rect 12298 1212 12332 1246
rect 12369 1212 12403 1246
rect 12440 1212 12474 1246
rect 12511 1212 12545 1246
rect 12582 1212 12616 1246
rect 12653 1212 12687 1246
rect 12724 1212 12758 1246
rect 12795 1212 12829 1246
rect 12866 1212 12900 1246
rect 12937 1212 12971 1246
rect 13008 1212 13042 1246
rect 13079 1212 13113 1246
rect 13150 1212 13184 1246
rect 13221 1212 13255 1246
rect 13292 1212 13326 1246
rect 13362 1212 13396 1246
rect 1561 1146 1595 1180
rect 1630 1146 1664 1180
rect 1699 1146 1733 1180
rect 1768 1146 1802 1180
rect 1837 1146 1871 1180
rect 1906 1146 1940 1180
rect 1975 1146 2009 1180
rect 2044 1146 2078 1180
rect 2113 1146 2147 1180
rect 2182 1146 2216 1180
rect 2251 1146 2285 1180
rect 2320 1146 2354 1180
rect 2389 1146 2423 1180
rect 2458 1146 2492 1180
rect 2527 1146 2561 1180
rect 2596 1146 2630 1180
rect 2665 1146 2699 1180
rect 2734 1146 2768 1180
rect 2803 1146 2837 1180
rect 2872 1146 2906 1180
rect 2941 1146 2975 1180
rect 3009 1146 3043 1180
rect 3077 1146 3111 1180
rect 3145 1146 3179 1180
rect 3213 1146 3247 1180
rect 3281 1146 3315 1180
rect 3349 1146 3383 1180
rect 3417 1146 3451 1180
rect 3485 1146 3519 1180
rect 3553 1146 3587 1180
rect 3621 1146 3655 1180
rect 3689 1146 3723 1180
rect 3757 1146 3791 1180
rect 3825 1146 3859 1180
rect 3893 1146 3927 1180
rect 3961 1146 3995 1180
rect 4029 1146 4063 1180
rect 4097 1146 4131 1180
rect 4165 1146 4199 1180
rect 4233 1146 4267 1180
rect 4301 1146 4335 1180
rect 4369 1146 4403 1180
rect 4437 1146 4471 1180
rect 4505 1146 4539 1180
rect 4573 1146 4607 1180
rect 4641 1146 4675 1180
rect 4709 1146 4743 1180
rect 4777 1146 4811 1180
rect 4845 1146 4879 1180
rect 4913 1146 4947 1180
rect 4981 1146 5015 1180
rect 5049 1146 5083 1180
rect 5117 1146 5151 1180
rect 5185 1146 5219 1180
rect 5253 1146 5287 1180
rect 5321 1146 5355 1180
rect 5389 1146 5423 1180
rect 5457 1146 5491 1180
rect 5525 1146 5559 1180
rect 5593 1146 5627 1180
rect 5661 1146 5695 1180
rect 5729 1146 5763 1180
rect 5797 1146 5831 1180
rect 5865 1146 5899 1180
rect 5933 1146 5967 1180
rect 6001 1146 6035 1180
rect 6069 1146 6103 1180
rect 6137 1146 6171 1180
rect 6205 1146 6239 1180
rect 6273 1146 6307 1180
rect 6341 1146 6375 1180
rect 6409 1146 6443 1180
rect 6477 1146 6511 1180
rect 6545 1146 6579 1180
rect 6613 1146 6647 1180
rect 6681 1146 6715 1180
rect 6749 1146 6783 1180
rect 6817 1146 6851 1180
rect 6885 1146 6919 1180
rect 6953 1146 6987 1180
rect 7021 1146 7055 1180
rect 7089 1146 7123 1180
rect 7157 1146 7191 1180
rect 7225 1146 7259 1180
rect 7293 1146 7327 1180
rect 7361 1146 7395 1180
rect 7429 1146 7463 1180
rect 7497 1146 7531 1180
rect 7565 1146 7599 1180
rect 7633 1146 7667 1180
rect 7701 1146 7735 1180
rect 7769 1146 7803 1180
rect 7837 1146 7871 1180
rect 7905 1146 7939 1180
rect 7973 1146 8007 1180
rect 8041 1146 8075 1180
rect 8109 1146 8143 1180
rect 8177 1146 8211 1180
rect 8245 1146 8279 1180
rect 8313 1146 8347 1180
rect 8381 1146 8415 1180
rect 8449 1146 8483 1180
rect 8517 1146 8551 1180
rect 8585 1146 8619 1180
rect 8653 1146 8687 1180
rect 8721 1146 8755 1180
rect 8789 1146 8823 1180
rect 8857 1146 8891 1180
rect 8925 1146 8959 1180
rect 8993 1146 9027 1180
rect 9061 1146 9095 1180
rect 9129 1146 9163 1180
rect 9197 1146 9231 1180
rect 9265 1146 9299 1180
rect 9333 1146 9367 1180
rect 9401 1146 9435 1180
rect 9469 1146 9503 1180
rect 9537 1146 9571 1180
rect 9605 1146 9639 1180
rect 9673 1146 9707 1180
rect 9741 1146 9775 1180
rect 9809 1146 9843 1180
rect 9877 1146 9911 1180
rect 9945 1146 9979 1180
rect 10013 1146 10047 1180
rect 10081 1146 10115 1180
rect 10149 1146 10183 1180
rect 10217 1146 10251 1180
rect 10285 1146 10319 1180
rect 10353 1146 10387 1180
rect 10421 1146 10455 1180
rect 10489 1146 10523 1180
rect 10557 1146 10591 1180
rect 10625 1146 10659 1180
rect 10693 1146 10727 1180
rect 10761 1146 10795 1180
rect 10829 1146 10863 1180
rect 10897 1146 10931 1180
rect 10965 1146 10999 1180
rect 11033 1146 11067 1180
rect 11101 1146 11135 1180
rect 11169 1146 11203 1180
rect 11237 1146 11271 1180
rect 11305 1146 11339 1180
rect 11373 1146 11407 1180
rect 11441 1146 11475 1180
rect 11509 1146 11543 1180
rect 11577 1146 11611 1180
rect 11645 1146 11679 1180
rect 11713 1146 11747 1180
rect 11781 1146 11815 1180
rect 11849 1146 11883 1180
rect 11917 1146 11951 1180
rect 11985 1146 12019 1180
rect 12053 1146 12087 1180
rect 12121 1146 12155 1180
rect 12189 1146 12223 1180
rect 12298 1114 12332 1148
rect 12369 1114 12403 1148
rect 12440 1114 12474 1148
rect 12511 1114 12545 1148
rect 12582 1114 12616 1148
rect 12653 1114 12687 1148
rect 12724 1114 12758 1148
rect 12795 1114 12829 1148
rect 12866 1114 12900 1148
rect 12937 1114 12971 1148
rect 13008 1114 13042 1148
rect 13079 1114 13113 1148
rect 13150 1114 13184 1148
rect 13221 1114 13255 1148
rect 13292 1114 13326 1148
rect 13362 1114 13396 1148
rect 12298 1016 12332 1050
rect 12369 1016 12403 1050
rect 12440 1016 12474 1050
rect 12511 1016 12545 1050
rect 12582 1016 12616 1050
rect 12653 1016 12687 1050
rect 12724 1016 12758 1050
rect 12795 1016 12829 1050
rect 12866 1016 12900 1050
rect 12937 1016 12971 1050
rect 13008 1016 13042 1050
rect 13079 1016 13113 1050
rect 13150 1016 13184 1050
rect 13221 1016 13255 1050
rect 13292 1016 13326 1050
rect 13362 1016 13396 1050
<< mvnsubdiffcont >>
rect -17 35671 17 35705
rect 55 35671 89 35705
rect 127 35671 161 35705
rect 199 35671 233 35705
rect 271 35671 305 35705
rect 343 35671 377 35705
rect 415 35671 449 35705
rect 487 35671 521 35705
rect 559 35671 593 35705
rect 631 35671 665 35705
rect 703 35671 737 35705
rect 775 35671 809 35705
rect 843 35695 877 35729
rect 915 35695 949 35729
rect -17 35603 17 35637
rect 55 35603 89 35637
rect 127 35603 161 35637
rect 199 35603 233 35637
rect 271 35603 305 35637
rect 343 35603 377 35637
rect 415 35603 449 35637
rect 487 35603 521 35637
rect 559 35603 593 35637
rect 631 35603 665 35637
rect 703 35603 737 35637
rect 775 35603 809 35637
rect 843 35611 877 35645
rect 915 35611 949 35645
rect -17 35535 17 35569
rect 55 35535 89 35569
rect 127 35535 161 35569
rect 199 35535 233 35569
rect 271 35535 305 35569
rect 343 35535 377 35569
rect 415 35535 449 35569
rect 487 35535 521 35569
rect 559 35535 593 35569
rect 631 35535 665 35569
rect 703 35535 737 35569
rect 775 35535 809 35569
rect 843 35527 877 35561
rect 915 35527 949 35561
rect -17 35467 17 35501
rect 55 35467 89 35501
rect 127 35467 161 35501
rect 199 35467 233 35501
rect 271 35467 305 35501
rect 343 35467 377 35501
rect 415 35467 449 35501
rect 487 35467 521 35501
rect 559 35467 593 35501
rect 631 35467 665 35501
rect 703 35467 737 35501
rect 775 35467 809 35501
rect 843 35443 877 35477
rect 915 35443 949 35477
rect -17 35399 17 35433
rect 55 35399 89 35433
rect 127 35399 161 35433
rect 199 35399 233 35433
rect 271 35399 305 35433
rect 343 35399 377 35433
rect 415 35399 449 35433
rect 487 35399 521 35433
rect 559 35399 593 35433
rect 631 35399 665 35433
rect 703 35399 737 35433
rect 775 35399 809 35433
rect -17 35331 17 35365
rect 55 35331 89 35365
rect 127 35331 161 35365
rect 199 35331 233 35365
rect 271 35331 305 35365
rect 343 35331 377 35365
rect 415 35331 449 35365
rect 487 35331 521 35365
rect 559 35331 593 35365
rect 631 35331 665 35365
rect 703 35331 737 35365
rect 775 35331 809 35365
rect 843 35359 877 35393
rect 915 35359 949 35393
rect -17 35263 17 35297
rect 55 35263 89 35297
rect 127 35263 161 35297
rect 199 35263 233 35297
rect 271 35263 305 35297
rect 343 35263 377 35297
rect 415 35263 449 35297
rect 487 35263 521 35297
rect 559 35263 593 35297
rect 631 35263 665 35297
rect 703 35263 737 35297
rect 775 35263 809 35297
rect 843 35275 877 35309
rect 915 35275 949 35309
rect -17 35195 17 35229
rect 55 35195 89 35229
rect 127 35195 161 35229
rect 199 35195 233 35229
rect 271 35195 305 35229
rect 343 35195 377 35229
rect 415 35195 449 35229
rect 487 35195 521 35229
rect 559 35195 593 35229
rect 631 35195 665 35229
rect 703 35195 737 35229
rect 775 35195 809 35229
rect 843 35191 877 35225
rect 915 35191 949 35225
rect -17 35127 17 35161
rect 55 35127 89 35161
rect 127 35127 161 35161
rect 199 35127 233 35161
rect 271 35127 305 35161
rect 343 35127 377 35161
rect 415 35127 449 35161
rect 487 35127 521 35161
rect 559 35127 593 35161
rect 631 35127 665 35161
rect 703 35127 737 35161
rect 775 35127 809 35161
rect 843 35107 877 35141
rect 915 35107 949 35141
rect -17 35059 17 35093
rect 55 35059 89 35093
rect 127 35059 161 35093
rect 199 35059 233 35093
rect 271 35059 305 35093
rect 343 35059 377 35093
rect 415 35059 449 35093
rect 487 35059 521 35093
rect 559 35059 593 35093
rect 631 35059 665 35093
rect 703 35059 737 35093
rect 775 35059 809 35093
rect -17 34991 17 35025
rect 55 34991 89 35025
rect 127 34991 161 35025
rect 199 34991 233 35025
rect 271 34991 305 35025
rect 343 34991 377 35025
rect 415 34991 449 35025
rect 487 34991 521 35025
rect 559 34991 593 35025
rect 631 34991 665 35025
rect 703 34991 737 35025
rect 775 34991 809 35025
rect 843 35023 877 35057
rect 915 35023 949 35057
rect -17 34923 17 34957
rect 55 34923 89 34957
rect 127 34923 161 34957
rect 199 34923 233 34957
rect 271 34923 305 34957
rect 343 34923 377 34957
rect 415 34923 449 34957
rect 487 34923 521 34957
rect 559 34923 593 34957
rect 631 34923 665 34957
rect 703 34923 737 34957
rect 775 34923 809 34957
rect 843 34939 877 34973
rect 915 34939 949 34973
rect -17 34855 17 34889
rect 55 34855 89 34889
rect 127 34855 161 34889
rect 199 34855 233 34889
rect 271 34855 305 34889
rect 343 34855 377 34889
rect 415 34855 449 34889
rect 487 34855 521 34889
rect 559 34855 593 34889
rect 631 34855 665 34889
rect 703 34855 737 34889
rect 775 34855 809 34889
rect 843 34855 877 34889
rect 915 34855 949 34889
rect -17 34787 17 34821
rect 55 34787 89 34821
rect 127 34787 161 34821
rect 199 34787 233 34821
rect 271 34787 305 34821
rect 343 34787 377 34821
rect 415 34787 449 34821
rect 487 34787 521 34821
rect 559 34787 593 34821
rect 631 34787 665 34821
rect 703 34787 737 34821
rect 775 34787 809 34821
rect 843 34771 877 34805
rect 915 34771 949 34805
rect -17 34719 17 34753
rect 55 34719 89 34753
rect 127 34719 161 34753
rect 199 34719 233 34753
rect 271 34719 305 34753
rect 343 34719 377 34753
rect 415 34719 449 34753
rect 487 34719 521 34753
rect 559 34719 593 34753
rect 631 34719 665 34753
rect 703 34719 737 34753
rect 775 34719 809 34753
rect 843 34687 877 34721
rect 915 34687 949 34721
rect -17 34651 17 34685
rect 55 34651 89 34685
rect 127 34651 161 34685
rect 199 34651 233 34685
rect 271 34651 305 34685
rect 343 34651 377 34685
rect 415 34651 449 34685
rect 487 34651 521 34685
rect 559 34651 593 34685
rect 631 34651 665 34685
rect 703 34651 737 34685
rect 775 34651 809 34685
rect -17 34583 17 34617
rect 55 34583 89 34617
rect 127 34583 161 34617
rect 199 34583 233 34617
rect 271 34583 305 34617
rect 343 34583 377 34617
rect 415 34583 449 34617
rect 487 34583 521 34617
rect 559 34583 593 34617
rect 631 34583 665 34617
rect 703 34583 737 34617
rect 775 34583 809 34617
rect 843 34603 877 34637
rect 915 34603 949 34637
rect -17 34515 17 34549
rect 55 34515 89 34549
rect 127 34515 161 34549
rect 199 34515 233 34549
rect 271 34515 305 34549
rect 343 34515 377 34549
rect 415 34515 449 34549
rect 487 34515 521 34549
rect 559 34515 593 34549
rect 631 34515 665 34549
rect 703 34515 737 34549
rect 775 34515 809 34549
rect 843 34519 877 34553
rect 915 34519 949 34553
rect -17 34447 17 34481
rect 55 34447 89 34481
rect 127 34447 161 34481
rect 199 34447 233 34481
rect 271 34447 305 34481
rect 343 34447 377 34481
rect 415 34447 449 34481
rect 487 34447 521 34481
rect 559 34447 593 34481
rect 631 34447 665 34481
rect 703 34447 737 34481
rect 775 34447 809 34481
rect 843 34435 877 34469
rect 915 34435 949 34469
rect -17 34379 17 34413
rect 55 34379 89 34413
rect 127 34379 161 34413
rect 199 34379 233 34413
rect 271 34379 305 34413
rect 343 34379 377 34413
rect 415 34379 449 34413
rect 487 34379 521 34413
rect 559 34379 593 34413
rect 631 34379 665 34413
rect 703 34379 737 34413
rect 775 34379 809 34413
rect 843 34351 877 34385
rect 915 34351 949 34385
rect -17 34311 17 34345
rect 55 34311 89 34345
rect 127 34311 161 34345
rect 199 34311 233 34345
rect 271 34311 305 34345
rect 343 34311 377 34345
rect 415 34311 449 34345
rect 487 34311 521 34345
rect 559 34311 593 34345
rect 631 34311 665 34345
rect 703 34311 737 34345
rect 775 34311 809 34345
rect -17 34243 17 34277
rect 55 34243 89 34277
rect 127 34243 161 34277
rect 199 34243 233 34277
rect 271 34243 305 34277
rect 343 34243 377 34277
rect 415 34243 449 34277
rect 487 34243 521 34277
rect 559 34243 593 34277
rect 631 34243 665 34277
rect 703 34243 737 34277
rect 775 34243 809 34277
rect 843 34267 877 34301
rect 915 34267 949 34301
rect -17 34175 17 34209
rect 55 34175 89 34209
rect 127 34175 161 34209
rect 199 34175 233 34209
rect 271 34175 305 34209
rect 343 34175 377 34209
rect 415 34175 449 34209
rect 487 34175 521 34209
rect 559 34175 593 34209
rect 631 34175 665 34209
rect 703 34175 737 34209
rect 775 34175 809 34209
rect 843 34183 877 34217
rect 915 34183 949 34217
rect -17 34107 17 34141
rect 55 34107 89 34141
rect 127 34107 161 34141
rect 199 34107 233 34141
rect 271 34107 305 34141
rect 343 34107 377 34141
rect 415 34107 449 34141
rect 487 34107 521 34141
rect 559 34107 593 34141
rect 631 34107 665 34141
rect 703 34107 737 34141
rect 775 34107 809 34141
rect 843 34099 877 34133
rect 915 34099 949 34133
rect -17 34039 17 34073
rect 55 34039 89 34073
rect 127 34039 161 34073
rect 199 34039 233 34073
rect 271 34039 305 34073
rect 343 34039 377 34073
rect 415 34039 449 34073
rect 487 34039 521 34073
rect 559 34039 593 34073
rect 631 34039 665 34073
rect 703 34039 737 34073
rect 775 34039 809 34073
rect 843 34015 877 34049
rect 915 34015 949 34049
rect -17 33971 17 34005
rect 55 33971 89 34005
rect 127 33971 161 34005
rect 199 33971 233 34005
rect 271 33971 305 34005
rect 343 33971 377 34005
rect 415 33971 449 34005
rect 487 33971 521 34005
rect 559 33971 593 34005
rect 631 33971 665 34005
rect 703 33971 737 34005
rect 775 33971 809 34005
rect -17 33903 17 33937
rect 55 33903 89 33937
rect 127 33903 161 33937
rect 199 33903 233 33937
rect 271 33903 305 33937
rect 343 33903 377 33937
rect 415 33903 449 33937
rect 487 33903 521 33937
rect 559 33903 593 33937
rect 631 33903 665 33937
rect 703 33903 737 33937
rect 775 33903 809 33937
rect 843 33931 877 33965
rect 915 33931 949 33965
rect -17 33835 17 33869
rect 55 33835 89 33869
rect 127 33835 161 33869
rect 199 33835 233 33869
rect 271 33835 305 33869
rect 343 33835 377 33869
rect 415 33835 449 33869
rect 487 33835 521 33869
rect 559 33835 593 33869
rect 631 33835 665 33869
rect 703 33835 737 33869
rect 775 33835 809 33869
rect 843 33847 877 33881
rect 915 33847 949 33881
rect -17 33767 17 33801
rect 55 33767 89 33801
rect 127 33767 161 33801
rect 199 33767 233 33801
rect 271 33767 305 33801
rect 343 33767 377 33801
rect 415 33767 449 33801
rect 487 33767 521 33801
rect 559 33767 593 33801
rect 631 33767 665 33801
rect 703 33767 737 33801
rect 775 33767 809 33801
rect 843 33763 877 33797
rect 915 33763 949 33797
rect -17 33699 17 33733
rect 55 33699 89 33733
rect 127 33699 161 33733
rect 199 33699 233 33733
rect 271 33699 305 33733
rect 343 33699 377 33733
rect 415 33699 449 33733
rect 487 33699 521 33733
rect 559 33699 593 33733
rect 631 33699 665 33733
rect 703 33699 737 33733
rect 775 33699 809 33733
rect 843 33679 877 33713
rect 915 33679 949 33713
rect -17 33631 17 33665
rect 55 33631 89 33665
rect 127 33631 161 33665
rect 199 33631 233 33665
rect 271 33631 305 33665
rect 343 33631 377 33665
rect 415 33631 449 33665
rect 487 33631 521 33665
rect 559 33631 593 33665
rect 631 33631 665 33665
rect 703 33631 737 33665
rect 775 33631 809 33665
rect -17 33563 17 33597
rect 55 33563 89 33597
rect 127 33563 161 33597
rect 199 33563 233 33597
rect 271 33563 305 33597
rect 343 33563 377 33597
rect 415 33563 449 33597
rect 487 33563 521 33597
rect 559 33563 593 33597
rect 631 33563 665 33597
rect 703 33563 737 33597
rect 775 33563 809 33597
rect 843 33595 877 33629
rect 915 33595 949 33629
rect -17 33495 17 33529
rect 55 33495 89 33529
rect 127 33495 161 33529
rect 199 33495 233 33529
rect 271 33495 305 33529
rect 343 33495 377 33529
rect 415 33495 449 33529
rect 487 33495 521 33529
rect 559 33495 593 33529
rect 631 33495 665 33529
rect 703 33495 737 33529
rect 775 33495 809 33529
rect 843 33511 877 33545
rect 915 33511 949 33545
rect -17 33427 17 33461
rect 55 33427 89 33461
rect 127 33427 161 33461
rect 199 33427 233 33461
rect 271 33427 305 33461
rect 343 33427 377 33461
rect 415 33427 449 33461
rect 487 33427 521 33461
rect 559 33427 593 33461
rect 631 33427 665 33461
rect 703 33427 737 33461
rect 775 33427 809 33461
rect 843 33427 877 33461
rect 915 33427 949 33461
rect -17 33359 17 33393
rect 55 33359 89 33393
rect 127 33359 161 33393
rect 199 33359 233 33393
rect 271 33359 305 33393
rect 343 33359 377 33393
rect 415 33359 449 33393
rect 487 33359 521 33393
rect 559 33359 593 33393
rect 631 33359 665 33393
rect 703 33359 737 33393
rect 775 33359 809 33393
rect 843 33343 877 33377
rect 915 33343 949 33377
rect -17 33291 17 33325
rect 55 33291 89 33325
rect 127 33291 161 33325
rect 199 33291 233 33325
rect 271 33291 305 33325
rect 343 33291 377 33325
rect 415 33291 449 33325
rect 487 33291 521 33325
rect 559 33291 593 33325
rect 631 33291 665 33325
rect 703 33291 737 33325
rect 775 33291 809 33325
rect 843 33259 877 33293
rect 915 33259 949 33293
rect -17 33223 17 33257
rect 55 33223 89 33257
rect 127 33223 161 33257
rect 199 33223 233 33257
rect 271 33223 305 33257
rect 343 33223 377 33257
rect 415 33223 449 33257
rect 487 33223 521 33257
rect 559 33223 593 33257
rect 631 33223 665 33257
rect 703 33223 737 33257
rect 775 33223 809 33257
rect -17 33155 17 33189
rect 55 33155 89 33189
rect 127 33155 161 33189
rect 199 33155 233 33189
rect 271 33155 305 33189
rect 343 33155 377 33189
rect 415 33155 449 33189
rect 487 33155 521 33189
rect 559 33155 593 33189
rect 631 33155 665 33189
rect 703 33155 737 33189
rect 775 33155 809 33189
rect 843 33175 877 33209
rect 915 33175 949 33209
rect -17 33087 17 33121
rect 55 33087 89 33121
rect 127 33087 161 33121
rect 199 33087 233 33121
rect 271 33087 305 33121
rect 343 33087 377 33121
rect 415 33087 449 33121
rect 487 33087 521 33121
rect 559 33087 593 33121
rect 631 33087 665 33121
rect 703 33087 737 33121
rect 775 33087 809 33121
rect 843 33091 877 33125
rect 915 33091 949 33125
rect -17 33019 17 33053
rect 55 33019 89 33053
rect 127 33019 161 33053
rect 199 33019 233 33053
rect 271 33019 305 33053
rect 343 33019 377 33053
rect 415 33019 449 33053
rect 487 33019 521 33053
rect 559 33019 593 33053
rect 631 33019 665 33053
rect 703 33019 737 33053
rect 775 33019 809 33053
rect 843 33007 877 33041
rect 915 33007 949 33041
rect -17 32951 17 32985
rect 55 32951 89 32985
rect 127 32951 161 32985
rect 199 32951 233 32985
rect 271 32951 305 32985
rect 343 32951 377 32985
rect 415 32951 449 32985
rect 487 32951 521 32985
rect 559 32951 593 32985
rect 631 32951 665 32985
rect 703 32951 737 32985
rect 775 32951 809 32985
rect 843 32923 877 32957
rect 915 32923 949 32957
rect -17 32883 17 32917
rect 55 32883 89 32917
rect 127 32883 161 32917
rect 199 32883 233 32917
rect 271 32883 305 32917
rect 343 32883 377 32917
rect 415 32883 449 32917
rect 487 32883 521 32917
rect 559 32883 593 32917
rect 631 32883 665 32917
rect 703 32883 737 32917
rect 775 32883 809 32917
rect -17 32815 17 32849
rect 55 32815 89 32849
rect 127 32815 161 32849
rect 199 32815 233 32849
rect 271 32815 305 32849
rect 343 32815 377 32849
rect 415 32815 449 32849
rect 487 32815 521 32849
rect 559 32815 593 32849
rect 631 32815 665 32849
rect 703 32815 737 32849
rect 775 32815 809 32849
rect 843 32839 877 32873
rect 915 32839 949 32873
rect -17 32747 17 32781
rect 55 32747 89 32781
rect 127 32747 161 32781
rect 199 32747 233 32781
rect 271 32747 305 32781
rect 343 32747 377 32781
rect 415 32747 449 32781
rect 487 32747 521 32781
rect 559 32747 593 32781
rect 631 32747 665 32781
rect 703 32747 737 32781
rect 775 32747 809 32781
rect 843 32755 877 32789
rect 915 32755 949 32789
rect -17 32679 17 32713
rect 55 32679 89 32713
rect 127 32679 161 32713
rect 199 32679 233 32713
rect 271 32679 305 32713
rect 343 32679 377 32713
rect 415 32679 449 32713
rect 487 32679 521 32713
rect 559 32679 593 32713
rect 631 32679 665 32713
rect 703 32679 737 32713
rect 775 32679 809 32713
rect 843 32671 877 32705
rect 915 32671 949 32705
rect -17 32611 17 32645
rect 55 32611 89 32645
rect 127 32611 161 32645
rect 199 32611 233 32645
rect 271 32611 305 32645
rect 343 32611 377 32645
rect 415 32611 449 32645
rect 487 32611 521 32645
rect 559 32611 593 32645
rect 631 32611 665 32645
rect 703 32611 737 32645
rect 775 32611 809 32645
rect 843 32587 877 32621
rect 915 32587 949 32621
rect -17 32543 17 32577
rect 55 32543 89 32577
rect 127 32543 161 32577
rect 199 32543 233 32577
rect 271 32543 305 32577
rect 343 32543 377 32577
rect 415 32543 449 32577
rect 487 32543 521 32577
rect 559 32543 593 32577
rect 631 32543 665 32577
rect 703 32543 737 32577
rect 775 32543 809 32577
rect -17 32475 17 32509
rect 55 32475 89 32509
rect 127 32475 161 32509
rect 199 32475 233 32509
rect 271 32475 305 32509
rect 343 32475 377 32509
rect 415 32475 449 32509
rect 487 32475 521 32509
rect 559 32475 593 32509
rect 631 32475 665 32509
rect 703 32475 737 32509
rect 775 32475 809 32509
rect 843 32503 877 32537
rect 915 32503 949 32537
rect -17 32407 17 32441
rect 55 32407 89 32441
rect 127 32407 161 32441
rect 199 32407 233 32441
rect 271 32407 305 32441
rect 343 32407 377 32441
rect 415 32407 449 32441
rect 487 32407 521 32441
rect 559 32407 593 32441
rect 631 32407 665 32441
rect 703 32407 737 32441
rect 775 32407 809 32441
rect 843 32419 877 32453
rect 915 32419 949 32453
rect -17 32339 17 32373
rect 55 32339 89 32373
rect 127 32339 161 32373
rect 199 32339 233 32373
rect 271 32339 305 32373
rect 343 32339 377 32373
rect 415 32339 449 32373
rect 487 32339 521 32373
rect 559 32339 593 32373
rect 631 32339 665 32373
rect 703 32339 737 32373
rect 775 32339 809 32373
rect 843 32335 877 32369
rect 915 32335 949 32369
rect -17 32271 17 32305
rect 55 32271 89 32305
rect 127 32271 161 32305
rect 199 32271 233 32305
rect 271 32271 305 32305
rect 343 32271 377 32305
rect 415 32271 449 32305
rect 487 32271 521 32305
rect 559 32271 593 32305
rect 631 32271 665 32305
rect 703 32271 737 32305
rect 775 32271 809 32305
rect 843 32251 877 32285
rect 915 32251 949 32285
rect -17 32203 17 32237
rect 55 32203 89 32237
rect 127 32203 161 32237
rect 199 32203 233 32237
rect 271 32203 305 32237
rect 343 32203 377 32237
rect 415 32203 449 32237
rect 487 32203 521 32237
rect 559 32203 593 32237
rect 631 32203 665 32237
rect 703 32203 737 32237
rect 775 32203 809 32237
rect -17 32135 17 32169
rect 55 32135 89 32169
rect 127 32135 161 32169
rect 199 32135 233 32169
rect 271 32135 305 32169
rect 343 32135 377 32169
rect 415 32135 449 32169
rect 487 32135 521 32169
rect 559 32135 593 32169
rect 631 32135 665 32169
rect 703 32135 737 32169
rect 775 32135 809 32169
rect 843 32167 877 32201
rect 915 32167 949 32201
rect -17 32067 17 32101
rect 55 32067 89 32101
rect 127 32067 161 32101
rect 199 32067 233 32101
rect 271 32067 305 32101
rect 343 32067 377 32101
rect 415 32067 449 32101
rect 487 32067 521 32101
rect 559 32067 593 32101
rect 631 32067 665 32101
rect 703 32067 737 32101
rect 775 32067 809 32101
rect 843 32083 877 32117
rect 915 32083 949 32117
rect -17 31999 17 32033
rect 55 31999 89 32033
rect 127 31999 161 32033
rect 199 31999 233 32033
rect 271 31999 305 32033
rect 343 31999 377 32033
rect 415 31999 449 32033
rect 487 31999 521 32033
rect 559 31999 593 32033
rect 631 31999 665 32033
rect 703 31999 737 32033
rect 775 31999 809 32033
rect 843 31999 877 32033
rect 915 31999 949 32033
rect -17 31931 17 31965
rect 55 31931 89 31965
rect 127 31931 161 31965
rect 199 31931 233 31965
rect 271 31931 305 31965
rect 343 31931 377 31965
rect 415 31931 449 31965
rect 487 31931 521 31965
rect 559 31931 593 31965
rect 631 31931 665 31965
rect 703 31931 737 31965
rect 775 31931 809 31965
rect 843 31915 877 31949
rect 915 31915 949 31949
rect -17 31863 17 31897
rect 55 31863 89 31897
rect 127 31863 161 31897
rect 199 31863 233 31897
rect 271 31863 305 31897
rect 343 31863 377 31897
rect 415 31863 449 31897
rect 487 31863 521 31897
rect 559 31863 593 31897
rect 631 31863 665 31897
rect 703 31863 737 31897
rect 775 31863 809 31897
rect 843 31831 877 31865
rect 915 31831 949 31865
rect -17 31795 17 31829
rect 55 31795 89 31829
rect 127 31795 161 31829
rect 199 31795 233 31829
rect 271 31795 305 31829
rect 343 31795 377 31829
rect 415 31795 449 31829
rect 487 31795 521 31829
rect 559 31795 593 31829
rect 631 31795 665 31829
rect 703 31795 737 31829
rect 775 31795 809 31829
rect -17 31727 17 31761
rect 55 31727 89 31761
rect 127 31727 161 31761
rect 199 31727 233 31761
rect 271 31727 305 31761
rect 343 31727 377 31761
rect 415 31727 449 31761
rect 487 31727 521 31761
rect 559 31727 593 31761
rect 631 31727 665 31761
rect 703 31727 737 31761
rect 775 31727 809 31761
rect 843 31747 877 31781
rect 915 31747 949 31781
rect -17 31659 17 31693
rect 55 31659 89 31693
rect 127 31659 161 31693
rect 199 31659 233 31693
rect 271 31659 305 31693
rect 343 31659 377 31693
rect 415 31659 449 31693
rect 487 31659 521 31693
rect 559 31659 593 31693
rect 631 31659 665 31693
rect 703 31659 737 31693
rect 775 31659 809 31693
rect 843 31663 877 31697
rect 915 31663 949 31697
rect -17 31591 17 31625
rect 55 31591 89 31625
rect 127 31591 161 31625
rect 199 31591 233 31625
rect 271 31591 305 31625
rect 343 31591 377 31625
rect 415 31591 449 31625
rect 487 31591 521 31625
rect 559 31591 593 31625
rect 631 31591 665 31625
rect 703 31591 737 31625
rect 775 31591 809 31625
rect 843 31579 877 31613
rect 915 31579 949 31613
rect -17 31523 17 31557
rect 55 31523 89 31557
rect 127 31523 161 31557
rect 199 31523 233 31557
rect 271 31523 305 31557
rect 343 31523 377 31557
rect 415 31523 449 31557
rect 487 31523 521 31557
rect 559 31523 593 31557
rect 631 31523 665 31557
rect 703 31523 737 31557
rect 775 31523 809 31557
rect 843 31495 877 31529
rect 915 31495 949 31529
rect -17 31455 17 31489
rect 55 31455 89 31489
rect 127 31455 161 31489
rect 199 31455 233 31489
rect 271 31455 305 31489
rect 343 31455 377 31489
rect 415 31455 449 31489
rect 487 31455 521 31489
rect 559 31455 593 31489
rect 631 31455 665 31489
rect 703 31455 737 31489
rect 775 31455 809 31489
rect -17 31387 17 31421
rect 55 31387 89 31421
rect 127 31387 161 31421
rect 199 31387 233 31421
rect 271 31387 305 31421
rect 343 31387 377 31421
rect 415 31387 449 31421
rect 487 31387 521 31421
rect 559 31387 593 31421
rect 631 31387 665 31421
rect 703 31387 737 31421
rect 775 31387 809 31421
rect 843 31411 877 31445
rect 915 31411 949 31445
rect -17 31319 17 31353
rect 55 31319 89 31353
rect 127 31319 161 31353
rect 199 31319 233 31353
rect 271 31319 305 31353
rect 343 31319 377 31353
rect 415 31319 449 31353
rect 487 31319 521 31353
rect 559 31319 593 31353
rect 631 31319 665 31353
rect 703 31319 737 31353
rect 775 31319 809 31353
rect 843 31327 877 31361
rect 915 31327 949 31361
rect -17 31251 17 31285
rect 55 31251 89 31285
rect 127 31251 161 31285
rect 199 31251 233 31285
rect 271 31251 305 31285
rect 343 31251 377 31285
rect 415 31251 449 31285
rect 487 31251 521 31285
rect 559 31251 593 31285
rect 631 31251 665 31285
rect 703 31251 737 31285
rect 775 31251 809 31285
rect 843 31243 877 31277
rect 915 31243 949 31277
rect -17 31183 17 31217
rect 55 31183 89 31217
rect 127 31183 161 31217
rect 199 31183 233 31217
rect 271 31183 305 31217
rect 343 31183 377 31217
rect 415 31183 449 31217
rect 487 31183 521 31217
rect 559 31183 593 31217
rect 631 31183 665 31217
rect 703 31183 737 31217
rect 775 31183 809 31217
rect 843 31159 877 31193
rect 915 31159 949 31193
rect -17 31115 17 31149
rect 55 31115 89 31149
rect 127 31115 161 31149
rect 199 31115 233 31149
rect 271 31115 305 31149
rect 343 31115 377 31149
rect 415 31115 449 31149
rect 487 31115 521 31149
rect 559 31115 593 31149
rect 631 31115 665 31149
rect 703 31115 737 31149
rect 775 31115 809 31149
rect -17 31047 17 31081
rect 55 31047 89 31081
rect 127 31047 161 31081
rect 199 31047 233 31081
rect 271 31047 305 31081
rect 343 31047 377 31081
rect 415 31047 449 31081
rect 487 31047 521 31081
rect 559 31047 593 31081
rect 631 31047 665 31081
rect 703 31047 737 31081
rect 775 31047 809 31081
rect 843 31075 877 31109
rect 915 31075 949 31109
rect -17 30979 17 31013
rect 55 30979 89 31013
rect 127 30979 161 31013
rect 199 30979 233 31013
rect 271 30979 305 31013
rect 343 30979 377 31013
rect 415 30979 449 31013
rect 487 30979 521 31013
rect 559 30979 593 31013
rect 631 30979 665 31013
rect 703 30979 737 31013
rect 775 30979 809 31013
rect 843 30991 877 31025
rect 915 30991 949 31025
rect -17 30911 17 30945
rect 55 30911 89 30945
rect 127 30911 161 30945
rect 199 30911 233 30945
rect 271 30911 305 30945
rect 343 30911 377 30945
rect 415 30911 449 30945
rect 487 30911 521 30945
rect 559 30911 593 30945
rect 631 30911 665 30945
rect 703 30911 737 30945
rect 775 30911 809 30945
rect 843 30907 877 30941
rect 915 30907 949 30941
rect -17 30843 17 30877
rect 55 30843 89 30877
rect 127 30843 161 30877
rect 199 30843 233 30877
rect 271 30843 305 30877
rect 343 30843 377 30877
rect 415 30843 449 30877
rect 487 30843 521 30877
rect 559 30843 593 30877
rect 631 30843 665 30877
rect 703 30843 737 30877
rect 775 30843 809 30877
rect 843 30823 877 30857
rect 915 30823 949 30857
rect -17 30775 17 30809
rect 55 30775 89 30809
rect 127 30775 161 30809
rect 199 30775 233 30809
rect 271 30775 305 30809
rect 343 30775 377 30809
rect 415 30775 449 30809
rect 487 30775 521 30809
rect 559 30775 593 30809
rect 631 30775 665 30809
rect 703 30775 737 30809
rect 775 30775 809 30809
rect -17 30707 17 30741
rect 55 30707 89 30741
rect 127 30707 161 30741
rect 199 30707 233 30741
rect 271 30707 305 30741
rect 343 30707 377 30741
rect 415 30707 449 30741
rect 487 30707 521 30741
rect 559 30707 593 30741
rect 631 30707 665 30741
rect 703 30707 737 30741
rect 775 30707 809 30741
rect 843 30739 877 30773
rect 915 30739 949 30773
rect -17 30639 17 30673
rect 55 30639 89 30673
rect 127 30639 161 30673
rect 199 30639 233 30673
rect 271 30639 305 30673
rect 343 30639 377 30673
rect 415 30639 449 30673
rect 487 30639 521 30673
rect 559 30639 593 30673
rect 631 30639 665 30673
rect 703 30639 737 30673
rect 775 30639 809 30673
rect 843 30655 877 30689
rect 915 30655 949 30689
rect -17 30571 17 30605
rect 55 30571 89 30605
rect 127 30571 161 30605
rect 199 30571 233 30605
rect 271 30571 305 30605
rect 343 30571 377 30605
rect 415 30571 449 30605
rect 487 30571 521 30605
rect 559 30571 593 30605
rect 631 30571 665 30605
rect 703 30571 737 30605
rect 775 30571 809 30605
rect 843 30571 877 30605
rect 915 30571 949 30605
rect -17 30503 17 30537
rect 55 30503 89 30537
rect 127 30503 161 30537
rect 199 30503 233 30537
rect 271 30503 305 30537
rect 343 30503 377 30537
rect 415 30503 449 30537
rect 487 30503 521 30537
rect 559 30503 593 30537
rect 631 30503 665 30537
rect 703 30503 737 30537
rect 775 30503 809 30537
rect 843 30487 877 30521
rect 915 30487 949 30521
rect -17 30435 17 30469
rect 55 30435 89 30469
rect 127 30435 161 30469
rect 199 30435 233 30469
rect 271 30435 305 30469
rect 343 30435 377 30469
rect 415 30435 449 30469
rect 487 30435 521 30469
rect 559 30435 593 30469
rect 631 30435 665 30469
rect 703 30435 737 30469
rect 775 30435 809 30469
rect 843 30402 877 30436
rect 915 30402 949 30436
rect -17 30367 17 30401
rect 55 30367 89 30401
rect 127 30367 161 30401
rect 199 30367 233 30401
rect 271 30367 305 30401
rect 343 30367 377 30401
rect 415 30367 449 30401
rect 487 30367 521 30401
rect 559 30367 593 30401
rect 631 30367 665 30401
rect 703 30367 737 30401
rect 775 30367 809 30401
rect -17 30299 17 30333
rect 55 30299 89 30333
rect 127 30299 161 30333
rect 199 30299 233 30333
rect 271 30299 305 30333
rect 343 30299 377 30333
rect 415 30299 449 30333
rect 487 30299 521 30333
rect 559 30299 593 30333
rect 631 30299 665 30333
rect 703 30299 737 30333
rect 775 30299 809 30333
rect 843 30317 877 30351
rect 915 30317 949 30351
rect -17 30231 17 30265
rect 55 30231 89 30265
rect 127 30231 161 30265
rect 199 30231 233 30265
rect 271 30231 305 30265
rect 343 30231 377 30265
rect 415 30231 449 30265
rect 487 30231 521 30265
rect 559 30231 593 30265
rect 631 30231 665 30265
rect 703 30231 737 30265
rect 775 30231 809 30265
rect 843 30232 877 30266
rect 915 30232 949 30266
rect -17 30163 17 30197
rect 55 30163 89 30197
rect 127 30163 161 30197
rect 199 30163 233 30197
rect 271 30163 305 30197
rect 343 30163 377 30197
rect 415 30163 449 30197
rect 487 30163 521 30197
rect 559 30163 593 30197
rect 631 30163 665 30197
rect 703 30163 737 30197
rect 775 30163 809 30197
rect 843 30147 877 30181
rect 915 30147 949 30181
rect -17 30095 17 30129
rect 55 30095 89 30129
rect 127 30095 161 30129
rect 199 30095 233 30129
rect 271 30095 305 30129
rect 343 30095 377 30129
rect 415 30095 449 30129
rect 487 30095 521 30129
rect 559 30095 593 30129
rect 631 30095 665 30129
rect 703 30095 737 30129
rect 775 30095 809 30129
rect 843 30062 877 30096
rect 915 30062 949 30096
rect -17 30027 17 30061
rect 55 30027 89 30061
rect 127 30027 161 30061
rect 199 30027 233 30061
rect 271 30027 305 30061
rect 343 30027 377 30061
rect 415 30027 449 30061
rect 487 30027 521 30061
rect 559 30027 593 30061
rect 631 30027 665 30061
rect 703 30027 737 30061
rect 775 30027 809 30061
rect -17 29959 17 29993
rect 55 29959 89 29993
rect 127 29959 161 29993
rect 199 29959 233 29993
rect 271 29959 305 29993
rect 343 29959 377 29993
rect 415 29959 449 29993
rect 487 29959 521 29993
rect 559 29959 593 29993
rect 631 29959 665 29993
rect 703 29959 737 29993
rect 775 29959 809 29993
rect 843 29977 877 30011
rect 915 29977 949 30011
rect -17 29891 17 29925
rect 55 29891 89 29925
rect 127 29891 161 29925
rect 199 29891 233 29925
rect 271 29891 305 29925
rect 343 29891 377 29925
rect 415 29891 449 29925
rect 487 29891 521 29925
rect 559 29891 593 29925
rect 631 29891 665 29925
rect 703 29891 737 29925
rect 775 29891 809 29925
rect 843 29892 877 29926
rect 915 29892 949 29926
rect -17 29823 17 29857
rect 55 29823 89 29857
rect 127 29823 161 29857
rect 199 29823 233 29857
rect 271 29823 305 29857
rect 343 29823 377 29857
rect 415 29823 449 29857
rect 487 29823 521 29857
rect 559 29823 593 29857
rect 631 29823 665 29857
rect 703 29823 737 29857
rect 775 29823 809 29857
rect 843 29807 877 29841
rect 915 29807 949 29841
rect -17 29755 17 29789
rect 55 29755 89 29789
rect 127 29755 161 29789
rect 199 29755 233 29789
rect 271 29755 305 29789
rect 343 29755 377 29789
rect 415 29755 449 29789
rect 487 29755 521 29789
rect 559 29755 593 29789
rect 631 29755 665 29789
rect 703 29755 737 29789
rect 775 29755 809 29789
rect 843 29722 877 29756
rect 915 29722 949 29756
rect -17 29687 17 29721
rect 55 29687 89 29721
rect 127 29687 161 29721
rect 199 29687 233 29721
rect 271 29687 305 29721
rect 343 29687 377 29721
rect 415 29687 449 29721
rect 487 29687 521 29721
rect 559 29687 593 29721
rect 631 29687 665 29721
rect 703 29687 737 29721
rect 775 29687 809 29721
rect -17 29618 17 29652
rect 55 29618 89 29652
rect 127 29618 161 29652
rect 199 29618 233 29652
rect 271 29618 305 29652
rect 343 29618 377 29652
rect 415 29618 449 29652
rect 487 29618 521 29652
rect 559 29618 593 29652
rect 631 29618 665 29652
rect 703 29618 737 29652
rect 775 29618 809 29652
rect 843 29637 877 29671
rect 915 29637 949 29671
rect -17 29549 17 29583
rect 55 29549 89 29583
rect 127 29549 161 29583
rect 199 29549 233 29583
rect 271 29549 305 29583
rect 343 29549 377 29583
rect 415 29549 449 29583
rect 487 29549 521 29583
rect 559 29549 593 29583
rect 631 29549 665 29583
rect 703 29549 737 29583
rect 775 29549 809 29583
rect 843 29552 877 29586
rect 915 29552 949 29586
rect -17 29480 17 29514
rect 55 29480 89 29514
rect 127 29480 161 29514
rect 199 29480 233 29514
rect 271 29480 305 29514
rect 343 29480 377 29514
rect 415 29480 449 29514
rect 487 29480 521 29514
rect 559 29480 593 29514
rect 631 29480 665 29514
rect 703 29480 737 29514
rect 775 29480 809 29514
rect 843 29467 877 29501
rect 915 29467 949 29501
rect -17 29411 17 29445
rect 55 29411 89 29445
rect 127 29411 161 29445
rect 199 29411 233 29445
rect 271 29411 305 29445
rect 343 29411 377 29445
rect 415 29411 449 29445
rect 487 29411 521 29445
rect 559 29411 593 29445
rect 631 29411 665 29445
rect 703 29411 737 29445
rect 775 29411 809 29445
rect 843 29382 877 29416
rect 915 29382 949 29416
rect -17 29342 17 29376
rect 55 29342 89 29376
rect 127 29342 161 29376
rect 199 29342 233 29376
rect 271 29342 305 29376
rect 343 29342 377 29376
rect 415 29342 449 29376
rect 487 29342 521 29376
rect 559 29342 593 29376
rect 631 29342 665 29376
rect 703 29342 737 29376
rect 775 29342 809 29376
rect -17 29273 17 29307
rect 55 29273 89 29307
rect 127 29273 161 29307
rect 199 29273 233 29307
rect 271 29273 305 29307
rect 343 29273 377 29307
rect 415 29273 449 29307
rect 487 29273 521 29307
rect 559 29273 593 29307
rect 631 29273 665 29307
rect 703 29273 737 29307
rect 775 29273 809 29307
rect 843 29297 877 29331
rect 915 29297 949 29331
rect -17 29204 17 29238
rect 55 29204 89 29238
rect 127 29204 161 29238
rect 199 29204 233 29238
rect 271 29204 305 29238
rect 343 29204 377 29238
rect 415 29204 449 29238
rect 487 29204 521 29238
rect 559 29204 593 29238
rect 631 29204 665 29238
rect 703 29204 737 29238
rect 775 29204 809 29238
rect 843 29212 877 29246
rect 915 29212 949 29246
rect -17 29135 17 29169
rect 55 29135 89 29169
rect 127 29135 161 29169
rect 199 29135 233 29169
rect 271 29135 305 29169
rect 343 29135 377 29169
rect 415 29135 449 29169
rect 487 29135 521 29169
rect 559 29135 593 29169
rect 631 29135 665 29169
rect 703 29135 737 29169
rect 775 29135 809 29169
rect 843 29127 877 29161
rect 915 29127 949 29161
rect -17 29066 17 29100
rect 55 29066 89 29100
rect 127 29066 161 29100
rect 199 29066 233 29100
rect 271 29066 305 29100
rect 343 29066 377 29100
rect 415 29066 449 29100
rect 487 29066 521 29100
rect 559 29066 593 29100
rect 631 29066 665 29100
rect 703 29066 737 29100
rect 775 29066 809 29100
rect 843 29042 877 29076
rect 915 29042 949 29076
rect -17 27952 17 27986
rect 55 27952 89 27986
rect 127 27952 161 27986
rect 199 27952 233 27986
rect 271 27952 305 27986
rect 343 27952 377 27986
rect 415 27952 449 27986
rect 487 27952 521 27986
rect 559 27952 593 27986
rect 631 27952 665 27986
rect 703 27952 737 27986
rect 775 27952 809 27986
rect 843 27976 877 28010
rect 915 27976 949 28010
rect -17 27883 17 27917
rect 55 27883 89 27917
rect 127 27883 161 27917
rect 199 27883 233 27917
rect 271 27883 305 27917
rect 343 27883 377 27917
rect 415 27883 449 27917
rect 487 27883 521 27917
rect 559 27883 593 27917
rect 631 27883 665 27917
rect 703 27883 737 27917
rect 775 27883 809 27917
rect 843 27908 877 27942
rect 915 27908 949 27942
rect -17 27814 17 27848
rect 55 27814 89 27848
rect 127 27814 161 27848
rect 199 27814 233 27848
rect 271 27814 305 27848
rect 343 27814 377 27848
rect 415 27814 449 27848
rect 487 27814 521 27848
rect 559 27814 593 27848
rect 631 27814 665 27848
rect 703 27814 737 27848
rect 775 27814 809 27848
rect 843 27840 877 27874
rect 915 27840 949 27874
rect -17 27745 17 27779
rect 55 27745 89 27779
rect 127 27745 161 27779
rect 199 27745 233 27779
rect 271 27745 305 27779
rect 343 27745 377 27779
rect 415 27745 449 27779
rect 487 27745 521 27779
rect 559 27745 593 27779
rect 631 27745 665 27779
rect 703 27745 737 27779
rect 775 27745 809 27779
rect 843 27772 877 27806
rect 915 27772 949 27806
rect -17 27676 17 27710
rect 55 27676 89 27710
rect 127 27676 161 27710
rect 199 27676 233 27710
rect 271 27676 305 27710
rect 343 27676 377 27710
rect 415 27676 449 27710
rect 487 27676 521 27710
rect 559 27676 593 27710
rect 631 27676 665 27710
rect 703 27676 737 27710
rect 775 27676 809 27710
rect 843 27704 877 27738
rect 915 27704 949 27738
rect -17 27607 17 27641
rect 55 27607 89 27641
rect 127 27607 161 27641
rect 199 27607 233 27641
rect 271 27607 305 27641
rect 343 27607 377 27641
rect 415 27607 449 27641
rect 487 27607 521 27641
rect 559 27607 593 27641
rect 631 27607 665 27641
rect 703 27607 737 27641
rect 775 27607 809 27641
rect 843 27636 877 27670
rect 915 27636 949 27670
rect -17 27538 17 27572
rect 55 27538 89 27572
rect 127 27538 161 27572
rect 199 27538 233 27572
rect 271 27538 305 27572
rect 343 27538 377 27572
rect 415 27538 449 27572
rect 487 27538 521 27572
rect 559 27538 593 27572
rect 631 27538 665 27572
rect 703 27538 737 27572
rect 775 27538 809 27572
rect 843 27568 877 27602
rect 915 27568 949 27602
rect -17 27469 17 27503
rect 55 27469 89 27503
rect 127 27469 161 27503
rect 199 27469 233 27503
rect 271 27469 305 27503
rect 343 27469 377 27503
rect 415 27469 449 27503
rect 487 27469 521 27503
rect 559 27469 593 27503
rect 631 27469 665 27503
rect 703 27469 737 27503
rect 775 27469 809 27503
rect 843 27500 877 27534
rect 915 27500 949 27534
rect -17 27400 17 27434
rect 55 27400 89 27434
rect 127 27400 161 27434
rect 199 27400 233 27434
rect 271 27400 305 27434
rect 343 27400 377 27434
rect 415 27400 449 27434
rect 487 27400 521 27434
rect 559 27400 593 27434
rect 631 27400 665 27434
rect 703 27400 737 27434
rect 775 27400 809 27434
rect 843 27432 877 27466
rect 915 27432 949 27466
rect -17 27331 17 27365
rect 55 27331 89 27365
rect 127 27331 161 27365
rect 199 27331 233 27365
rect 271 27331 305 27365
rect 343 27331 377 27365
rect 415 27331 449 27365
rect 487 27331 521 27365
rect 559 27331 593 27365
rect 631 27331 665 27365
rect 703 27331 737 27365
rect 775 27331 809 27365
rect 843 27364 877 27398
rect 915 27364 949 27398
rect 843 27296 877 27330
rect 915 27296 949 27330
rect -17 27262 17 27296
rect 55 27262 89 27296
rect 127 27262 161 27296
rect 199 27262 233 27296
rect 271 27262 305 27296
rect 343 27262 377 27296
rect 415 27262 449 27296
rect 487 27262 521 27296
rect 559 27262 593 27296
rect 631 27262 665 27296
rect 703 27262 737 27296
rect 775 27262 809 27296
rect 843 27228 877 27262
rect 915 27228 949 27262
rect -17 27193 17 27227
rect 55 27193 89 27227
rect 127 27193 161 27227
rect 199 27193 233 27227
rect 271 27193 305 27227
rect 343 27193 377 27227
rect 415 27193 449 27227
rect 487 27193 521 27227
rect 559 27193 593 27227
rect 631 27193 665 27227
rect 703 27193 737 27227
rect 775 27193 809 27227
rect 843 27160 877 27194
rect 915 27160 949 27194
rect -17 27124 17 27158
rect 55 27124 89 27158
rect 127 27124 161 27158
rect 199 27124 233 27158
rect 271 27124 305 27158
rect 343 27124 377 27158
rect 415 27124 449 27158
rect 487 27124 521 27158
rect 559 27124 593 27158
rect 631 27124 665 27158
rect 703 27124 737 27158
rect 775 27124 809 27158
rect 843 27092 877 27126
rect 915 27092 949 27126
rect -17 27055 17 27089
rect 55 27055 89 27089
rect 127 27055 161 27089
rect 199 27055 233 27089
rect 271 27055 305 27089
rect 343 27055 377 27089
rect 415 27055 449 27089
rect 487 27055 521 27089
rect 559 27055 593 27089
rect 631 27055 665 27089
rect 703 27055 737 27089
rect 775 27055 809 27089
rect 843 27024 877 27058
rect 915 27024 949 27058
rect -17 26986 17 27020
rect 55 26986 89 27020
rect 127 26986 161 27020
rect 199 26986 233 27020
rect 271 26986 305 27020
rect 343 26986 377 27020
rect 415 26986 449 27020
rect 487 26986 521 27020
rect 559 26986 593 27020
rect 631 26986 665 27020
rect 703 26986 737 27020
rect 775 26986 809 27020
rect 843 26956 877 26990
rect 915 26956 949 26990
rect -17 26917 17 26951
rect 55 26917 89 26951
rect 127 26917 161 26951
rect 199 26917 233 26951
rect 271 26917 305 26951
rect 343 26917 377 26951
rect 415 26917 449 26951
rect 487 26917 521 26951
rect 559 26917 593 26951
rect 631 26917 665 26951
rect 703 26917 737 26951
rect 775 26917 809 26951
rect 843 26888 877 26922
rect 915 26888 949 26922
rect -17 26848 17 26882
rect 55 26848 89 26882
rect 127 26848 161 26882
rect 199 26848 233 26882
rect 271 26848 305 26882
rect 343 26848 377 26882
rect 415 26848 449 26882
rect 487 26848 521 26882
rect 559 26848 593 26882
rect 631 26848 665 26882
rect 703 26848 737 26882
rect 775 26848 809 26882
rect 843 26820 877 26854
rect 915 26820 949 26854
rect -17 26779 17 26813
rect 55 26779 89 26813
rect 127 26779 161 26813
rect 199 26779 233 26813
rect 271 26779 305 26813
rect 343 26779 377 26813
rect 415 26779 449 26813
rect 487 26779 521 26813
rect 559 26779 593 26813
rect 631 26779 665 26813
rect 703 26779 737 26813
rect 775 26779 809 26813
rect 843 26751 877 26785
rect 915 26751 949 26785
rect -17 26710 17 26744
rect 55 26710 89 26744
rect 127 26710 161 26744
rect 199 26710 233 26744
rect 271 26710 305 26744
rect 343 26710 377 26744
rect 415 26710 449 26744
rect 487 26710 521 26744
rect 559 26710 593 26744
rect 631 26710 665 26744
rect 703 26710 737 26744
rect 775 26710 809 26744
rect 843 26682 877 26716
rect 915 26682 949 26716
rect -17 26641 17 26675
rect 55 26641 89 26675
rect 127 26641 161 26675
rect 199 26641 233 26675
rect 271 26641 305 26675
rect 343 26641 377 26675
rect 415 26641 449 26675
rect 487 26641 521 26675
rect 559 26641 593 26675
rect 631 26641 665 26675
rect 703 26641 737 26675
rect 775 26641 809 26675
rect 843 26613 877 26647
rect 915 26613 949 26647
rect -17 26572 17 26606
rect 55 26572 89 26606
rect 127 26572 161 26606
rect 199 26572 233 26606
rect 271 26572 305 26606
rect 343 26572 377 26606
rect 415 26572 449 26606
rect 487 26572 521 26606
rect 559 26572 593 26606
rect 631 26572 665 26606
rect 703 26572 737 26606
rect 775 26572 809 26606
rect 843 26544 877 26578
rect 915 26544 949 26578
rect -17 26503 17 26537
rect 55 26503 89 26537
rect 127 26503 161 26537
rect 199 26503 233 26537
rect 271 26503 305 26537
rect 343 26503 377 26537
rect 415 26503 449 26537
rect 487 26503 521 26537
rect 559 26503 593 26537
rect 631 26503 665 26537
rect 703 26503 737 26537
rect 775 26503 809 26537
rect 843 26475 877 26509
rect 915 26475 949 26509
rect -17 26433 17 26467
rect 55 26433 89 26467
rect 127 26433 161 26467
rect 199 26433 233 26467
rect 271 26433 305 26467
rect 343 26433 377 26467
rect 415 26433 449 26467
rect 487 26433 521 26467
rect 559 26433 593 26467
rect 631 26433 665 26467
rect 703 26433 737 26467
rect 775 26433 809 26467
rect 843 26406 877 26440
rect 915 26406 949 26440
rect -17 26363 17 26397
rect 55 26363 89 26397
rect 127 26363 161 26397
rect 199 26363 233 26397
rect 271 26363 305 26397
rect 343 26363 377 26397
rect 415 26363 449 26397
rect 487 26363 521 26397
rect 559 26363 593 26397
rect 631 26363 665 26397
rect 703 26363 737 26397
rect 775 26363 809 26397
rect 843 26337 877 26371
rect 915 26337 949 26371
rect -17 26293 17 26327
rect 55 26293 89 26327
rect 127 26293 161 26327
rect 199 26293 233 26327
rect 271 26293 305 26327
rect 343 26293 377 26327
rect 415 26293 449 26327
rect 487 26293 521 26327
rect 559 26293 593 26327
rect 631 26293 665 26327
rect 703 26293 737 26327
rect 775 26293 809 26327
rect 843 26268 877 26302
rect 915 26268 949 26302
rect -17 26223 17 26257
rect 55 26223 89 26257
rect 127 26223 161 26257
rect 199 26223 233 26257
rect 271 26223 305 26257
rect 343 26223 377 26257
rect 415 26223 449 26257
rect 487 26223 521 26257
rect 559 26223 593 26257
rect 631 26223 665 26257
rect 703 26223 737 26257
rect 775 26223 809 26257
rect 843 26199 877 26233
rect 915 26199 949 26233
rect 15983 7087 16017 7121
rect 15983 7018 16017 7052
rect 15983 6949 16017 6983
rect 15983 6880 16017 6914
rect 15983 6811 16017 6845
rect 15983 6742 16017 6776
rect 15983 6673 16017 6707
rect 15983 6604 16017 6638
rect 15983 6535 16017 6569
rect 15983 6466 16017 6500
rect 15983 6397 16017 6431
rect 15983 6327 16017 6361
rect 15983 6257 16017 6291
rect 15983 6187 16017 6221
rect 15983 6117 16017 6151
rect 15983 6047 16017 6081
rect 15983 4945 16017 4979
rect 15983 4877 16017 4911
rect 15983 4809 16017 4843
rect 15983 4741 16017 4775
rect 15983 4673 16017 4707
rect 15983 4605 16017 4639
rect 15983 4537 16017 4571
rect 15983 4469 16017 4503
rect 15983 4401 16017 4435
rect 15983 4333 16017 4367
rect 15983 4265 16017 4299
rect 15983 4197 16017 4231
rect 15983 4128 16017 4162
rect 15983 4059 16017 4093
rect 15983 3990 16017 4024
rect 15983 3921 16017 3955
<< locali >>
rect 8771 36041 8900 36074
rect 11345 36041 11461 36074
rect 3146 35996 13785 36041
rect 13925 35996 15577 36041
rect 3146 35981 3157 35996
rect 3191 35981 3230 35996
rect 3264 35981 3303 35996
rect 3337 35981 3376 35996
rect 3410 35981 3449 35996
rect 3483 35981 3522 35996
rect 3556 35981 3595 35996
rect 3191 35962 3215 35981
rect 3264 35962 3284 35981
rect 3337 35962 3353 35981
rect 3410 35962 3422 35981
rect 3483 35962 3491 35981
rect 3556 35962 3560 35981
rect 3180 35947 3215 35962
rect 3249 35947 3284 35962
rect 3318 35947 3353 35962
rect 3387 35947 3422 35962
rect 3456 35947 3491 35962
rect 3525 35947 3560 35962
rect 3594 35962 3595 35981
rect 3629 35981 3668 35996
rect 3702 35981 3741 35996
rect 3775 35981 3814 35996
rect 3848 35981 3887 35996
rect 3921 35981 3960 35996
rect 3994 35981 4033 35996
rect 4067 35981 4106 35996
rect 4140 35981 4179 35996
rect 4213 35981 4252 35996
rect 4286 35981 4325 35996
rect 4359 35981 4398 35996
rect 4432 35981 4471 35996
rect 4505 35981 4544 35996
rect 4578 35981 4617 35996
rect 4651 35981 4690 35996
rect 4724 35981 4763 35996
rect 4797 35981 4836 35996
rect 3594 35947 3629 35962
rect 3663 35962 3668 35981
rect 3732 35962 3741 35981
rect 3801 35962 3814 35981
rect 3870 35962 3887 35981
rect 3939 35962 3960 35981
rect 4008 35962 4033 35981
rect 4077 35962 4106 35981
rect 4146 35962 4179 35981
rect 3663 35947 3698 35962
rect 3732 35947 3767 35962
rect 3801 35947 3836 35962
rect 3870 35947 3905 35962
rect 3939 35947 3974 35962
rect 4008 35947 4043 35962
rect 4077 35947 4112 35962
rect 4146 35947 4181 35962
rect 4215 35947 4250 35981
rect 4286 35962 4319 35981
rect 4359 35962 4388 35981
rect 4432 35962 4457 35981
rect 4505 35962 4526 35981
rect 4578 35962 4595 35981
rect 4651 35962 4664 35981
rect 4724 35962 4733 35981
rect 4797 35962 4802 35981
rect 4284 35947 4319 35962
rect 4353 35947 4388 35962
rect 4422 35947 4457 35962
rect 4491 35947 4526 35962
rect 4560 35947 4595 35962
rect 4629 35947 4664 35962
rect 4698 35947 4733 35962
rect 4767 35947 4802 35962
rect 4870 35981 4909 35996
rect 4943 35981 4982 35996
rect 5016 35981 5055 35996
rect 15529 35981 15577 35996
rect 4870 35962 4871 35981
rect 4836 35947 4871 35962
rect 4905 35962 4909 35981
rect 4974 35962 4982 35981
rect 4905 35947 4940 35962
rect 4974 35947 5009 35962
rect 5043 35947 5055 35981
rect 15529 35947 15543 35981
rect 3146 35924 5055 35947
rect 3146 35890 3157 35924
rect 3191 35890 3230 35924
rect 3264 35890 3303 35924
rect 3337 35890 3376 35924
rect 3410 35890 3449 35924
rect 3483 35890 3522 35924
rect 3556 35890 3595 35924
rect 3629 35890 3668 35924
rect 3702 35890 3741 35924
rect 3775 35890 3814 35924
rect 3848 35890 3887 35924
rect 3921 35890 3960 35924
rect 3994 35890 4033 35924
rect 4067 35890 4106 35924
rect 4140 35890 4179 35924
rect 4213 35890 4252 35924
rect 4286 35890 4325 35924
rect 4359 35890 4398 35924
rect 4432 35890 4471 35924
rect 4505 35890 4544 35924
rect 4578 35890 4617 35924
rect 4651 35890 4690 35924
rect 4724 35890 4763 35924
rect 4797 35890 4836 35924
rect 4870 35890 4909 35924
rect 4943 35890 4982 35924
rect 5016 35890 5055 35924
rect 15529 35890 15577 35947
rect 3146 35887 13785 35890
rect 13925 35887 15577 35890
rect -17 35705 843 35729
rect 17 35671 55 35705
rect 89 35671 127 35705
rect 161 35671 199 35705
rect 233 35671 271 35705
rect 305 35671 343 35705
rect 377 35671 415 35705
rect 449 35671 487 35705
rect 521 35671 559 35705
rect 593 35671 631 35705
rect 665 35671 703 35705
rect 737 35671 775 35705
rect 809 35695 843 35705
rect 877 35695 915 35729
rect 949 35695 983 35729
rect 809 35671 983 35695
rect -17 35648 983 35671
rect -17 35637 463 35648
rect 929 35645 983 35648
rect 17 35603 55 35637
rect 89 35603 127 35637
rect 161 35603 199 35637
rect 233 35603 271 35637
rect 305 35603 343 35637
rect 377 35603 415 35637
rect 449 35603 463 35637
rect 949 35611 983 35645
rect -17 35569 463 35603
rect 17 35535 55 35569
rect 89 35535 127 35569
rect 161 35535 199 35569
rect 233 35535 271 35569
rect 305 35535 343 35569
rect 377 35535 415 35569
rect 449 35535 463 35569
rect 929 35561 983 35611
rect -17 35501 463 35535
rect 949 35527 983 35561
rect 17 35467 55 35501
rect 89 35467 127 35501
rect 161 35467 199 35501
rect 233 35467 271 35501
rect 305 35467 343 35501
rect 377 35467 415 35501
rect 449 35467 463 35501
rect 929 35477 983 35527
rect -17 35433 463 35467
rect 949 35443 983 35477
rect 17 35399 55 35433
rect 89 35399 127 35433
rect 161 35399 199 35433
rect 233 35399 271 35433
rect 305 35399 343 35433
rect 377 35399 415 35433
rect 449 35399 463 35433
rect -17 35365 463 35399
rect 929 35393 983 35443
rect 17 35331 55 35365
rect 89 35331 127 35365
rect 161 35331 199 35365
rect 233 35331 271 35365
rect 305 35331 343 35365
rect 377 35331 415 35365
rect 449 35331 463 35365
rect 949 35359 983 35393
rect -17 35297 463 35331
rect 929 35309 983 35359
rect 17 35263 55 35297
rect 89 35263 127 35297
rect 161 35263 199 35297
rect 233 35263 271 35297
rect 305 35263 343 35297
rect 377 35263 415 35297
rect 449 35263 463 35297
rect 949 35275 983 35309
rect -17 35229 463 35263
rect 17 35195 55 35229
rect 89 35195 127 35229
rect 161 35195 199 35229
rect 233 35195 271 35229
rect 305 35195 343 35229
rect 377 35195 415 35229
rect 449 35195 463 35229
rect 929 35225 983 35275
rect -17 35161 463 35195
rect 949 35191 983 35225
rect 17 35127 55 35161
rect 89 35127 127 35161
rect 161 35127 199 35161
rect 233 35127 271 35161
rect 305 35127 343 35161
rect 377 35127 415 35161
rect 449 35127 463 35161
rect 929 35141 983 35191
rect -17 35093 463 35127
rect 949 35107 983 35141
rect 17 35059 55 35093
rect 89 35059 127 35093
rect 161 35059 199 35093
rect 233 35059 271 35093
rect 305 35059 343 35093
rect 377 35059 415 35093
rect 449 35059 463 35093
rect -17 35025 463 35059
rect 929 35057 983 35107
rect 17 34991 55 35025
rect 89 34991 127 35025
rect 161 34991 199 35025
rect 233 34991 271 35025
rect 305 34991 343 35025
rect 377 34991 415 35025
rect 449 34991 463 35025
rect 949 35023 983 35057
rect -17 34957 463 34991
rect 929 34973 983 35023
rect 17 34923 55 34957
rect 89 34923 127 34957
rect 161 34923 199 34957
rect 233 34923 271 34957
rect 305 34923 343 34957
rect 377 34923 415 34957
rect 449 34923 463 34957
rect 949 34939 983 34973
rect -17 34889 463 34923
rect 929 34889 983 34939
rect 17 34855 55 34889
rect 89 34855 127 34889
rect 161 34855 199 34889
rect 233 34855 271 34889
rect 305 34855 343 34889
rect 377 34855 415 34889
rect 449 34855 463 34889
rect 949 34855 983 34889
rect -17 34821 463 34855
rect 17 34787 55 34821
rect 89 34787 127 34821
rect 161 34787 199 34821
rect 233 34787 271 34821
rect 305 34787 343 34821
rect 377 34787 415 34821
rect 449 34787 463 34821
rect 929 34805 983 34855
rect -17 34753 463 34787
rect 949 34771 983 34805
rect 17 34719 55 34753
rect 89 34719 127 34753
rect 161 34719 199 34753
rect 233 34719 271 34753
rect 305 34719 343 34753
rect 377 34719 415 34753
rect 449 34719 463 34753
rect 929 34721 983 34771
rect -17 34685 463 34719
rect 949 34687 983 34721
rect 17 34651 55 34685
rect 89 34651 127 34685
rect 161 34651 199 34685
rect 233 34651 271 34685
rect 305 34651 343 34685
rect 377 34651 415 34685
rect 449 34651 463 34685
rect -17 34617 463 34651
rect 929 34637 983 34687
rect 17 34583 55 34617
rect 89 34583 127 34617
rect 161 34583 199 34617
rect 233 34583 271 34617
rect 305 34583 343 34617
rect 377 34583 415 34617
rect 449 34583 463 34617
rect 949 34603 983 34637
rect -17 34549 463 34583
rect 929 34553 983 34603
rect 17 34515 55 34549
rect 89 34515 127 34549
rect 161 34515 199 34549
rect 233 34515 271 34549
rect 305 34515 343 34549
rect 377 34515 415 34549
rect 449 34515 463 34549
rect 949 34519 983 34553
rect -17 34481 463 34515
rect 17 34447 55 34481
rect 89 34447 127 34481
rect 161 34447 199 34481
rect 233 34447 271 34481
rect 305 34447 343 34481
rect 377 34447 415 34481
rect 449 34447 463 34481
rect 929 34469 983 34519
rect -17 34413 463 34447
rect 949 34435 983 34469
rect 17 34379 55 34413
rect 89 34379 127 34413
rect 161 34379 199 34413
rect 233 34379 271 34413
rect 305 34379 343 34413
rect 377 34379 415 34413
rect 449 34379 463 34413
rect 929 34385 983 34435
rect -17 34345 463 34379
rect 949 34351 983 34385
rect 17 34311 55 34345
rect 89 34311 127 34345
rect 161 34311 199 34345
rect 233 34311 271 34345
rect 305 34311 343 34345
rect 377 34311 415 34345
rect 449 34311 463 34345
rect -17 34277 463 34311
rect 929 34301 983 34351
rect 17 34243 55 34277
rect 89 34243 127 34277
rect 161 34243 199 34277
rect 233 34243 271 34277
rect 305 34243 343 34277
rect 377 34243 415 34277
rect 449 34246 463 34277
rect 949 34267 983 34301
rect 929 34246 983 34267
rect 449 34243 487 34246
rect 521 34243 559 34246
rect 593 34243 631 34246
rect 665 34243 703 34246
rect 737 34243 775 34246
rect 809 34243 983 34246
rect -17 34217 983 34243
rect -17 34209 843 34217
rect 17 34175 55 34209
rect 89 34175 127 34209
rect 161 34175 199 34209
rect 233 34175 271 34209
rect 305 34175 343 34209
rect 377 34175 415 34209
rect 449 34207 487 34209
rect 521 34207 559 34209
rect 593 34207 631 34209
rect 665 34207 703 34209
rect 737 34207 775 34209
rect 809 34207 843 34209
rect 877 34207 915 34217
rect 449 34175 463 34207
rect 521 34175 535 34207
rect 593 34175 607 34207
rect 665 34175 679 34207
rect 737 34175 751 34207
rect 809 34175 823 34207
rect 877 34183 895 34207
rect 949 34183 983 34217
rect -17 34173 463 34175
rect 497 34173 535 34175
rect 569 34173 607 34175
rect 641 34173 679 34175
rect 713 34173 751 34175
rect 785 34173 823 34175
rect 857 34173 895 34183
rect 929 34173 983 34183
rect -17 34141 983 34173
rect 17 34107 55 34141
rect 89 34107 127 34141
rect 161 34107 199 34141
rect 233 34107 271 34141
rect 305 34107 343 34141
rect 377 34107 415 34141
rect 449 34134 487 34141
rect 521 34134 559 34141
rect 593 34134 631 34141
rect 665 34134 703 34141
rect 737 34134 775 34141
rect 809 34134 983 34141
rect 449 34107 463 34134
rect 521 34107 535 34134
rect 593 34107 607 34134
rect 665 34107 679 34134
rect 737 34107 751 34134
rect 809 34107 823 34134
rect 857 34133 895 34134
rect 929 34133 983 34134
rect -17 34100 463 34107
rect 497 34100 535 34107
rect 569 34100 607 34107
rect 641 34100 679 34107
rect 713 34100 751 34107
rect 785 34100 823 34107
rect 877 34100 895 34133
rect -17 34099 843 34100
rect 877 34099 915 34100
rect 949 34099 983 34133
rect -17 34073 983 34099
rect 17 34039 55 34073
rect 89 34039 127 34073
rect 161 34039 199 34073
rect 233 34039 271 34073
rect 305 34039 343 34073
rect 377 34039 415 34073
rect 449 34061 487 34073
rect 521 34061 559 34073
rect 593 34061 631 34073
rect 665 34061 703 34073
rect 737 34061 775 34073
rect 809 34061 983 34073
rect 449 34039 463 34061
rect 521 34039 535 34061
rect 593 34039 607 34061
rect 665 34039 679 34061
rect 737 34039 751 34061
rect 809 34039 823 34061
rect 857 34049 895 34061
rect 929 34049 983 34061
rect -17 34027 463 34039
rect 497 34027 535 34039
rect 569 34027 607 34039
rect 641 34027 679 34039
rect 713 34027 751 34039
rect 785 34027 823 34039
rect 877 34027 895 34049
rect -17 34018 843 34027
rect -23 34015 843 34018
rect 877 34015 915 34027
rect 949 34015 983 34049
rect -23 34005 983 34015
rect -23 33952 -17 34005
rect 17 33971 55 34005
rect 89 33986 127 34005
rect 109 33971 127 33986
rect 161 33986 199 34005
rect 233 33986 271 34005
rect 161 33971 167 33986
rect 233 33971 259 33986
rect 305 33971 343 34005
rect 377 33971 415 34005
rect 449 33988 487 34005
rect 521 33988 559 34005
rect 593 33988 631 34005
rect 665 33988 703 34005
rect 737 33988 775 34005
rect 809 33988 983 34005
rect 449 33971 463 33988
rect 521 33971 535 33988
rect 593 33971 607 33988
rect 665 33971 679 33988
rect 737 33971 751 33988
rect 809 33971 823 33988
rect 17 33952 75 33971
rect 109 33952 167 33971
rect 201 33952 259 33971
rect 293 33954 463 33971
rect 497 33954 535 33971
rect 569 33954 607 33971
rect 641 33954 679 33971
rect 713 33954 751 33971
rect 785 33954 823 33971
rect 857 33965 895 33988
rect 929 33965 983 33988
rect 877 33954 895 33965
rect 293 33952 843 33954
rect -23 33937 843 33952
rect -23 33880 -17 33937
rect 17 33903 55 33937
rect 89 33914 127 33937
rect 109 33903 127 33914
rect 161 33914 199 33937
rect 233 33914 271 33937
rect 161 33903 167 33914
rect 233 33903 259 33914
rect 305 33903 343 33937
rect 377 33903 415 33937
rect 449 33915 487 33937
rect 521 33915 559 33937
rect 593 33915 631 33937
rect 665 33915 703 33937
rect 737 33915 775 33937
rect 809 33931 843 33937
rect 877 33931 915 33954
rect 949 33931 983 33965
rect 809 33915 983 33931
rect 449 33903 463 33915
rect 521 33903 535 33915
rect 593 33903 607 33915
rect 665 33903 679 33915
rect 737 33903 751 33915
rect 809 33903 823 33915
rect 17 33880 75 33903
rect 109 33880 167 33903
rect 201 33880 259 33903
rect 293 33881 463 33903
rect 497 33881 535 33903
rect 569 33881 607 33903
rect 641 33881 679 33903
rect 713 33881 751 33903
rect 785 33881 823 33903
rect 857 33881 895 33915
rect 929 33881 983 33915
rect 293 33880 843 33881
rect -23 33869 843 33880
rect -23 33808 -17 33869
rect 17 33835 55 33869
rect 89 33842 127 33869
rect 109 33835 127 33842
rect 161 33842 199 33869
rect 233 33842 271 33869
rect 161 33835 167 33842
rect 233 33835 259 33842
rect 305 33835 343 33869
rect 377 33835 415 33869
rect 449 33842 487 33869
rect 521 33842 559 33869
rect 593 33842 631 33869
rect 665 33842 703 33869
rect 737 33842 775 33869
rect 809 33847 843 33869
rect 877 33847 915 33881
rect 949 33847 983 33881
rect 809 33842 983 33847
rect 449 33835 463 33842
rect 521 33835 535 33842
rect 593 33835 607 33842
rect 665 33835 679 33842
rect 737 33835 751 33842
rect 809 33835 823 33842
rect 17 33808 75 33835
rect 109 33808 167 33835
rect 201 33808 259 33835
rect 293 33808 463 33835
rect 497 33808 535 33835
rect 569 33808 607 33835
rect 641 33808 679 33835
rect 713 33808 751 33835
rect 785 33808 823 33835
rect 857 33808 895 33842
rect 929 33808 983 33842
rect -23 33801 983 33808
rect -23 33735 -17 33801
rect 17 33767 55 33801
rect 89 33769 127 33801
rect 109 33767 127 33769
rect 161 33769 199 33801
rect 233 33769 271 33801
rect 161 33767 167 33769
rect 233 33767 259 33769
rect 305 33767 343 33801
rect 377 33767 415 33801
rect 449 33769 487 33801
rect 521 33769 559 33801
rect 593 33769 631 33801
rect 665 33769 703 33801
rect 737 33769 775 33801
rect 809 33797 983 33801
rect 809 33769 843 33797
rect 877 33769 915 33797
rect 449 33767 463 33769
rect 521 33767 535 33769
rect 593 33767 607 33769
rect 665 33767 679 33769
rect 737 33767 751 33769
rect 809 33767 823 33769
rect 17 33735 75 33767
rect 109 33735 167 33767
rect 201 33735 259 33767
rect 293 33735 463 33767
rect 497 33735 535 33767
rect 569 33735 607 33767
rect 641 33735 679 33767
rect 713 33735 751 33767
rect 785 33735 823 33767
rect 877 33763 895 33769
rect 949 33763 983 33797
rect 857 33735 895 33763
rect 929 33735 983 33763
rect -23 33733 983 33735
rect -23 33699 -17 33733
rect 17 33699 55 33733
rect 89 33699 127 33733
rect 161 33699 199 33733
rect 233 33699 271 33733
rect 305 33699 343 33733
rect 377 33699 415 33733
rect 449 33699 487 33733
rect 521 33699 559 33733
rect 593 33699 631 33733
rect 665 33699 703 33733
rect 737 33699 775 33733
rect 809 33713 983 33733
rect 809 33699 843 33713
rect -23 33696 843 33699
rect 877 33696 915 33713
rect -23 33631 -17 33696
rect 17 33665 75 33696
rect 109 33665 167 33696
rect 201 33665 259 33696
rect 293 33665 463 33696
rect 497 33665 535 33696
rect 569 33665 607 33696
rect 641 33665 679 33696
rect 713 33665 751 33696
rect 785 33665 823 33696
rect 877 33679 895 33696
rect 949 33679 983 33713
rect 17 33631 55 33665
rect 109 33662 127 33665
rect 89 33631 127 33662
rect 161 33662 167 33665
rect 233 33662 259 33665
rect 161 33631 199 33662
rect 233 33631 271 33662
rect 305 33631 343 33665
rect 377 33631 415 33665
rect 449 33662 463 33665
rect 521 33662 535 33665
rect 593 33662 607 33665
rect 665 33662 679 33665
rect 737 33662 751 33665
rect 809 33662 823 33665
rect 857 33662 895 33679
rect 929 33662 983 33679
rect 449 33631 487 33662
rect 521 33631 559 33662
rect 593 33631 631 33662
rect 665 33631 703 33662
rect 737 33631 775 33662
rect 809 33631 983 33662
rect -23 33629 983 33631
rect -23 33623 843 33629
rect 877 33623 915 33629
rect -23 33563 -17 33623
rect 17 33597 75 33623
rect 109 33597 167 33623
rect 201 33597 259 33623
rect 293 33597 463 33623
rect 497 33597 535 33623
rect 569 33597 607 33623
rect 641 33597 679 33623
rect 713 33597 751 33623
rect 785 33597 823 33623
rect 17 33563 55 33597
rect 109 33589 127 33597
rect 89 33563 127 33589
rect 161 33589 167 33597
rect 233 33589 259 33597
rect 161 33563 199 33589
rect 233 33563 271 33589
rect 305 33563 343 33597
rect 377 33563 415 33597
rect 449 33589 463 33597
rect 521 33589 535 33597
rect 593 33589 607 33597
rect 665 33589 679 33597
rect 737 33589 751 33597
rect 809 33589 823 33597
rect 877 33595 895 33623
rect 949 33595 983 33629
rect 857 33589 895 33595
rect 929 33589 983 33595
rect 449 33563 487 33589
rect 521 33563 559 33589
rect 593 33563 631 33589
rect 665 33563 703 33589
rect 737 33563 775 33589
rect 809 33563 983 33589
rect -23 33550 983 33563
rect -23 33495 -17 33550
rect 17 33529 75 33550
rect 109 33529 167 33550
rect 201 33529 259 33550
rect 293 33529 463 33550
rect 497 33529 535 33550
rect 569 33529 607 33550
rect 641 33529 679 33550
rect 713 33529 751 33550
rect 785 33529 823 33550
rect 857 33545 895 33550
rect 929 33545 983 33550
rect 17 33495 55 33529
rect 109 33516 127 33529
rect 89 33495 127 33516
rect 161 33516 167 33529
rect 233 33516 259 33529
rect 161 33495 199 33516
rect 233 33495 271 33516
rect 305 33495 343 33529
rect 377 33495 415 33529
rect 449 33516 463 33529
rect 521 33516 535 33529
rect 593 33516 607 33529
rect 665 33516 679 33529
rect 737 33516 751 33529
rect 809 33516 823 33529
rect 877 33516 895 33545
rect 449 33495 487 33516
rect 521 33495 559 33516
rect 593 33495 631 33516
rect 665 33495 703 33516
rect 737 33495 775 33516
rect 809 33511 843 33516
rect 877 33511 915 33516
rect 949 33511 983 33545
rect 809 33495 983 33511
rect -23 33477 983 33495
rect -23 33427 -17 33477
rect 17 33461 75 33477
rect 109 33461 167 33477
rect 201 33461 259 33477
rect 293 33461 463 33477
rect 497 33461 535 33477
rect 569 33461 607 33477
rect 641 33461 679 33477
rect 713 33461 751 33477
rect 785 33461 823 33477
rect 857 33461 895 33477
rect 929 33461 983 33477
rect 17 33427 55 33461
rect 109 33443 127 33461
rect 89 33427 127 33443
rect 161 33443 167 33461
rect 233 33443 259 33461
rect 161 33427 199 33443
rect 233 33427 271 33443
rect 305 33427 343 33461
rect 377 33427 415 33461
rect 449 33443 463 33461
rect 521 33443 535 33461
rect 593 33443 607 33461
rect 665 33443 679 33461
rect 737 33443 751 33461
rect 809 33443 823 33461
rect 877 33443 895 33461
rect 449 33427 487 33443
rect 521 33427 559 33443
rect 593 33427 631 33443
rect 665 33427 703 33443
rect 737 33427 775 33443
rect 809 33427 843 33443
rect 877 33427 915 33443
rect 949 33427 983 33461
rect -23 33404 983 33427
rect -23 33359 -17 33404
rect 17 33393 75 33404
rect 109 33393 167 33404
rect 201 33393 259 33404
rect 293 33393 463 33404
rect 497 33393 535 33404
rect 569 33393 607 33404
rect 641 33393 679 33404
rect 713 33393 751 33404
rect 785 33393 823 33404
rect 17 33359 55 33393
rect 109 33370 127 33393
rect 89 33359 127 33370
rect 161 33370 167 33393
rect 233 33370 259 33393
rect 161 33359 199 33370
rect 233 33359 271 33370
rect 305 33359 343 33393
rect 377 33359 415 33393
rect 449 33370 463 33393
rect 521 33370 535 33393
rect 593 33370 607 33393
rect 665 33370 679 33393
rect 737 33370 751 33393
rect 809 33370 823 33393
rect 857 33377 895 33404
rect 929 33377 983 33404
rect 877 33370 895 33377
rect 449 33359 487 33370
rect 521 33359 559 33370
rect 593 33359 631 33370
rect 665 33359 703 33370
rect 737 33359 775 33370
rect 809 33359 843 33370
rect -23 33343 843 33359
rect 877 33343 915 33370
rect 949 33343 983 33377
rect -23 33331 983 33343
rect -23 33291 -17 33331
rect 17 33325 75 33331
rect 109 33325 167 33331
rect 201 33325 259 33331
rect 293 33325 463 33331
rect 497 33325 535 33331
rect 569 33325 607 33331
rect 641 33325 679 33331
rect 713 33325 751 33331
rect 785 33325 823 33331
rect 17 33291 55 33325
rect 109 33297 127 33325
rect 89 33291 127 33297
rect 161 33297 167 33325
rect 233 33297 259 33325
rect 161 33291 199 33297
rect 233 33291 271 33297
rect 305 33291 343 33325
rect 377 33291 415 33325
rect 449 33297 463 33325
rect 521 33297 535 33325
rect 593 33297 607 33325
rect 665 33297 679 33325
rect 737 33297 751 33325
rect 809 33297 823 33325
rect 857 33297 895 33331
rect 929 33297 983 33331
rect 449 33291 487 33297
rect 521 33291 559 33297
rect 593 33291 631 33297
rect 665 33291 703 33297
rect 737 33291 775 33297
rect 809 33293 983 33297
rect 809 33291 843 33293
rect -23 33259 843 33291
rect 877 33259 915 33293
rect 949 33259 983 33293
rect -23 33258 983 33259
rect -23 33223 -17 33258
rect 17 33257 75 33258
rect 109 33257 167 33258
rect 201 33257 259 33258
rect 293 33257 463 33258
rect 497 33257 535 33258
rect 569 33257 607 33258
rect 641 33257 679 33258
rect 713 33257 751 33258
rect 785 33257 823 33258
rect 17 33223 55 33257
rect 109 33224 127 33257
rect 89 33223 127 33224
rect 161 33224 167 33257
rect 233 33224 259 33257
rect 161 33223 199 33224
rect 233 33223 271 33224
rect 305 33223 343 33257
rect 377 33223 415 33257
rect 449 33224 463 33257
rect 521 33224 535 33257
rect 593 33224 607 33257
rect 665 33224 679 33257
rect 737 33224 751 33257
rect 809 33224 823 33257
rect 857 33224 895 33258
rect 929 33224 983 33258
rect 449 33223 487 33224
rect 521 33223 559 33224
rect 593 33223 631 33224
rect 665 33223 703 33224
rect 737 33223 775 33224
rect 809 33223 983 33224
rect -23 33209 983 33223
rect -23 33189 843 33209
rect -23 33151 -17 33189
rect 17 33155 55 33189
rect 89 33185 127 33189
rect 109 33155 127 33185
rect 161 33185 199 33189
rect 233 33185 271 33189
rect 161 33155 167 33185
rect 233 33155 259 33185
rect 305 33155 343 33189
rect 377 33155 415 33189
rect 449 33185 487 33189
rect 521 33185 559 33189
rect 593 33185 631 33189
rect 665 33185 703 33189
rect 737 33185 775 33189
rect 809 33185 843 33189
rect 877 33185 915 33209
rect 449 33155 463 33185
rect 521 33155 535 33185
rect 593 33155 607 33185
rect 665 33155 679 33185
rect 737 33155 751 33185
rect 809 33155 823 33185
rect 877 33175 895 33185
rect 949 33175 983 33209
rect 17 33151 75 33155
rect 109 33151 167 33155
rect 201 33151 259 33155
rect 293 33151 463 33155
rect 497 33151 535 33155
rect 569 33151 607 33155
rect 641 33151 679 33155
rect 713 33151 751 33155
rect 785 33151 823 33155
rect 857 33151 895 33175
rect 929 33151 983 33175
rect -23 33125 983 33151
rect -23 33121 843 33125
rect -23 33078 -17 33121
rect 17 33087 55 33121
rect 89 33112 127 33121
rect 109 33087 127 33112
rect 161 33112 199 33121
rect 233 33112 271 33121
rect 161 33087 167 33112
rect 233 33087 259 33112
rect 305 33087 343 33121
rect 377 33087 415 33121
rect 449 33112 487 33121
rect 521 33112 559 33121
rect 593 33112 631 33121
rect 665 33112 703 33121
rect 737 33112 775 33121
rect 809 33112 843 33121
rect 877 33112 915 33125
rect 449 33087 463 33112
rect 521 33087 535 33112
rect 593 33087 607 33112
rect 665 33087 679 33112
rect 737 33087 751 33112
rect 809 33087 823 33112
rect 877 33091 895 33112
rect 949 33091 983 33125
rect 17 33078 75 33087
rect 109 33078 167 33087
rect 201 33078 259 33087
rect 293 33078 463 33087
rect 497 33078 535 33087
rect 569 33078 607 33087
rect 641 33078 679 33087
rect 713 33078 751 33087
rect 785 33078 823 33087
rect 857 33078 895 33091
rect 929 33078 983 33091
rect -23 33053 983 33078
rect -23 33005 -17 33053
rect 17 33019 55 33053
rect 89 33039 127 33053
rect 109 33019 127 33039
rect 161 33039 199 33053
rect 233 33039 271 33053
rect 161 33019 167 33039
rect 233 33019 259 33039
rect 305 33019 343 33053
rect 377 33019 415 33053
rect 449 33039 487 33053
rect 521 33039 559 33053
rect 593 33039 631 33053
rect 665 33039 703 33053
rect 737 33039 775 33053
rect 809 33041 983 33053
rect 809 33039 843 33041
rect 877 33039 915 33041
rect 449 33019 463 33039
rect 521 33019 535 33039
rect 593 33019 607 33039
rect 665 33019 679 33039
rect 737 33019 751 33039
rect 809 33019 823 33039
rect 17 33005 75 33019
rect 109 33005 167 33019
rect 201 33005 259 33019
rect 293 33005 463 33019
rect 497 33005 535 33019
rect 569 33005 607 33019
rect 641 33005 679 33019
rect 713 33005 751 33019
rect 785 33005 823 33019
rect 877 33007 895 33039
rect 949 33007 983 33041
rect 857 33005 895 33007
rect 929 33005 983 33007
rect -23 32985 983 33005
rect -23 32932 -17 32985
rect 17 32951 55 32985
rect 89 32966 127 32985
rect 109 32951 127 32966
rect 161 32966 199 32985
rect 233 32966 271 32985
rect 161 32951 167 32966
rect 233 32951 259 32966
rect 305 32951 343 32985
rect 377 32951 415 32985
rect 449 32966 487 32985
rect 521 32966 559 32985
rect 593 32966 631 32985
rect 665 32966 703 32985
rect 737 32966 775 32985
rect 809 32966 983 32985
rect 449 32951 463 32966
rect 521 32951 535 32966
rect 593 32951 607 32966
rect 665 32951 679 32966
rect 737 32951 751 32966
rect 809 32951 823 32966
rect 857 32957 895 32966
rect 929 32957 983 32966
rect 17 32932 75 32951
rect 109 32932 167 32951
rect 201 32932 259 32951
rect 293 32932 463 32951
rect 497 32932 535 32951
rect 569 32932 607 32951
rect 641 32932 679 32951
rect 713 32932 751 32951
rect 785 32932 823 32951
rect 877 32932 895 32957
rect -23 32923 843 32932
rect 877 32923 915 32932
rect 949 32923 983 32957
rect -23 32917 983 32923
rect -23 32859 -17 32917
rect 17 32883 55 32917
rect 89 32893 127 32917
rect 109 32883 127 32893
rect 161 32893 199 32917
rect 233 32893 271 32917
rect 161 32883 167 32893
rect 233 32883 259 32893
rect 305 32883 343 32917
rect 377 32883 415 32917
rect 449 32893 487 32917
rect 521 32893 559 32917
rect 593 32893 631 32917
rect 665 32893 703 32917
rect 737 32893 775 32917
rect 809 32893 983 32917
rect 449 32883 463 32893
rect 521 32883 535 32893
rect 593 32883 607 32893
rect 665 32883 679 32893
rect 737 32883 751 32893
rect 809 32883 823 32893
rect 17 32859 75 32883
rect 109 32859 167 32883
rect 201 32859 259 32883
rect 293 32859 463 32883
rect 497 32859 535 32883
rect 569 32859 607 32883
rect 641 32859 679 32883
rect 713 32859 751 32883
rect 785 32859 823 32883
rect 857 32873 895 32893
rect 929 32873 983 32893
rect 877 32859 895 32873
rect -23 32849 843 32859
rect -23 32786 -17 32849
rect 17 32815 55 32849
rect 89 32820 127 32849
rect 109 32815 127 32820
rect 161 32820 199 32849
rect 233 32820 271 32849
rect 161 32815 167 32820
rect 233 32815 259 32820
rect 305 32815 343 32849
rect 377 32815 415 32849
rect 449 32820 487 32849
rect 521 32820 559 32849
rect 593 32820 631 32849
rect 665 32820 703 32849
rect 737 32820 775 32849
rect 809 32839 843 32849
rect 877 32839 915 32859
rect 949 32839 983 32873
rect 809 32820 983 32839
rect 449 32815 463 32820
rect 521 32815 535 32820
rect 593 32815 607 32820
rect 665 32815 679 32820
rect 737 32815 751 32820
rect 809 32815 823 32820
rect 17 32786 75 32815
rect 109 32786 167 32815
rect 201 32786 259 32815
rect 293 32786 463 32815
rect 497 32786 535 32815
rect 569 32786 607 32815
rect 641 32786 679 32815
rect 713 32786 751 32815
rect 785 32786 823 32815
rect 857 32789 895 32820
rect 929 32789 983 32820
rect 877 32786 895 32789
rect -23 32781 843 32786
rect -23 32679 -17 32781
rect 17 32747 55 32781
rect 89 32747 127 32781
rect 161 32747 199 32781
rect 233 32747 271 32781
rect 305 32747 343 32781
rect 377 32747 415 32781
rect 449 32747 487 32781
rect 521 32747 559 32781
rect 593 32747 631 32781
rect 665 32747 703 32781
rect 737 32747 775 32781
rect 809 32755 843 32781
rect 877 32755 915 32786
rect 949 32755 983 32789
rect 809 32747 983 32755
rect 17 32713 75 32747
rect 109 32713 167 32747
rect 201 32713 259 32747
rect 293 32713 463 32747
rect 497 32713 535 32747
rect 569 32713 607 32747
rect 641 32713 679 32747
rect 713 32713 751 32747
rect 785 32713 823 32747
rect 857 32713 895 32747
rect 929 32713 983 32747
rect 17 32679 55 32713
rect 89 32679 127 32713
rect 161 32679 199 32713
rect 233 32679 271 32713
rect 305 32679 343 32713
rect 377 32679 415 32713
rect 449 32679 487 32713
rect 521 32679 559 32713
rect 593 32679 631 32713
rect 665 32679 703 32713
rect 737 32679 775 32713
rect 809 32705 983 32713
rect 809 32679 843 32705
rect -23 32674 843 32679
rect 877 32674 915 32705
rect -23 32611 -17 32674
rect 17 32645 75 32674
rect 109 32645 167 32674
rect 201 32645 259 32674
rect 293 32645 463 32674
rect 497 32645 535 32674
rect 569 32645 607 32674
rect 641 32645 679 32674
rect 713 32645 751 32674
rect 785 32645 823 32674
rect 877 32671 895 32674
rect 949 32671 983 32705
rect 17 32611 55 32645
rect 109 32640 127 32645
rect 89 32611 127 32640
rect 161 32640 167 32645
rect 233 32640 259 32645
rect 161 32611 199 32640
rect 233 32611 271 32640
rect 305 32611 343 32645
rect 377 32611 415 32645
rect 449 32640 463 32645
rect 521 32640 535 32645
rect 593 32640 607 32645
rect 665 32640 679 32645
rect 737 32640 751 32645
rect 809 32640 823 32645
rect 857 32640 895 32671
rect 929 32640 983 32671
rect 449 32611 487 32640
rect 521 32611 559 32640
rect 593 32611 631 32640
rect 665 32611 703 32640
rect 737 32611 775 32640
rect 809 32621 983 32640
rect 809 32611 843 32621
rect -23 32601 843 32611
rect 877 32601 915 32621
rect -23 32543 -17 32601
rect 17 32577 75 32601
rect 109 32577 167 32601
rect 201 32577 259 32601
rect 293 32577 463 32601
rect 497 32577 535 32601
rect 569 32577 607 32601
rect 641 32577 679 32601
rect 713 32577 751 32601
rect 785 32577 823 32601
rect 877 32587 895 32601
rect 949 32587 983 32621
rect 17 32543 55 32577
rect 109 32567 127 32577
rect 89 32543 127 32567
rect 161 32567 167 32577
rect 233 32567 259 32577
rect 161 32543 199 32567
rect 233 32543 271 32567
rect 305 32543 343 32577
rect 377 32543 415 32577
rect 449 32567 463 32577
rect 521 32567 535 32577
rect 593 32567 607 32577
rect 665 32567 679 32577
rect 737 32567 751 32577
rect 809 32567 823 32577
rect 857 32567 895 32587
rect 929 32567 983 32587
rect 449 32543 487 32567
rect 521 32543 559 32567
rect 593 32543 631 32567
rect 665 32543 703 32567
rect 737 32543 775 32567
rect 809 32543 983 32567
rect -23 32537 983 32543
rect -23 32528 843 32537
rect 877 32528 915 32537
rect -23 32475 -17 32528
rect 17 32509 75 32528
rect 109 32509 167 32528
rect 201 32509 259 32528
rect 293 32509 463 32528
rect 497 32509 535 32528
rect 569 32509 607 32528
rect 641 32509 679 32528
rect 713 32509 751 32528
rect 785 32509 823 32528
rect 17 32475 55 32509
rect 109 32494 127 32509
rect 89 32475 127 32494
rect 161 32494 167 32509
rect 233 32494 259 32509
rect 161 32475 199 32494
rect 233 32475 271 32494
rect 305 32475 343 32509
rect 377 32475 415 32509
rect 449 32494 463 32509
rect 521 32494 535 32509
rect 593 32494 607 32509
rect 665 32494 679 32509
rect 737 32494 751 32509
rect 809 32494 823 32509
rect 877 32503 895 32528
rect 949 32503 983 32537
rect 857 32494 895 32503
rect 929 32494 983 32503
rect 449 32475 487 32494
rect 521 32475 559 32494
rect 593 32475 631 32494
rect 665 32475 703 32494
rect 737 32475 775 32494
rect 809 32475 983 32494
rect -23 32455 983 32475
rect -23 32407 -17 32455
rect 17 32441 75 32455
rect 109 32441 167 32455
rect 201 32441 259 32455
rect 293 32441 463 32455
rect 497 32441 535 32455
rect 569 32441 607 32455
rect 641 32441 679 32455
rect 713 32441 751 32455
rect 785 32441 823 32455
rect 857 32453 895 32455
rect 929 32453 983 32455
rect 17 32407 55 32441
rect 109 32421 127 32441
rect 89 32407 127 32421
rect 161 32421 167 32441
rect 233 32421 259 32441
rect 161 32407 199 32421
rect 233 32407 271 32421
rect 305 32407 343 32441
rect 377 32407 415 32441
rect 449 32421 463 32441
rect 521 32421 535 32441
rect 593 32421 607 32441
rect 665 32421 679 32441
rect 737 32421 751 32441
rect 809 32421 823 32441
rect 877 32421 895 32453
rect 449 32407 487 32421
rect 521 32407 559 32421
rect 593 32407 631 32421
rect 665 32407 703 32421
rect 737 32407 775 32421
rect 809 32419 843 32421
rect 877 32419 915 32421
rect 949 32419 983 32453
rect 809 32407 983 32419
rect -23 32382 983 32407
rect -23 32339 -17 32382
rect 17 32373 75 32382
rect 109 32373 167 32382
rect 201 32373 259 32382
rect 293 32373 463 32382
rect 497 32373 535 32382
rect 569 32373 607 32382
rect 641 32373 679 32382
rect 713 32373 751 32382
rect 785 32373 823 32382
rect 17 32339 55 32373
rect 109 32348 127 32373
rect 89 32339 127 32348
rect 161 32348 167 32373
rect 233 32348 259 32373
rect 161 32339 199 32348
rect 233 32339 271 32348
rect 305 32339 343 32373
rect 377 32339 415 32373
rect 449 32348 463 32373
rect 521 32348 535 32373
rect 593 32348 607 32373
rect 665 32348 679 32373
rect 737 32348 751 32373
rect 809 32348 823 32373
rect 857 32369 895 32382
rect 929 32369 983 32382
rect 877 32348 895 32369
rect 449 32339 487 32348
rect 521 32339 559 32348
rect 593 32339 631 32348
rect 665 32339 703 32348
rect 737 32339 775 32348
rect 809 32339 843 32348
rect -23 32335 843 32339
rect 877 32335 915 32348
rect 949 32335 983 32369
rect -23 32309 983 32335
rect -23 32271 -17 32309
rect 17 32305 75 32309
rect 109 32305 167 32309
rect 201 32305 259 32309
rect 293 32305 463 32309
rect 497 32305 535 32309
rect 569 32305 607 32309
rect 641 32305 679 32309
rect 713 32305 751 32309
rect 785 32305 823 32309
rect 17 32271 55 32305
rect 109 32275 127 32305
rect 89 32271 127 32275
rect 161 32275 167 32305
rect 233 32275 259 32305
rect 161 32271 199 32275
rect 233 32271 271 32275
rect 305 32271 343 32305
rect 377 32271 415 32305
rect 449 32275 463 32305
rect 521 32275 535 32305
rect 593 32275 607 32305
rect 665 32275 679 32305
rect 737 32275 751 32305
rect 809 32275 823 32305
rect 857 32285 895 32309
rect 929 32285 983 32309
rect 877 32275 895 32285
rect 449 32271 487 32275
rect 521 32271 559 32275
rect 593 32271 631 32275
rect 665 32271 703 32275
rect 737 32271 775 32275
rect 809 32271 843 32275
rect -23 32251 843 32271
rect 877 32251 915 32275
rect 949 32251 983 32285
rect -23 32237 983 32251
rect -23 32202 -17 32237
rect 17 32203 55 32237
rect 89 32236 127 32237
rect 109 32203 127 32236
rect 161 32236 199 32237
rect 233 32236 271 32237
rect 161 32203 167 32236
rect 233 32203 259 32236
rect 305 32203 343 32237
rect 377 32203 415 32237
rect 449 32236 487 32237
rect 521 32236 559 32237
rect 593 32236 631 32237
rect 665 32236 703 32237
rect 737 32236 775 32237
rect 809 32236 983 32237
rect 449 32203 463 32236
rect 521 32203 535 32236
rect 593 32203 607 32236
rect 665 32203 679 32236
rect 737 32203 751 32236
rect 809 32203 823 32236
rect 17 32202 75 32203
rect 109 32202 167 32203
rect 201 32202 259 32203
rect 293 32202 463 32203
rect 497 32202 535 32203
rect 569 32202 607 32203
rect 641 32202 679 32203
rect 713 32202 751 32203
rect 785 32202 823 32203
rect 857 32202 895 32236
rect 929 32202 983 32236
rect -23 32201 983 32202
rect -23 32169 843 32201
rect -23 32129 -17 32169
rect 17 32135 55 32169
rect 89 32163 127 32169
rect 109 32135 127 32163
rect 161 32163 199 32169
rect 233 32163 271 32169
rect 161 32135 167 32163
rect 233 32135 259 32163
rect 305 32135 343 32169
rect 377 32135 415 32169
rect 449 32163 487 32169
rect 521 32163 559 32169
rect 593 32163 631 32169
rect 665 32163 703 32169
rect 737 32163 775 32169
rect 809 32167 843 32169
rect 877 32167 915 32201
rect 949 32167 983 32201
rect 809 32163 983 32167
rect 449 32135 463 32163
rect 521 32135 535 32163
rect 593 32135 607 32163
rect 665 32135 679 32163
rect 737 32135 751 32163
rect 809 32135 823 32163
rect 17 32129 75 32135
rect 109 32129 167 32135
rect 201 32129 259 32135
rect 293 32129 463 32135
rect 497 32129 535 32135
rect 569 32129 607 32135
rect 641 32129 679 32135
rect 713 32129 751 32135
rect 785 32129 823 32135
rect 857 32129 895 32163
rect 929 32129 983 32163
rect -23 32117 983 32129
rect -23 32101 843 32117
rect -23 32056 -17 32101
rect 17 32067 55 32101
rect 89 32090 127 32101
rect 109 32067 127 32090
rect 161 32090 199 32101
rect 233 32090 271 32101
rect 161 32067 167 32090
rect 233 32067 259 32090
rect 305 32067 343 32101
rect 377 32067 415 32101
rect 449 32090 487 32101
rect 521 32090 559 32101
rect 593 32090 631 32101
rect 665 32090 703 32101
rect 737 32090 775 32101
rect 809 32090 843 32101
rect 877 32090 915 32117
rect 449 32067 463 32090
rect 521 32067 535 32090
rect 593 32067 607 32090
rect 665 32067 679 32090
rect 737 32067 751 32090
rect 809 32067 823 32090
rect 877 32083 895 32090
rect 949 32083 983 32117
rect 17 32056 75 32067
rect 109 32056 167 32067
rect 201 32056 259 32067
rect 293 32056 463 32067
rect 497 32056 535 32067
rect 569 32056 607 32067
rect 641 32056 679 32067
rect 713 32056 751 32067
rect 785 32056 823 32067
rect 857 32056 895 32083
rect 929 32056 983 32083
rect -23 32033 983 32056
rect -23 31983 -17 32033
rect 17 31999 55 32033
rect 89 32017 127 32033
rect 109 31999 127 32017
rect 161 32017 199 32033
rect 233 32017 271 32033
rect 161 31999 167 32017
rect 233 31999 259 32017
rect 305 31999 343 32033
rect 377 31999 415 32033
rect 449 32017 487 32033
rect 521 32017 559 32033
rect 593 32017 631 32033
rect 665 32017 703 32033
rect 737 32017 775 32033
rect 809 32017 843 32033
rect 877 32017 915 32033
rect 449 31999 463 32017
rect 521 31999 535 32017
rect 593 31999 607 32017
rect 665 31999 679 32017
rect 737 31999 751 32017
rect 809 31999 823 32017
rect 877 31999 895 32017
rect 949 31999 983 32033
rect 17 31983 75 31999
rect 109 31983 167 31999
rect 201 31983 259 31999
rect 293 31983 463 31999
rect 497 31983 535 31999
rect 569 31983 607 31999
rect 641 31983 679 31999
rect 713 31983 751 31999
rect 785 31983 823 31999
rect 857 31983 895 31999
rect 929 31983 983 31999
rect -23 31965 983 31983
rect -23 31910 -17 31965
rect 17 31931 55 31965
rect 89 31944 127 31965
rect 109 31931 127 31944
rect 161 31944 199 31965
rect 233 31944 271 31965
rect 161 31931 167 31944
rect 233 31931 259 31944
rect 305 31931 343 31965
rect 377 31931 415 31965
rect 449 31944 487 31965
rect 521 31944 559 31965
rect 593 31944 631 31965
rect 665 31944 703 31965
rect 737 31944 775 31965
rect 809 31949 983 31965
rect 809 31944 843 31949
rect 877 31944 915 31949
rect 449 31931 463 31944
rect 521 31931 535 31944
rect 593 31931 607 31944
rect 665 31931 679 31944
rect 737 31931 751 31944
rect 809 31931 823 31944
rect 17 31910 75 31931
rect 109 31910 167 31931
rect 201 31910 259 31931
rect 293 31910 463 31931
rect 497 31910 535 31931
rect 569 31910 607 31931
rect 641 31910 679 31931
rect 713 31910 751 31931
rect 785 31910 823 31931
rect 877 31915 895 31944
rect 949 31915 983 31949
rect 857 31910 895 31915
rect 929 31910 983 31915
rect -23 31897 983 31910
rect -23 31837 -17 31897
rect 17 31863 55 31897
rect 89 31871 127 31897
rect 109 31863 127 31871
rect 161 31871 199 31897
rect 233 31871 271 31897
rect 161 31863 167 31871
rect 233 31863 259 31871
rect 305 31863 343 31897
rect 377 31863 415 31897
rect 449 31871 487 31897
rect 521 31871 559 31897
rect 593 31871 631 31897
rect 665 31871 703 31897
rect 737 31871 775 31897
rect 809 31871 983 31897
rect 449 31863 463 31871
rect 521 31863 535 31871
rect 593 31863 607 31871
rect 665 31863 679 31871
rect 737 31863 751 31871
rect 809 31863 823 31871
rect 857 31865 895 31871
rect 929 31865 983 31871
rect 17 31837 75 31863
rect 109 31837 167 31863
rect 201 31837 259 31863
rect 293 31837 463 31863
rect 497 31837 535 31863
rect 569 31837 607 31863
rect 641 31837 679 31863
rect 713 31837 751 31863
rect 785 31837 823 31863
rect 877 31837 895 31865
rect -23 31831 843 31837
rect 877 31831 915 31837
rect 949 31831 983 31865
rect -23 31829 983 31831
rect -23 31764 -17 31829
rect 17 31795 55 31829
rect 89 31798 127 31829
rect 109 31795 127 31798
rect 161 31798 199 31829
rect 233 31798 271 31829
rect 161 31795 167 31798
rect 233 31795 259 31798
rect 305 31795 343 31829
rect 377 31795 415 31829
rect 449 31798 487 31829
rect 521 31798 559 31829
rect 593 31798 631 31829
rect 665 31798 703 31829
rect 737 31798 775 31829
rect 809 31798 983 31829
rect 449 31795 463 31798
rect 521 31795 535 31798
rect 593 31795 607 31798
rect 665 31795 679 31798
rect 737 31795 751 31798
rect 809 31795 823 31798
rect 17 31764 75 31795
rect 109 31764 167 31795
rect 201 31764 259 31795
rect 293 31764 463 31795
rect 497 31764 535 31795
rect 569 31764 607 31795
rect 641 31764 679 31795
rect 713 31764 751 31795
rect 785 31764 823 31795
rect 857 31781 895 31798
rect 929 31781 983 31798
rect 877 31764 895 31781
rect -23 31761 843 31764
rect -23 31727 -17 31761
rect 17 31727 55 31761
rect 89 31727 127 31761
rect 161 31727 199 31761
rect 233 31727 271 31761
rect 305 31727 343 31761
rect 377 31727 415 31761
rect 449 31727 487 31761
rect 521 31727 559 31761
rect 593 31727 631 31761
rect 665 31727 703 31761
rect 737 31727 775 31761
rect 809 31747 843 31761
rect 877 31747 915 31764
rect 949 31747 983 31781
rect 809 31727 983 31747
rect -23 31725 983 31727
rect -23 31659 -17 31725
rect 17 31693 75 31725
rect 109 31693 167 31725
rect 201 31693 259 31725
rect 293 31693 463 31725
rect 497 31693 535 31725
rect 569 31693 607 31725
rect 641 31693 679 31725
rect 713 31693 751 31725
rect 785 31693 823 31725
rect 857 31697 895 31725
rect 929 31697 983 31725
rect 17 31659 55 31693
rect 109 31691 127 31693
rect 89 31659 127 31691
rect 161 31691 167 31693
rect 233 31691 259 31693
rect 161 31659 199 31691
rect 233 31659 271 31691
rect 305 31659 343 31693
rect 377 31659 415 31693
rect 449 31691 463 31693
rect 521 31691 535 31693
rect 593 31691 607 31693
rect 665 31691 679 31693
rect 737 31691 751 31693
rect 809 31691 823 31693
rect 877 31691 895 31697
rect 449 31659 487 31691
rect 521 31659 559 31691
rect 593 31659 631 31691
rect 665 31659 703 31691
rect 737 31659 775 31691
rect 809 31663 843 31691
rect 877 31663 915 31691
rect 949 31663 983 31697
rect 809 31659 983 31663
rect -23 31652 983 31659
rect -23 31591 -17 31652
rect 17 31625 75 31652
rect 109 31625 167 31652
rect 201 31625 259 31652
rect 293 31625 463 31652
rect 497 31625 535 31652
rect 569 31625 607 31652
rect 641 31625 679 31652
rect 713 31625 751 31652
rect 785 31625 823 31652
rect 17 31591 55 31625
rect 109 31618 127 31625
rect 89 31591 127 31618
rect 161 31618 167 31625
rect 233 31618 259 31625
rect 161 31591 199 31618
rect 233 31591 271 31618
rect 305 31591 343 31625
rect 377 31591 415 31625
rect 449 31618 463 31625
rect 521 31618 535 31625
rect 593 31618 607 31625
rect 665 31618 679 31625
rect 737 31618 751 31625
rect 809 31618 823 31625
rect 857 31618 895 31652
rect 929 31618 983 31652
rect 449 31591 487 31618
rect 521 31591 559 31618
rect 593 31591 631 31618
rect 665 31591 703 31618
rect 737 31591 775 31618
rect 809 31613 983 31618
rect 809 31591 843 31613
rect -23 31579 843 31591
rect 877 31579 915 31613
rect 949 31579 983 31613
rect -23 31523 -17 31579
rect 17 31557 75 31579
rect 109 31557 167 31579
rect 201 31557 259 31579
rect 293 31557 463 31579
rect 497 31557 535 31579
rect 569 31557 607 31579
rect 641 31557 679 31579
rect 713 31557 751 31579
rect 785 31557 823 31579
rect 17 31523 55 31557
rect 109 31545 127 31557
rect 89 31523 127 31545
rect 161 31545 167 31557
rect 233 31545 259 31557
rect 161 31523 199 31545
rect 233 31523 271 31545
rect 305 31523 343 31557
rect 377 31523 415 31557
rect 449 31545 463 31557
rect 521 31545 535 31557
rect 593 31545 607 31557
rect 665 31545 679 31557
rect 737 31545 751 31557
rect 809 31545 823 31557
rect 857 31545 895 31579
rect 929 31545 983 31579
rect 449 31523 487 31545
rect 521 31523 559 31545
rect 593 31523 631 31545
rect 665 31523 703 31545
rect 737 31523 775 31545
rect 809 31529 983 31545
rect 809 31523 843 31529
rect -23 31506 843 31523
rect 877 31506 915 31529
rect -23 31455 -17 31506
rect 17 31489 75 31506
rect 109 31489 167 31506
rect 201 31489 259 31506
rect 293 31489 463 31506
rect 497 31489 535 31506
rect 569 31489 607 31506
rect 641 31489 679 31506
rect 713 31489 751 31506
rect 785 31489 823 31506
rect 877 31495 895 31506
rect 949 31495 983 31529
rect 17 31455 55 31489
rect 109 31472 127 31489
rect 89 31455 127 31472
rect 161 31472 167 31489
rect 233 31472 259 31489
rect 161 31455 199 31472
rect 233 31455 271 31472
rect 305 31455 343 31489
rect 377 31455 415 31489
rect 449 31472 463 31489
rect 521 31472 535 31489
rect 593 31472 607 31489
rect 665 31472 679 31489
rect 737 31472 751 31489
rect 809 31472 823 31489
rect 857 31472 895 31495
rect 929 31472 983 31495
rect 449 31455 487 31472
rect 521 31455 559 31472
rect 593 31455 631 31472
rect 665 31455 703 31472
rect 737 31455 775 31472
rect 809 31455 983 31472
rect -23 31445 983 31455
rect -23 31433 843 31445
rect 877 31433 915 31445
rect -23 31387 -17 31433
rect 17 31421 75 31433
rect 109 31421 167 31433
rect 201 31421 259 31433
rect 293 31421 463 31433
rect 497 31421 535 31433
rect 569 31421 607 31433
rect 641 31421 679 31433
rect 713 31421 751 31433
rect 785 31421 823 31433
rect 17 31387 55 31421
rect 109 31399 127 31421
rect 89 31387 127 31399
rect 161 31399 167 31421
rect 233 31399 259 31421
rect 161 31387 199 31399
rect 233 31387 271 31399
rect 305 31387 343 31421
rect 377 31387 415 31421
rect 449 31399 463 31421
rect 521 31399 535 31421
rect 593 31399 607 31421
rect 665 31399 679 31421
rect 737 31399 751 31421
rect 809 31399 823 31421
rect 877 31411 895 31433
rect 949 31411 983 31445
rect 857 31399 895 31411
rect 929 31399 983 31411
rect 449 31387 487 31399
rect 521 31387 559 31399
rect 593 31387 631 31399
rect 665 31387 703 31399
rect 737 31387 775 31399
rect 809 31387 983 31399
rect -23 31361 983 31387
rect -23 31360 843 31361
rect 877 31360 915 31361
rect -23 31319 -17 31360
rect 17 31353 75 31360
rect 109 31353 167 31360
rect 201 31353 259 31360
rect 293 31353 463 31360
rect 497 31353 535 31360
rect 569 31353 607 31360
rect 641 31353 679 31360
rect 713 31353 751 31360
rect 785 31353 823 31360
rect 17 31319 55 31353
rect 109 31326 127 31353
rect 89 31319 127 31326
rect 161 31326 167 31353
rect 233 31326 259 31353
rect 161 31319 199 31326
rect 233 31319 271 31326
rect 305 31319 343 31353
rect 377 31319 415 31353
rect 449 31326 463 31353
rect 521 31326 535 31353
rect 593 31326 607 31353
rect 665 31326 679 31353
rect 737 31326 751 31353
rect 809 31326 823 31353
rect 877 31327 895 31360
rect 949 31327 983 31361
rect 857 31326 895 31327
rect 929 31326 983 31327
rect 449 31319 487 31326
rect 521 31319 559 31326
rect 593 31319 631 31326
rect 665 31319 703 31326
rect 737 31319 775 31326
rect 809 31319 983 31326
rect -23 31287 983 31319
rect -23 31251 -17 31287
rect 17 31285 75 31287
rect 109 31285 167 31287
rect 201 31285 259 31287
rect 293 31285 463 31287
rect 497 31285 535 31287
rect 569 31285 607 31287
rect 641 31285 679 31287
rect 713 31285 751 31287
rect 785 31285 823 31287
rect 17 31251 55 31285
rect 109 31253 127 31285
rect 89 31251 127 31253
rect 161 31253 167 31285
rect 233 31253 259 31285
rect 161 31251 199 31253
rect 233 31251 271 31253
rect 305 31251 343 31285
rect 377 31251 415 31285
rect 449 31253 463 31285
rect 521 31253 535 31285
rect 593 31253 607 31285
rect 665 31253 679 31285
rect 737 31253 751 31285
rect 809 31253 823 31285
rect 857 31277 895 31287
rect 929 31277 983 31287
rect 877 31253 895 31277
rect 449 31251 487 31253
rect 521 31251 559 31253
rect 593 31251 631 31253
rect 665 31251 703 31253
rect 737 31251 775 31253
rect 809 31251 843 31253
rect -23 31243 843 31251
rect 877 31243 915 31253
rect 949 31243 983 31277
rect -23 31217 983 31243
rect -23 31180 -17 31217
rect 17 31183 55 31217
rect 89 31214 127 31217
rect 109 31183 127 31214
rect 161 31214 199 31217
rect 233 31214 271 31217
rect 161 31183 167 31214
rect 233 31183 259 31214
rect 305 31183 343 31217
rect 377 31183 415 31217
rect 449 31214 487 31217
rect 521 31214 559 31217
rect 593 31214 631 31217
rect 665 31214 703 31217
rect 737 31214 775 31217
rect 809 31214 983 31217
rect 449 31183 463 31214
rect 521 31183 535 31214
rect 593 31183 607 31214
rect 665 31183 679 31214
rect 737 31183 751 31214
rect 809 31183 823 31214
rect 857 31193 895 31214
rect 929 31193 983 31214
rect 17 31180 75 31183
rect 109 31180 167 31183
rect 201 31180 259 31183
rect 293 31180 463 31183
rect 497 31180 535 31183
rect 569 31180 607 31183
rect 641 31180 679 31183
rect 713 31180 751 31183
rect 785 31180 823 31183
rect 877 31180 895 31193
rect -23 31159 843 31180
rect 877 31159 915 31180
rect 949 31159 983 31193
rect -23 31149 983 31159
rect -23 31107 -17 31149
rect 17 31115 55 31149
rect 89 31141 127 31149
rect 109 31115 127 31141
rect 161 31141 199 31149
rect 233 31141 271 31149
rect 161 31115 167 31141
rect 233 31115 259 31141
rect 305 31115 343 31149
rect 377 31115 415 31149
rect 449 31141 487 31149
rect 521 31141 559 31149
rect 593 31141 631 31149
rect 665 31141 703 31149
rect 737 31141 775 31149
rect 809 31141 983 31149
rect 449 31115 463 31141
rect 521 31115 535 31141
rect 593 31115 607 31141
rect 665 31115 679 31141
rect 737 31115 751 31141
rect 809 31115 823 31141
rect 17 31107 75 31115
rect 109 31107 167 31115
rect 201 31107 259 31115
rect 293 31107 463 31115
rect 497 31107 535 31115
rect 569 31107 607 31115
rect 641 31107 679 31115
rect 713 31107 751 31115
rect 785 31107 823 31115
rect 857 31109 895 31141
rect 929 31109 983 31141
rect 877 31107 895 31109
rect -23 31081 843 31107
rect -23 31034 -17 31081
rect 17 31047 55 31081
rect 89 31068 127 31081
rect 109 31047 127 31068
rect 161 31068 199 31081
rect 233 31068 271 31081
rect 161 31047 167 31068
rect 233 31047 259 31068
rect 305 31047 343 31081
rect 377 31047 415 31081
rect 449 31068 487 31081
rect 521 31068 559 31081
rect 593 31068 631 31081
rect 665 31068 703 31081
rect 737 31068 775 31081
rect 809 31075 843 31081
rect 877 31075 915 31107
rect 949 31075 983 31109
rect 809 31068 983 31075
rect 449 31047 463 31068
rect 521 31047 535 31068
rect 593 31047 607 31068
rect 665 31047 679 31068
rect 737 31047 751 31068
rect 809 31047 823 31068
rect 17 31034 75 31047
rect 109 31034 167 31047
rect 201 31034 259 31047
rect 293 31034 463 31047
rect 497 31034 535 31047
rect 569 31034 607 31047
rect 641 31034 679 31047
rect 713 31034 751 31047
rect 785 31034 823 31047
rect 857 31034 895 31068
rect 929 31034 983 31068
rect -23 31025 983 31034
rect -23 31013 843 31025
rect -23 30961 -17 31013
rect 17 30979 55 31013
rect 89 30995 127 31013
rect 109 30979 127 30995
rect 161 30995 199 31013
rect 233 30995 271 31013
rect 161 30979 167 30995
rect 233 30979 259 30995
rect 305 30979 343 31013
rect 377 30979 415 31013
rect 449 30995 487 31013
rect 521 30995 559 31013
rect 593 30995 631 31013
rect 665 30995 703 31013
rect 737 30995 775 31013
rect 809 30995 843 31013
rect 877 30995 915 31025
rect 449 30979 463 30995
rect 521 30979 535 30995
rect 593 30979 607 30995
rect 665 30979 679 30995
rect 737 30979 751 30995
rect 809 30979 823 30995
rect 877 30991 895 30995
rect 949 30991 983 31025
rect 17 30961 75 30979
rect 109 30961 167 30979
rect 201 30961 259 30979
rect 293 30961 463 30979
rect 497 30961 535 30979
rect 569 30961 607 30979
rect 641 30961 679 30979
rect 713 30961 751 30979
rect 785 30961 823 30979
rect 857 30961 895 30991
rect 929 30961 983 30991
rect -23 30945 983 30961
rect -23 30888 -17 30945
rect 17 30911 55 30945
rect 89 30922 127 30945
rect 109 30911 127 30922
rect 161 30922 199 30945
rect 233 30922 271 30945
rect 161 30911 167 30922
rect 233 30911 259 30922
rect 305 30911 343 30945
rect 377 30911 415 30945
rect 449 30922 487 30945
rect 521 30922 559 30945
rect 593 30922 631 30945
rect 665 30922 703 30945
rect 737 30922 775 30945
rect 809 30941 983 30945
rect 809 30922 843 30941
rect 877 30922 915 30941
rect 449 30911 463 30922
rect 521 30911 535 30922
rect 593 30911 607 30922
rect 665 30911 679 30922
rect 737 30911 751 30922
rect 809 30911 823 30922
rect 17 30888 75 30911
rect 109 30888 167 30911
rect 201 30888 259 30911
rect 293 30888 463 30911
rect 497 30888 535 30911
rect 569 30888 607 30911
rect 641 30888 679 30911
rect 713 30888 751 30911
rect 785 30888 823 30911
rect 877 30907 895 30922
rect 949 30907 983 30941
rect 857 30888 895 30907
rect 929 30888 983 30907
rect -23 30877 983 30888
rect -23 30815 -17 30877
rect 17 30843 55 30877
rect 89 30849 127 30877
rect 109 30843 127 30849
rect 161 30849 199 30877
rect 233 30849 271 30877
rect 161 30843 167 30849
rect 233 30843 259 30849
rect 305 30843 343 30877
rect 377 30843 415 30877
rect 449 30849 487 30877
rect 521 30849 559 30877
rect 593 30849 631 30877
rect 665 30849 703 30877
rect 737 30849 775 30877
rect 809 30857 983 30877
rect 809 30849 843 30857
rect 877 30849 915 30857
rect 449 30843 463 30849
rect 521 30843 535 30849
rect 593 30843 607 30849
rect 665 30843 679 30849
rect 737 30843 751 30849
rect 809 30843 823 30849
rect 17 30815 75 30843
rect 109 30815 167 30843
rect 201 30815 259 30843
rect 293 30815 463 30843
rect 497 30815 535 30843
rect 569 30815 607 30843
rect 641 30815 679 30843
rect 713 30815 751 30843
rect 785 30815 823 30843
rect 877 30823 895 30849
rect 949 30823 983 30857
rect 857 30815 895 30823
rect 929 30815 983 30823
rect -23 30809 983 30815
rect -23 30742 -17 30809
rect 17 30775 55 30809
rect 89 30776 127 30809
rect 109 30775 127 30776
rect 161 30776 199 30809
rect 233 30776 271 30809
rect 161 30775 167 30776
rect 233 30775 259 30776
rect 305 30775 343 30809
rect 377 30775 415 30809
rect 449 30776 487 30809
rect 521 30776 559 30809
rect 593 30776 631 30809
rect 665 30776 703 30809
rect 737 30776 775 30809
rect 809 30776 983 30809
rect 449 30775 463 30776
rect 521 30775 535 30776
rect 593 30775 607 30776
rect 665 30775 679 30776
rect 737 30775 751 30776
rect 809 30775 823 30776
rect 17 30742 75 30775
rect 109 30742 167 30775
rect 201 30742 259 30775
rect 293 30742 463 30775
rect 497 30742 535 30775
rect 569 30742 607 30775
rect 641 30742 679 30775
rect 713 30742 751 30775
rect 785 30742 823 30775
rect 857 30773 895 30776
rect 929 30773 983 30776
rect 877 30742 895 30773
rect -23 30741 843 30742
rect -23 30707 -17 30741
rect 17 30707 55 30741
rect 89 30707 127 30741
rect 161 30707 199 30741
rect 233 30707 271 30741
rect 305 30707 343 30741
rect 377 30707 415 30741
rect 449 30707 487 30741
rect 521 30707 559 30741
rect 593 30707 631 30741
rect 665 30707 703 30741
rect 737 30707 775 30741
rect 809 30739 843 30741
rect 877 30739 915 30742
rect 949 30739 983 30773
rect 809 30707 983 30739
rect -23 30703 983 30707
rect -23 30639 -17 30703
rect 17 30673 75 30703
rect 109 30673 167 30703
rect 201 30673 259 30703
rect 293 30673 463 30703
rect 497 30673 535 30703
rect 569 30673 607 30703
rect 641 30673 679 30703
rect 713 30673 751 30703
rect 785 30673 823 30703
rect 857 30689 895 30703
rect 929 30689 983 30703
rect 17 30639 55 30673
rect 109 30669 127 30673
rect 89 30639 127 30669
rect 161 30669 167 30673
rect 233 30669 259 30673
rect 161 30639 199 30669
rect 233 30639 271 30669
rect 305 30639 343 30673
rect 377 30639 415 30673
rect 449 30669 463 30673
rect 521 30669 535 30673
rect 593 30669 607 30673
rect 665 30669 679 30673
rect 737 30669 751 30673
rect 809 30669 823 30673
rect 877 30669 895 30689
rect 449 30639 487 30669
rect 521 30639 559 30669
rect 593 30639 631 30669
rect 665 30639 703 30669
rect 737 30639 775 30669
rect 809 30655 843 30669
rect 877 30655 915 30669
rect 949 30655 983 30689
rect 809 30639 983 30655
rect -23 30630 983 30639
rect -23 30571 -17 30630
rect 17 30605 75 30630
rect 109 30605 167 30630
rect 201 30605 259 30630
rect 293 30605 463 30630
rect 497 30605 535 30630
rect 569 30605 607 30630
rect 641 30605 679 30630
rect 713 30605 751 30630
rect 785 30605 823 30630
rect 857 30605 895 30630
rect 929 30605 983 30630
rect 17 30571 55 30605
rect 109 30596 127 30605
rect 89 30571 127 30596
rect 161 30596 167 30605
rect 233 30596 259 30605
rect 161 30571 199 30596
rect 233 30571 271 30596
rect 305 30571 343 30605
rect 377 30571 415 30605
rect 449 30596 463 30605
rect 521 30596 535 30605
rect 593 30596 607 30605
rect 665 30596 679 30605
rect 737 30596 751 30605
rect 809 30596 823 30605
rect 877 30596 895 30605
rect 449 30571 487 30596
rect 521 30571 559 30596
rect 593 30571 631 30596
rect 665 30571 703 30596
rect 737 30571 775 30596
rect 809 30571 843 30596
rect 877 30571 915 30596
rect 949 30571 983 30605
rect -23 30557 983 30571
rect -23 30503 -17 30557
rect 17 30537 75 30557
rect 109 30537 167 30557
rect 201 30537 259 30557
rect 293 30537 463 30557
rect 497 30537 535 30557
rect 569 30537 607 30557
rect 641 30537 679 30557
rect 713 30537 751 30557
rect 785 30537 823 30557
rect 17 30503 55 30537
rect 109 30523 127 30537
rect 89 30503 127 30523
rect 161 30523 167 30537
rect 233 30523 259 30537
rect 161 30503 199 30523
rect 233 30503 271 30523
rect 305 30503 343 30537
rect 377 30503 415 30537
rect 449 30523 463 30537
rect 521 30523 535 30537
rect 593 30523 607 30537
rect 665 30523 679 30537
rect 737 30523 751 30537
rect 809 30523 823 30537
rect 857 30523 895 30557
rect 929 30523 983 30557
rect 449 30503 487 30523
rect 521 30503 559 30523
rect 593 30503 631 30523
rect 665 30503 703 30523
rect 737 30503 775 30523
rect 809 30521 983 30523
rect 809 30503 843 30521
rect -23 30487 843 30503
rect 877 30487 915 30521
rect 949 30487 983 30521
rect -23 30484 983 30487
rect -23 30435 -17 30484
rect 17 30469 75 30484
rect 109 30469 167 30484
rect 201 30469 259 30484
rect 293 30469 463 30484
rect 497 30469 535 30484
rect 569 30469 607 30484
rect 641 30469 679 30484
rect 713 30469 751 30484
rect 785 30469 823 30484
rect 17 30435 55 30469
rect 109 30450 127 30469
rect 89 30435 127 30450
rect 161 30450 167 30469
rect 233 30450 259 30469
rect 161 30435 199 30450
rect 233 30435 271 30450
rect 305 30435 343 30469
rect 377 30435 415 30469
rect 449 30450 463 30469
rect 521 30450 535 30469
rect 593 30450 607 30469
rect 665 30450 679 30469
rect 737 30450 751 30469
rect 809 30450 823 30469
rect 857 30450 895 30484
rect 929 30450 983 30484
rect 449 30435 487 30450
rect 521 30435 559 30450
rect 593 30435 631 30450
rect 665 30435 703 30450
rect 737 30435 775 30450
rect 809 30436 983 30450
rect 809 30435 843 30436
rect -23 30411 843 30435
rect 877 30411 915 30436
rect -23 30367 -17 30411
rect 17 30401 75 30411
rect 109 30401 167 30411
rect 201 30401 259 30411
rect 293 30401 463 30411
rect 497 30401 535 30411
rect 569 30401 607 30411
rect 641 30401 679 30411
rect 713 30401 751 30411
rect 785 30401 823 30411
rect 877 30402 895 30411
rect 949 30402 983 30436
rect 17 30367 55 30401
rect 109 30377 127 30401
rect 89 30367 127 30377
rect 161 30377 167 30401
rect 233 30377 259 30401
rect 161 30367 199 30377
rect 233 30367 271 30377
rect 305 30367 343 30401
rect 377 30367 415 30401
rect 449 30377 463 30401
rect 521 30377 535 30401
rect 593 30377 607 30401
rect 665 30377 679 30401
rect 737 30377 751 30401
rect 809 30377 823 30401
rect 857 30377 895 30402
rect 929 30377 983 30402
rect 449 30367 487 30377
rect 521 30367 559 30377
rect 593 30367 631 30377
rect 665 30367 703 30377
rect 737 30367 775 30377
rect 809 30367 983 30377
rect -23 30351 983 30367
rect -23 30338 843 30351
rect 877 30338 915 30351
rect -23 30299 -17 30338
rect 17 30333 75 30338
rect 109 30333 167 30338
rect 201 30333 259 30338
rect 293 30333 463 30338
rect 497 30333 535 30338
rect 569 30333 607 30338
rect 641 30333 679 30338
rect 713 30333 751 30338
rect 785 30333 823 30338
rect 17 30299 55 30333
rect 109 30304 127 30333
rect 89 30299 127 30304
rect 161 30304 167 30333
rect 233 30304 259 30333
rect 161 30299 199 30304
rect 233 30299 271 30304
rect 305 30299 343 30333
rect 377 30299 415 30333
rect 449 30304 463 30333
rect 521 30304 535 30333
rect 593 30304 607 30333
rect 665 30304 679 30333
rect 737 30304 751 30333
rect 809 30304 823 30333
rect 877 30317 895 30338
rect 949 30317 983 30351
rect 857 30304 895 30317
rect 929 30304 983 30317
rect 449 30299 487 30304
rect 521 30299 559 30304
rect 593 30299 631 30304
rect 665 30299 703 30304
rect 737 30299 775 30304
rect 809 30299 983 30304
rect -23 30266 983 30299
rect -23 30265 843 30266
rect 877 30265 915 30266
rect -23 30231 -17 30265
rect 17 30231 55 30265
rect 109 30231 127 30265
rect 161 30231 167 30265
rect 233 30231 259 30265
rect 305 30231 343 30265
rect 377 30231 415 30265
rect 449 30231 463 30265
rect 521 30231 535 30265
rect 593 30231 607 30265
rect 665 30231 679 30265
rect 737 30231 751 30265
rect 809 30231 823 30265
rect 877 30232 895 30265
rect 949 30232 983 30266
rect 857 30231 895 30232
rect 929 30231 983 30232
rect -23 30197 983 30231
rect -23 30158 -17 30197
rect 17 30163 55 30197
rect 89 30192 127 30197
rect 109 30163 127 30192
rect 161 30192 199 30197
rect 233 30192 271 30197
rect 161 30163 167 30192
rect 233 30163 259 30192
rect 305 30163 343 30197
rect 377 30163 415 30197
rect 449 30192 487 30197
rect 521 30192 559 30197
rect 593 30192 631 30197
rect 665 30192 703 30197
rect 737 30192 775 30197
rect 809 30192 983 30197
rect 449 30163 463 30192
rect 521 30163 535 30192
rect 593 30163 607 30192
rect 665 30163 679 30192
rect 737 30163 751 30192
rect 809 30163 823 30192
rect 857 30181 895 30192
rect 929 30181 983 30192
rect 17 30158 75 30163
rect 109 30158 167 30163
rect 201 30158 259 30163
rect 293 30158 463 30163
rect 497 30158 535 30163
rect 569 30158 607 30163
rect 641 30158 679 30163
rect 713 30158 751 30163
rect 785 30158 823 30163
rect 877 30158 895 30181
rect -23 30147 843 30158
rect 877 30147 915 30158
rect 949 30147 983 30181
rect -23 30129 983 30147
rect -23 30085 -17 30129
rect 17 30095 55 30129
rect 89 30119 127 30129
rect 109 30095 127 30119
rect 161 30119 199 30129
rect 233 30119 271 30129
rect 161 30095 167 30119
rect 233 30095 259 30119
rect 305 30095 343 30129
rect 377 30095 415 30129
rect 449 30119 487 30129
rect 521 30119 559 30129
rect 593 30119 631 30129
rect 665 30119 703 30129
rect 737 30119 775 30129
rect 809 30119 983 30129
rect 449 30095 463 30119
rect 521 30095 535 30119
rect 593 30095 607 30119
rect 665 30095 679 30119
rect 737 30095 751 30119
rect 809 30095 823 30119
rect 857 30096 895 30119
rect 929 30096 983 30119
rect 17 30085 75 30095
rect 109 30085 167 30095
rect 201 30085 259 30095
rect 293 30085 463 30095
rect 497 30085 535 30095
rect 569 30085 607 30095
rect 641 30085 679 30095
rect 713 30085 751 30095
rect 785 30085 823 30095
rect 877 30085 895 30096
rect -23 30062 843 30085
rect 877 30062 915 30085
rect 949 30062 983 30096
rect -23 30061 983 30062
rect -23 30012 -17 30061
rect 17 30027 55 30061
rect 89 30046 127 30061
rect 109 30027 127 30046
rect 161 30046 199 30061
rect 233 30046 271 30061
rect 161 30027 167 30046
rect 233 30027 259 30046
rect 305 30027 343 30061
rect 377 30027 415 30061
rect 449 30046 487 30061
rect 521 30046 559 30061
rect 593 30046 631 30061
rect 665 30046 703 30061
rect 737 30046 775 30061
rect 809 30046 983 30061
rect 449 30027 463 30046
rect 521 30027 535 30046
rect 593 30027 607 30046
rect 665 30027 679 30046
rect 737 30027 751 30046
rect 809 30027 823 30046
rect 17 30012 75 30027
rect 109 30012 167 30027
rect 201 30012 259 30027
rect 293 30012 463 30027
rect 497 30012 535 30027
rect 569 30012 607 30027
rect 641 30012 679 30027
rect 713 30012 751 30027
rect 785 30012 823 30027
rect 857 30012 895 30046
rect 929 30012 983 30046
rect -23 30011 983 30012
rect -23 29993 843 30011
rect -23 29939 -17 29993
rect 17 29959 55 29993
rect 89 29973 127 29993
rect 109 29959 127 29973
rect 161 29973 199 29993
rect 233 29973 271 29993
rect 161 29959 167 29973
rect 233 29959 259 29973
rect 305 29959 343 29993
rect 377 29959 415 29993
rect 449 29973 487 29993
rect 521 29973 559 29993
rect 593 29973 631 29993
rect 665 29973 703 29993
rect 737 29973 775 29993
rect 809 29977 843 29993
rect 877 29977 915 30011
rect 949 29977 983 30011
rect 809 29973 983 29977
rect 449 29959 463 29973
rect 521 29959 535 29973
rect 593 29959 607 29973
rect 665 29959 679 29973
rect 737 29959 751 29973
rect 809 29959 823 29973
rect 17 29939 75 29959
rect 109 29939 167 29959
rect 201 29939 259 29959
rect 293 29939 463 29959
rect 497 29939 535 29959
rect 569 29939 607 29959
rect 641 29939 679 29959
rect 713 29939 751 29959
rect 785 29939 823 29959
rect 857 29939 895 29973
rect 929 29939 983 29973
rect -23 29926 983 29939
rect -23 29925 843 29926
rect -23 29866 -17 29925
rect 17 29891 55 29925
rect 89 29900 127 29925
rect 109 29891 127 29900
rect 161 29900 199 29925
rect 233 29900 271 29925
rect 161 29891 167 29900
rect 233 29891 259 29900
rect 305 29891 343 29925
rect 377 29891 415 29925
rect 449 29900 487 29925
rect 521 29900 559 29925
rect 593 29900 631 29925
rect 665 29900 703 29925
rect 737 29900 775 29925
rect 809 29900 843 29925
rect 877 29900 915 29926
rect 449 29891 463 29900
rect 521 29891 535 29900
rect 593 29891 607 29900
rect 665 29891 679 29900
rect 737 29891 751 29900
rect 809 29891 823 29900
rect 877 29892 895 29900
rect 949 29892 983 29926
rect 17 29866 75 29891
rect 109 29866 167 29891
rect 201 29866 259 29891
rect 293 29866 463 29891
rect 497 29866 535 29891
rect 569 29866 607 29891
rect 641 29866 679 29891
rect 713 29866 751 29891
rect 785 29866 823 29891
rect 857 29866 895 29892
rect 929 29866 983 29892
rect -23 29857 983 29866
rect -23 29793 -17 29857
rect 17 29823 55 29857
rect 89 29827 127 29857
rect 109 29823 127 29827
rect 161 29827 199 29857
rect 233 29827 271 29857
rect 161 29823 167 29827
rect 233 29823 259 29827
rect 305 29823 343 29857
rect 377 29823 415 29857
rect 449 29827 487 29857
rect 521 29827 559 29857
rect 593 29827 631 29857
rect 665 29827 703 29857
rect 737 29827 775 29857
rect 809 29841 983 29857
rect 809 29827 843 29841
rect 877 29827 915 29841
rect 449 29823 463 29827
rect 521 29823 535 29827
rect 593 29823 607 29827
rect 665 29823 679 29827
rect 737 29823 751 29827
rect 809 29823 823 29827
rect 17 29793 75 29823
rect 109 29793 167 29823
rect 201 29793 259 29823
rect 293 29793 463 29823
rect 497 29793 535 29823
rect 569 29793 607 29823
rect 641 29793 679 29823
rect 713 29793 751 29823
rect 785 29793 823 29823
rect 877 29807 895 29827
rect 949 29807 983 29841
rect 857 29793 895 29807
rect 929 29793 983 29807
rect -23 29789 983 29793
rect -23 29755 -17 29789
rect 17 29755 55 29789
rect 89 29755 127 29789
rect 161 29755 199 29789
rect 233 29755 271 29789
rect 305 29755 343 29789
rect 377 29755 415 29789
rect 449 29755 487 29789
rect 521 29755 559 29789
rect 593 29755 631 29789
rect 665 29755 703 29789
rect 737 29755 775 29789
rect 809 29756 983 29789
rect 809 29755 843 29756
rect -23 29754 843 29755
rect 877 29754 915 29756
rect -23 29687 -17 29754
rect 17 29721 75 29754
rect 109 29721 167 29754
rect 201 29721 259 29754
rect 293 29721 463 29754
rect 497 29721 535 29754
rect 569 29721 607 29754
rect 641 29721 679 29754
rect 713 29721 751 29754
rect 785 29721 823 29754
rect 877 29722 895 29754
rect 949 29722 983 29756
rect 17 29687 55 29721
rect 109 29720 127 29721
rect 89 29687 127 29720
rect 161 29720 167 29721
rect 233 29720 259 29721
rect 161 29687 199 29720
rect 233 29687 271 29720
rect 305 29687 343 29721
rect 377 29687 415 29721
rect 449 29720 463 29721
rect 521 29720 535 29721
rect 593 29720 607 29721
rect 665 29720 679 29721
rect 737 29720 751 29721
rect 809 29720 823 29721
rect 857 29720 895 29722
rect 929 29720 983 29722
rect 449 29687 487 29720
rect 521 29687 559 29720
rect 593 29687 631 29720
rect 665 29687 703 29720
rect 737 29687 775 29720
rect 809 29687 983 29720
rect -23 29681 983 29687
rect -23 29618 -17 29681
rect 17 29652 75 29681
rect 109 29652 167 29681
rect 201 29652 259 29681
rect 293 29652 463 29681
rect 497 29652 535 29681
rect 569 29652 607 29681
rect 641 29652 679 29681
rect 713 29652 751 29681
rect 785 29652 823 29681
rect 857 29671 895 29681
rect 929 29671 983 29681
rect 17 29618 55 29652
rect 109 29647 127 29652
rect 89 29618 127 29647
rect 161 29647 167 29652
rect 233 29647 259 29652
rect 161 29618 199 29647
rect 233 29618 271 29647
rect 305 29618 343 29652
rect 377 29618 415 29652
rect 449 29647 463 29652
rect 521 29647 535 29652
rect 593 29647 607 29652
rect 665 29647 679 29652
rect 737 29647 751 29652
rect 809 29647 823 29652
rect 877 29647 895 29671
rect 449 29618 487 29647
rect 521 29618 559 29647
rect 593 29618 631 29647
rect 665 29618 703 29647
rect 737 29618 775 29647
rect 809 29637 843 29647
rect 877 29637 915 29647
rect 949 29637 983 29671
rect 809 29618 983 29637
rect -23 29608 983 29618
rect -23 29549 -17 29608
rect 17 29583 75 29608
rect 109 29583 167 29608
rect 201 29583 259 29608
rect 293 29583 463 29608
rect 497 29583 535 29608
rect 569 29583 607 29608
rect 641 29583 679 29608
rect 713 29583 751 29608
rect 785 29583 823 29608
rect 857 29586 895 29608
rect 929 29586 983 29608
rect 17 29549 55 29583
rect 109 29574 127 29583
rect 89 29549 127 29574
rect 161 29574 167 29583
rect 233 29574 259 29583
rect 161 29549 199 29574
rect 233 29549 271 29574
rect 305 29549 343 29583
rect 377 29549 415 29583
rect 449 29574 463 29583
rect 521 29574 535 29583
rect 593 29574 607 29583
rect 665 29574 679 29583
rect 737 29574 751 29583
rect 809 29574 823 29583
rect 877 29574 895 29586
rect 449 29549 487 29574
rect 521 29549 559 29574
rect 593 29549 631 29574
rect 665 29549 703 29574
rect 737 29549 775 29574
rect 809 29552 843 29574
rect 877 29552 915 29574
rect 949 29552 983 29586
rect 809 29549 983 29552
rect -23 29535 983 29549
rect -23 29480 -17 29535
rect 17 29514 75 29535
rect 109 29514 167 29535
rect 201 29514 259 29535
rect 293 29514 463 29535
rect 497 29514 535 29535
rect 569 29514 607 29535
rect 641 29514 679 29535
rect 713 29514 751 29535
rect 785 29514 823 29535
rect 17 29480 55 29514
rect 109 29501 127 29514
rect 89 29480 127 29501
rect 161 29501 167 29514
rect 233 29501 259 29514
rect 161 29480 199 29501
rect 233 29480 271 29501
rect 305 29480 343 29514
rect 377 29480 415 29514
rect 449 29501 463 29514
rect 521 29501 535 29514
rect 593 29501 607 29514
rect 665 29501 679 29514
rect 737 29501 751 29514
rect 809 29501 823 29514
rect 857 29501 895 29535
rect 929 29501 983 29535
rect 449 29480 487 29501
rect 521 29480 559 29501
rect 593 29480 631 29501
rect 665 29480 703 29501
rect 737 29480 775 29501
rect 809 29480 843 29501
rect -23 29467 843 29480
rect 877 29467 915 29501
rect 949 29467 983 29501
rect -23 29462 983 29467
rect -23 29411 -17 29462
rect 17 29445 75 29462
rect 109 29445 167 29462
rect 201 29445 259 29462
rect 293 29445 463 29462
rect 497 29445 535 29462
rect 569 29445 607 29462
rect 641 29445 679 29462
rect 713 29445 751 29462
rect 785 29445 823 29462
rect 17 29411 55 29445
rect 109 29428 127 29445
rect 89 29411 127 29428
rect 161 29428 167 29445
rect 233 29428 259 29445
rect 161 29411 199 29428
rect 233 29411 271 29428
rect 305 29411 343 29445
rect 377 29411 415 29445
rect 449 29428 463 29445
rect 521 29428 535 29445
rect 593 29428 607 29445
rect 665 29428 679 29445
rect 737 29428 751 29445
rect 809 29428 823 29445
rect 857 29428 895 29462
rect 929 29428 983 29462
rect 449 29411 487 29428
rect 521 29411 559 29428
rect 593 29411 631 29428
rect 665 29411 703 29428
rect 737 29411 775 29428
rect 809 29416 983 29428
rect 809 29411 843 29416
rect -23 29389 843 29411
rect 877 29389 915 29416
rect -23 29342 -17 29389
rect 17 29376 75 29389
rect 109 29376 167 29389
rect 201 29376 259 29389
rect 293 29376 463 29389
rect 497 29376 535 29389
rect 569 29376 607 29389
rect 641 29376 679 29389
rect 713 29376 751 29389
rect 785 29376 823 29389
rect 877 29382 895 29389
rect 949 29382 983 29416
rect 17 29342 55 29376
rect 109 29355 127 29376
rect 89 29342 127 29355
rect 161 29355 167 29376
rect 233 29355 259 29376
rect 161 29342 199 29355
rect 233 29342 271 29355
rect 305 29342 343 29376
rect 377 29342 415 29376
rect 449 29355 463 29376
rect 521 29355 535 29376
rect 593 29355 607 29376
rect 665 29355 679 29376
rect 737 29355 751 29376
rect 809 29355 823 29376
rect 857 29355 895 29382
rect 929 29355 983 29382
rect 449 29342 487 29355
rect 521 29342 559 29355
rect 593 29342 631 29355
rect 665 29342 703 29355
rect 737 29342 775 29355
rect 809 29342 983 29355
rect -23 29331 983 29342
rect -23 29316 843 29331
rect 877 29316 915 29331
rect -23 29273 -17 29316
rect 17 29307 75 29316
rect 109 29307 167 29316
rect 201 29307 259 29316
rect 293 29307 463 29316
rect 497 29307 535 29316
rect 569 29307 607 29316
rect 641 29307 679 29316
rect 713 29307 751 29316
rect 785 29307 823 29316
rect 17 29273 55 29307
rect 109 29282 127 29307
rect 89 29273 127 29282
rect 161 29282 167 29307
rect 233 29282 259 29307
rect 161 29273 199 29282
rect 233 29273 271 29282
rect 305 29273 343 29307
rect 377 29273 415 29307
rect 449 29282 463 29307
rect 521 29282 535 29307
rect 593 29282 607 29307
rect 665 29282 679 29307
rect 737 29282 751 29307
rect 809 29282 823 29307
rect 877 29297 895 29316
rect 949 29297 983 29331
rect 857 29282 895 29297
rect 929 29282 983 29297
rect 449 29273 487 29282
rect 521 29273 559 29282
rect 593 29273 631 29282
rect 665 29273 703 29282
rect 737 29273 775 29282
rect 809 29273 983 29282
rect -23 29246 983 29273
rect -23 29243 843 29246
rect 877 29243 915 29246
rect -23 29204 -17 29243
rect 17 29238 75 29243
rect 109 29238 167 29243
rect 201 29238 259 29243
rect 293 29238 463 29243
rect 497 29238 535 29243
rect 569 29238 607 29243
rect 641 29238 679 29243
rect 713 29238 751 29243
rect 785 29238 823 29243
rect 17 29204 55 29238
rect 109 29209 127 29238
rect 89 29204 127 29209
rect 161 29209 167 29238
rect 233 29209 259 29238
rect 161 29204 199 29209
rect 233 29204 271 29209
rect 305 29204 343 29238
rect 377 29204 415 29238
rect 449 29209 463 29238
rect 521 29209 535 29238
rect 593 29209 607 29238
rect 665 29209 679 29238
rect 737 29209 751 29238
rect 809 29209 823 29238
rect 877 29212 895 29243
rect 949 29212 983 29246
rect 857 29209 895 29212
rect 929 29209 983 29212
rect 449 29204 487 29209
rect 521 29204 559 29209
rect 593 29204 631 29209
rect 665 29204 703 29209
rect 737 29204 775 29209
rect 809 29204 983 29209
rect -23 29170 983 29204
rect -23 29135 -17 29170
rect 17 29169 75 29170
rect 109 29169 167 29170
rect 201 29169 259 29170
rect 293 29169 463 29170
rect 497 29169 535 29170
rect 569 29169 607 29170
rect 641 29169 679 29170
rect 713 29169 751 29170
rect 785 29169 823 29170
rect 17 29135 55 29169
rect 109 29136 127 29169
rect 89 29135 127 29136
rect 161 29136 167 29169
rect 233 29136 259 29169
rect 161 29135 199 29136
rect 233 29135 271 29136
rect 305 29135 343 29169
rect 377 29135 415 29169
rect 449 29136 463 29169
rect 521 29136 535 29169
rect 593 29136 607 29169
rect 665 29136 679 29169
rect 737 29136 751 29169
rect 809 29136 823 29169
rect 857 29161 895 29170
rect 929 29161 983 29170
rect 877 29136 895 29161
rect 449 29135 487 29136
rect 521 29135 559 29136
rect 593 29135 631 29136
rect 665 29135 703 29136
rect 737 29135 775 29136
rect 809 29135 843 29136
rect -23 29127 843 29135
rect 877 29127 915 29136
rect 949 29127 983 29161
rect -23 29100 983 29127
rect -23 29063 -17 29100
rect 17 29066 55 29100
rect 89 29097 127 29100
rect 109 29066 127 29097
rect 161 29097 199 29100
rect 233 29097 271 29100
rect 161 29066 167 29097
rect 233 29066 259 29097
rect 305 29066 343 29100
rect 377 29066 415 29100
rect 449 29097 487 29100
rect 521 29097 559 29100
rect 593 29097 631 29100
rect 665 29097 703 29100
rect 737 29097 775 29100
rect 809 29097 983 29100
rect 449 29066 463 29097
rect 521 29066 535 29097
rect 593 29066 607 29097
rect 665 29066 679 29097
rect 737 29066 751 29097
rect 809 29066 823 29097
rect 857 29076 895 29097
rect 929 29076 983 29097
rect 17 29063 75 29066
rect 109 29063 167 29066
rect 201 29063 259 29066
rect 293 29063 463 29066
rect 497 29063 535 29066
rect 569 29063 607 29066
rect 641 29063 679 29066
rect 713 29063 751 29066
rect 785 29063 823 29066
rect 877 29063 895 29076
rect -23 29042 843 29063
rect 877 29042 915 29063
rect 949 29042 983 29076
rect -23 29031 299 29042
rect 452 29031 940 29042
rect -23 28010 299 28030
rect -23 27998 843 28010
rect -23 27952 -17 27998
rect 17 27986 75 27998
rect 109 27986 167 27998
rect 201 27986 259 27998
rect 293 27986 843 27998
rect 17 27952 55 27986
rect 109 27964 127 27986
rect 89 27952 127 27964
rect 161 27964 167 27986
rect 233 27964 259 27986
rect 161 27952 199 27964
rect 233 27952 271 27964
rect 305 27952 343 27986
rect 377 27952 415 27986
rect 449 27978 487 27986
rect 521 27978 559 27986
rect 593 27978 631 27986
rect 665 27978 703 27986
rect 737 27978 775 27986
rect 809 27978 843 27986
rect 877 27978 915 28010
rect 449 27952 463 27978
rect 521 27952 535 27978
rect 593 27952 607 27978
rect 665 27952 679 27978
rect 737 27952 751 27978
rect 809 27952 823 27978
rect 877 27976 895 27978
rect 949 27976 983 28010
rect -23 27944 463 27952
rect 497 27944 535 27952
rect 569 27944 607 27952
rect 641 27944 679 27952
rect 713 27944 751 27952
rect 785 27944 823 27952
rect 857 27944 895 27976
rect 929 27944 983 27976
rect -23 27942 983 27944
rect -23 27925 843 27942
rect -23 27883 -17 27925
rect 17 27917 75 27925
rect 109 27917 167 27925
rect 201 27917 259 27925
rect 293 27917 843 27925
rect 17 27883 55 27917
rect 109 27891 127 27917
rect 89 27883 127 27891
rect 161 27891 167 27917
rect 233 27891 259 27917
rect 161 27883 199 27891
rect 233 27883 271 27891
rect 305 27883 343 27917
rect 377 27883 415 27917
rect 449 27903 487 27917
rect 521 27903 559 27917
rect 593 27903 631 27917
rect 665 27903 703 27917
rect 737 27903 775 27917
rect 809 27908 843 27917
rect 877 27908 915 27942
rect 949 27908 983 27942
rect 809 27903 983 27908
rect 449 27883 463 27903
rect 521 27883 535 27903
rect 593 27883 607 27903
rect 665 27883 679 27903
rect 737 27883 751 27903
rect 809 27883 823 27903
rect -23 27869 463 27883
rect 497 27869 535 27883
rect 569 27869 607 27883
rect 641 27869 679 27883
rect 713 27869 751 27883
rect 785 27869 823 27883
rect 857 27874 895 27903
rect 929 27874 983 27903
rect 877 27869 895 27874
rect -23 27852 843 27869
rect -23 27814 -17 27852
rect 17 27848 75 27852
rect 109 27848 167 27852
rect 201 27848 259 27852
rect 293 27848 843 27852
rect 17 27814 55 27848
rect 109 27818 127 27848
rect 89 27814 127 27818
rect 161 27818 167 27848
rect 233 27818 259 27848
rect 161 27814 199 27818
rect 233 27814 271 27818
rect 305 27814 343 27848
rect 377 27814 415 27848
rect 449 27828 487 27848
rect 521 27828 559 27848
rect 593 27828 631 27848
rect 665 27828 703 27848
rect 737 27828 775 27848
rect 809 27840 843 27848
rect 877 27840 915 27869
rect 949 27840 983 27874
rect 809 27828 983 27840
rect 449 27814 463 27828
rect 521 27814 535 27828
rect 593 27814 607 27828
rect 665 27814 679 27828
rect 737 27814 751 27828
rect 809 27814 823 27828
rect -23 27794 463 27814
rect 497 27794 535 27814
rect 569 27794 607 27814
rect 641 27794 679 27814
rect 713 27794 751 27814
rect 785 27794 823 27814
rect 857 27806 895 27828
rect 929 27806 983 27828
rect 877 27794 895 27806
rect -23 27779 843 27794
rect -23 27745 -17 27779
rect 17 27745 55 27779
rect 109 27745 127 27779
rect 161 27745 167 27779
rect 233 27745 259 27779
rect 305 27745 343 27779
rect 377 27745 415 27779
rect 449 27753 487 27779
rect 521 27753 559 27779
rect 593 27753 631 27779
rect 665 27753 703 27779
rect 737 27753 775 27779
rect 809 27772 843 27779
rect 877 27772 915 27794
rect 949 27772 983 27806
rect 809 27753 983 27772
rect 449 27745 463 27753
rect 521 27745 535 27753
rect 593 27745 607 27753
rect 665 27745 679 27753
rect 737 27745 751 27753
rect 809 27745 823 27753
rect -23 27719 463 27745
rect 497 27719 535 27745
rect 569 27719 607 27745
rect 641 27719 679 27745
rect 713 27719 751 27745
rect 785 27719 823 27745
rect 857 27738 895 27753
rect 929 27738 983 27753
rect 877 27719 895 27738
rect -23 27710 843 27719
rect -23 27672 -17 27710
rect 17 27676 55 27710
rect 89 27706 127 27710
rect 109 27676 127 27706
rect 161 27706 199 27710
rect 233 27706 271 27710
rect 161 27676 167 27706
rect 233 27676 259 27706
rect 305 27676 343 27710
rect 377 27676 415 27710
rect 449 27678 487 27710
rect 521 27678 559 27710
rect 593 27678 631 27710
rect 665 27678 703 27710
rect 737 27678 775 27710
rect 809 27704 843 27710
rect 877 27704 915 27719
rect 949 27704 983 27738
rect 809 27678 983 27704
rect 449 27676 463 27678
rect 521 27676 535 27678
rect 593 27676 607 27678
rect 665 27676 679 27678
rect 737 27676 751 27678
rect 809 27676 823 27678
rect 17 27672 75 27676
rect 109 27672 167 27676
rect 201 27672 259 27676
rect 293 27672 463 27676
rect -23 27644 463 27672
rect 497 27644 535 27676
rect 569 27644 607 27676
rect 641 27644 679 27676
rect 713 27644 751 27676
rect 785 27644 823 27676
rect 857 27670 895 27678
rect 929 27670 983 27678
rect 877 27644 895 27670
rect -23 27641 843 27644
rect -23 27599 -17 27641
rect 17 27607 55 27641
rect 89 27633 127 27641
rect 109 27607 127 27633
rect 161 27633 199 27641
rect 233 27633 271 27641
rect 161 27607 167 27633
rect 233 27607 259 27633
rect 305 27607 343 27641
rect 377 27607 415 27641
rect 449 27607 487 27641
rect 521 27607 559 27641
rect 593 27607 631 27641
rect 665 27607 703 27641
rect 737 27607 775 27641
rect 809 27636 843 27641
rect 877 27636 915 27644
rect 949 27636 983 27670
rect 809 27607 983 27636
rect 17 27599 75 27607
rect 109 27599 167 27607
rect 201 27599 259 27607
rect 293 27603 983 27607
rect 293 27599 463 27603
rect -23 27572 463 27599
rect 497 27572 535 27603
rect 569 27572 607 27603
rect 641 27572 679 27603
rect 713 27572 751 27603
rect 785 27572 823 27603
rect 857 27602 895 27603
rect 929 27602 983 27603
rect -23 27526 -17 27572
rect 17 27538 55 27572
rect 89 27560 127 27572
rect 109 27538 127 27560
rect 161 27560 199 27572
rect 233 27560 271 27572
rect 161 27538 167 27560
rect 233 27538 259 27560
rect 305 27538 343 27572
rect 377 27538 415 27572
rect 449 27569 463 27572
rect 521 27569 535 27572
rect 593 27569 607 27572
rect 665 27569 679 27572
rect 737 27569 751 27572
rect 809 27569 823 27572
rect 877 27569 895 27602
rect 449 27538 487 27569
rect 521 27538 559 27569
rect 593 27538 631 27569
rect 665 27538 703 27569
rect 737 27538 775 27569
rect 809 27568 843 27569
rect 877 27568 915 27569
rect 949 27568 983 27602
rect 809 27538 983 27568
rect 17 27526 75 27538
rect 109 27526 167 27538
rect 201 27526 259 27538
rect 293 27534 983 27538
rect 293 27528 843 27534
rect 877 27528 915 27534
rect 293 27526 463 27528
rect -23 27503 463 27526
rect 497 27503 535 27528
rect 569 27503 607 27528
rect 641 27503 679 27528
rect 713 27503 751 27528
rect 785 27503 823 27528
rect -23 27453 -17 27503
rect 17 27469 55 27503
rect 89 27487 127 27503
rect 109 27469 127 27487
rect 161 27487 199 27503
rect 233 27487 271 27503
rect 161 27469 167 27487
rect 233 27469 259 27487
rect 305 27469 343 27503
rect 377 27469 415 27503
rect 449 27494 463 27503
rect 521 27494 535 27503
rect 593 27494 607 27503
rect 665 27494 679 27503
rect 737 27494 751 27503
rect 809 27494 823 27503
rect 877 27500 895 27528
rect 949 27500 983 27534
rect 857 27494 895 27500
rect 929 27494 983 27500
rect 449 27469 487 27494
rect 521 27469 559 27494
rect 593 27469 631 27494
rect 665 27469 703 27494
rect 737 27469 775 27494
rect 809 27469 983 27494
rect 17 27453 75 27469
rect 109 27453 167 27469
rect 201 27453 259 27469
rect 293 27466 983 27469
rect 293 27453 843 27466
rect 877 27453 915 27466
rect -23 27434 463 27453
rect 497 27434 535 27453
rect 569 27434 607 27453
rect 641 27434 679 27453
rect 713 27434 751 27453
rect 785 27434 823 27453
rect -23 27380 -17 27434
rect 17 27400 55 27434
rect 89 27414 127 27434
rect 109 27400 127 27414
rect 161 27414 199 27434
rect 233 27414 271 27434
rect 161 27400 167 27414
rect 233 27400 259 27414
rect 305 27400 343 27434
rect 377 27400 415 27434
rect 449 27419 463 27434
rect 521 27419 535 27434
rect 593 27419 607 27434
rect 665 27419 679 27434
rect 737 27419 751 27434
rect 809 27419 823 27434
rect 877 27432 895 27453
rect 949 27432 983 27466
rect 857 27419 895 27432
rect 929 27419 983 27432
rect 449 27400 487 27419
rect 521 27400 559 27419
rect 593 27400 631 27419
rect 665 27400 703 27419
rect 737 27400 775 27419
rect 809 27400 983 27419
rect 17 27380 75 27400
rect 109 27380 167 27400
rect 201 27380 259 27400
rect 293 27398 983 27400
rect 293 27380 843 27398
rect -23 27378 843 27380
rect 877 27378 915 27398
rect -23 27365 463 27378
rect 497 27365 535 27378
rect 569 27365 607 27378
rect 641 27365 679 27378
rect 713 27365 751 27378
rect 785 27365 823 27378
rect -23 27307 -17 27365
rect 17 27331 55 27365
rect 89 27341 127 27365
rect 109 27331 127 27341
rect 161 27341 199 27365
rect 233 27341 271 27365
rect 161 27331 167 27341
rect 233 27331 259 27341
rect 305 27331 343 27365
rect 377 27331 415 27365
rect 449 27344 463 27365
rect 521 27344 535 27365
rect 593 27344 607 27365
rect 665 27344 679 27365
rect 737 27344 751 27365
rect 809 27344 823 27365
rect 877 27364 895 27378
rect 949 27364 983 27398
rect 857 27344 895 27364
rect 929 27344 983 27364
rect 449 27331 487 27344
rect 521 27331 559 27344
rect 593 27331 631 27344
rect 665 27331 703 27344
rect 737 27331 775 27344
rect 809 27331 983 27344
rect 17 27307 75 27331
rect 109 27307 167 27331
rect 201 27307 259 27331
rect 293 27330 983 27331
rect 293 27307 843 27330
rect -23 27303 843 27307
rect 877 27303 915 27330
rect -23 27296 463 27303
rect 497 27296 535 27303
rect 569 27296 607 27303
rect 641 27296 679 27303
rect 713 27296 751 27303
rect 785 27296 823 27303
rect 877 27296 895 27303
rect 949 27296 983 27330
rect -23 27234 -17 27296
rect 17 27262 55 27296
rect 89 27268 127 27296
rect 109 27262 127 27268
rect 161 27268 199 27296
rect 233 27268 271 27296
rect 161 27262 167 27268
rect 233 27262 259 27268
rect 305 27262 343 27296
rect 377 27262 415 27296
rect 449 27269 463 27296
rect 521 27269 535 27296
rect 593 27269 607 27296
rect 665 27269 679 27296
rect 737 27269 751 27296
rect 809 27269 823 27296
rect 857 27269 895 27296
rect 929 27269 983 27296
rect 449 27262 487 27269
rect 521 27262 559 27269
rect 593 27262 631 27269
rect 665 27262 703 27269
rect 737 27262 775 27269
rect 809 27262 983 27269
rect 17 27234 75 27262
rect 109 27234 167 27262
rect 201 27234 259 27262
rect 293 27234 843 27262
rect -23 27228 843 27234
rect 877 27228 915 27262
rect 949 27228 983 27262
rect -23 27227 463 27228
rect 497 27227 535 27228
rect 569 27227 607 27228
rect 641 27227 679 27228
rect 713 27227 751 27228
rect 785 27227 823 27228
rect -23 27161 -17 27227
rect 17 27193 55 27227
rect 89 27195 127 27227
rect 109 27193 127 27195
rect 161 27195 199 27227
rect 233 27195 271 27227
rect 161 27193 167 27195
rect 233 27193 259 27195
rect 305 27193 343 27227
rect 377 27193 415 27227
rect 449 27194 463 27227
rect 521 27194 535 27227
rect 593 27194 607 27227
rect 665 27194 679 27227
rect 737 27194 751 27227
rect 809 27194 823 27227
rect 857 27194 895 27228
rect 929 27194 983 27228
rect 449 27193 487 27194
rect 521 27193 559 27194
rect 593 27193 631 27194
rect 665 27193 703 27194
rect 737 27193 775 27194
rect 809 27193 843 27194
rect 17 27161 75 27193
rect 109 27161 167 27193
rect 201 27161 259 27193
rect 293 27161 843 27193
rect -23 27160 843 27161
rect 877 27160 915 27194
rect 949 27160 983 27194
rect -23 27158 983 27160
rect -23 27124 -17 27158
rect 17 27124 55 27158
rect 89 27124 127 27158
rect 161 27124 199 27158
rect 233 27124 271 27158
rect 305 27124 343 27158
rect 377 27124 415 27158
rect 449 27153 487 27158
rect 521 27153 559 27158
rect 593 27153 631 27158
rect 665 27153 703 27158
rect 737 27153 775 27158
rect 809 27153 983 27158
rect 449 27124 463 27153
rect 521 27124 535 27153
rect 593 27124 607 27153
rect 665 27124 679 27153
rect 737 27124 751 27153
rect 809 27124 823 27153
rect 857 27126 895 27153
rect 929 27126 983 27153
rect -23 27122 463 27124
rect -23 27055 -17 27122
rect 17 27089 75 27122
rect 109 27089 167 27122
rect 201 27089 259 27122
rect 293 27119 463 27122
rect 497 27119 535 27124
rect 569 27119 607 27124
rect 641 27119 679 27124
rect 713 27119 751 27124
rect 785 27119 823 27124
rect 877 27119 895 27126
rect 293 27092 843 27119
rect 877 27092 915 27119
rect 949 27092 983 27126
rect 293 27089 983 27092
rect 17 27055 55 27089
rect 109 27088 127 27089
rect 89 27055 127 27088
rect 161 27088 167 27089
rect 233 27088 259 27089
rect 161 27055 199 27088
rect 233 27055 271 27088
rect 305 27055 343 27089
rect 377 27055 415 27089
rect 449 27079 487 27089
rect 521 27079 559 27089
rect 593 27079 631 27089
rect 665 27079 703 27089
rect 737 27079 775 27089
rect 809 27079 983 27089
rect 449 27055 463 27079
rect 521 27055 535 27079
rect 593 27055 607 27079
rect 665 27055 679 27079
rect 737 27055 751 27079
rect 809 27055 823 27079
rect 857 27058 895 27079
rect 929 27058 983 27079
rect -23 27049 463 27055
rect -23 26986 -17 27049
rect 17 27020 75 27049
rect 109 27020 167 27049
rect 201 27020 259 27049
rect 293 27045 463 27049
rect 497 27045 535 27055
rect 569 27045 607 27055
rect 641 27045 679 27055
rect 713 27045 751 27055
rect 785 27045 823 27055
rect 877 27045 895 27058
rect 293 27024 843 27045
rect 877 27024 915 27045
rect 949 27024 983 27058
rect 293 27020 983 27024
rect 17 26986 55 27020
rect 109 27015 127 27020
rect 89 26986 127 27015
rect 161 27015 167 27020
rect 233 27015 259 27020
rect 161 26986 199 27015
rect 233 26986 271 27015
rect 305 26986 343 27020
rect 377 26986 415 27020
rect 449 27005 487 27020
rect 521 27005 559 27020
rect 593 27005 631 27020
rect 665 27005 703 27020
rect 737 27005 775 27020
rect 809 27005 983 27020
rect 449 26986 463 27005
rect 521 26986 535 27005
rect 593 26986 607 27005
rect 665 26986 679 27005
rect 737 26986 751 27005
rect 809 26986 823 27005
rect 857 26990 895 27005
rect 929 26990 983 27005
rect -23 26976 463 26986
rect -23 26917 -17 26976
rect 17 26951 75 26976
rect 109 26951 167 26976
rect 201 26951 259 26976
rect 293 26971 463 26976
rect 497 26971 535 26986
rect 569 26971 607 26986
rect 641 26971 679 26986
rect 713 26971 751 26986
rect 785 26971 823 26986
rect 877 26971 895 26990
rect 293 26956 843 26971
rect 877 26956 915 26971
rect 949 26956 983 26990
rect 293 26951 983 26956
rect 17 26917 55 26951
rect 109 26942 127 26951
rect 89 26917 127 26942
rect 161 26942 167 26951
rect 233 26942 259 26951
rect 161 26917 199 26942
rect 233 26917 271 26942
rect 305 26917 343 26951
rect 377 26917 415 26951
rect 449 26931 487 26951
rect 521 26931 559 26951
rect 593 26931 631 26951
rect 665 26931 703 26951
rect 737 26931 775 26951
rect 809 26931 983 26951
rect 449 26917 463 26931
rect 521 26917 535 26931
rect 593 26917 607 26931
rect 665 26917 679 26931
rect 737 26917 751 26931
rect 809 26917 823 26931
rect 857 26922 895 26931
rect 929 26922 983 26931
rect -23 26903 463 26917
rect -23 26848 -17 26903
rect 17 26882 75 26903
rect 109 26882 167 26903
rect 201 26882 259 26903
rect 293 26897 463 26903
rect 497 26897 535 26917
rect 569 26897 607 26917
rect 641 26897 679 26917
rect 713 26897 751 26917
rect 785 26897 823 26917
rect 877 26897 895 26922
rect 293 26888 843 26897
rect 877 26888 915 26897
rect 949 26888 983 26922
rect 293 26882 983 26888
rect 17 26848 55 26882
rect 109 26869 127 26882
rect 89 26848 127 26869
rect 161 26869 167 26882
rect 233 26869 259 26882
rect 161 26848 199 26869
rect 233 26848 271 26869
rect 305 26848 343 26882
rect 377 26848 415 26882
rect 449 26857 487 26882
rect 521 26857 559 26882
rect 593 26857 631 26882
rect 665 26857 703 26882
rect 737 26857 775 26882
rect 809 26857 983 26882
rect 449 26848 463 26857
rect 521 26848 535 26857
rect 593 26848 607 26857
rect 665 26848 679 26857
rect 737 26848 751 26857
rect 809 26848 823 26857
rect 857 26854 895 26857
rect 929 26854 983 26857
rect -23 26830 463 26848
rect -23 26779 -17 26830
rect 17 26813 75 26830
rect 109 26813 167 26830
rect 201 26813 259 26830
rect 293 26823 463 26830
rect 497 26823 535 26848
rect 569 26823 607 26848
rect 641 26823 679 26848
rect 713 26823 751 26848
rect 785 26823 823 26848
rect 877 26823 895 26854
rect 293 26820 843 26823
rect 877 26820 915 26823
rect 949 26820 983 26854
rect 293 26813 983 26820
rect 17 26779 55 26813
rect 109 26796 127 26813
rect 89 26779 127 26796
rect 161 26796 167 26813
rect 233 26796 259 26813
rect 161 26779 199 26796
rect 233 26779 271 26796
rect 305 26779 343 26813
rect 377 26779 415 26813
rect 449 26783 487 26813
rect 521 26783 559 26813
rect 593 26783 631 26813
rect 665 26783 703 26813
rect 737 26783 775 26813
rect 809 26785 983 26813
rect 809 26783 843 26785
rect 877 26783 915 26785
rect 449 26779 463 26783
rect 521 26779 535 26783
rect 593 26779 607 26783
rect 665 26779 679 26783
rect 737 26779 751 26783
rect 809 26779 823 26783
rect -23 26757 463 26779
rect -23 26710 -17 26757
rect 17 26744 75 26757
rect 109 26744 167 26757
rect 201 26744 259 26757
rect 293 26749 463 26757
rect 497 26749 535 26779
rect 569 26749 607 26779
rect 641 26749 679 26779
rect 713 26749 751 26779
rect 785 26749 823 26779
rect 877 26751 895 26783
rect 949 26751 983 26785
rect 857 26749 895 26751
rect 929 26749 983 26751
rect 293 26744 983 26749
rect 17 26710 55 26744
rect 109 26723 127 26744
rect 89 26710 127 26723
rect 161 26723 167 26744
rect 233 26723 259 26744
rect 161 26710 199 26723
rect 233 26710 271 26723
rect 305 26710 343 26744
rect 377 26710 415 26744
rect 449 26710 487 26744
rect 521 26710 559 26744
rect 593 26710 631 26744
rect 665 26710 703 26744
rect 737 26710 775 26744
rect 809 26716 983 26744
rect 809 26710 843 26716
rect -23 26709 843 26710
rect 877 26709 915 26716
rect -23 26684 463 26709
rect -23 26641 -17 26684
rect 17 26675 75 26684
rect 109 26675 167 26684
rect 201 26675 259 26684
rect 293 26675 463 26684
rect 497 26675 535 26709
rect 569 26675 607 26709
rect 641 26675 679 26709
rect 713 26675 751 26709
rect 785 26675 823 26709
rect 877 26682 895 26709
rect 949 26682 983 26716
rect 857 26675 895 26682
rect 929 26675 983 26682
rect 17 26641 55 26675
rect 109 26650 127 26675
rect 89 26641 127 26650
rect 161 26650 167 26675
rect 233 26650 259 26675
rect 161 26641 199 26650
rect 233 26641 271 26650
rect 305 26641 343 26675
rect 377 26641 415 26675
rect 449 26641 487 26675
rect 521 26641 559 26675
rect 593 26641 631 26675
rect 665 26641 703 26675
rect 737 26641 775 26675
rect 809 26647 983 26675
rect 809 26641 843 26647
rect -23 26635 843 26641
rect 877 26635 915 26647
rect -23 26611 463 26635
rect -23 26572 -17 26611
rect 17 26606 75 26611
rect 109 26606 167 26611
rect 201 26606 259 26611
rect 293 26606 463 26611
rect 497 26606 535 26635
rect 569 26606 607 26635
rect 641 26606 679 26635
rect 713 26606 751 26635
rect 785 26606 823 26635
rect 877 26613 895 26635
rect 949 26613 983 26647
rect 17 26572 55 26606
rect 109 26577 127 26606
rect 89 26572 127 26577
rect 161 26577 167 26606
rect 233 26577 259 26606
rect 161 26572 199 26577
rect 233 26572 271 26577
rect 305 26572 343 26606
rect 377 26572 415 26606
rect 449 26601 463 26606
rect 521 26601 535 26606
rect 593 26601 607 26606
rect 665 26601 679 26606
rect 737 26601 751 26606
rect 809 26601 823 26606
rect 857 26601 895 26613
rect 929 26601 983 26613
rect 449 26572 487 26601
rect 521 26572 559 26601
rect 593 26572 631 26601
rect 665 26572 703 26601
rect 737 26572 775 26601
rect 809 26578 983 26601
rect 809 26572 843 26578
rect -23 26561 843 26572
rect 877 26561 915 26578
rect -23 26538 463 26561
rect -23 26503 -17 26538
rect 17 26537 75 26538
rect 109 26537 167 26538
rect 201 26537 259 26538
rect 293 26537 463 26538
rect 497 26537 535 26561
rect 569 26537 607 26561
rect 641 26537 679 26561
rect 713 26537 751 26561
rect 785 26537 823 26561
rect 877 26544 895 26561
rect 949 26544 983 26578
rect 17 26503 55 26537
rect 109 26504 127 26537
rect 89 26503 127 26504
rect 161 26504 167 26537
rect 233 26504 259 26537
rect 161 26503 199 26504
rect 233 26503 271 26504
rect 305 26503 343 26537
rect 377 26503 415 26537
rect 449 26527 463 26537
rect 521 26527 535 26537
rect 593 26527 607 26537
rect 665 26527 679 26537
rect 737 26527 751 26537
rect 809 26527 823 26537
rect 857 26527 895 26544
rect 929 26527 983 26544
rect 449 26503 487 26527
rect 521 26503 559 26527
rect 593 26503 631 26527
rect 665 26503 703 26527
rect 737 26503 775 26527
rect 809 26509 983 26527
rect 809 26503 843 26509
rect -23 26487 843 26503
rect 877 26487 915 26509
rect -23 26467 463 26487
rect 497 26467 535 26487
rect 569 26467 607 26487
rect 641 26467 679 26487
rect 713 26467 751 26487
rect 785 26467 823 26487
rect 877 26475 895 26487
rect 949 26475 983 26509
rect -23 26431 -17 26467
rect 17 26433 55 26467
rect 89 26465 127 26467
rect 109 26433 127 26465
rect 161 26465 199 26467
rect 233 26465 271 26467
rect 161 26433 167 26465
rect 233 26433 259 26465
rect 305 26433 343 26467
rect 377 26433 415 26467
rect 449 26453 463 26467
rect 521 26453 535 26467
rect 593 26453 607 26467
rect 665 26453 679 26467
rect 737 26453 751 26467
rect 809 26453 823 26467
rect 857 26453 895 26475
rect 929 26453 983 26475
rect 449 26433 487 26453
rect 521 26433 559 26453
rect 593 26433 631 26453
rect 665 26433 703 26453
rect 737 26433 775 26453
rect 809 26440 983 26453
rect 809 26433 843 26440
rect 17 26431 75 26433
rect 109 26431 167 26433
rect 201 26431 259 26433
rect 293 26431 843 26433
rect -23 26413 843 26431
rect 877 26413 915 26440
rect -23 26397 463 26413
rect 497 26397 535 26413
rect 569 26397 607 26413
rect 641 26397 679 26413
rect 713 26397 751 26413
rect 785 26397 823 26413
rect 877 26406 895 26413
rect 949 26406 983 26440
rect -23 26359 -17 26397
rect 17 26363 55 26397
rect 89 26393 127 26397
rect 109 26363 127 26393
rect 161 26393 199 26397
rect 233 26393 271 26397
rect 161 26363 167 26393
rect 233 26363 259 26393
rect 305 26363 343 26397
rect 377 26363 415 26397
rect 449 26379 463 26397
rect 521 26379 535 26397
rect 593 26379 607 26397
rect 665 26379 679 26397
rect 737 26379 751 26397
rect 809 26379 823 26397
rect 857 26379 895 26406
rect 929 26379 983 26406
rect 449 26363 487 26379
rect 521 26363 559 26379
rect 593 26363 631 26379
rect 665 26363 703 26379
rect 737 26363 775 26379
rect 809 26371 983 26379
rect 809 26363 843 26371
rect 17 26359 75 26363
rect 109 26359 167 26363
rect 201 26359 259 26363
rect 293 26359 843 26363
rect -23 26339 843 26359
rect 877 26339 915 26371
rect -23 26327 463 26339
rect 497 26327 535 26339
rect 569 26327 607 26339
rect 641 26327 679 26339
rect 713 26327 751 26339
rect 785 26327 823 26339
rect 877 26337 895 26339
rect 949 26337 983 26371
rect -23 26287 -17 26327
rect 17 26293 55 26327
rect 89 26321 127 26327
rect 109 26293 127 26321
rect 161 26321 199 26327
rect 233 26321 271 26327
rect 161 26293 167 26321
rect 233 26293 259 26321
rect 305 26293 343 26327
rect 377 26293 415 26327
rect 449 26305 463 26327
rect 521 26305 535 26327
rect 593 26305 607 26327
rect 665 26305 679 26327
rect 737 26305 751 26327
rect 809 26305 823 26327
rect 857 26305 895 26337
rect 929 26305 983 26337
rect 449 26293 487 26305
rect 521 26293 559 26305
rect 593 26293 631 26305
rect 665 26293 703 26305
rect 737 26293 775 26305
rect 809 26302 983 26305
rect 809 26293 843 26302
rect 17 26287 75 26293
rect 109 26287 167 26293
rect 201 26287 259 26293
rect 293 26287 843 26293
rect -23 26268 843 26287
rect 877 26268 915 26302
rect 949 26268 983 26302
rect -23 26265 983 26268
rect -23 26257 463 26265
rect 497 26257 535 26265
rect 569 26257 607 26265
rect 641 26257 679 26265
rect 713 26257 751 26265
rect 785 26257 823 26265
rect -23 26255 -17 26257
rect 17 26223 55 26257
rect 89 26223 127 26257
rect 161 26223 199 26257
rect 233 26223 271 26257
rect 305 26223 343 26257
rect 377 26223 415 26257
rect 449 26231 463 26257
rect 521 26231 535 26257
rect 593 26231 607 26257
rect 665 26231 679 26257
rect 737 26231 751 26257
rect 809 26231 823 26257
rect 857 26233 895 26265
rect 929 26233 983 26265
rect 877 26231 895 26233
rect 449 26223 487 26231
rect 521 26223 559 26231
rect 593 26223 631 26231
rect 665 26223 703 26231
rect 737 26223 775 26231
rect 809 26223 843 26231
rect -17 26199 843 26223
rect 877 26199 915 26231
rect 949 26199 983 26233
rect -17 26044 843 26045
rect -23 26021 843 26044
rect -23 25978 -17 26021
rect 17 25987 55 26021
rect 89 26012 127 26021
rect 109 25987 127 26012
rect 161 26012 199 26021
rect 233 26012 271 26021
rect 161 25987 167 26012
rect 233 25987 259 26012
rect 305 25987 343 26021
rect 377 25987 415 26021
rect 449 26012 487 26021
rect 521 26012 559 26021
rect 593 26012 631 26021
rect 665 26012 703 26021
rect 737 26012 775 26021
rect 449 25987 459 26012
rect 521 25987 537 26012
rect 593 25987 615 26012
rect 665 25987 693 26012
rect 737 25987 771 26012
rect 809 26011 843 26021
rect 877 26011 915 26045
rect 949 26011 983 26045
rect 809 25988 983 26011
rect 809 25987 863 25988
rect 17 25978 75 25987
rect 109 25978 167 25987
rect 201 25978 259 25987
rect 293 25978 459 25987
rect 493 25978 537 25987
rect 571 25978 615 25987
rect 649 25978 693 25987
rect 727 25978 771 25987
rect 805 25978 863 25987
rect -23 25972 863 25978
rect 897 25972 983 25988
rect -23 25952 843 25972
rect 897 25954 915 25972
rect -23 25906 -17 25952
rect 17 25918 55 25952
rect 89 25940 127 25952
rect 109 25918 127 25940
rect 161 25940 199 25952
rect 233 25940 271 25952
rect 161 25918 167 25940
rect 233 25918 259 25940
rect 305 25918 343 25952
rect 377 25918 415 25952
rect 449 25940 487 25952
rect 521 25940 559 25952
rect 593 25940 631 25952
rect 665 25940 703 25952
rect 737 25940 775 25952
rect 449 25918 459 25940
rect 521 25918 537 25940
rect 593 25918 615 25940
rect 665 25918 693 25940
rect 737 25918 771 25940
rect 809 25938 843 25952
rect 877 25938 915 25954
rect 949 25938 983 25972
rect 809 25918 983 25938
rect 17 25906 75 25918
rect 109 25906 167 25918
rect 201 25906 259 25918
rect 293 25906 459 25918
rect 493 25906 537 25918
rect 571 25906 615 25918
rect 649 25906 693 25918
rect 727 25906 771 25918
rect 805 25915 983 25918
rect 805 25906 863 25915
rect -23 25899 863 25906
rect 897 25899 983 25915
rect -23 25883 843 25899
rect -23 25834 -17 25883
rect 17 25849 55 25883
rect 89 25868 127 25883
rect 109 25849 127 25868
rect 161 25868 199 25883
rect 233 25868 271 25883
rect 161 25849 167 25868
rect 233 25849 259 25868
rect 305 25849 343 25883
rect 377 25849 415 25883
rect 449 25868 487 25883
rect 521 25868 559 25883
rect 593 25868 631 25883
rect 665 25868 703 25883
rect 737 25868 775 25883
rect 449 25849 459 25868
rect 521 25849 537 25868
rect 593 25849 615 25868
rect 665 25849 693 25868
rect 737 25849 771 25868
rect 809 25865 843 25883
rect 897 25881 915 25899
rect 877 25865 915 25881
rect 949 25865 983 25899
rect 809 25849 983 25865
rect 17 25834 75 25849
rect 109 25834 167 25849
rect 201 25834 259 25849
rect 293 25834 459 25849
rect 493 25834 537 25849
rect 571 25834 615 25849
rect 649 25834 693 25849
rect 727 25834 771 25849
rect 805 25842 983 25849
rect 805 25834 863 25842
rect -23 25826 863 25834
rect 897 25826 983 25842
rect -23 25814 843 25826
rect -23 25762 -17 25814
rect 17 25780 55 25814
rect 89 25796 127 25814
rect 109 25780 127 25796
rect 161 25796 199 25814
rect 233 25796 271 25814
rect 161 25780 167 25796
rect 233 25780 259 25796
rect 305 25780 343 25814
rect 377 25780 415 25814
rect 449 25796 487 25814
rect 521 25796 559 25814
rect 593 25796 631 25814
rect 665 25796 703 25814
rect 737 25796 775 25814
rect 449 25780 459 25796
rect 521 25780 537 25796
rect 593 25780 615 25796
rect 665 25780 693 25796
rect 737 25780 771 25796
rect 809 25792 843 25814
rect 897 25808 915 25826
rect 877 25792 915 25808
rect 949 25792 983 25826
rect 809 25780 983 25792
rect 17 25762 75 25780
rect 109 25762 167 25780
rect 201 25762 259 25780
rect 293 25762 459 25780
rect 493 25762 537 25780
rect 571 25762 615 25780
rect 649 25762 693 25780
rect 727 25762 771 25780
rect 805 25769 983 25780
rect 805 25762 863 25769
rect -23 25753 863 25762
rect 897 25753 983 25769
rect -23 25745 843 25753
rect -23 25690 -17 25745
rect 17 25711 55 25745
rect 89 25724 127 25745
rect 109 25711 127 25724
rect 161 25724 199 25745
rect 233 25724 271 25745
rect 161 25711 167 25724
rect 233 25711 259 25724
rect 305 25711 343 25745
rect 377 25711 415 25745
rect 449 25724 487 25745
rect 521 25724 559 25745
rect 593 25724 631 25745
rect 665 25724 703 25745
rect 737 25724 775 25745
rect 449 25711 459 25724
rect 521 25711 537 25724
rect 593 25711 615 25724
rect 665 25711 693 25724
rect 737 25711 771 25724
rect 809 25719 843 25745
rect 897 25735 915 25753
rect 877 25719 915 25735
rect 949 25719 983 25753
rect 809 25711 983 25719
rect 17 25690 75 25711
rect 109 25690 167 25711
rect 201 25690 259 25711
rect 293 25690 459 25711
rect 493 25690 537 25711
rect 571 25690 615 25711
rect 649 25690 693 25711
rect 727 25690 771 25711
rect 805 25696 983 25711
rect 805 25690 863 25696
rect -23 25680 863 25690
rect 897 25680 983 25696
rect 13833 26021 15917 26023
rect 13867 25987 13906 26021
rect 13940 25987 13979 26021
rect 14013 25987 14052 26021
rect 14086 25987 14125 26021
rect 14159 25987 14198 26021
rect 14232 25987 14271 26021
rect 14305 25987 14344 26021
rect 14378 25987 14417 26021
rect 14451 25987 14490 26021
rect 14524 25987 14563 26021
rect 14597 25987 14636 26021
rect 14670 25987 14709 26021
rect 14743 25987 14782 26021
rect 14816 25987 14855 26021
rect 14889 25987 14928 26021
rect 14962 25987 15001 26021
rect 15035 25987 15074 26021
rect 15108 25987 15147 26021
rect 15181 25987 15220 26021
rect 15254 25987 15293 26021
rect 15327 25987 15366 26021
rect 15400 25987 15439 26021
rect 15473 25987 15513 26021
rect 15547 25987 15587 26021
rect 15621 25987 15661 26021
rect 15695 25987 15735 26021
rect 15769 25987 15809 26021
rect 15843 25987 15883 26021
rect 13833 25947 15917 25987
rect 13867 25913 13906 25947
rect 13940 25913 13979 25947
rect 14013 25913 14052 25947
rect 14086 25913 14125 25947
rect 14159 25913 14198 25947
rect 14232 25913 14271 25947
rect 14305 25913 14344 25947
rect 14378 25913 14417 25947
rect 14451 25913 14490 25947
rect 14524 25913 14563 25947
rect 14597 25913 14636 25947
rect 14670 25913 14709 25947
rect 14743 25913 14782 25947
rect 14816 25913 14855 25947
rect 14889 25913 14928 25947
rect 14962 25913 15001 25947
rect 15035 25913 15074 25947
rect 15108 25913 15147 25947
rect 15181 25913 15220 25947
rect 15254 25913 15293 25947
rect 15327 25913 15366 25947
rect 15400 25913 15439 25947
rect 15473 25913 15513 25947
rect 15547 25913 15587 25947
rect 15621 25913 15661 25947
rect 15695 25913 15735 25947
rect 15769 25913 15809 25947
rect 15843 25913 15883 25947
rect 13833 25873 15917 25913
rect 13867 25839 13906 25873
rect 13940 25839 13979 25873
rect 14013 25839 14052 25873
rect 14086 25839 14125 25873
rect 14159 25839 14198 25873
rect 14232 25839 14271 25873
rect 14305 25839 14344 25873
rect 14378 25839 14417 25873
rect 14451 25839 14490 25873
rect 14524 25839 14563 25873
rect 14597 25839 14636 25873
rect 14670 25839 14709 25873
rect 14743 25839 14782 25873
rect 14816 25839 14855 25873
rect 14889 25839 14928 25873
rect 14962 25839 15001 25873
rect 15035 25839 15074 25873
rect 15108 25839 15147 25873
rect 15181 25839 15220 25873
rect 15254 25839 15293 25873
rect 15327 25839 15366 25873
rect 15400 25839 15439 25873
rect 15473 25839 15513 25873
rect 15547 25839 15587 25873
rect 15621 25839 15661 25873
rect 15695 25839 15735 25873
rect 15769 25839 15809 25873
rect 15843 25839 15883 25873
rect 13833 25799 15917 25839
rect 13867 25765 13906 25799
rect 13940 25765 13979 25799
rect 14013 25765 14052 25799
rect 14086 25765 14125 25799
rect 14159 25765 14198 25799
rect 14232 25765 14271 25799
rect 14305 25765 14344 25799
rect 14378 25765 14417 25799
rect 14451 25765 14490 25799
rect 14524 25765 14563 25799
rect 14597 25765 14636 25799
rect 14670 25765 14709 25799
rect 14743 25765 14782 25799
rect 14816 25765 14855 25799
rect 14889 25765 14928 25799
rect 14962 25765 15001 25799
rect 15035 25765 15074 25799
rect 15108 25765 15147 25799
rect 15181 25765 15220 25799
rect 15254 25765 15293 25799
rect 15327 25765 15366 25799
rect 15400 25765 15439 25799
rect 15473 25765 15513 25799
rect 15547 25765 15587 25799
rect 15621 25765 15661 25799
rect 15695 25765 15735 25799
rect 15769 25765 15809 25799
rect 15843 25765 15883 25799
rect 13833 25725 15917 25765
rect 13867 25691 13906 25725
rect 13940 25691 13979 25725
rect 14013 25691 14052 25725
rect 14086 25691 14125 25725
rect 14159 25691 14198 25725
rect 14232 25691 14271 25725
rect 14305 25691 14344 25725
rect 14378 25691 14417 25725
rect 14451 25691 14490 25725
rect 14524 25691 14563 25725
rect 14597 25691 14636 25725
rect 14670 25691 14709 25725
rect 14743 25691 14782 25725
rect 14816 25691 14855 25725
rect 14889 25691 14928 25725
rect 14962 25691 15001 25725
rect 15035 25691 15074 25725
rect 15108 25691 15147 25725
rect 15181 25691 15220 25725
rect 15254 25691 15293 25725
rect 15327 25691 15366 25725
rect 15400 25691 15439 25725
rect 15473 25691 15513 25725
rect 15547 25691 15587 25725
rect 15621 25691 15661 25725
rect 15695 25691 15735 25725
rect 15769 25691 15809 25725
rect 15843 25691 15883 25725
rect 13833 25689 15917 25691
rect -23 25676 843 25680
rect -23 25618 -17 25676
rect 17 25642 55 25676
rect 89 25652 127 25676
rect 109 25642 127 25652
rect 161 25652 199 25676
rect 233 25652 271 25676
rect 161 25642 167 25652
rect 233 25642 259 25652
rect 305 25642 343 25676
rect 377 25642 415 25676
rect 449 25652 487 25676
rect 521 25652 559 25676
rect 593 25652 631 25676
rect 665 25652 703 25676
rect 737 25652 775 25676
rect 449 25642 459 25652
rect 521 25642 537 25652
rect 593 25642 615 25652
rect 665 25642 693 25652
rect 737 25642 771 25652
rect 809 25646 843 25676
rect 897 25662 915 25680
rect 877 25646 915 25662
rect 949 25646 983 25680
rect 809 25642 983 25646
rect 17 25618 75 25642
rect 109 25618 167 25642
rect 201 25618 259 25642
rect 293 25618 459 25642
rect 493 25618 537 25642
rect 571 25618 615 25642
rect 649 25618 693 25642
rect 727 25618 771 25642
rect 805 25623 983 25642
rect 805 25618 863 25623
rect -23 25607 863 25618
rect 897 25607 983 25623
rect -23 25546 -17 25607
rect 17 25573 55 25607
rect 89 25580 127 25607
rect 109 25573 127 25580
rect 161 25580 199 25607
rect 233 25580 271 25607
rect 161 25573 167 25580
rect 233 25573 259 25580
rect 305 25573 343 25607
rect 377 25573 415 25607
rect 449 25580 487 25607
rect 521 25580 559 25607
rect 593 25580 631 25607
rect 665 25580 703 25607
rect 737 25580 775 25607
rect 449 25573 459 25580
rect 521 25573 537 25580
rect 593 25573 615 25580
rect 665 25573 693 25580
rect 737 25573 771 25580
rect 809 25573 843 25607
rect 897 25589 915 25607
rect 877 25573 915 25589
rect 949 25573 983 25607
rect 17 25546 75 25573
rect 109 25546 167 25573
rect 201 25546 259 25573
rect 293 25546 459 25573
rect 493 25546 537 25573
rect 571 25546 615 25573
rect 649 25546 693 25573
rect 727 25546 771 25573
rect 805 25550 983 25573
rect 805 25546 863 25550
rect -23 25539 863 25546
rect -23 25474 -17 25539
rect 17 25505 55 25539
rect 89 25508 127 25539
rect 109 25505 127 25508
rect 161 25508 199 25539
rect 233 25508 271 25539
rect 161 25505 167 25508
rect 233 25505 259 25508
rect 305 25505 343 25539
rect 377 25505 415 25539
rect 449 25508 487 25539
rect 521 25508 559 25539
rect 593 25508 631 25539
rect 665 25508 703 25539
rect 737 25508 775 25539
rect 809 25534 863 25539
rect 897 25534 983 25550
rect 449 25505 459 25508
rect 521 25505 537 25508
rect 593 25505 615 25508
rect 665 25505 693 25508
rect 737 25505 771 25508
rect 809 25505 843 25534
rect 897 25516 915 25534
rect 17 25474 75 25505
rect 109 25474 167 25505
rect 201 25474 259 25505
rect 293 25474 459 25505
rect 493 25474 537 25505
rect 571 25474 615 25505
rect 649 25474 693 25505
rect 727 25474 771 25505
rect 805 25500 843 25505
rect 877 25500 915 25516
rect 949 25500 983 25534
rect 805 25476 983 25500
rect 805 25474 863 25476
rect -23 25471 863 25474
rect -23 25437 -17 25471
rect 17 25437 55 25471
rect 89 25437 127 25471
rect 161 25437 199 25471
rect 233 25437 271 25471
rect 305 25437 343 25471
rect 377 25437 415 25471
rect 449 25437 487 25471
rect 521 25437 559 25471
rect 593 25437 631 25471
rect 665 25437 703 25471
rect 737 25437 775 25471
rect 809 25461 863 25471
rect 897 25461 983 25476
rect 809 25437 843 25461
rect 897 25442 915 25461
rect -23 25436 843 25437
rect -23 25369 -17 25436
rect 17 25403 75 25436
rect 109 25403 167 25436
rect 201 25403 259 25436
rect 293 25403 459 25436
rect 493 25403 537 25436
rect 571 25403 615 25436
rect 649 25403 693 25436
rect 727 25403 771 25436
rect 805 25427 843 25436
rect 877 25427 915 25442
rect 949 25427 983 25461
rect 805 25403 983 25427
rect 17 25369 55 25403
rect 109 25402 127 25403
rect 89 25369 127 25402
rect 161 25402 167 25403
rect 233 25402 259 25403
rect 161 25369 199 25402
rect 233 25369 271 25402
rect 305 25369 343 25403
rect 377 25369 415 25403
rect 449 25402 459 25403
rect 521 25402 537 25403
rect 593 25402 615 25403
rect 665 25402 693 25403
rect 737 25402 771 25403
rect 809 25402 983 25403
rect 449 25369 487 25402
rect 521 25369 559 25402
rect 593 25369 631 25402
rect 665 25369 703 25402
rect 737 25369 775 25402
rect 809 25388 863 25402
rect 897 25388 983 25402
rect 809 25369 843 25388
rect -23 25364 843 25369
rect 897 25368 915 25388
rect -23 25301 -17 25364
rect 17 25335 75 25364
rect 109 25335 167 25364
rect 201 25335 259 25364
rect 293 25335 459 25364
rect 493 25335 537 25364
rect 571 25335 615 25364
rect 649 25335 693 25364
rect 727 25335 771 25364
rect 805 25354 843 25364
rect 877 25354 915 25368
rect 949 25354 983 25388
rect 805 25335 983 25354
rect 17 25301 55 25335
rect 109 25330 127 25335
rect 89 25301 127 25330
rect 161 25330 167 25335
rect 233 25330 259 25335
rect 161 25301 199 25330
rect 233 25301 271 25330
rect 305 25301 343 25335
rect 377 25301 415 25335
rect 449 25330 459 25335
rect 521 25330 537 25335
rect 593 25330 615 25335
rect 665 25330 693 25335
rect 737 25330 771 25335
rect 449 25301 487 25330
rect 521 25301 559 25330
rect 593 25301 631 25330
rect 665 25301 703 25330
rect 737 25301 775 25330
rect 809 25328 983 25335
rect 809 25316 863 25328
rect 897 25316 983 25328
rect 809 25301 843 25316
rect -23 25292 843 25301
rect 897 25294 915 25316
rect -23 25233 -17 25292
rect 17 25267 75 25292
rect 109 25267 167 25292
rect 201 25267 259 25292
rect 293 25267 459 25292
rect 493 25267 537 25292
rect 571 25267 615 25292
rect 649 25267 693 25292
rect 727 25267 771 25292
rect 805 25282 843 25292
rect 877 25282 915 25294
rect 949 25282 983 25316
rect 805 25267 983 25282
rect 17 25233 55 25267
rect 109 25258 127 25267
rect 89 25233 127 25258
rect 161 25258 167 25267
rect 233 25258 259 25267
rect 161 25233 199 25258
rect 233 25233 271 25258
rect 305 25233 343 25267
rect 377 25233 415 25267
rect 449 25258 459 25267
rect 521 25258 537 25267
rect 593 25258 615 25267
rect 665 25258 693 25267
rect 737 25258 771 25267
rect 449 25233 487 25258
rect 521 25233 559 25258
rect 593 25233 631 25258
rect 665 25233 703 25258
rect 737 25233 775 25258
rect 809 25233 983 25267
rect -23 25220 983 25233
rect -23 25165 -17 25220
rect 17 25199 75 25220
rect 109 25199 167 25220
rect 201 25199 259 25220
rect 293 25199 459 25220
rect 493 25199 537 25220
rect 571 25199 615 25220
rect 649 25199 693 25220
rect 727 25199 771 25220
rect 805 25199 983 25220
rect 17 25165 55 25199
rect 109 25186 127 25199
rect 89 25165 127 25186
rect 161 25186 167 25199
rect 233 25186 259 25199
rect 161 25165 199 25186
rect 233 25165 271 25186
rect 305 25165 343 25199
rect 377 25165 415 25199
rect 449 25186 459 25199
rect 521 25186 537 25199
rect 593 25186 615 25199
rect 665 25186 693 25199
rect 737 25186 771 25199
rect 449 25165 487 25186
rect 521 25165 559 25186
rect 593 25165 631 25186
rect 665 25165 703 25186
rect 737 25165 775 25186
rect 809 25165 983 25199
rect -23 25148 983 25165
rect -23 25097 -17 25148
rect 17 25131 75 25148
rect 109 25131 167 25148
rect 201 25131 259 25148
rect 293 25131 459 25148
rect 493 25131 537 25148
rect 571 25131 615 25148
rect 649 25131 693 25148
rect 727 25131 771 25148
rect 805 25131 983 25148
rect 17 25097 55 25131
rect 109 25114 127 25131
rect 89 25097 127 25114
rect 161 25114 167 25131
rect 233 25114 259 25131
rect 161 25097 199 25114
rect 233 25097 271 25114
rect 305 25097 343 25131
rect 377 25097 415 25131
rect 449 25114 459 25131
rect 521 25114 537 25131
rect 593 25114 615 25131
rect 665 25114 693 25131
rect 737 25114 771 25131
rect 449 25097 487 25114
rect 521 25097 559 25114
rect 593 25097 631 25114
rect 665 25097 703 25114
rect 737 25097 775 25114
rect 809 25097 983 25131
rect -23 25076 983 25097
rect -23 25029 -17 25076
rect 17 25063 75 25076
rect 109 25063 167 25076
rect 201 25063 259 25076
rect 293 25063 459 25076
rect 493 25063 537 25076
rect 571 25063 615 25076
rect 649 25063 693 25076
rect 727 25063 771 25076
rect 805 25063 983 25076
rect 17 25029 55 25063
rect 109 25042 127 25063
rect 89 25029 127 25042
rect 161 25042 167 25063
rect 233 25042 259 25063
rect 161 25029 199 25042
rect 233 25029 271 25042
rect 305 25029 343 25063
rect 377 25029 415 25063
rect 449 25042 459 25063
rect 521 25042 537 25063
rect 593 25042 615 25063
rect 665 25042 693 25063
rect 737 25042 771 25063
rect 449 25029 487 25042
rect 521 25029 559 25042
rect 593 25029 631 25042
rect 665 25029 703 25042
rect 737 25029 775 25042
rect 809 25029 983 25063
rect -23 25004 983 25029
rect -23 24961 -17 25004
rect 17 24995 75 25004
rect 109 24995 167 25004
rect 201 24995 259 25004
rect 293 24995 459 25004
rect 493 24995 537 25004
rect 571 24995 615 25004
rect 649 24995 693 25004
rect 727 24995 771 25004
rect 805 24995 983 25004
rect 17 24961 55 24995
rect 109 24970 127 24995
rect 89 24961 127 24970
rect 161 24970 167 24995
rect 233 24970 259 24995
rect 161 24961 199 24970
rect 233 24961 271 24970
rect 305 24961 343 24995
rect 377 24961 415 24995
rect 449 24970 459 24995
rect 521 24970 537 24995
rect 593 24970 615 24995
rect 665 24970 693 24995
rect 737 24970 771 24995
rect 449 24961 487 24970
rect 521 24961 559 24970
rect 593 24961 631 24970
rect 665 24961 703 24970
rect 737 24961 775 24970
rect 809 24961 983 24995
rect -23 24932 983 24961
rect -23 24893 -17 24932
rect 17 24927 75 24932
rect 109 24927 167 24932
rect 201 24927 259 24932
rect 293 24927 459 24932
rect 493 24927 537 24932
rect 571 24927 615 24932
rect 649 24927 693 24932
rect 727 24927 771 24932
rect 805 24927 983 24932
rect 17 24893 55 24927
rect 109 24898 127 24927
rect 89 24893 127 24898
rect 161 24898 167 24927
rect 233 24898 259 24927
rect 161 24893 199 24898
rect 233 24893 271 24898
rect 305 24893 343 24927
rect 377 24893 415 24927
rect 449 24898 459 24927
rect 521 24898 537 24927
rect 593 24898 615 24927
rect 665 24898 693 24927
rect 737 24898 771 24927
rect 449 24893 487 24898
rect 521 24893 559 24898
rect 593 24893 631 24898
rect 665 24893 703 24898
rect 737 24893 775 24898
rect 809 24893 983 24927
rect -23 24860 983 24893
rect -23 24825 -17 24860
rect 17 24859 75 24860
rect 109 24859 167 24860
rect 201 24859 259 24860
rect 293 24859 459 24860
rect 493 24859 537 24860
rect 571 24859 615 24860
rect 649 24859 693 24860
rect 727 24859 771 24860
rect 805 24859 983 24860
rect 17 24825 55 24859
rect 109 24826 127 24859
rect 89 24825 127 24826
rect 161 24826 167 24859
rect 233 24826 259 24859
rect 161 24825 199 24826
rect 233 24825 271 24826
rect 305 24825 343 24859
rect 377 24825 415 24859
rect 449 24826 459 24859
rect 521 24826 537 24859
rect 593 24826 615 24859
rect 665 24826 693 24859
rect 737 24826 771 24859
rect 449 24825 487 24826
rect 521 24825 559 24826
rect 593 24825 631 24826
rect 665 24825 703 24826
rect 737 24825 775 24826
rect 809 24825 983 24859
rect -23 24791 983 24825
rect -23 24754 -17 24791
rect 17 24757 55 24791
rect 89 24788 127 24791
rect 109 24757 127 24788
rect 161 24788 199 24791
rect 233 24788 271 24791
rect 161 24757 167 24788
rect 233 24757 259 24788
rect 305 24757 343 24791
rect 377 24757 415 24791
rect 449 24788 487 24791
rect 521 24788 559 24791
rect 593 24788 631 24791
rect 665 24788 703 24791
rect 737 24788 775 24791
rect 449 24757 459 24788
rect 521 24757 537 24788
rect 593 24757 615 24788
rect 665 24757 693 24788
rect 737 24757 771 24788
rect 809 24757 983 24791
rect 17 24754 75 24757
rect 109 24754 167 24757
rect 201 24754 259 24757
rect 293 24754 459 24757
rect 493 24754 537 24757
rect 571 24754 615 24757
rect 649 24754 693 24757
rect 727 24754 771 24757
rect 805 24754 983 24757
rect -23 24723 983 24754
rect -23 24682 -17 24723
rect 17 24689 55 24723
rect 89 24716 127 24723
rect 109 24689 127 24716
rect 161 24716 199 24723
rect 233 24716 271 24723
rect 161 24689 167 24716
rect 233 24689 259 24716
rect 305 24689 343 24723
rect 377 24689 415 24723
rect 449 24716 487 24723
rect 521 24716 559 24723
rect 593 24716 631 24723
rect 665 24716 703 24723
rect 737 24716 775 24723
rect 449 24689 459 24716
rect 521 24689 537 24716
rect 593 24689 615 24716
rect 665 24689 693 24716
rect 737 24689 771 24716
rect 809 24689 983 24723
rect 17 24682 75 24689
rect 109 24682 167 24689
rect 201 24682 259 24689
rect 293 24682 459 24689
rect 493 24682 537 24689
rect 571 24682 615 24689
rect 649 24682 693 24689
rect 727 24682 771 24689
rect 805 24682 983 24689
rect -23 24655 983 24682
rect -23 24610 -17 24655
rect 17 24621 55 24655
rect 89 24644 127 24655
rect 109 24621 127 24644
rect 161 24644 199 24655
rect 233 24644 271 24655
rect 161 24621 167 24644
rect 233 24621 259 24644
rect 305 24621 343 24655
rect 377 24621 415 24655
rect 449 24644 487 24655
rect 521 24644 559 24655
rect 593 24644 631 24655
rect 665 24644 703 24655
rect 737 24644 775 24655
rect 449 24621 459 24644
rect 521 24621 537 24644
rect 593 24621 615 24644
rect 665 24621 693 24644
rect 737 24621 771 24644
rect 809 24621 983 24655
rect 17 24610 75 24621
rect 109 24610 167 24621
rect 201 24610 259 24621
rect 293 24610 459 24621
rect 493 24610 537 24621
rect 571 24610 615 24621
rect 649 24610 693 24621
rect 727 24610 771 24621
rect 805 24610 983 24621
rect -23 24587 983 24610
rect -23 24538 -17 24587
rect 17 24553 55 24587
rect 89 24572 127 24587
rect 109 24553 127 24572
rect 161 24572 199 24587
rect 233 24572 271 24587
rect 161 24553 167 24572
rect 233 24553 259 24572
rect 305 24553 343 24587
rect 377 24553 415 24587
rect 449 24572 487 24587
rect 521 24572 559 24587
rect 593 24572 631 24587
rect 665 24572 703 24587
rect 737 24572 775 24587
rect 449 24553 459 24572
rect 521 24553 537 24572
rect 593 24553 615 24572
rect 665 24553 693 24572
rect 737 24553 771 24572
rect 809 24553 983 24587
rect 17 24538 75 24553
rect 109 24538 167 24553
rect 201 24538 259 24553
rect 293 24538 459 24553
rect 493 24538 537 24553
rect 571 24538 615 24553
rect 649 24538 693 24553
rect 727 24538 771 24553
rect 805 24538 983 24553
rect -23 24519 983 24538
rect -23 24466 -17 24519
rect 17 24485 55 24519
rect 89 24500 127 24519
rect 109 24485 127 24500
rect 161 24500 199 24519
rect 233 24500 271 24519
rect 161 24485 167 24500
rect 233 24485 259 24500
rect 305 24485 343 24519
rect 377 24485 415 24519
rect 449 24500 487 24519
rect 521 24500 559 24519
rect 593 24500 631 24519
rect 665 24500 703 24519
rect 737 24500 775 24519
rect 449 24485 459 24500
rect 521 24485 537 24500
rect 593 24485 615 24500
rect 665 24485 693 24500
rect 737 24485 771 24500
rect 809 24485 983 24519
rect 17 24466 75 24485
rect 109 24466 167 24485
rect 201 24466 259 24485
rect 293 24466 459 24485
rect 493 24466 537 24485
rect 571 24466 615 24485
rect 649 24466 693 24485
rect 727 24466 771 24485
rect 805 24466 983 24485
rect -23 24451 983 24466
rect -23 24394 -17 24451
rect 17 24417 55 24451
rect 89 24428 127 24451
rect 109 24417 127 24428
rect 161 24428 199 24451
rect 233 24428 271 24451
rect 161 24417 167 24428
rect 233 24417 259 24428
rect 305 24417 343 24451
rect 377 24417 415 24451
rect 449 24428 487 24451
rect 521 24428 559 24451
rect 593 24428 631 24451
rect 665 24428 703 24451
rect 737 24428 775 24451
rect 449 24417 459 24428
rect 521 24417 537 24428
rect 593 24417 615 24428
rect 665 24417 693 24428
rect 737 24417 771 24428
rect 809 24417 983 24451
rect 17 24394 75 24417
rect 109 24394 167 24417
rect 201 24394 259 24417
rect 293 24394 459 24417
rect 493 24394 537 24417
rect 571 24394 615 24417
rect 649 24394 693 24417
rect 727 24394 771 24417
rect 805 24394 983 24417
rect -23 24383 983 24394
rect -23 24321 -17 24383
rect 17 24349 55 24383
rect 89 24355 127 24383
rect 109 24349 127 24355
rect 161 24355 199 24383
rect 233 24355 271 24383
rect 161 24349 167 24355
rect 233 24349 259 24355
rect 305 24349 343 24383
rect 377 24349 415 24383
rect 449 24355 487 24383
rect 521 24355 559 24383
rect 593 24355 631 24383
rect 665 24355 703 24383
rect 737 24355 775 24383
rect 449 24349 459 24355
rect 521 24349 537 24355
rect 593 24349 615 24355
rect 665 24349 693 24355
rect 737 24349 771 24355
rect 809 24349 983 24383
rect 17 24321 75 24349
rect 109 24321 167 24349
rect 201 24321 259 24349
rect 293 24321 459 24349
rect 493 24321 537 24349
rect 571 24321 615 24349
rect 649 24321 693 24349
rect 727 24321 771 24349
rect 805 24321 983 24349
rect -23 24315 983 24321
rect -23 24248 -17 24315
rect 17 24281 55 24315
rect 89 24282 127 24315
rect 109 24281 127 24282
rect 161 24282 199 24315
rect 233 24282 271 24315
rect 161 24281 167 24282
rect 233 24281 259 24282
rect 305 24281 343 24315
rect 377 24281 415 24315
rect 449 24282 487 24315
rect 521 24282 559 24315
rect 593 24282 631 24315
rect 665 24282 703 24315
rect 737 24282 775 24315
rect 449 24281 459 24282
rect 521 24281 537 24282
rect 593 24281 615 24282
rect 665 24281 693 24282
rect 737 24281 771 24282
rect 809 24281 983 24315
rect 17 24248 75 24281
rect 109 24248 167 24281
rect 201 24248 259 24281
rect 293 24248 459 24281
rect 493 24248 537 24281
rect 571 24248 615 24281
rect 649 24248 693 24281
rect 727 24248 771 24281
rect 805 24248 983 24281
rect -23 24247 983 24248
rect -23 24213 -17 24247
rect 17 24213 55 24247
rect 89 24213 127 24247
rect 161 24213 199 24247
rect 233 24213 271 24247
rect 305 24213 343 24247
rect 377 24213 415 24247
rect 449 24213 487 24247
rect 521 24213 559 24247
rect 593 24213 631 24247
rect 665 24213 703 24247
rect 737 24213 775 24247
rect 809 24213 983 24247
rect -23 24209 983 24213
rect -23 24145 -17 24209
rect 17 24179 75 24209
rect 109 24179 167 24209
rect 201 24179 259 24209
rect 293 24179 459 24209
rect 493 24179 537 24209
rect 571 24179 615 24209
rect 649 24179 693 24209
rect 727 24179 771 24209
rect 805 24179 983 24209
rect 17 24145 55 24179
rect 109 24175 127 24179
rect 89 24145 127 24175
rect 161 24175 167 24179
rect 233 24175 259 24179
rect 161 24145 199 24175
rect 233 24145 271 24175
rect 305 24145 343 24179
rect 377 24145 415 24179
rect 449 24175 459 24179
rect 521 24175 537 24179
rect 593 24175 615 24179
rect 665 24175 693 24179
rect 737 24175 771 24179
rect 449 24145 487 24175
rect 521 24145 559 24175
rect 593 24145 631 24175
rect 665 24145 703 24175
rect 737 24145 775 24175
rect 809 24145 983 24179
rect -23 24136 983 24145
rect -23 24077 -17 24136
rect 17 24111 75 24136
rect 109 24111 167 24136
rect 201 24111 259 24136
rect 293 24111 459 24136
rect 493 24111 537 24136
rect 571 24111 615 24136
rect 649 24111 693 24136
rect 727 24111 771 24136
rect 805 24111 983 24136
rect 17 24077 55 24111
rect 109 24102 127 24111
rect 89 24077 127 24102
rect 161 24102 167 24111
rect 233 24102 259 24111
rect 161 24077 199 24102
rect 233 24077 271 24102
rect 305 24077 343 24111
rect 377 24077 415 24111
rect 449 24102 459 24111
rect 521 24102 537 24111
rect 593 24102 615 24111
rect 665 24102 693 24111
rect 737 24102 771 24111
rect 449 24077 487 24102
rect 521 24077 559 24102
rect 593 24077 631 24102
rect 665 24077 703 24102
rect 737 24077 775 24102
rect 809 24077 983 24111
rect -23 24063 983 24077
rect -23 24009 -17 24063
rect 17 24043 75 24063
rect 109 24043 167 24063
rect 201 24043 259 24063
rect 293 24043 459 24063
rect 493 24043 537 24063
rect 571 24043 615 24063
rect 649 24043 693 24063
rect 727 24043 771 24063
rect 805 24043 983 24063
rect 17 24009 55 24043
rect 109 24029 127 24043
rect 89 24009 127 24029
rect 161 24029 167 24043
rect 233 24029 259 24043
rect 161 24009 199 24029
rect 233 24009 271 24029
rect 305 24009 343 24043
rect 377 24009 415 24043
rect 449 24029 459 24043
rect 521 24029 537 24043
rect 593 24029 615 24043
rect 665 24029 693 24043
rect 737 24029 771 24043
rect 449 24009 487 24029
rect 521 24009 559 24029
rect 593 24009 631 24029
rect 665 24009 703 24029
rect 737 24009 775 24029
rect 809 24009 983 24043
rect -23 23990 983 24009
rect -23 23941 -17 23990
rect 17 23975 75 23990
rect 109 23975 167 23990
rect 201 23975 259 23990
rect 293 23975 459 23990
rect 493 23975 537 23990
rect 571 23975 615 23990
rect 649 23975 693 23990
rect 727 23975 771 23990
rect 805 23975 983 23990
rect 17 23941 55 23975
rect 109 23956 127 23975
rect 89 23941 127 23956
rect 161 23956 167 23975
rect 233 23956 259 23975
rect 161 23941 199 23956
rect 233 23941 271 23956
rect 305 23941 343 23975
rect 377 23941 415 23975
rect 449 23956 459 23975
rect 521 23956 537 23975
rect 593 23956 615 23975
rect 665 23956 693 23975
rect 737 23956 771 23975
rect 449 23941 487 23956
rect 521 23941 559 23956
rect 593 23941 631 23956
rect 665 23941 703 23956
rect 737 23941 775 23956
rect 809 23941 983 23975
rect -23 23917 983 23941
rect -23 23873 -17 23917
rect 17 23907 75 23917
rect 109 23907 167 23917
rect 201 23907 259 23917
rect 293 23907 459 23917
rect 493 23907 537 23917
rect 571 23907 615 23917
rect 649 23907 693 23917
rect 727 23907 771 23917
rect 805 23907 983 23917
rect 17 23873 55 23907
rect 109 23883 127 23907
rect 89 23873 127 23883
rect 161 23883 167 23907
rect 233 23883 259 23907
rect 161 23873 199 23883
rect 233 23873 271 23883
rect 305 23873 343 23907
rect 377 23873 415 23907
rect 449 23883 459 23907
rect 521 23883 537 23907
rect 593 23883 615 23907
rect 665 23883 693 23907
rect 737 23883 771 23907
rect 449 23873 487 23883
rect 521 23873 559 23883
rect 593 23873 631 23883
rect 665 23873 703 23883
rect 737 23873 775 23883
rect 809 23873 983 23907
rect -23 23844 983 23873
rect -23 23805 -17 23844
rect 17 23839 75 23844
rect 109 23839 167 23844
rect 201 23839 259 23844
rect 293 23839 459 23844
rect 493 23839 537 23844
rect 571 23839 615 23844
rect 649 23839 693 23844
rect 727 23839 771 23844
rect 805 23839 983 23844
rect 17 23805 55 23839
rect 109 23810 127 23839
rect 89 23805 127 23810
rect 161 23810 167 23839
rect 233 23810 259 23839
rect 161 23805 199 23810
rect 233 23805 271 23810
rect 305 23805 343 23839
rect 377 23805 415 23839
rect 449 23810 459 23839
rect 521 23810 537 23839
rect 593 23810 615 23839
rect 665 23810 693 23839
rect 737 23810 771 23839
rect 449 23805 487 23810
rect 521 23805 559 23810
rect 593 23805 631 23810
rect 665 23805 703 23810
rect 737 23805 775 23810
rect 809 23805 983 23839
rect -23 23771 983 23805
rect -23 23737 -17 23771
rect 17 23737 55 23771
rect 109 23737 127 23771
rect 161 23737 167 23771
rect 233 23737 259 23771
rect 305 23737 343 23771
rect 377 23737 415 23771
rect 449 23737 459 23771
rect 521 23737 537 23771
rect 593 23737 615 23771
rect 665 23737 693 23771
rect 737 23737 771 23771
rect 809 23737 983 23771
rect -23 23703 983 23737
rect -23 23664 -17 23703
rect 17 23669 55 23703
rect 89 23698 127 23703
rect 109 23669 127 23698
rect 161 23698 199 23703
rect 233 23698 271 23703
rect 161 23669 167 23698
rect 233 23669 259 23698
rect 305 23669 343 23703
rect 377 23669 415 23703
rect 449 23698 487 23703
rect 521 23698 559 23703
rect 593 23698 631 23703
rect 665 23698 703 23703
rect 737 23698 775 23703
rect 449 23669 459 23698
rect 521 23669 537 23698
rect 593 23669 615 23698
rect 665 23669 693 23698
rect 737 23669 771 23698
rect 809 23669 983 23703
rect 17 23664 75 23669
rect 109 23664 167 23669
rect 201 23664 259 23669
rect 293 23664 459 23669
rect 493 23664 537 23669
rect 571 23664 615 23669
rect 649 23664 693 23669
rect 727 23664 771 23669
rect 805 23664 983 23669
rect -23 23635 983 23664
rect -23 23591 -17 23635
rect 17 23601 55 23635
rect 89 23625 127 23635
rect 109 23601 127 23625
rect 161 23625 199 23635
rect 233 23625 271 23635
rect 161 23601 167 23625
rect 233 23601 259 23625
rect 305 23601 343 23635
rect 377 23601 415 23635
rect 449 23625 487 23635
rect 521 23625 559 23635
rect 593 23625 631 23635
rect 665 23625 703 23635
rect 737 23625 775 23635
rect 449 23601 459 23625
rect 521 23601 537 23625
rect 593 23601 615 23625
rect 665 23601 693 23625
rect 737 23601 771 23625
rect 809 23601 983 23635
rect 17 23591 75 23601
rect 109 23591 167 23601
rect 201 23591 259 23601
rect 293 23591 459 23601
rect 493 23591 537 23601
rect 571 23591 615 23601
rect 649 23591 693 23601
rect 727 23591 771 23601
rect 805 23591 983 23601
rect -23 23567 983 23591
rect -23 23518 -17 23567
rect 17 23533 55 23567
rect 89 23552 127 23567
rect 109 23533 127 23552
rect 161 23552 199 23567
rect 233 23552 271 23567
rect 161 23533 167 23552
rect 233 23533 259 23552
rect 305 23533 343 23567
rect 377 23533 415 23567
rect 449 23552 487 23567
rect 521 23552 559 23567
rect 593 23552 631 23567
rect 665 23552 703 23567
rect 737 23552 775 23567
rect 449 23533 459 23552
rect 521 23533 537 23552
rect 593 23533 615 23552
rect 665 23533 693 23552
rect 737 23533 771 23552
rect 809 23533 983 23567
rect 17 23518 75 23533
rect 109 23518 167 23533
rect 201 23518 259 23533
rect 293 23518 459 23533
rect 493 23518 537 23533
rect 571 23518 615 23533
rect 649 23518 693 23533
rect 727 23518 771 23533
rect 805 23518 983 23533
rect -23 23499 983 23518
rect -23 23445 -17 23499
rect 17 23465 55 23499
rect 89 23479 127 23499
rect 109 23465 127 23479
rect 161 23479 199 23499
rect 233 23479 271 23499
rect 161 23465 167 23479
rect 233 23465 259 23479
rect 305 23465 343 23499
rect 377 23465 415 23499
rect 449 23479 487 23499
rect 521 23479 559 23499
rect 593 23479 631 23499
rect 665 23479 703 23499
rect 737 23479 775 23499
rect 449 23465 459 23479
rect 521 23465 537 23479
rect 593 23465 615 23479
rect 665 23465 693 23479
rect 737 23465 771 23479
rect 809 23465 983 23499
rect 17 23445 75 23465
rect 109 23445 167 23465
rect 201 23445 259 23465
rect 293 23445 459 23465
rect 493 23445 537 23465
rect 571 23445 615 23465
rect 649 23445 693 23465
rect 727 23445 771 23465
rect 805 23445 983 23465
rect -23 23431 983 23445
rect -23 23372 -17 23431
rect 17 23397 55 23431
rect 89 23406 127 23431
rect 109 23397 127 23406
rect 161 23406 199 23431
rect 233 23406 271 23431
rect 161 23397 167 23406
rect 233 23397 259 23406
rect 305 23397 343 23431
rect 377 23397 415 23431
rect 449 23406 487 23431
rect 521 23406 559 23431
rect 593 23406 631 23431
rect 665 23406 703 23431
rect 737 23406 775 23431
rect 449 23397 459 23406
rect 521 23397 537 23406
rect 593 23397 615 23406
rect 665 23397 693 23406
rect 737 23397 771 23406
rect 809 23397 983 23431
rect 17 23372 75 23397
rect 109 23372 167 23397
rect 201 23372 259 23397
rect 293 23372 459 23397
rect 493 23372 537 23397
rect 571 23372 615 23397
rect 649 23372 693 23397
rect 727 23372 771 23397
rect 805 23372 983 23397
rect -23 23363 983 23372
rect -23 23299 -17 23363
rect 17 23329 55 23363
rect 89 23333 127 23363
rect 109 23329 127 23333
rect 161 23333 199 23363
rect 233 23333 271 23363
rect 161 23329 167 23333
rect 233 23329 259 23333
rect 305 23329 343 23363
rect 377 23329 415 23363
rect 449 23333 487 23363
rect 521 23333 559 23363
rect 593 23333 631 23363
rect 665 23333 703 23363
rect 737 23333 775 23363
rect 449 23329 459 23333
rect 521 23329 537 23333
rect 593 23329 615 23333
rect 665 23329 693 23333
rect 737 23329 771 23333
rect 809 23329 983 23363
rect 17 23299 75 23329
rect 109 23299 167 23329
rect 201 23299 259 23329
rect 293 23299 459 23329
rect 493 23299 537 23329
rect 571 23299 615 23329
rect 649 23299 693 23329
rect 727 23299 771 23329
rect 805 23299 983 23329
rect -23 23295 983 23299
rect -23 23261 -17 23295
rect 17 23261 55 23295
rect 89 23261 127 23295
rect 161 23261 199 23295
rect 233 23261 271 23295
rect 305 23261 343 23295
rect 377 23261 415 23295
rect 449 23261 487 23295
rect 521 23261 559 23295
rect 593 23261 631 23295
rect 665 23261 703 23295
rect 737 23261 775 23295
rect 809 23261 983 23295
rect -23 23260 983 23261
rect -23 23193 -17 23260
rect 17 23227 75 23260
rect 109 23227 167 23260
rect 201 23227 259 23260
rect 293 23227 459 23260
rect 493 23227 537 23260
rect 571 23227 615 23260
rect 649 23227 693 23260
rect 727 23227 771 23260
rect 805 23227 983 23260
rect 17 23193 55 23227
rect 109 23226 127 23227
rect 89 23193 127 23226
rect 161 23226 167 23227
rect 233 23226 259 23227
rect 161 23193 199 23226
rect 233 23193 271 23226
rect 305 23193 343 23227
rect 377 23193 415 23227
rect 449 23226 459 23227
rect 521 23226 537 23227
rect 593 23226 615 23227
rect 665 23226 693 23227
rect 737 23226 771 23227
rect 449 23193 487 23226
rect 521 23193 559 23226
rect 593 23193 631 23226
rect 665 23193 703 23226
rect 737 23193 775 23226
rect 809 23193 983 23227
rect -23 23187 983 23193
rect -23 23125 -17 23187
rect 17 23159 75 23187
rect 109 23159 167 23187
rect 201 23159 259 23187
rect 293 23159 459 23187
rect 493 23159 537 23187
rect 571 23159 615 23187
rect 649 23159 693 23187
rect 727 23159 771 23187
rect 805 23159 983 23187
rect 17 23125 55 23159
rect 109 23153 127 23159
rect 89 23125 127 23153
rect 161 23153 167 23159
rect 233 23153 259 23159
rect 161 23125 199 23153
rect 233 23125 271 23153
rect 305 23125 343 23159
rect 377 23125 415 23159
rect 449 23153 459 23159
rect 521 23153 537 23159
rect 593 23153 615 23159
rect 665 23153 693 23159
rect 737 23153 771 23159
rect 449 23125 487 23153
rect 521 23125 559 23153
rect 593 23125 631 23153
rect 665 23125 703 23153
rect 737 23125 775 23153
rect 809 23125 983 23159
rect -23 23114 983 23125
rect -23 23057 -17 23114
rect 17 23091 75 23114
rect 109 23091 167 23114
rect 201 23091 259 23114
rect 293 23091 459 23114
rect 493 23091 537 23114
rect 571 23091 615 23114
rect 649 23091 693 23114
rect 727 23091 771 23114
rect 805 23091 983 23114
rect 17 23057 55 23091
rect 109 23080 127 23091
rect 89 23057 127 23080
rect 161 23080 167 23091
rect 233 23080 259 23091
rect 161 23057 199 23080
rect 233 23057 271 23080
rect 305 23057 343 23091
rect 377 23057 415 23091
rect 449 23080 459 23091
rect 521 23080 537 23091
rect 593 23080 615 23091
rect 665 23080 693 23091
rect 737 23080 771 23091
rect 449 23057 487 23080
rect 521 23057 559 23080
rect 593 23057 631 23080
rect 665 23057 703 23080
rect 737 23057 775 23080
rect 809 23057 983 23091
rect -23 23041 983 23057
rect -23 22989 -17 23041
rect 17 23023 75 23041
rect 109 23023 167 23041
rect 201 23023 259 23041
rect 293 23023 459 23041
rect 493 23023 537 23041
rect 571 23023 615 23041
rect 649 23023 693 23041
rect 727 23023 771 23041
rect 805 23023 983 23041
rect 17 22989 55 23023
rect 109 23007 127 23023
rect 89 22989 127 23007
rect 161 23007 167 23023
rect 233 23007 259 23023
rect 161 22989 199 23007
rect 233 22989 271 23007
rect 305 22989 343 23023
rect 377 22989 415 23023
rect 449 23007 459 23023
rect 521 23007 537 23023
rect 593 23007 615 23023
rect 665 23007 693 23023
rect 737 23007 771 23023
rect 449 22989 487 23007
rect 521 22989 559 23007
rect 593 22989 631 23007
rect 665 22989 703 23007
rect 737 22989 775 23007
rect 809 22989 983 23023
rect -23 22968 983 22989
rect -23 22921 -17 22968
rect 17 22955 75 22968
rect 109 22955 167 22968
rect 201 22955 259 22968
rect 293 22955 459 22968
rect 493 22955 537 22968
rect 571 22955 615 22968
rect 649 22955 693 22968
rect 727 22955 771 22968
rect 805 22955 983 22968
rect 17 22921 55 22955
rect 109 22934 127 22955
rect 89 22921 127 22934
rect 161 22934 167 22955
rect 233 22934 259 22955
rect 161 22921 199 22934
rect 233 22921 271 22934
rect 305 22921 343 22955
rect 377 22921 415 22955
rect 449 22934 459 22955
rect 521 22934 537 22955
rect 593 22934 615 22955
rect 665 22934 693 22955
rect 737 22934 771 22955
rect 449 22921 487 22934
rect 521 22921 559 22934
rect 593 22921 631 22934
rect 665 22921 703 22934
rect 737 22921 775 22934
rect 809 22921 983 22955
rect -23 22895 983 22921
rect -23 22853 -17 22895
rect 17 22887 75 22895
rect 109 22887 167 22895
rect 201 22887 259 22895
rect 293 22887 459 22895
rect 493 22887 537 22895
rect 571 22887 615 22895
rect 649 22887 693 22895
rect 727 22887 771 22895
rect 805 22887 983 22895
rect 17 22853 55 22887
rect 109 22861 127 22887
rect 89 22853 127 22861
rect 161 22861 167 22887
rect 233 22861 259 22887
rect 161 22853 199 22861
rect 233 22853 271 22861
rect 305 22853 343 22887
rect 377 22853 415 22887
rect 449 22861 459 22887
rect 521 22861 537 22887
rect 593 22861 615 22887
rect 665 22861 693 22887
rect 737 22861 771 22887
rect 449 22853 487 22861
rect 521 22853 559 22861
rect 593 22853 631 22861
rect 665 22853 703 22861
rect 737 22853 775 22861
rect 809 22853 983 22887
rect -23 22822 983 22853
rect -23 22785 -17 22822
rect 17 22819 75 22822
rect 109 22819 167 22822
rect 201 22819 259 22822
rect 293 22819 459 22822
rect 493 22819 537 22822
rect 571 22819 615 22822
rect 649 22819 693 22822
rect 727 22819 771 22822
rect 805 22819 983 22822
rect 17 22785 55 22819
rect 109 22788 127 22819
rect 89 22785 127 22788
rect 161 22788 167 22819
rect 233 22788 259 22819
rect 161 22785 199 22788
rect 233 22785 271 22788
rect 305 22785 343 22819
rect 377 22785 415 22819
rect 449 22788 459 22819
rect 521 22788 537 22819
rect 593 22788 615 22819
rect 665 22788 693 22819
rect 737 22788 771 22819
rect 449 22785 487 22788
rect 521 22785 559 22788
rect 593 22785 631 22788
rect 665 22785 703 22788
rect 737 22785 775 22788
rect 809 22785 983 22819
rect -23 22751 983 22785
rect -23 22715 -17 22751
rect 17 22717 55 22751
rect 89 22749 127 22751
rect 109 22717 127 22749
rect 161 22749 199 22751
rect 233 22749 271 22751
rect 161 22717 167 22749
rect 233 22717 259 22749
rect 305 22717 343 22751
rect 377 22717 415 22751
rect 449 22749 487 22751
rect 521 22749 559 22751
rect 593 22749 631 22751
rect 665 22749 703 22751
rect 737 22749 775 22751
rect 449 22717 459 22749
rect 521 22717 537 22749
rect 593 22717 615 22749
rect 665 22717 693 22749
rect 737 22717 771 22749
rect 809 22717 983 22751
rect 17 22715 75 22717
rect 109 22715 167 22717
rect 201 22715 259 22717
rect 293 22715 459 22717
rect 493 22715 537 22717
rect 571 22715 615 22717
rect 649 22715 693 22717
rect 727 22715 771 22717
rect 805 22715 983 22717
rect -23 22683 983 22715
rect -23 22642 -17 22683
rect 17 22649 55 22683
rect 89 22676 127 22683
rect 109 22649 127 22676
rect 161 22676 199 22683
rect 233 22676 271 22683
rect 161 22649 167 22676
rect 233 22649 259 22676
rect 305 22649 343 22683
rect 377 22649 415 22683
rect 449 22676 487 22683
rect 521 22676 559 22683
rect 593 22676 631 22683
rect 665 22676 703 22683
rect 737 22676 775 22683
rect 449 22649 459 22676
rect 521 22649 537 22676
rect 593 22649 615 22676
rect 665 22649 693 22676
rect 737 22649 771 22676
rect 809 22649 983 22683
rect 17 22642 75 22649
rect 109 22642 167 22649
rect 201 22642 259 22649
rect 293 22642 459 22649
rect 493 22642 537 22649
rect 571 22642 615 22649
rect 649 22642 693 22649
rect 727 22642 771 22649
rect 805 22642 983 22649
rect -23 22615 983 22642
rect -23 22569 -17 22615
rect 17 22581 55 22615
rect 89 22603 127 22615
rect 109 22581 127 22603
rect 161 22603 199 22615
rect 233 22603 271 22615
rect 161 22581 167 22603
rect 233 22581 259 22603
rect 305 22581 343 22615
rect 377 22581 415 22615
rect 449 22603 487 22615
rect 521 22603 559 22615
rect 593 22603 631 22615
rect 665 22603 703 22615
rect 737 22603 775 22615
rect 449 22581 459 22603
rect 521 22581 537 22603
rect 593 22581 615 22603
rect 665 22581 693 22603
rect 737 22581 771 22603
rect 809 22581 983 22615
rect 17 22569 75 22581
rect 109 22569 167 22581
rect 201 22569 259 22581
rect 293 22569 459 22581
rect 493 22569 537 22581
rect 571 22569 615 22581
rect 649 22569 693 22581
rect 727 22569 771 22581
rect 805 22569 983 22581
rect -23 22547 983 22569
rect -23 22496 -17 22547
rect 17 22513 55 22547
rect 89 22530 127 22547
rect 109 22513 127 22530
rect 161 22530 199 22547
rect 233 22530 271 22547
rect 161 22513 167 22530
rect 233 22513 259 22530
rect 305 22513 343 22547
rect 377 22513 415 22547
rect 449 22530 487 22547
rect 521 22530 559 22547
rect 593 22530 631 22547
rect 665 22530 703 22547
rect 737 22530 775 22547
rect 449 22513 459 22530
rect 521 22513 537 22530
rect 593 22513 615 22530
rect 665 22513 693 22530
rect 737 22513 771 22530
rect 809 22513 983 22547
rect 17 22496 75 22513
rect 109 22496 167 22513
rect 201 22496 259 22513
rect 293 22496 459 22513
rect 493 22496 537 22513
rect 571 22496 615 22513
rect 649 22496 693 22513
rect 727 22496 771 22513
rect 805 22496 983 22513
rect -23 22479 983 22496
rect -23 22423 -17 22479
rect 17 22445 55 22479
rect 89 22457 127 22479
rect 109 22445 127 22457
rect 161 22457 199 22479
rect 233 22457 271 22479
rect 161 22445 167 22457
rect 233 22445 259 22457
rect 305 22445 343 22479
rect 377 22445 415 22479
rect 449 22457 487 22479
rect 521 22457 559 22479
rect 593 22457 631 22479
rect 665 22457 703 22479
rect 737 22457 775 22479
rect 449 22445 459 22457
rect 521 22445 537 22457
rect 593 22445 615 22457
rect 665 22445 693 22457
rect 737 22445 771 22457
rect 809 22445 983 22479
rect 17 22423 75 22445
rect 109 22423 167 22445
rect 201 22423 259 22445
rect 293 22423 459 22445
rect 493 22423 537 22445
rect 571 22423 615 22445
rect 649 22423 693 22445
rect 727 22423 771 22445
rect 805 22423 983 22445
rect -23 22411 983 22423
rect -23 22350 -17 22411
rect 17 22377 55 22411
rect 89 22384 127 22411
rect 109 22377 127 22384
rect 161 22384 199 22411
rect 233 22384 271 22411
rect 161 22377 167 22384
rect 233 22377 259 22384
rect 305 22377 343 22411
rect 377 22377 415 22411
rect 449 22384 487 22411
rect 521 22384 559 22411
rect 593 22384 631 22411
rect 665 22384 703 22411
rect 737 22384 775 22411
rect 449 22377 459 22384
rect 521 22377 537 22384
rect 593 22377 615 22384
rect 665 22377 693 22384
rect 737 22377 771 22384
rect 809 22377 983 22411
rect 17 22350 75 22377
rect 109 22350 167 22377
rect 201 22350 259 22377
rect 293 22350 459 22377
rect 493 22350 537 22377
rect 571 22350 615 22377
rect 649 22350 693 22377
rect 727 22350 771 22377
rect 805 22350 983 22377
rect -23 22343 983 22350
rect -23 22277 -17 22343
rect 17 22309 55 22343
rect 89 22311 127 22343
rect 109 22309 127 22311
rect 161 22311 199 22343
rect 233 22311 271 22343
rect 161 22309 167 22311
rect 233 22309 259 22311
rect 305 22309 343 22343
rect 377 22309 415 22343
rect 449 22311 487 22343
rect 521 22311 559 22343
rect 593 22311 631 22343
rect 665 22311 703 22343
rect 737 22311 775 22343
rect 449 22309 459 22311
rect 521 22309 537 22311
rect 593 22309 615 22311
rect 665 22309 693 22311
rect 737 22309 771 22311
rect 809 22309 983 22343
rect 17 22277 75 22309
rect 109 22277 167 22309
rect 201 22277 259 22309
rect 293 22277 459 22309
rect 493 22277 537 22309
rect 571 22277 615 22309
rect 649 22277 693 22309
rect 727 22277 771 22309
rect 805 22277 983 22309
rect -23 22275 983 22277
rect -23 22241 -17 22275
rect 17 22241 55 22275
rect 89 22241 127 22275
rect 161 22241 199 22275
rect 233 22241 271 22275
rect 305 22241 343 22275
rect 377 22241 415 22275
rect 449 22241 487 22275
rect 521 22241 559 22275
rect 593 22241 631 22275
rect 665 22241 703 22275
rect 737 22241 775 22275
rect 809 22241 983 22275
rect -23 22238 983 22241
rect -23 22173 -17 22238
rect 17 22207 75 22238
rect 109 22207 167 22238
rect 201 22207 259 22238
rect 293 22207 459 22238
rect 493 22207 537 22238
rect 571 22207 615 22238
rect 649 22207 693 22238
rect 727 22207 771 22238
rect 805 22207 983 22238
rect 17 22173 55 22207
rect 109 22204 127 22207
rect 89 22173 127 22204
rect 161 22204 167 22207
rect 233 22204 259 22207
rect 161 22173 199 22204
rect 233 22173 271 22204
rect 305 22173 343 22207
rect 377 22173 415 22207
rect 449 22204 459 22207
rect 521 22204 537 22207
rect 593 22204 615 22207
rect 665 22204 693 22207
rect 737 22204 771 22207
rect 449 22173 487 22204
rect 521 22173 559 22204
rect 593 22173 631 22204
rect 665 22173 703 22204
rect 737 22173 775 22204
rect 809 22173 983 22207
rect -23 22165 983 22173
rect -23 22105 -17 22165
rect 17 22139 75 22165
rect 109 22139 167 22165
rect 201 22139 259 22165
rect 293 22139 459 22165
rect 493 22139 537 22165
rect 571 22139 615 22165
rect 649 22139 693 22165
rect 727 22139 771 22165
rect 805 22139 983 22165
rect 17 22105 55 22139
rect 109 22131 127 22139
rect 89 22105 127 22131
rect 161 22131 167 22139
rect 233 22131 259 22139
rect 161 22105 199 22131
rect 233 22105 271 22131
rect 305 22105 343 22139
rect 377 22105 415 22139
rect 449 22131 459 22139
rect 521 22131 537 22139
rect 593 22131 615 22139
rect 665 22131 693 22139
rect 737 22131 771 22139
rect 449 22105 487 22131
rect 521 22105 559 22131
rect 593 22105 631 22131
rect 665 22105 703 22131
rect 737 22105 775 22131
rect 809 22105 983 22139
rect -23 22092 983 22105
rect -23 22037 -17 22092
rect 17 22071 75 22092
rect 109 22071 167 22092
rect 201 22071 259 22092
rect 293 22071 459 22092
rect 493 22071 537 22092
rect 571 22071 615 22092
rect 649 22071 693 22092
rect 727 22071 771 22092
rect 805 22071 983 22092
rect 17 22037 55 22071
rect 109 22058 127 22071
rect 89 22037 127 22058
rect 161 22058 167 22071
rect 233 22058 259 22071
rect 161 22037 199 22058
rect 233 22037 271 22058
rect 305 22037 343 22071
rect 377 22037 415 22071
rect 449 22058 459 22071
rect 521 22058 537 22071
rect 593 22058 615 22071
rect 665 22058 693 22071
rect 737 22058 771 22071
rect 449 22037 487 22058
rect 521 22037 559 22058
rect 593 22037 631 22058
rect 665 22037 703 22058
rect 737 22037 775 22058
rect 809 22037 983 22071
rect -23 22019 983 22037
rect -23 21969 -17 22019
rect 17 22003 75 22019
rect 109 22003 167 22019
rect 201 22003 259 22019
rect 293 22003 459 22019
rect 493 22003 537 22019
rect 571 22003 615 22019
rect 649 22003 693 22019
rect 727 22003 771 22019
rect 805 22003 983 22019
rect 17 21969 55 22003
rect 109 21985 127 22003
rect 89 21969 127 21985
rect 161 21985 167 22003
rect 233 21985 259 22003
rect 161 21969 199 21985
rect 233 21969 271 21985
rect 305 21969 343 22003
rect 377 21969 415 22003
rect 449 21985 459 22003
rect 521 21985 537 22003
rect 593 21985 615 22003
rect 665 21985 693 22003
rect 737 21985 771 22003
rect 449 21969 487 21985
rect 521 21969 559 21985
rect 593 21969 631 21985
rect 665 21969 703 21985
rect 737 21969 775 21985
rect 809 21969 983 22003
rect -23 21946 983 21969
rect -23 21901 -17 21946
rect 17 21935 75 21946
rect 109 21935 167 21946
rect 201 21935 259 21946
rect 293 21935 459 21946
rect 493 21935 537 21946
rect 571 21935 615 21946
rect 649 21935 693 21946
rect 727 21935 771 21946
rect 805 21935 983 21946
rect 17 21901 55 21935
rect 109 21912 127 21935
rect 89 21901 127 21912
rect 161 21912 167 21935
rect 233 21912 259 21935
rect 161 21901 199 21912
rect 233 21901 271 21912
rect 305 21901 343 21935
rect 377 21901 415 21935
rect 449 21912 459 21935
rect 521 21912 537 21935
rect 593 21912 615 21935
rect 665 21912 693 21935
rect 737 21912 771 21935
rect 449 21901 487 21912
rect 521 21901 559 21912
rect 593 21901 631 21912
rect 665 21901 703 21912
rect 737 21901 775 21912
rect 809 21901 983 21935
rect -23 21873 983 21901
rect -23 21833 -17 21873
rect 17 21867 75 21873
rect 109 21867 167 21873
rect 201 21867 259 21873
rect 293 21867 459 21873
rect 493 21867 537 21873
rect 571 21867 615 21873
rect 649 21867 693 21873
rect 727 21867 771 21873
rect 805 21867 983 21873
rect 17 21833 55 21867
rect 109 21839 127 21867
rect 89 21833 127 21839
rect 161 21839 167 21867
rect 233 21839 259 21867
rect 161 21833 199 21839
rect 233 21833 271 21839
rect 305 21833 343 21867
rect 377 21833 415 21867
rect 449 21839 459 21867
rect 521 21839 537 21867
rect 593 21839 615 21867
rect 665 21839 693 21867
rect 737 21839 771 21867
rect 449 21833 487 21839
rect 521 21833 559 21839
rect 593 21833 631 21839
rect 665 21833 703 21839
rect 737 21833 775 21839
rect 809 21833 983 21867
rect -23 21800 983 21833
rect -23 21765 -17 21800
rect 17 21799 75 21800
rect 109 21799 167 21800
rect 201 21799 259 21800
rect 293 21799 459 21800
rect 493 21799 537 21800
rect 571 21799 615 21800
rect 649 21799 693 21800
rect 727 21799 771 21800
rect 805 21799 983 21800
rect 17 21765 55 21799
rect 109 21766 127 21799
rect 89 21765 127 21766
rect 161 21766 167 21799
rect 233 21766 259 21799
rect 161 21765 199 21766
rect 233 21765 271 21766
rect 305 21765 343 21799
rect 377 21765 415 21799
rect 449 21766 459 21799
rect 521 21766 537 21799
rect 593 21766 615 21799
rect 665 21766 693 21799
rect 737 21766 771 21799
rect 449 21765 487 21766
rect 521 21765 559 21766
rect 593 21765 631 21766
rect 665 21765 703 21766
rect 737 21765 775 21766
rect 809 21765 983 21799
rect -23 21731 983 21765
rect -23 21693 -17 21731
rect 17 21697 55 21731
rect 89 21727 127 21731
rect 109 21697 127 21727
rect 161 21727 199 21731
rect 233 21727 271 21731
rect 161 21697 167 21727
rect 233 21697 259 21727
rect 305 21697 343 21731
rect 377 21697 415 21731
rect 449 21727 487 21731
rect 521 21727 559 21731
rect 593 21727 631 21731
rect 665 21727 703 21731
rect 737 21727 775 21731
rect 449 21697 459 21727
rect 521 21697 537 21727
rect 593 21697 615 21727
rect 665 21697 693 21727
rect 737 21697 771 21727
rect 809 21697 983 21731
rect 17 21693 75 21697
rect 109 21693 167 21697
rect 201 21693 259 21697
rect 293 21693 459 21697
rect 493 21693 537 21697
rect 571 21693 615 21697
rect 649 21693 693 21697
rect 727 21693 771 21697
rect 805 21693 983 21697
rect -23 21663 983 21693
rect -23 21620 -17 21663
rect 17 21629 55 21663
rect 89 21654 127 21663
rect 109 21629 127 21654
rect 161 21654 199 21663
rect 233 21654 271 21663
rect 161 21629 167 21654
rect 233 21629 259 21654
rect 305 21629 343 21663
rect 377 21629 415 21663
rect 449 21654 487 21663
rect 521 21654 559 21663
rect 593 21654 631 21663
rect 665 21654 703 21663
rect 737 21654 775 21663
rect 449 21629 459 21654
rect 521 21629 537 21654
rect 593 21629 615 21654
rect 665 21629 693 21654
rect 737 21629 771 21654
rect 809 21629 983 21663
rect 17 21620 75 21629
rect 109 21620 167 21629
rect 201 21620 259 21629
rect 293 21620 459 21629
rect 493 21620 537 21629
rect 571 21620 615 21629
rect 649 21620 693 21629
rect 727 21620 771 21629
rect 805 21620 983 21629
rect -23 21595 983 21620
rect -23 21547 -17 21595
rect 17 21561 55 21595
rect 89 21581 127 21595
rect 109 21561 127 21581
rect 161 21581 199 21595
rect 233 21581 271 21595
rect 161 21561 167 21581
rect 233 21561 259 21581
rect 305 21561 343 21595
rect 377 21561 415 21595
rect 449 21581 487 21595
rect 521 21581 559 21595
rect 593 21581 631 21595
rect 665 21581 703 21595
rect 737 21581 775 21595
rect 449 21561 459 21581
rect 521 21561 537 21581
rect 593 21561 615 21581
rect 665 21561 693 21581
rect 737 21561 771 21581
rect 809 21561 983 21595
rect 17 21547 75 21561
rect 109 21547 167 21561
rect 201 21547 259 21561
rect 293 21547 459 21561
rect 493 21547 537 21561
rect 571 21547 615 21561
rect 649 21547 693 21561
rect 727 21547 771 21561
rect 805 21547 983 21561
rect -23 21527 983 21547
rect -23 21474 -17 21527
rect 17 21493 55 21527
rect 89 21508 127 21527
rect 109 21493 127 21508
rect 161 21508 199 21527
rect 233 21508 271 21527
rect 161 21493 167 21508
rect 233 21493 259 21508
rect 305 21493 343 21527
rect 377 21493 415 21527
rect 449 21508 487 21527
rect 521 21508 559 21527
rect 593 21508 631 21527
rect 665 21508 703 21527
rect 737 21508 775 21527
rect 449 21493 459 21508
rect 521 21493 537 21508
rect 593 21493 615 21508
rect 665 21493 693 21508
rect 737 21493 771 21508
rect 809 21493 983 21527
rect 17 21474 75 21493
rect 109 21474 167 21493
rect 201 21474 259 21493
rect 293 21474 459 21493
rect 493 21474 537 21493
rect 571 21474 615 21493
rect 649 21474 693 21493
rect 727 21474 771 21493
rect 805 21474 983 21493
rect -23 21459 983 21474
rect -23 21401 -17 21459
rect 17 21425 55 21459
rect 89 21435 127 21459
rect 109 21425 127 21435
rect 161 21435 199 21459
rect 233 21435 271 21459
rect 161 21425 167 21435
rect 233 21425 259 21435
rect 305 21425 343 21459
rect 377 21425 415 21459
rect 449 21435 487 21459
rect 521 21435 559 21459
rect 593 21435 631 21459
rect 665 21435 703 21459
rect 737 21435 775 21459
rect 449 21425 459 21435
rect 521 21425 537 21435
rect 593 21425 615 21435
rect 665 21425 693 21435
rect 737 21425 771 21435
rect 809 21425 983 21459
rect 17 21401 75 21425
rect 109 21401 167 21425
rect 201 21401 259 21425
rect 293 21401 459 21425
rect 493 21401 537 21425
rect 571 21401 615 21425
rect 649 21401 693 21425
rect 727 21401 771 21425
rect 805 21401 983 21425
rect -23 21391 983 21401
rect -23 21328 -17 21391
rect 17 21357 55 21391
rect 89 21362 127 21391
rect 109 21357 127 21362
rect 161 21362 199 21391
rect 233 21362 271 21391
rect 161 21357 167 21362
rect 233 21357 259 21362
rect 305 21357 343 21391
rect 377 21357 415 21391
rect 449 21362 487 21391
rect 521 21362 559 21391
rect 593 21362 631 21391
rect 665 21362 703 21391
rect 737 21362 775 21391
rect 449 21357 459 21362
rect 521 21357 537 21362
rect 593 21357 615 21362
rect 665 21357 693 21362
rect 737 21357 771 21362
rect 809 21357 983 21391
rect 17 21328 75 21357
rect 109 21328 167 21357
rect 201 21328 259 21357
rect 293 21328 459 21357
rect 493 21328 537 21357
rect 571 21328 615 21357
rect 649 21328 693 21357
rect 727 21328 771 21357
rect 805 21328 983 21357
rect -23 21323 983 21328
rect -23 21221 -17 21323
rect 17 21289 55 21323
rect 89 21289 127 21323
rect 161 21289 199 21323
rect 233 21289 271 21323
rect 305 21289 343 21323
rect 377 21289 415 21323
rect 449 21289 487 21323
rect 521 21289 559 21323
rect 593 21289 631 21323
rect 665 21289 703 21323
rect 737 21289 775 21323
rect 809 21289 983 21323
rect 17 21255 75 21289
rect 109 21255 167 21289
rect 201 21255 259 21289
rect 293 21255 459 21289
rect 493 21255 537 21289
rect 571 21255 615 21289
rect 649 21255 693 21289
rect 727 21255 771 21289
rect 805 21255 983 21289
rect 17 21221 55 21255
rect 89 21221 127 21255
rect 161 21221 199 21255
rect 233 21221 271 21255
rect 305 21221 343 21255
rect 377 21221 415 21255
rect 449 21221 487 21255
rect 521 21221 559 21255
rect 593 21221 631 21255
rect 665 21221 703 21255
rect 737 21221 775 21255
rect 809 21221 983 21255
rect -23 21216 983 21221
rect -23 21153 -17 21216
rect 17 21187 75 21216
rect 109 21187 167 21216
rect 201 21187 259 21216
rect 293 21187 459 21216
rect 493 21187 537 21216
rect 571 21187 615 21216
rect 649 21187 693 21216
rect 727 21187 771 21216
rect 805 21187 983 21216
rect 17 21153 55 21187
rect 109 21182 127 21187
rect 89 21153 127 21182
rect 161 21182 167 21187
rect 233 21182 259 21187
rect 161 21153 199 21182
rect 233 21153 271 21182
rect 305 21153 343 21187
rect 377 21153 415 21187
rect 449 21182 459 21187
rect 521 21182 537 21187
rect 593 21182 615 21187
rect 665 21182 693 21187
rect 737 21182 771 21187
rect 449 21153 487 21182
rect 521 21153 559 21182
rect 593 21153 631 21182
rect 665 21153 703 21182
rect 737 21153 775 21182
rect 809 21153 983 21187
rect -23 21143 983 21153
rect -23 21085 -17 21143
rect 17 21119 75 21143
rect 109 21119 167 21143
rect 201 21119 259 21143
rect 293 21119 459 21143
rect 493 21119 537 21143
rect 571 21119 615 21143
rect 649 21119 693 21143
rect 727 21119 771 21143
rect 805 21119 983 21143
rect 17 21085 55 21119
rect 109 21109 127 21119
rect 89 21085 127 21109
rect 161 21109 167 21119
rect 233 21109 259 21119
rect 161 21085 199 21109
rect 233 21085 271 21109
rect 305 21085 343 21119
rect 377 21085 415 21119
rect 449 21109 459 21119
rect 521 21109 537 21119
rect 593 21109 615 21119
rect 665 21109 693 21119
rect 737 21109 771 21119
rect 449 21085 487 21109
rect 521 21085 559 21109
rect 593 21085 631 21109
rect 665 21085 703 21109
rect 737 21085 775 21109
rect 809 21085 983 21119
rect -23 21070 983 21085
rect -23 21017 -17 21070
rect 17 21051 75 21070
rect 109 21051 167 21070
rect 201 21051 259 21070
rect 293 21051 459 21070
rect 493 21051 537 21070
rect 571 21051 615 21070
rect 649 21051 693 21070
rect 727 21051 771 21070
rect 805 21051 983 21070
rect 17 21017 55 21051
rect 109 21036 127 21051
rect 89 21017 127 21036
rect 161 21036 167 21051
rect 233 21036 259 21051
rect 161 21017 199 21036
rect 233 21017 271 21036
rect 305 21017 343 21051
rect 377 21017 415 21051
rect 449 21036 459 21051
rect 521 21036 537 21051
rect 593 21036 615 21051
rect 665 21036 693 21051
rect 737 21036 771 21051
rect 449 21017 487 21036
rect 521 21017 559 21036
rect 593 21017 631 21036
rect 665 21017 703 21036
rect 737 21017 775 21036
rect 809 21017 983 21051
rect -23 20997 983 21017
rect -23 20949 -17 20997
rect 17 20983 75 20997
rect 109 20983 167 20997
rect 201 20983 259 20997
rect 293 20983 459 20997
rect 493 20983 537 20997
rect 571 20983 615 20997
rect 649 20983 693 20997
rect 727 20983 771 20997
rect 805 20983 983 20997
rect 17 20949 55 20983
rect 109 20963 127 20983
rect 89 20949 127 20963
rect 161 20963 167 20983
rect 233 20963 259 20983
rect 161 20949 199 20963
rect 233 20949 271 20963
rect 305 20949 343 20983
rect 377 20949 415 20983
rect 449 20963 459 20983
rect 521 20963 537 20983
rect 593 20963 615 20983
rect 665 20963 693 20983
rect 737 20963 771 20983
rect 449 20949 487 20963
rect 521 20949 559 20963
rect 593 20949 631 20963
rect 665 20949 703 20963
rect 737 20949 775 20963
rect 809 20949 983 20983
rect -23 20924 983 20949
rect -23 20881 -17 20924
rect 17 20915 75 20924
rect 109 20915 167 20924
rect 201 20915 259 20924
rect 293 20915 459 20924
rect 493 20915 537 20924
rect 571 20915 615 20924
rect 649 20915 693 20924
rect 727 20915 771 20924
rect 805 20915 983 20924
rect 17 20881 55 20915
rect 109 20890 127 20915
rect 89 20881 127 20890
rect 161 20890 167 20915
rect 233 20890 259 20915
rect 161 20881 199 20890
rect 233 20881 271 20890
rect 305 20881 343 20915
rect 377 20881 415 20915
rect 449 20890 459 20915
rect 521 20890 537 20915
rect 593 20890 615 20915
rect 665 20890 693 20915
rect 737 20890 771 20915
rect 449 20881 487 20890
rect 521 20881 559 20890
rect 593 20881 631 20890
rect 665 20881 703 20890
rect 737 20881 775 20890
rect 809 20881 983 20915
rect -23 20851 983 20881
rect -23 20813 -17 20851
rect 17 20847 75 20851
rect 109 20847 167 20851
rect 201 20847 259 20851
rect 293 20847 459 20851
rect 493 20847 537 20851
rect 571 20847 615 20851
rect 649 20847 693 20851
rect 727 20847 771 20851
rect 805 20847 983 20851
rect 17 20813 55 20847
rect 109 20817 127 20847
rect 89 20813 127 20817
rect 161 20817 167 20847
rect 233 20817 259 20847
rect 161 20813 199 20817
rect 233 20813 271 20817
rect 305 20813 343 20847
rect 377 20813 415 20847
rect 449 20817 459 20847
rect 521 20817 537 20847
rect 593 20817 615 20847
rect 665 20817 693 20847
rect 737 20817 771 20847
rect 449 20813 487 20817
rect 521 20813 559 20817
rect 593 20813 631 20817
rect 665 20813 703 20817
rect 737 20813 775 20817
rect 809 20813 983 20847
rect -23 20779 983 20813
rect -23 20744 -17 20779
rect 17 20745 55 20779
rect 89 20778 127 20779
rect 109 20745 127 20778
rect 161 20778 199 20779
rect 233 20778 271 20779
rect 161 20745 167 20778
rect 233 20745 259 20778
rect 305 20745 343 20779
rect 377 20745 415 20779
rect 449 20778 487 20779
rect 521 20778 559 20779
rect 593 20778 631 20779
rect 665 20778 703 20779
rect 737 20778 775 20779
rect 449 20745 459 20778
rect 521 20745 537 20778
rect 593 20745 615 20778
rect 665 20745 693 20778
rect 737 20745 771 20778
rect 809 20745 983 20779
rect 17 20744 75 20745
rect 109 20744 167 20745
rect 201 20744 259 20745
rect 293 20744 459 20745
rect 493 20744 537 20745
rect 571 20744 615 20745
rect 649 20744 693 20745
rect 727 20744 771 20745
rect 805 20744 983 20745
rect -23 20711 983 20744
rect -23 20671 -17 20711
rect 17 20677 55 20711
rect 89 20705 127 20711
rect 109 20677 127 20705
rect 161 20705 199 20711
rect 233 20705 271 20711
rect 161 20677 167 20705
rect 233 20677 259 20705
rect 305 20677 343 20711
rect 377 20677 415 20711
rect 449 20705 487 20711
rect 521 20705 559 20711
rect 593 20705 631 20711
rect 665 20705 703 20711
rect 737 20705 775 20711
rect 449 20677 459 20705
rect 521 20677 537 20705
rect 593 20677 615 20705
rect 665 20677 693 20705
rect 737 20677 771 20705
rect 809 20677 983 20711
rect 17 20671 75 20677
rect 109 20671 167 20677
rect 201 20671 259 20677
rect 293 20671 459 20677
rect 493 20671 537 20677
rect 571 20671 615 20677
rect 649 20671 693 20677
rect 727 20671 771 20677
rect 805 20671 983 20677
rect -23 20643 983 20671
rect -23 20598 -17 20643
rect 17 20609 55 20643
rect 89 20632 127 20643
rect 109 20609 127 20632
rect 161 20632 199 20643
rect 233 20632 271 20643
rect 161 20609 167 20632
rect 233 20609 259 20632
rect 305 20609 343 20643
rect 377 20609 415 20643
rect 449 20632 487 20643
rect 521 20632 559 20643
rect 593 20632 631 20643
rect 665 20632 703 20643
rect 737 20632 775 20643
rect 449 20609 459 20632
rect 521 20609 537 20632
rect 593 20609 615 20632
rect 665 20609 693 20632
rect 737 20609 771 20632
rect 809 20609 983 20643
rect 17 20598 75 20609
rect 109 20598 167 20609
rect 201 20598 259 20609
rect 293 20598 459 20609
rect 493 20598 537 20609
rect 571 20598 615 20609
rect 649 20598 693 20609
rect 727 20598 771 20609
rect 805 20598 983 20609
rect -23 20575 983 20598
rect -23 20525 -17 20575
rect 17 20541 55 20575
rect 89 20559 127 20575
rect 109 20541 127 20559
rect 161 20559 199 20575
rect 233 20559 271 20575
rect 161 20541 167 20559
rect 233 20541 259 20559
rect 305 20541 343 20575
rect 377 20541 415 20575
rect 449 20559 487 20575
rect 521 20559 559 20575
rect 593 20559 631 20575
rect 665 20559 703 20575
rect 737 20559 775 20575
rect 449 20541 459 20559
rect 521 20541 537 20559
rect 593 20541 615 20559
rect 665 20541 693 20559
rect 737 20541 771 20559
rect 809 20541 983 20575
rect 17 20525 75 20541
rect 109 20525 167 20541
rect 201 20525 259 20541
rect 293 20525 459 20541
rect 493 20525 537 20541
rect 571 20525 615 20541
rect 649 20525 693 20541
rect 727 20525 771 20541
rect 805 20525 983 20541
rect -23 20507 983 20525
rect -23 20452 -17 20507
rect 17 20473 55 20507
rect 89 20486 127 20507
rect 109 20473 127 20486
rect 161 20486 199 20507
rect 233 20486 271 20507
rect 161 20473 167 20486
rect 233 20473 259 20486
rect 305 20473 343 20507
rect 377 20473 415 20507
rect 449 20486 487 20507
rect 521 20486 559 20507
rect 593 20486 631 20507
rect 665 20486 703 20507
rect 737 20486 775 20507
rect 449 20473 459 20486
rect 521 20473 537 20486
rect 593 20473 615 20486
rect 665 20473 693 20486
rect 737 20473 771 20486
rect 809 20484 983 20507
rect 809 20473 843 20484
rect 17 20452 75 20473
rect 109 20452 167 20473
rect 201 20452 259 20473
rect 293 20452 459 20473
rect 493 20452 537 20473
rect 571 20452 615 20473
rect 649 20452 693 20473
rect 727 20452 771 20473
rect 805 20452 843 20473
rect -23 20450 843 20452
rect 877 20450 915 20484
rect 949 20450 983 20484
rect -23 20439 983 20450
rect -23 20379 -17 20439
rect 17 20405 55 20439
rect 89 20413 127 20439
rect 109 20405 127 20413
rect 161 20413 199 20439
rect 233 20413 271 20439
rect 161 20405 167 20413
rect 233 20405 259 20413
rect 305 20405 343 20439
rect 377 20405 415 20439
rect 449 20413 487 20439
rect 521 20413 559 20439
rect 593 20413 631 20439
rect 665 20413 703 20439
rect 737 20413 775 20439
rect 809 20418 983 20439
rect 809 20415 868 20418
rect 902 20415 983 20418
rect 449 20405 459 20413
rect 521 20405 537 20413
rect 593 20405 615 20413
rect 665 20405 693 20413
rect 737 20405 771 20413
rect 17 20379 75 20405
rect 109 20379 167 20405
rect 201 20379 259 20405
rect 293 20379 459 20405
rect 493 20379 537 20405
rect 571 20379 615 20405
rect 649 20379 693 20405
rect 727 20379 771 20405
rect 902 20384 915 20415
rect 877 20381 915 20384
rect 949 20381 983 20415
rect -23 20371 775 20379
rect -23 20306 -17 20371
rect 17 20337 55 20371
rect 89 20340 127 20371
rect 109 20337 127 20340
rect 161 20340 199 20371
rect 233 20340 271 20371
rect 161 20337 167 20340
rect 233 20337 259 20340
rect 305 20337 343 20371
rect 377 20337 415 20371
rect 449 20340 487 20371
rect 521 20340 559 20371
rect 593 20340 631 20371
rect 665 20340 703 20371
rect 737 20340 775 20371
rect 877 20347 983 20381
rect 877 20343 915 20347
rect 449 20337 459 20340
rect 521 20337 537 20340
rect 593 20337 615 20340
rect 665 20337 693 20340
rect 737 20337 771 20340
rect 17 20306 75 20337
rect 109 20306 167 20337
rect 201 20306 259 20337
rect 293 20306 459 20337
rect 493 20306 537 20337
rect 571 20306 615 20337
rect 649 20306 693 20337
rect 727 20306 771 20337
rect 902 20313 915 20343
rect 949 20313 983 20347
rect 902 20309 983 20313
rect -23 20303 775 20306
rect -23 20269 -17 20303
rect 17 20269 55 20303
rect 89 20269 127 20303
rect 161 20269 199 20303
rect 233 20269 271 20303
rect 305 20269 343 20303
rect 377 20269 415 20303
rect 449 20269 487 20303
rect 521 20269 559 20303
rect 593 20269 631 20303
rect 665 20269 703 20303
rect 737 20269 775 20303
rect -23 20267 775 20269
rect 877 20279 983 20309
rect 877 20268 915 20279
rect -23 20201 -17 20267
rect 17 20235 75 20267
rect 109 20235 167 20267
rect 201 20235 259 20267
rect 293 20235 459 20267
rect 493 20235 537 20267
rect 571 20235 615 20267
rect 649 20235 693 20267
rect 727 20235 771 20267
rect 17 20201 55 20235
rect 109 20233 127 20235
rect 89 20201 127 20233
rect 161 20233 167 20235
rect 233 20233 259 20235
rect 161 20201 199 20233
rect 233 20201 271 20233
rect 305 20201 343 20235
rect 377 20201 415 20235
rect 449 20233 459 20235
rect 521 20233 537 20235
rect 593 20233 615 20235
rect 665 20233 693 20235
rect 737 20233 771 20235
rect 902 20245 915 20268
rect 949 20245 983 20279
rect 902 20234 983 20245
rect 449 20201 487 20233
rect 521 20201 559 20233
rect 593 20201 631 20233
rect 665 20201 703 20233
rect 737 20201 775 20233
rect -23 20194 775 20201
rect 877 20211 983 20234
rect -23 20133 -17 20194
rect 17 20167 75 20194
rect 109 20167 167 20194
rect 201 20167 259 20194
rect 293 20167 459 20194
rect 493 20167 537 20194
rect 571 20167 615 20194
rect 649 20167 693 20194
rect 727 20167 771 20194
rect 17 20133 55 20167
rect 109 20160 127 20167
rect 89 20133 127 20160
rect 161 20160 167 20167
rect 233 20160 259 20167
rect 161 20133 199 20160
rect 233 20133 271 20160
rect 305 20133 343 20167
rect 377 20133 415 20167
rect 449 20160 459 20167
rect 521 20160 537 20167
rect 593 20160 615 20167
rect 665 20160 693 20167
rect 737 20160 771 20167
rect 877 20193 915 20211
rect 449 20133 487 20160
rect 521 20133 559 20160
rect 593 20133 631 20160
rect 665 20133 703 20160
rect 737 20133 775 20160
rect 902 20177 915 20193
rect 949 20177 983 20211
rect 902 20159 983 20177
rect -23 20121 775 20133
rect 877 20143 983 20159
rect -23 20065 -17 20121
rect 17 20099 75 20121
rect 109 20099 167 20121
rect 201 20099 259 20121
rect 293 20099 459 20121
rect 493 20099 537 20121
rect 571 20099 615 20121
rect 649 20099 693 20121
rect 727 20099 771 20121
rect 17 20065 55 20099
rect 109 20087 127 20099
rect 89 20065 127 20087
rect 161 20087 167 20099
rect 233 20087 259 20099
rect 161 20065 199 20087
rect 233 20065 271 20087
rect 305 20065 343 20099
rect 377 20065 415 20099
rect 449 20087 459 20099
rect 521 20087 537 20099
rect 593 20087 615 20099
rect 665 20087 693 20099
rect 737 20087 771 20099
rect 877 20117 915 20143
rect 449 20065 487 20087
rect 521 20065 559 20087
rect 593 20065 631 20087
rect 665 20065 703 20087
rect 737 20065 775 20087
rect 902 20109 915 20117
rect 949 20109 983 20143
rect 902 20083 983 20109
rect -23 20048 775 20065
rect 877 20075 983 20083
rect -23 19997 -17 20048
rect 17 20031 75 20048
rect 109 20031 167 20048
rect 201 20031 259 20048
rect 293 20031 459 20048
rect 493 20031 537 20048
rect 571 20031 615 20048
rect 649 20031 693 20048
rect 727 20031 771 20048
rect 17 19997 55 20031
rect 109 20014 127 20031
rect 89 19997 127 20014
rect 161 20014 167 20031
rect 233 20014 259 20031
rect 161 19997 199 20014
rect 233 19997 271 20014
rect 305 19997 343 20031
rect 377 19997 415 20031
rect 449 20014 459 20031
rect 521 20014 537 20031
rect 593 20014 615 20031
rect 665 20014 693 20031
rect 737 20014 771 20031
rect 877 20041 915 20075
rect 949 20041 983 20075
rect 449 19997 487 20014
rect 521 19997 559 20014
rect 593 19997 631 20014
rect 665 19997 703 20014
rect 737 19997 775 20014
rect 902 20007 983 20041
rect -23 19975 775 19997
rect -23 19929 -17 19975
rect 17 19963 75 19975
rect 109 19963 167 19975
rect 201 19963 259 19975
rect 293 19963 459 19975
rect 493 19963 537 19975
rect 571 19963 615 19975
rect 649 19963 693 19975
rect 727 19963 771 19975
rect 17 19929 55 19963
rect 109 19941 127 19963
rect 89 19929 127 19941
rect 161 19941 167 19963
rect 233 19941 259 19963
rect 161 19929 199 19941
rect 233 19929 271 19941
rect 305 19929 343 19963
rect 377 19929 415 19963
rect 449 19941 459 19963
rect 521 19941 537 19963
rect 593 19941 615 19963
rect 665 19941 693 19963
rect 737 19941 771 19963
rect 877 19973 915 20007
rect 949 19973 983 20007
rect 877 19965 983 19973
rect 449 19929 487 19941
rect 521 19929 559 19941
rect 593 19929 631 19941
rect 665 19929 703 19941
rect 737 19929 775 19941
rect 902 19939 983 19965
rect 902 19931 915 19939
rect -23 19902 775 19929
rect 877 19905 915 19931
rect 949 19905 983 19939
rect -23 19861 -17 19902
rect 17 19895 75 19902
rect 109 19895 167 19902
rect 201 19895 259 19902
rect 293 19895 459 19902
rect 493 19895 537 19902
rect 571 19895 615 19902
rect 649 19895 693 19902
rect 727 19895 771 19902
rect 17 19861 55 19895
rect 109 19868 127 19895
rect 89 19861 127 19868
rect 161 19868 167 19895
rect 233 19868 259 19895
rect 161 19861 199 19868
rect 233 19861 271 19868
rect 305 19861 343 19895
rect 377 19861 415 19895
rect 449 19868 459 19895
rect 521 19868 537 19895
rect 593 19868 615 19895
rect 665 19868 693 19895
rect 737 19868 771 19895
rect 877 19889 983 19905
rect 449 19861 487 19868
rect 521 19861 559 19868
rect 593 19861 631 19868
rect 665 19861 703 19868
rect 737 19861 775 19868
rect -23 19829 775 19861
rect 902 19871 983 19889
rect 902 19855 915 19871
rect 877 19837 915 19855
rect 949 19837 983 19871
rect -23 19793 -17 19829
rect 17 19827 75 19829
rect 109 19827 167 19829
rect 201 19827 259 19829
rect 293 19827 459 19829
rect 493 19827 537 19829
rect 571 19827 615 19829
rect 649 19827 693 19829
rect 727 19827 771 19829
rect 17 19793 55 19827
rect 109 19795 127 19827
rect 89 19793 127 19795
rect 161 19795 167 19827
rect 233 19795 259 19827
rect 161 19793 199 19795
rect 233 19793 271 19795
rect 305 19793 343 19827
rect 377 19793 415 19827
rect 449 19795 459 19827
rect 521 19795 537 19827
rect 593 19795 615 19827
rect 665 19795 693 19827
rect 737 19795 771 19827
rect 877 19813 983 19837
rect 449 19793 487 19795
rect 521 19793 559 19795
rect 593 19793 631 19795
rect 665 19793 703 19795
rect 737 19793 775 19795
rect -23 19759 775 19793
rect 902 19803 983 19813
rect 902 19779 915 19803
rect -23 19722 -17 19759
rect 17 19725 55 19759
rect 89 19756 127 19759
rect 109 19725 127 19756
rect 161 19756 199 19759
rect 233 19756 271 19759
rect 161 19725 167 19756
rect 233 19725 259 19756
rect 305 19725 343 19759
rect 377 19725 415 19759
rect 449 19756 487 19759
rect 521 19756 559 19759
rect 593 19756 631 19759
rect 665 19756 703 19759
rect 737 19756 775 19759
rect 877 19769 915 19779
rect 949 19769 983 19803
rect 449 19725 459 19756
rect 521 19725 537 19756
rect 593 19725 615 19756
rect 665 19725 693 19756
rect 737 19725 771 19756
rect 17 19722 75 19725
rect 109 19722 167 19725
rect 201 19722 259 19725
rect 293 19722 459 19725
rect 493 19722 537 19725
rect 571 19722 615 19725
rect 649 19722 693 19725
rect 727 19722 771 19725
rect 877 19737 983 19769
rect -23 19691 775 19722
rect 902 19735 983 19737
rect 902 19703 915 19735
rect -23 19649 -17 19691
rect 17 19657 55 19691
rect 89 19683 127 19691
rect 109 19657 127 19683
rect 161 19683 199 19691
rect 233 19683 271 19691
rect 161 19657 167 19683
rect 233 19657 259 19683
rect 305 19657 343 19691
rect 377 19657 415 19691
rect 449 19683 487 19691
rect 521 19683 559 19691
rect 593 19683 631 19691
rect 665 19683 703 19691
rect 737 19683 775 19691
rect 877 19701 915 19703
rect 949 19701 983 19735
rect 449 19657 459 19683
rect 521 19657 537 19683
rect 593 19657 615 19683
rect 665 19657 693 19683
rect 737 19657 771 19683
rect 17 19649 75 19657
rect 109 19649 167 19657
rect 201 19649 259 19657
rect 293 19649 459 19657
rect 493 19649 537 19657
rect 571 19649 615 19657
rect 649 19649 693 19657
rect 727 19649 771 19657
rect 877 19667 983 19701
rect 877 19661 915 19667
rect -23 19623 775 19649
rect 902 19633 915 19661
rect 949 19633 983 19667
rect 902 19627 983 19633
rect -23 19576 -17 19623
rect 17 19589 55 19623
rect 89 19610 127 19623
rect 109 19589 127 19610
rect 161 19610 199 19623
rect 233 19610 271 19623
rect 161 19589 167 19610
rect 233 19589 259 19610
rect 305 19589 343 19623
rect 377 19589 415 19623
rect 449 19610 487 19623
rect 521 19610 559 19623
rect 593 19610 631 19623
rect 665 19610 703 19623
rect 737 19610 775 19623
rect 449 19589 459 19610
rect 521 19589 537 19610
rect 593 19589 615 19610
rect 665 19589 693 19610
rect 737 19589 771 19610
rect 17 19576 75 19589
rect 109 19576 167 19589
rect 201 19576 259 19589
rect 293 19576 459 19589
rect 493 19576 537 19589
rect 571 19576 615 19589
rect 649 19576 693 19589
rect 727 19576 771 19589
rect 877 19599 983 19627
rect 877 19585 915 19599
rect -23 19555 775 19576
rect -23 19503 -17 19555
rect 17 19521 55 19555
rect 89 19537 127 19555
rect 109 19521 127 19537
rect 161 19537 199 19555
rect 233 19537 271 19555
rect 161 19521 167 19537
rect 233 19521 259 19537
rect 305 19521 343 19555
rect 377 19521 415 19555
rect 449 19537 487 19555
rect 521 19537 559 19555
rect 593 19537 631 19555
rect 665 19537 703 19555
rect 737 19537 775 19555
rect 902 19565 915 19585
rect 949 19565 983 19599
rect 902 19551 983 19565
rect 449 19521 459 19537
rect 521 19521 537 19537
rect 593 19521 615 19537
rect 665 19521 693 19537
rect 737 19521 771 19537
rect 17 19503 75 19521
rect 109 19503 167 19521
rect 201 19503 259 19521
rect 293 19503 459 19521
rect 493 19503 537 19521
rect 571 19503 615 19521
rect 649 19503 693 19521
rect 727 19503 771 19521
rect 877 19531 983 19551
rect 877 19509 915 19531
rect -23 19487 775 19503
rect -23 19430 -17 19487
rect 17 19453 55 19487
rect 89 19464 127 19487
rect 109 19453 127 19464
rect 161 19464 199 19487
rect 233 19464 271 19487
rect 161 19453 167 19464
rect 233 19453 259 19464
rect 305 19453 343 19487
rect 377 19453 415 19487
rect 449 19464 487 19487
rect 521 19464 559 19487
rect 593 19464 631 19487
rect 665 19464 703 19487
rect 737 19464 775 19487
rect 902 19497 915 19509
rect 949 19497 983 19531
rect 902 19475 983 19497
rect 449 19453 459 19464
rect 521 19453 537 19464
rect 593 19453 615 19464
rect 665 19453 693 19464
rect 737 19453 771 19464
rect 17 19430 75 19453
rect 109 19430 167 19453
rect 201 19430 259 19453
rect 293 19430 459 19453
rect 493 19430 537 19453
rect 571 19430 615 19453
rect 649 19430 693 19453
rect 727 19430 771 19453
rect 877 19463 983 19475
rect 877 19433 915 19463
rect -23 19419 775 19430
rect -23 19357 -17 19419
rect 17 19385 55 19419
rect 89 19391 127 19419
rect 109 19385 127 19391
rect 161 19391 199 19419
rect 233 19391 271 19419
rect 161 19385 167 19391
rect 233 19385 259 19391
rect 305 19385 343 19419
rect 377 19385 415 19419
rect 449 19391 487 19419
rect 521 19391 559 19419
rect 593 19391 631 19419
rect 665 19391 703 19419
rect 737 19391 775 19419
rect 902 19429 915 19433
rect 949 19429 983 19463
rect 902 19399 983 19429
rect 877 19395 983 19399
rect 449 19385 459 19391
rect 521 19385 537 19391
rect 593 19385 615 19391
rect 665 19385 693 19391
rect 737 19385 771 19391
rect 17 19357 75 19385
rect 109 19357 167 19385
rect 201 19357 259 19385
rect 293 19357 459 19385
rect 493 19357 537 19385
rect 571 19357 615 19385
rect 649 19357 693 19385
rect 727 19357 771 19385
rect 877 19361 915 19395
rect 949 19361 983 19395
rect 877 19357 983 19361
rect -23 19351 775 19357
rect -23 19284 -17 19351
rect 17 19317 55 19351
rect 89 19318 127 19351
rect 109 19317 127 19318
rect 161 19318 199 19351
rect 233 19318 271 19351
rect 161 19317 167 19318
rect 233 19317 259 19318
rect 305 19317 343 19351
rect 377 19317 415 19351
rect 449 19318 487 19351
rect 521 19318 559 19351
rect 593 19318 631 19351
rect 665 19318 703 19351
rect 737 19318 775 19351
rect 902 19327 983 19357
rect 902 19323 915 19327
rect 449 19317 459 19318
rect 521 19317 537 19318
rect 593 19317 615 19318
rect 665 19317 693 19318
rect 737 19317 771 19318
rect 17 19284 75 19317
rect 109 19284 167 19317
rect 201 19284 259 19317
rect 293 19284 459 19317
rect 493 19284 537 19317
rect 571 19284 615 19317
rect 649 19284 693 19317
rect 727 19284 771 19317
rect 877 19293 915 19323
rect 949 19293 983 19327
rect -23 19283 775 19284
rect -23 19249 -17 19283
rect 17 19249 55 19283
rect 89 19249 127 19283
rect 161 19249 199 19283
rect 233 19249 271 19283
rect 305 19249 343 19283
rect 377 19249 415 19283
rect 449 19249 487 19283
rect 521 19249 559 19283
rect 593 19249 631 19283
rect 665 19249 703 19283
rect 737 19249 775 19283
rect 877 19281 983 19293
rect -23 19245 775 19249
rect 902 19259 983 19281
rect 902 19247 915 19259
rect -23 19181 -17 19245
rect 17 19215 75 19245
rect 109 19215 167 19245
rect 201 19215 259 19245
rect 293 19215 459 19245
rect 493 19215 537 19245
rect 571 19215 615 19245
rect 649 19215 693 19245
rect 727 19215 771 19245
rect 17 19181 55 19215
rect 109 19211 127 19215
rect 89 19181 127 19211
rect 161 19211 167 19215
rect 233 19211 259 19215
rect 161 19181 199 19211
rect 233 19181 271 19211
rect 305 19181 343 19215
rect 377 19181 415 19215
rect 449 19211 459 19215
rect 521 19211 537 19215
rect 593 19211 615 19215
rect 665 19211 693 19215
rect 737 19211 771 19215
rect 877 19225 915 19247
rect 949 19225 983 19259
rect 449 19181 487 19211
rect 521 19181 559 19211
rect 593 19181 631 19211
rect 665 19181 703 19211
rect 737 19181 775 19211
rect -23 19179 775 19181
rect -17 19153 775 19179
rect 877 19191 983 19225
rect 7937 19191 9142 19221
rect 877 19153 915 19191
rect 949 19157 9142 19191
rect 1017 19153 1058 19157
rect 1092 19153 1133 19157
rect 1167 19153 1208 19157
rect 1242 19153 1283 19157
rect 1317 19153 1358 19157
rect 1392 19153 1433 19157
rect 1467 19153 1508 19157
rect 1542 19153 1583 19157
rect 1617 19153 1658 19157
rect 1692 19153 9142 19157
rect -17 19147 472 19153
rect 506 19147 545 19153
rect 579 19147 618 19153
rect 652 19147 691 19153
rect 725 19147 764 19153
rect 17 19113 55 19147
rect 89 19113 127 19147
rect 161 19113 199 19147
rect 233 19113 271 19147
rect 305 19113 343 19147
rect 377 19113 415 19147
rect 449 19119 472 19147
rect 521 19119 545 19147
rect 593 19119 618 19147
rect 665 19119 691 19147
rect 737 19119 764 19147
rect 877 19119 910 19153
rect 1017 19119 1056 19153
rect 1092 19123 1129 19153
rect 1167 19123 1202 19153
rect 1242 19123 1275 19153
rect 1317 19123 1348 19153
rect 1392 19123 1420 19153
rect 1467 19123 1492 19153
rect 1542 19123 1564 19153
rect 1617 19123 1636 19153
rect 1692 19123 1708 19153
rect 1090 19119 1129 19123
rect 1163 19119 1202 19123
rect 1236 19119 1275 19123
rect 1309 19119 1348 19123
rect 1382 19119 1420 19123
rect 1454 19119 1492 19123
rect 1526 19119 1564 19123
rect 1598 19119 1636 19123
rect 1670 19119 1708 19123
rect 1763 19138 9142 19153
rect 1763 19119 1800 19138
rect 449 19113 487 19119
rect 521 19113 559 19119
rect 593 19113 631 19119
rect 665 19113 703 19119
rect 737 19113 775 19119
rect -17 19079 775 19113
rect 17 19045 55 19079
rect 89 19045 127 19079
rect 161 19045 199 19079
rect 233 19045 271 19079
rect 305 19045 343 19079
rect 377 19045 415 19079
rect 449 19063 487 19079
rect 521 19063 559 19079
rect 593 19063 631 19079
rect 665 19063 703 19079
rect 737 19063 775 19079
rect 877 19063 915 19119
rect 1017 19104 1800 19119
rect 1834 19104 1869 19138
rect 1903 19104 1938 19138
rect 1972 19104 2007 19138
rect 2041 19104 2076 19138
rect 2110 19104 2145 19138
rect 2179 19104 2214 19138
rect 2248 19104 2283 19138
rect 2317 19104 2352 19138
rect 2386 19104 2421 19138
rect 2455 19104 2490 19138
rect 2524 19104 2559 19138
rect 2593 19104 2628 19138
rect 2662 19104 2697 19138
rect 2731 19104 2766 19138
rect 2800 19104 2835 19138
rect 2869 19104 2904 19138
rect 2938 19104 2973 19138
rect 3007 19104 3042 19138
rect 3076 19104 3111 19138
rect 3145 19104 3180 19138
rect 3214 19104 3249 19138
rect 3283 19104 3318 19138
rect 3352 19104 3387 19138
rect 3421 19104 3456 19138
rect 3490 19104 3525 19138
rect 3559 19104 3594 19138
rect 3628 19104 3663 19138
rect 3697 19104 3732 19138
rect 3766 19104 3801 19138
rect 3835 19104 3870 19138
rect 3904 19104 3939 19138
rect 3973 19104 4008 19138
rect 4042 19104 4076 19138
rect 4110 19104 4144 19138
rect 4178 19104 4212 19138
rect 4246 19104 4280 19138
rect 4314 19104 4348 19138
rect 4382 19104 4416 19138
rect 4450 19104 4484 19138
rect 4518 19104 4552 19138
rect 4586 19104 4620 19138
rect 4654 19104 4688 19138
rect 4722 19104 4756 19138
rect 4790 19104 4824 19138
rect 4858 19104 4892 19138
rect 4926 19104 4960 19138
rect 4994 19104 5028 19138
rect 5062 19104 5096 19138
rect 5130 19104 5164 19138
rect 5198 19104 5232 19138
rect 5266 19104 5300 19138
rect 5334 19104 5368 19138
rect 5402 19104 5436 19138
rect 5470 19104 5504 19138
rect 5538 19104 5572 19138
rect 5606 19104 5640 19138
rect 5674 19104 5708 19138
rect 5742 19104 5776 19138
rect 5810 19104 5844 19138
rect 5878 19104 5912 19138
rect 5946 19104 5980 19138
rect 6014 19104 6048 19138
rect 6082 19104 6116 19138
rect 6150 19104 6184 19138
rect 6218 19104 6252 19138
rect 6286 19104 6320 19138
rect 6354 19104 6388 19138
rect 6422 19104 6456 19138
rect 6490 19104 6524 19138
rect 6558 19104 6592 19138
rect 6626 19104 6660 19138
rect 6694 19104 6728 19138
rect 6762 19104 6796 19138
rect 6830 19104 6864 19138
rect 6898 19104 6932 19138
rect 6966 19104 7000 19138
rect 7034 19104 7068 19138
rect 7102 19104 7136 19138
rect 7170 19104 7204 19138
rect 7238 19104 7272 19138
rect 7306 19104 7340 19138
rect 7374 19104 7408 19138
rect 7442 19104 7476 19138
rect 7510 19104 7544 19138
rect 7578 19104 7612 19138
rect 7646 19104 7680 19138
rect 7714 19104 7748 19138
rect 7782 19104 7816 19138
rect 7850 19104 7884 19138
rect 7918 19104 7952 19138
rect 7986 19104 8020 19138
rect 8054 19104 8088 19138
rect 8122 19104 8156 19138
rect 8190 19104 8224 19138
rect 8258 19104 8292 19138
rect 8326 19104 8360 19138
rect 8394 19104 8428 19138
rect 8462 19104 8496 19138
rect 8530 19104 8564 19138
rect 8598 19104 8632 19138
rect 8666 19104 8700 19138
rect 8734 19104 8768 19138
rect 8802 19104 8836 19138
rect 8870 19104 8904 19138
rect 8938 19104 8972 19138
rect 9006 19104 9040 19138
rect 9074 19104 9108 19138
rect 1017 19089 9142 19104
rect 1017 19063 1058 19089
rect 1092 19063 1133 19089
rect 1167 19063 1208 19089
rect 1242 19063 1283 19089
rect 1317 19063 1358 19089
rect 1392 19063 1433 19089
rect 1467 19063 1508 19089
rect 1542 19063 1583 19089
rect 1617 19063 1658 19089
rect 1692 19081 9142 19089
rect 1692 19063 1729 19081
rect 449 19045 472 19063
rect 521 19045 545 19063
rect 593 19045 618 19063
rect 665 19045 691 19063
rect 737 19045 764 19063
rect -17 19029 472 19045
rect 506 19029 545 19045
rect 579 19029 618 19045
rect 652 19029 691 19045
rect 725 19029 764 19045
rect 877 19029 910 19063
rect 1017 19029 1056 19063
rect 1092 19055 1129 19063
rect 1167 19055 1202 19063
rect 1242 19055 1275 19063
rect 1317 19055 1348 19063
rect 1392 19055 1420 19063
rect 1467 19055 1492 19063
rect 1542 19055 1564 19063
rect 1617 19055 1636 19063
rect 1692 19055 1708 19063
rect 1090 19029 1129 19055
rect 1163 19029 1202 19055
rect 1236 19029 1275 19055
rect 1309 19029 1348 19055
rect 1382 19029 1420 19055
rect 1454 19029 1492 19055
rect 1526 19029 1564 19055
rect 1598 19029 1636 19055
rect 1670 19029 1708 19055
rect 1763 19051 9142 19081
rect 1763 19047 1800 19051
rect 1742 19029 1800 19047
rect -17 19011 775 19029
rect 17 18977 55 19011
rect 89 18977 127 19011
rect 161 18977 199 19011
rect 233 18977 271 19011
rect 305 18977 343 19011
rect 377 18977 415 19011
rect 449 18977 487 19011
rect 521 18977 559 19011
rect 593 18977 631 19011
rect 665 18977 703 19011
rect 737 18977 775 19011
rect -17 18943 775 18977
rect 17 18909 55 18943
rect 89 18909 127 18943
rect 161 18909 199 18943
rect 233 18909 271 18943
rect 305 18909 343 18943
rect 377 18909 415 18943
rect 449 18909 487 18943
rect 521 18909 559 18943
rect 593 18909 631 18943
rect 665 18909 703 18943
rect 737 18909 775 18943
rect -17 18875 775 18909
rect 17 18841 55 18875
rect 89 18841 127 18875
rect 161 18841 199 18875
rect 233 18841 271 18875
rect 305 18841 343 18875
rect 377 18841 415 18875
rect 449 18841 487 18875
rect 521 18841 559 18875
rect 593 18841 631 18875
rect 665 18841 703 18875
rect 737 18841 775 18875
rect -17 18807 775 18841
rect 17 18773 55 18807
rect 89 18773 127 18807
rect 161 18773 199 18807
rect 233 18773 271 18807
rect 305 18773 343 18807
rect 377 18773 415 18807
rect 449 18773 487 18807
rect 521 18773 559 18807
rect 593 18773 631 18807
rect 665 18773 703 18807
rect 737 18773 775 18807
rect -17 18739 775 18773
rect 17 18705 55 18739
rect 89 18705 127 18739
rect 161 18705 199 18739
rect 233 18705 271 18739
rect 305 18705 343 18739
rect 377 18705 415 18739
rect 449 18705 487 18739
rect 521 18705 559 18739
rect 593 18705 631 18739
rect 665 18705 703 18739
rect 737 18705 775 18739
rect -17 18671 775 18705
rect 17 18637 55 18671
rect 89 18637 127 18671
rect 161 18637 199 18671
rect 233 18637 271 18671
rect 305 18637 343 18671
rect 377 18637 415 18671
rect 449 18637 487 18671
rect 521 18637 559 18671
rect 593 18637 631 18671
rect 665 18637 703 18671
rect 737 18637 775 18671
rect -17 18613 843 18637
rect 877 18613 915 19029
rect 1017 19021 1800 19029
rect 5772 19025 9142 19051
rect 1017 18987 1058 19021
rect 1092 18987 1133 19021
rect 1167 18987 1208 19021
rect 1242 18987 1283 19021
rect 1317 18987 1358 19021
rect 1392 18987 1433 19021
rect 1467 18987 1508 19021
rect 1542 18987 1583 19021
rect 1617 18987 1658 19021
rect 1692 19009 1800 19021
rect 1692 18987 1729 19009
rect 1017 18975 1729 18987
rect 1763 18975 1800 19009
rect 1017 18953 1800 18975
rect 1017 18919 1058 18953
rect 1092 18919 1133 18953
rect 1167 18919 1208 18953
rect 1242 18919 1283 18953
rect 1317 18919 1358 18953
rect 1392 18919 1433 18953
rect 1467 18919 1508 18953
rect 1542 18919 1583 18953
rect 1617 18919 1658 18953
rect 1692 18937 1800 18953
rect 1692 18919 1729 18937
rect 1017 18903 1729 18919
rect 1763 18903 1800 18937
rect 1017 18885 1800 18903
rect 1017 18851 1058 18885
rect 1092 18851 1133 18885
rect 1167 18851 1208 18885
rect 1242 18851 1283 18885
rect 1317 18851 1358 18885
rect 1392 18851 1433 18885
rect 1467 18851 1508 18885
rect 1542 18851 1583 18885
rect 1617 18851 1658 18885
rect 1692 18865 1800 18885
rect 1692 18851 1729 18865
rect 1017 18831 1729 18851
rect 1763 18831 1800 18865
rect 1017 18817 1800 18831
rect 1017 18783 1058 18817
rect 1092 18783 1133 18817
rect 1167 18783 1208 18817
rect 1242 18783 1283 18817
rect 1317 18783 1358 18817
rect 1392 18783 1433 18817
rect 1467 18783 1508 18817
rect 1542 18783 1583 18817
rect 1617 18783 1658 18817
rect 1692 18793 1800 18817
rect 1692 18783 1729 18793
rect 1017 18759 1729 18783
rect 1763 18759 1800 18793
rect 1017 18749 1800 18759
rect 1017 18715 1058 18749
rect 1092 18715 1133 18749
rect 1167 18715 1208 18749
rect 1242 18715 1283 18749
rect 1317 18715 1358 18749
rect 1392 18715 1433 18749
rect 1467 18715 1508 18749
rect 1542 18715 1583 18749
rect 1617 18715 1658 18749
rect 1692 18720 1800 18749
rect 1692 18715 1729 18720
rect 1017 18686 1729 18715
rect 1763 18686 1800 18720
rect 1017 18681 1800 18686
rect 1017 18647 1058 18681
rect 1092 18647 1133 18681
rect 1167 18647 1208 18681
rect 1242 18647 1283 18681
rect 1317 18647 1358 18681
rect 1392 18647 1433 18681
rect 1467 18647 1508 18681
rect 1542 18647 1583 18681
rect 1617 18647 1658 18681
rect 1692 18647 1800 18681
rect 949 18613 1729 18647
rect 1763 18613 1800 18647
rect 1298 18577 1800 18613
rect 1298 18543 1332 18577
rect 1366 18543 1412 18577
rect 1446 18543 1492 18577
rect 1526 18543 1572 18577
rect 1606 18543 1652 18577
rect 1686 18543 1732 18577
rect 1766 18543 1800 18577
rect 1298 18509 1800 18543
rect 1298 18475 1332 18509
rect 1366 18475 1412 18509
rect 1446 18475 1492 18509
rect 1526 18475 1572 18509
rect 1606 18475 1652 18509
rect 1686 18475 1732 18509
rect 1766 18475 1800 18509
rect 1298 18441 1800 18475
rect 1298 18407 1332 18441
rect 1366 18407 1412 18441
rect 1446 18407 1492 18441
rect 1526 18407 1572 18441
rect 1606 18407 1652 18441
rect 1686 18407 1732 18441
rect 1766 18407 1800 18441
rect 1298 18373 1800 18407
rect 1298 18339 1332 18373
rect 1366 18339 1412 18373
rect 1446 18339 1492 18373
rect 1526 18339 1572 18373
rect 1606 18339 1652 18373
rect 1686 18339 1732 18373
rect 1766 18339 1800 18373
rect 1298 18305 1800 18339
rect 1298 18271 1332 18305
rect 1366 18271 1412 18305
rect 1446 18271 1492 18305
rect 1526 18271 1572 18305
rect 1606 18271 1652 18305
rect 1686 18271 1732 18305
rect 1766 18271 1800 18305
rect 1298 18237 1800 18271
rect 1298 18203 1332 18237
rect 1366 18203 1412 18237
rect 1446 18203 1492 18237
rect 1526 18203 1572 18237
rect 1606 18203 1652 18237
rect 1686 18203 1732 18237
rect 1766 18203 1800 18237
rect 1298 18169 1800 18203
rect 1298 18135 1332 18169
rect 1366 18135 1412 18169
rect 1446 18135 1492 18169
rect 1526 18135 1572 18169
rect 1606 18158 1652 18169
rect 1686 18158 1732 18169
rect 1766 18135 1800 18169
rect 1298 18100 1584 18135
rect 1762 18100 1800 18135
rect 1298 18066 1332 18100
rect 1366 18066 1412 18100
rect 1446 18066 1492 18100
rect 1526 18066 1572 18100
rect 1766 18066 1800 18100
rect 1298 18031 1584 18066
rect 1762 18031 1800 18066
rect 1298 17997 1332 18031
rect 1366 17997 1412 18031
rect 1446 17997 1492 18031
rect 1526 17997 1572 18031
rect 1766 17997 1800 18031
rect 1298 17962 1584 17997
rect 1762 17962 1800 17997
rect 1298 17928 1332 17962
rect 1366 17928 1412 17962
rect 1446 17928 1492 17962
rect 1526 17928 1572 17962
rect 1766 17928 1800 17962
rect 1298 17908 1584 17928
rect 1762 17908 1800 17928
rect 1298 17893 1800 17908
rect 1298 17859 1332 17893
rect 1366 17859 1412 17893
rect 1446 17859 1492 17893
rect 1526 17859 1572 17893
rect 1606 17869 1652 17893
rect 1686 17869 1732 17893
rect 1618 17859 1652 17869
rect 1298 17835 1584 17859
rect 1618 17835 1656 17859
rect 1690 17835 1728 17869
rect 1766 17859 1800 17893
rect 1762 17835 1800 17859
rect 1298 17824 1800 17835
rect 1298 17790 1332 17824
rect 1366 17790 1412 17824
rect 1446 17790 1492 17824
rect 1526 17790 1572 17824
rect 1606 17790 1652 17824
rect 1686 17790 1732 17824
rect 1766 17790 1800 17824
rect 5569 13855 5608 13889
rect 5642 13855 5681 13889
rect 5715 13855 5754 13889
rect 5788 13855 5827 13889
rect 5861 13855 5900 13889
rect 5535 13781 5934 13855
rect 5569 13747 5608 13781
rect 5642 13747 5681 13781
rect 5715 13747 5754 13781
rect 5788 13747 5827 13781
rect 5861 13747 5900 13781
rect 5339 13529 5380 13563
rect 5414 13529 5455 13563
rect 5489 13529 5530 13563
rect 5564 13529 5604 13563
rect 5638 13529 5678 13563
rect 5712 13529 5752 13563
rect 5786 13529 5826 13563
rect 5860 13529 5900 13563
rect 5305 13455 5934 13529
rect 5339 13421 5380 13455
rect 5414 13421 5455 13455
rect 5489 13421 5530 13455
rect 5564 13421 5604 13455
rect 5638 13421 5678 13455
rect 5712 13421 5752 13455
rect 5786 13421 5826 13455
rect 5860 13421 5900 13455
rect 5532 12876 5581 12910
rect 5615 12876 5664 12910
rect 5698 12876 5747 12910
rect 5781 12876 5829 12910
rect 5498 12828 5863 12876
rect 5532 12794 5581 12828
rect 5615 12794 5664 12828
rect 5698 12794 5747 12828
rect 5781 12794 5829 12828
rect 5220 11991 5266 12025
rect 5300 11991 5346 12025
rect 5380 11991 5426 12025
rect 5460 11991 5506 12025
rect 5540 11991 5586 12025
rect 5186 11939 5620 11991
rect 5220 11905 5266 11939
rect 5300 11905 5346 11939
rect 5380 11905 5426 11939
rect 5460 11905 5506 11939
rect 5540 11905 5586 11939
rect 5186 11853 5620 11905
rect 5220 11819 5266 11853
rect 5300 11819 5346 11853
rect 5380 11819 5426 11853
rect 5460 11819 5506 11853
rect 5540 11819 5586 11853
rect 5668 11870 5702 11908
rect 5221 11739 5260 11773
rect 5294 11739 5333 11773
rect 5367 11739 5406 11773
rect 5440 11739 5479 11773
rect 5513 11739 5552 11773
rect 5586 11739 5624 11773
rect 5658 11739 5696 11773
rect 5730 11739 5768 11773
rect 5802 11739 5840 11773
rect 5187 11699 5874 11739
rect 5221 11665 5260 11699
rect 5294 11665 5333 11699
rect 5367 11665 5406 11699
rect 5440 11665 5479 11699
rect 5513 11665 5552 11699
rect 5586 11665 5624 11699
rect 5658 11665 5696 11699
rect 5730 11665 5768 11699
rect 5802 11665 5840 11699
rect 5187 11625 5874 11665
rect 5221 11591 5260 11625
rect 5294 11591 5333 11625
rect 5367 11591 5406 11625
rect 5440 11591 5479 11625
rect 5513 11591 5552 11625
rect 5586 11591 5624 11625
rect 5658 11591 5696 11625
rect 5730 11591 5768 11625
rect 5802 11591 5840 11625
rect 5187 11551 5874 11591
rect 5221 11517 5260 11551
rect 5294 11517 5333 11551
rect 5367 11517 5406 11551
rect 5440 11517 5479 11551
rect 5513 11517 5552 11551
rect 5586 11517 5624 11551
rect 5658 11517 5696 11551
rect 5730 11517 5768 11551
rect 5802 11517 5840 11551
rect 338 9109 359 9143
rect 396 9109 433 9143
rect 477 9109 504 9143
rect 561 9109 575 9143
rect 609 9109 611 9143
rect 645 9109 646 9143
rect 680 9109 694 9143
rect 751 9109 777 9143
rect 822 9109 859 9143
rect 894 9109 917 9143
rect 1860 6400 1932 7350
rect 2066 6400 2138 7350
rect 2282 6400 2333 7452
rect 2388 6222 2473 7353
rect 2522 6400 2628 7452
rect 2834 7350 2861 7452
rect 2678 6400 2784 7350
rect 2834 6400 2940 7350
rect 2991 6400 3097 7452
rect 3146 6400 3252 7350
rect 3302 6400 3390 7452
rect 3442 6400 3530 7350
rect 3628 6412 3726 7350
rect 3810 6400 3916 7350
rect 4128 6400 4234 7350
rect 4434 6400 4540 7351
rect 4745 6400 4851 7351
rect 5135 6450 5218 7400
rect 5277 6450 5373 7466
rect 5409 6450 5515 7400
rect 5566 6449 5672 7466
rect 5721 6450 5827 7401
rect 5878 6450 5984 7466
rect 6033 6450 6139 7400
rect 6190 6450 6275 7466
rect 6332 6450 6417 7401
rect 6482 6412 6614 7350
rect 6700 6398 6786 7416
rect 6861 6395 6973 7350
rect 7012 6398 7098 7416
rect 7173 6395 7285 7350
rect 7324 6398 7410 7416
rect 7485 6395 7597 7350
rect 7636 6398 7722 7416
rect 7797 6395 7909 7350
rect 7943 6398 8018 7350
rect 8116 6431 8180 7342
rect 8840 6654 8878 7302
rect 9062 7268 9272 7394
rect 15976 7133 16024 7145
rect 15976 7087 15983 7133
rect 16017 7087 16024 7133
rect 15976 7061 16024 7087
rect 15976 7018 15983 7061
rect 16017 7018 16024 7061
rect 15976 6989 16024 7018
rect 15976 6949 15983 6989
rect 16017 6949 16024 6989
rect 15976 6917 16024 6949
rect 15976 6880 15983 6917
rect 16017 6880 16024 6917
rect 15976 6845 16024 6880
rect 15976 6811 15983 6845
rect 16017 6811 16024 6845
rect 15976 6776 16024 6811
rect 15976 6739 15983 6776
rect 16017 6739 16024 6776
rect 10221 6489 10352 6738
rect 9868 6413 10352 6489
rect 15976 6707 16024 6739
rect 15976 6667 15983 6707
rect 16017 6667 16024 6707
rect 15976 6638 16024 6667
rect 15976 6595 15983 6638
rect 16017 6595 16024 6638
rect 15976 6569 16024 6595
rect 15976 6523 15983 6569
rect 16017 6523 16024 6569
rect 15976 6500 16024 6523
rect 15976 6451 15983 6500
rect 16017 6451 16024 6500
rect 15976 6431 16024 6451
rect 15976 6379 15983 6431
rect 16017 6379 16024 6431
rect 15976 6361 16024 6379
rect 15976 6307 15983 6361
rect 16017 6307 16024 6361
rect 15976 6291 16024 6307
rect 15976 6235 15983 6291
rect 16017 6235 16024 6291
rect 15976 6221 16024 6235
rect 15976 6163 15983 6221
rect 16017 6163 16024 6221
rect 15976 6151 16024 6163
rect 15976 6091 15983 6151
rect 16017 6091 16024 6151
rect 15976 6081 16024 6091
rect 2864 5914 2898 6022
rect 2864 5894 2934 5914
rect 2864 5352 2900 5894
rect 3021 5352 3127 5938
rect 3177 5352 3283 5894
rect 3334 5352 3440 5938
rect 3607 5352 3690 5894
rect 3808 5352 3891 5894
rect 3958 5352 4064 5894
rect 4338 5352 4426 5894
rect 4760 5352 4832 5894
rect 4868 5181 4967 5938
rect 5003 5352 5109 5894
rect 5278 5352 5350 5938
rect 5502 5298 5618 6072
rect 15976 6047 15983 6081
rect 16017 6047 16024 6081
rect 15976 6023 16024 6047
rect 7174 5377 7261 5647
rect 7854 5377 7938 5647
rect 4868 5116 5266 5181
rect 8676 4970 8774 5512
rect 10410 4971 10516 5513
rect 10694 4971 10800 5513
rect 10974 4971 11080 5513
rect 15976 4991 16024 5003
rect 15976 4945 15983 4991
rect 16017 4945 16024 4991
rect 15976 4919 16024 4945
rect 15976 4877 15983 4919
rect 16017 4877 16024 4919
rect 224 4465 262 4499
rect 196 4293 262 4327
rect 230 4121 262 4155
rect 230 3949 262 3983
rect 5245 3919 5334 4875
rect 5395 3920 5484 4873
rect 15976 4847 16024 4877
rect 15976 4809 15983 4847
rect 16017 4809 16024 4847
rect 15976 4775 16024 4809
rect 190 3777 262 3811
rect 5736 3799 5842 4750
rect 5878 3793 6016 4749
rect 6054 3799 6160 4749
rect 6364 3799 6470 4749
rect 15976 4741 15983 4775
rect 16017 4741 16024 4775
rect 15976 4707 16024 4741
rect 15976 4669 15983 4707
rect 16017 4669 16024 4707
rect 15976 4639 16024 4669
rect 15976 4597 15983 4639
rect 16017 4597 16024 4639
rect 15976 4571 16024 4597
rect 15976 4525 15983 4571
rect 16017 4525 16024 4571
rect 15976 4503 16024 4525
rect 15976 4453 15983 4503
rect 16017 4453 16024 4503
rect 15976 4435 16024 4453
rect 15976 4381 15983 4435
rect 16017 4381 16024 4435
rect 15976 4367 16024 4381
rect 15976 4309 15983 4367
rect 16017 4309 16024 4367
rect 15976 4299 16024 4309
rect 15976 4237 15983 4299
rect 16017 4237 16024 4299
rect 15976 4231 16024 4237
rect 15976 4165 15983 4231
rect 16017 4165 16024 4231
rect 15976 4162 16024 4165
rect 15976 4128 15983 4162
rect 16017 4128 16024 4162
rect 15976 4127 16024 4128
rect 15976 4059 15983 4127
rect 16017 4059 16024 4127
rect 15976 4055 16024 4059
rect 15976 3990 15983 4055
rect 16017 3990 16024 4055
rect 15976 3983 16024 3990
rect 15976 3921 15983 3983
rect 16017 3921 16024 3983
rect 15976 3897 16024 3921
rect 13933 2251 14330 2285
rect 13967 2217 14006 2251
rect 14040 2217 14079 2251
rect 14113 2217 14152 2251
rect 14186 2217 14224 2251
rect 14258 2217 14296 2251
rect 13933 2173 14330 2217
rect 13967 2139 14006 2173
rect 14040 2139 14079 2173
rect 14113 2139 14152 2173
rect 14186 2139 14224 2173
rect 14258 2139 14296 2173
rect 13933 2095 14330 2139
rect 13967 2068 14006 2095
rect 14040 2068 14079 2095
rect 13983 2061 14006 2068
rect 14065 2061 14079 2068
rect 14113 2068 14152 2095
rect 13933 2037 13949 2061
rect 13278 2003 13312 2037
rect 13346 2003 13382 2037
rect 13416 2003 13451 2037
rect 13485 2003 13520 2037
rect 13554 2003 13589 2037
rect 13623 2003 13658 2037
rect 13692 2003 13727 2037
rect 13761 2024 13796 2037
rect 13830 2024 13865 2037
rect 13899 2034 13949 2037
rect 13983 2034 14031 2061
rect 14065 2034 14113 2061
rect 14147 2061 14152 2068
rect 14186 2068 14224 2095
rect 14258 2068 14296 2095
rect 14186 2061 14195 2068
rect 14258 2061 14277 2068
rect 14147 2034 14195 2061
rect 14229 2034 14277 2061
rect 14311 2034 14330 2061
rect 13761 2003 13782 2024
rect 13830 2003 13854 2024
rect 13899 2017 14330 2034
rect 13899 2003 13933 2017
rect 13278 1990 13782 2003
rect 13816 1990 13854 2003
rect 13888 1990 13933 2003
rect 13278 1983 13933 1990
rect 13967 1983 14006 2017
rect 14040 1983 14079 2017
rect 14113 1983 14152 2017
rect 14186 1983 14224 2017
rect 14258 1983 14296 2017
rect 13278 1949 14330 1983
rect 13278 1915 13312 1949
rect 13346 1915 13382 1949
rect 13416 1915 13451 1949
rect 13485 1915 13520 1949
rect 13563 1915 13589 1949
rect 13641 1915 13658 1949
rect 13719 1915 13727 1949
rect 13761 1915 13762 1949
rect 13830 1915 13839 1949
rect 13899 1915 13933 1949
rect 13278 1914 13420 1915
rect 13132 1880 13420 1914
rect 13132 1846 13133 1880
rect 13167 1846 13217 1880
rect 13251 1846 13301 1880
rect 13335 1873 13385 1880
rect 13335 1846 13379 1873
rect 13419 1846 13420 1880
rect 13132 1839 13379 1846
rect 13413 1839 13420 1846
rect 13132 1810 13420 1839
rect 13132 1776 13133 1810
rect 13167 1776 13217 1810
rect 13251 1776 13301 1810
rect 13335 1797 13385 1810
rect 13335 1776 13379 1797
rect 13419 1776 13420 1810
rect 13132 1763 13379 1776
rect 13413 1763 13420 1776
rect 13132 1740 13420 1763
rect 13132 1706 13133 1740
rect 13167 1706 13217 1740
rect 13251 1706 13301 1740
rect 13335 1721 13385 1740
rect 13335 1706 13379 1721
rect 13419 1706 13420 1740
rect 13132 1687 13379 1706
rect 13413 1687 13420 1706
rect 13132 1669 13420 1687
rect 13132 1635 13133 1669
rect 13167 1635 13217 1669
rect 13251 1635 13301 1669
rect 13335 1635 13385 1669
rect 13419 1635 13420 1669
rect 13132 1598 13420 1635
rect 14616 1616 14982 1766
rect 13132 1564 13133 1598
rect 13167 1564 13217 1598
rect 13251 1564 13301 1598
rect 13335 1564 13385 1598
rect 13419 1564 13420 1598
rect 15482 1564 15886 1616
rect 13132 1527 13420 1564
rect 13132 1493 13133 1527
rect 13167 1493 13217 1527
rect 13251 1493 13301 1527
rect 13335 1493 13385 1527
rect 13419 1493 13420 1527
rect 13132 1456 13420 1493
rect 13132 1422 13133 1456
rect 13167 1422 13217 1456
rect 13251 1422 13301 1456
rect 13335 1422 13385 1456
rect 13419 1422 13420 1456
rect 13132 1385 13420 1422
rect 13132 1351 13133 1385
rect 13167 1351 13217 1385
rect 13251 1351 13301 1385
rect 13335 1351 13385 1385
rect 13419 1351 13420 1385
rect 13132 1314 13420 1351
rect 1175 1188 1281 1293
rect 13132 1280 13133 1314
rect 13167 1280 13217 1314
rect 13251 1280 13301 1314
rect 13335 1280 13385 1314
rect 13419 1280 13420 1314
rect 13132 1246 13420 1280
rect 1561 1212 12298 1246
rect 12332 1212 12369 1246
rect 12403 1212 12440 1246
rect 12474 1212 12511 1246
rect 12545 1212 12582 1246
rect 12616 1212 12653 1246
rect 12687 1212 12724 1246
rect 12758 1212 12795 1246
rect 12829 1212 12866 1246
rect 12900 1212 12937 1246
rect 12971 1212 13008 1246
rect 13042 1212 13079 1246
rect 13113 1212 13150 1246
rect 13184 1212 13221 1246
rect 13255 1212 13292 1246
rect 13326 1212 13362 1246
rect 13396 1212 13420 1246
rect 1561 1180 13420 1212
rect 1595 1146 1630 1180
rect 1664 1146 1699 1180
rect 1733 1146 1768 1180
rect 1802 1146 1837 1180
rect 1871 1146 1906 1180
rect 1940 1146 1975 1180
rect 2009 1146 2044 1180
rect 2078 1146 2113 1180
rect 2147 1146 2182 1180
rect 2216 1146 2251 1180
rect 2285 1146 2320 1180
rect 2354 1146 2389 1180
rect 2423 1146 2458 1180
rect 2492 1146 2527 1180
rect 2561 1146 2596 1180
rect 2630 1146 2665 1180
rect 2699 1146 2734 1180
rect 2768 1146 2803 1180
rect 2837 1146 2872 1180
rect 2906 1146 2941 1180
rect 2975 1146 3009 1180
rect 3043 1146 3077 1180
rect 3111 1146 3145 1180
rect 3179 1146 3213 1180
rect 3247 1146 3281 1180
rect 3315 1146 3349 1180
rect 3383 1146 3417 1180
rect 3451 1146 3485 1180
rect 3519 1146 3553 1180
rect 3587 1146 3621 1180
rect 3655 1146 3689 1180
rect 3723 1146 3757 1180
rect 3791 1146 3825 1180
rect 3859 1146 3893 1180
rect 3927 1146 3961 1180
rect 3995 1146 4029 1180
rect 4063 1146 4097 1180
rect 4131 1146 4165 1180
rect 4199 1146 4233 1180
rect 4267 1146 4301 1180
rect 4335 1146 4369 1180
rect 4403 1146 4437 1180
rect 4471 1146 4505 1180
rect 4539 1146 4573 1180
rect 4607 1146 4641 1180
rect 4675 1146 4709 1180
rect 4743 1146 4777 1180
rect 4811 1146 4845 1180
rect 4879 1146 4913 1180
rect 4947 1146 4981 1180
rect 5015 1146 5049 1180
rect 5083 1146 5117 1180
rect 5151 1146 5185 1180
rect 5219 1146 5253 1180
rect 5287 1146 5321 1180
rect 5355 1146 5389 1180
rect 5423 1146 5457 1180
rect 5491 1146 5525 1180
rect 5559 1146 5593 1180
rect 5627 1146 5661 1180
rect 5695 1146 5729 1180
rect 5763 1146 5797 1180
rect 5831 1146 5865 1180
rect 5899 1146 5933 1180
rect 5967 1146 6001 1180
rect 6035 1146 6069 1180
rect 6103 1146 6137 1180
rect 6171 1146 6205 1180
rect 6239 1146 6273 1180
rect 6307 1146 6341 1180
rect 6375 1146 6409 1180
rect 6443 1146 6477 1180
rect 6511 1146 6545 1180
rect 6579 1146 6613 1180
rect 6647 1146 6681 1180
rect 6715 1146 6749 1180
rect 6783 1146 6817 1180
rect 6851 1146 6885 1180
rect 6919 1146 6953 1180
rect 6987 1146 7021 1180
rect 7055 1146 7089 1180
rect 7123 1146 7157 1180
rect 7191 1146 7225 1180
rect 7259 1146 7293 1180
rect 7327 1146 7361 1180
rect 7395 1146 7429 1180
rect 7463 1146 7497 1180
rect 7531 1146 7565 1180
rect 7599 1146 7633 1180
rect 7667 1146 7701 1180
rect 7735 1146 7769 1180
rect 7803 1146 7837 1180
rect 7871 1146 7905 1180
rect 7939 1146 7973 1180
rect 8007 1146 8041 1180
rect 8075 1146 8109 1180
rect 8143 1146 8177 1180
rect 8211 1146 8245 1180
rect 8279 1146 8313 1180
rect 8347 1146 8381 1180
rect 8415 1146 8449 1180
rect 8483 1146 8517 1180
rect 8551 1146 8585 1180
rect 8619 1146 8653 1180
rect 8687 1146 8721 1180
rect 8755 1146 8789 1180
rect 8823 1146 8857 1180
rect 8891 1146 8925 1180
rect 8959 1146 8993 1180
rect 9027 1146 9061 1180
rect 9095 1146 9129 1180
rect 9163 1146 9197 1180
rect 9231 1146 9265 1180
rect 9299 1146 9333 1180
rect 9367 1146 9401 1180
rect 9435 1146 9469 1180
rect 9503 1146 9537 1180
rect 9571 1146 9605 1180
rect 9639 1146 9673 1180
rect 9707 1146 9741 1180
rect 9775 1146 9809 1180
rect 9843 1146 9877 1180
rect 9911 1146 9945 1180
rect 9979 1146 10013 1180
rect 10047 1146 10081 1180
rect 10115 1146 10149 1180
rect 10183 1146 10217 1180
rect 10251 1146 10285 1180
rect 10319 1146 10353 1180
rect 10387 1146 10421 1180
rect 10455 1146 10489 1180
rect 10523 1146 10557 1180
rect 10591 1146 10625 1180
rect 10659 1146 10693 1180
rect 10727 1146 10761 1180
rect 10795 1146 10829 1180
rect 10863 1146 10897 1180
rect 10931 1146 10965 1180
rect 10999 1146 11033 1180
rect 11067 1146 11101 1180
rect 11135 1146 11169 1180
rect 11203 1146 11237 1180
rect 11271 1146 11305 1180
rect 11339 1146 11373 1180
rect 11407 1146 11441 1180
rect 11475 1146 11509 1180
rect 11543 1146 11577 1180
rect 11611 1146 11645 1180
rect 11679 1146 11713 1180
rect 11747 1146 11781 1180
rect 11815 1146 11849 1180
rect 11883 1146 11917 1180
rect 11951 1146 11985 1180
rect 12019 1146 12053 1180
rect 12087 1146 12121 1180
rect 12155 1146 12189 1180
rect 12223 1148 13420 1180
rect 12223 1146 12298 1148
rect 1561 1114 12298 1146
rect 12332 1114 12369 1148
rect 12403 1114 12440 1148
rect 12474 1114 12511 1148
rect 12545 1114 12582 1148
rect 12616 1114 12653 1148
rect 12687 1114 12724 1148
rect 12758 1114 12795 1148
rect 12829 1114 12866 1148
rect 12900 1114 12937 1148
rect 12971 1114 13008 1148
rect 13042 1114 13079 1148
rect 13113 1114 13150 1148
rect 13184 1114 13221 1148
rect 13255 1114 13292 1148
rect 13326 1114 13362 1148
rect 13396 1114 13420 1148
rect 1561 1080 13420 1114
rect 12223 1069 13420 1080
rect 14982 1160 15886 1564
rect 12223 1050 12312 1069
rect 12346 1050 12387 1069
rect 12421 1050 12462 1069
rect 12496 1050 12536 1069
rect 12570 1050 12610 1069
rect 12644 1050 12684 1069
rect 12718 1050 12758 1069
rect 12223 1046 12298 1050
rect 12274 1016 12298 1046
rect 12346 1035 12369 1050
rect 12421 1035 12440 1050
rect 12496 1035 12511 1050
rect 12570 1035 12582 1050
rect 12644 1035 12653 1050
rect 12718 1035 12724 1050
rect 12332 1016 12369 1035
rect 12403 1016 12440 1035
rect 12474 1016 12511 1035
rect 12545 1016 12582 1035
rect 12616 1016 12653 1035
rect 12687 1016 12724 1035
rect 12792 1050 12832 1069
rect 12792 1035 12795 1050
rect 12758 1016 12795 1035
rect 12829 1035 12832 1050
rect 12866 1050 12906 1069
rect 12940 1050 12980 1069
rect 13014 1050 13054 1069
rect 13088 1050 13128 1069
rect 13162 1050 13202 1069
rect 13236 1050 13276 1069
rect 13310 1050 13350 1069
rect 13384 1050 13424 1069
rect 12829 1016 12866 1035
rect 12900 1035 12906 1050
rect 12971 1035 12980 1050
rect 13042 1035 13054 1050
rect 13113 1035 13128 1050
rect 13184 1035 13202 1050
rect 13255 1035 13276 1050
rect 13326 1035 13350 1050
rect 13396 1035 13424 1050
rect 12900 1016 12937 1035
rect 12971 1016 13008 1035
rect 13042 1016 13079 1035
rect 13113 1016 13150 1035
rect 13184 1016 13221 1035
rect 13255 1016 13292 1035
rect 13326 1016 13362 1035
rect 13396 1016 13458 1035
rect 14982 1034 15386 1160
rect 12312 987 13458 1016
rect 12346 953 12387 987
rect 12421 953 12462 987
rect 12496 953 12536 987
rect 12570 953 12610 987
rect 12644 953 12684 987
rect 12718 953 12758 987
rect 12792 953 12832 987
rect 12866 953 12906 987
rect 12940 953 12980 987
rect 13014 953 13054 987
rect 13088 953 13128 987
rect 13162 953 13202 987
rect 13236 953 13276 987
rect 13310 953 13350 987
rect 13384 953 13424 987
rect 15473 1000 15521 1034
rect 15439 948 15555 1000
rect 15473 914 15521 948
rect 15439 884 15555 914
rect 13658 784 13851 792
rect 11872 558 11944 686
rect 11872 524 11899 558
rect 11933 524 11944 558
rect 11872 486 11944 524
rect 11872 452 11899 486
rect 11933 452 11944 486
rect 13658 606 13664 784
rect 13770 606 13851 784
rect 13658 567 13851 606
rect 13658 533 13664 567
rect 13698 533 13736 567
rect 13770 533 13851 567
rect 13658 494 13851 533
rect 13658 460 13664 494
rect 13698 460 13736 494
rect 13770 460 13851 494
rect 13658 388 13851 460
rect 14463 388 14867 884
rect 15439 862 15886 884
rect 15473 828 15521 862
rect 15555 828 15886 862
rect 15439 775 15886 828
rect 15473 741 15521 775
rect 15555 741 15886 775
rect 15482 740 15886 741
rect 12875 176 13215 200
rect 12909 171 12977 176
rect 13011 171 13079 176
rect 13113 171 13181 176
rect 12875 137 12887 142
rect 12921 137 12960 171
rect 13011 142 13033 171
rect 12994 137 13033 142
rect 13067 142 13079 171
rect 13067 137 13105 142
rect 13139 137 13177 171
rect 13211 137 13215 142
rect 12875 108 13215 137
rect 12909 93 12977 108
rect 13011 93 13079 108
rect 13113 93 13181 108
rect 12875 59 12887 74
rect 12921 59 12960 93
rect 13011 74 13033 93
rect 12994 59 13033 74
rect 13067 74 13079 93
rect 13067 59 13105 74
rect 13139 59 13177 93
rect 13211 59 13215 74
rect 12875 50 13215 59
<< viali >>
rect 3157 35981 3191 35996
rect 3230 35981 3264 35996
rect 3303 35981 3337 35996
rect 3376 35981 3410 35996
rect 3449 35981 3483 35996
rect 3522 35981 3556 35996
rect 3157 35962 3180 35981
rect 3180 35962 3191 35981
rect 3230 35962 3249 35981
rect 3249 35962 3264 35981
rect 3303 35962 3318 35981
rect 3318 35962 3337 35981
rect 3376 35962 3387 35981
rect 3387 35962 3410 35981
rect 3449 35962 3456 35981
rect 3456 35962 3483 35981
rect 3522 35962 3525 35981
rect 3525 35962 3556 35981
rect 3595 35962 3629 35996
rect 3668 35981 3702 35996
rect 3741 35981 3775 35996
rect 3814 35981 3848 35996
rect 3887 35981 3921 35996
rect 3960 35981 3994 35996
rect 4033 35981 4067 35996
rect 4106 35981 4140 35996
rect 4179 35981 4213 35996
rect 4252 35981 4286 35996
rect 4325 35981 4359 35996
rect 4398 35981 4432 35996
rect 4471 35981 4505 35996
rect 4544 35981 4578 35996
rect 4617 35981 4651 35996
rect 4690 35981 4724 35996
rect 4763 35981 4797 35996
rect 3668 35962 3698 35981
rect 3698 35962 3702 35981
rect 3741 35962 3767 35981
rect 3767 35962 3775 35981
rect 3814 35962 3836 35981
rect 3836 35962 3848 35981
rect 3887 35962 3905 35981
rect 3905 35962 3921 35981
rect 3960 35962 3974 35981
rect 3974 35962 3994 35981
rect 4033 35962 4043 35981
rect 4043 35962 4067 35981
rect 4106 35962 4112 35981
rect 4112 35962 4140 35981
rect 4179 35962 4181 35981
rect 4181 35962 4213 35981
rect 4252 35962 4284 35981
rect 4284 35962 4286 35981
rect 4325 35962 4353 35981
rect 4353 35962 4359 35981
rect 4398 35962 4422 35981
rect 4422 35962 4432 35981
rect 4471 35962 4491 35981
rect 4491 35962 4505 35981
rect 4544 35962 4560 35981
rect 4560 35962 4578 35981
rect 4617 35962 4629 35981
rect 4629 35962 4651 35981
rect 4690 35962 4698 35981
rect 4698 35962 4724 35981
rect 4763 35962 4767 35981
rect 4767 35962 4797 35981
rect 4836 35962 4870 35996
rect 4909 35981 4943 35996
rect 4982 35981 5016 35996
rect 5055 35981 15529 35996
rect 4909 35962 4940 35981
rect 4940 35962 4943 35981
rect 4982 35962 5009 35981
rect 5009 35962 5016 35981
rect 5055 35947 5078 35981
rect 5078 35947 5112 35981
rect 5112 35947 5147 35981
rect 5147 35947 5181 35981
rect 5181 35947 5216 35981
rect 5216 35947 5250 35981
rect 5250 35947 5285 35981
rect 5285 35947 5319 35981
rect 5319 35947 5354 35981
rect 5354 35947 5388 35981
rect 5388 35947 5423 35981
rect 5423 35947 5457 35981
rect 5457 35947 5492 35981
rect 5492 35947 5526 35981
rect 5526 35947 5561 35981
rect 5561 35947 5595 35981
rect 5595 35947 5630 35981
rect 5630 35947 5664 35981
rect 5664 35947 5699 35981
rect 5699 35947 5733 35981
rect 5733 35947 5768 35981
rect 5768 35947 5802 35981
rect 5802 35947 5837 35981
rect 5837 35947 5871 35981
rect 5871 35947 5906 35981
rect 5906 35947 5940 35981
rect 5940 35947 5975 35981
rect 5975 35947 6009 35981
rect 6009 35947 6044 35981
rect 6044 35947 6078 35981
rect 6078 35947 6113 35981
rect 6113 35947 6147 35981
rect 6147 35947 6182 35981
rect 6182 35947 6216 35981
rect 6216 35947 6251 35981
rect 6251 35947 6285 35981
rect 6285 35947 6320 35981
rect 6320 35947 6354 35981
rect 6354 35947 6389 35981
rect 6389 35947 6423 35981
rect 6423 35947 6458 35981
rect 6458 35947 6492 35981
rect 6492 35947 6527 35981
rect 6527 35947 6561 35981
rect 6561 35947 6596 35981
rect 6596 35947 6630 35981
rect 6630 35947 6665 35981
rect 6665 35947 6699 35981
rect 6699 35947 6734 35981
rect 6734 35947 6768 35981
rect 6768 35947 6803 35981
rect 6803 35947 6837 35981
rect 6837 35947 6872 35981
rect 6872 35947 6906 35981
rect 6906 35947 6941 35981
rect 6941 35947 6975 35981
rect 6975 35947 7010 35981
rect 7010 35947 7044 35981
rect 7044 35947 7079 35981
rect 7079 35947 7113 35981
rect 7113 35947 7148 35981
rect 7148 35947 7182 35981
rect 7182 35947 7217 35981
rect 7217 35947 7251 35981
rect 7251 35947 7286 35981
rect 7286 35947 7320 35981
rect 7320 35947 7355 35981
rect 7355 35947 7389 35981
rect 7389 35947 7424 35981
rect 7424 35947 7458 35981
rect 7458 35947 7493 35981
rect 7493 35947 7527 35981
rect 7527 35947 7562 35981
rect 7562 35947 7596 35981
rect 7596 35947 7631 35981
rect 7631 35947 7665 35981
rect 7665 35947 7699 35981
rect 7699 35947 7733 35981
rect 7733 35947 7767 35981
rect 7767 35947 7801 35981
rect 7801 35947 7835 35981
rect 7835 35947 7869 35981
rect 7869 35947 7903 35981
rect 7903 35947 7937 35981
rect 7937 35947 7971 35981
rect 7971 35947 8005 35981
rect 8005 35947 8039 35981
rect 8039 35947 8073 35981
rect 8073 35947 8107 35981
rect 8107 35947 8141 35981
rect 8141 35947 8175 35981
rect 8175 35947 8209 35981
rect 8209 35947 8243 35981
rect 8243 35947 8277 35981
rect 8277 35947 8311 35981
rect 8311 35947 8345 35981
rect 8345 35947 8379 35981
rect 8379 35947 8413 35981
rect 8413 35947 8447 35981
rect 8447 35947 8481 35981
rect 8481 35947 8515 35981
rect 8515 35947 8549 35981
rect 8549 35947 8583 35981
rect 8583 35947 8617 35981
rect 8617 35947 8651 35981
rect 8651 35947 8685 35981
rect 8685 35947 8719 35981
rect 8719 35947 8753 35981
rect 8753 35947 8787 35981
rect 8787 35947 8821 35981
rect 8821 35947 8855 35981
rect 8855 35947 8889 35981
rect 8889 35947 8923 35981
rect 8923 35947 8957 35981
rect 8957 35947 8991 35981
rect 8991 35947 9025 35981
rect 9025 35947 9059 35981
rect 9059 35947 9093 35981
rect 9093 35947 9127 35981
rect 9127 35947 9161 35981
rect 9161 35947 9195 35981
rect 9195 35947 9229 35981
rect 9229 35947 9263 35981
rect 9263 35947 9297 35981
rect 9297 35947 9331 35981
rect 9331 35947 9365 35981
rect 9365 35947 9399 35981
rect 9399 35947 9433 35981
rect 9433 35947 9467 35981
rect 9467 35947 9501 35981
rect 9501 35947 9535 35981
rect 9535 35947 9569 35981
rect 9569 35947 9603 35981
rect 9603 35947 9637 35981
rect 9637 35947 9671 35981
rect 9671 35947 9705 35981
rect 9705 35947 9739 35981
rect 9739 35947 9773 35981
rect 9773 35947 9807 35981
rect 9807 35947 9841 35981
rect 9841 35947 9875 35981
rect 9875 35947 9909 35981
rect 9909 35947 9943 35981
rect 9943 35947 9977 35981
rect 9977 35947 10011 35981
rect 10011 35947 10045 35981
rect 10045 35947 10079 35981
rect 10079 35947 10113 35981
rect 10113 35947 10147 35981
rect 10147 35947 10181 35981
rect 10181 35947 10215 35981
rect 10215 35947 10249 35981
rect 10249 35947 10283 35981
rect 10283 35947 10317 35981
rect 10317 35947 10351 35981
rect 10351 35947 10385 35981
rect 10385 35947 10419 35981
rect 10419 35947 10453 35981
rect 10453 35947 10487 35981
rect 10487 35947 10521 35981
rect 10521 35947 10555 35981
rect 10555 35947 10589 35981
rect 10589 35947 10623 35981
rect 10623 35947 10657 35981
rect 10657 35947 10691 35981
rect 10691 35947 10725 35981
rect 10725 35947 10759 35981
rect 10759 35947 10793 35981
rect 10793 35947 10827 35981
rect 10827 35947 10861 35981
rect 10861 35947 10895 35981
rect 10895 35947 10929 35981
rect 10929 35947 10963 35981
rect 10963 35947 10997 35981
rect 10997 35947 11031 35981
rect 11031 35947 11065 35981
rect 11065 35947 11099 35981
rect 11099 35947 11133 35981
rect 11133 35947 11167 35981
rect 11167 35947 11201 35981
rect 11201 35947 11235 35981
rect 11235 35947 11269 35981
rect 11269 35947 11303 35981
rect 11303 35947 11337 35981
rect 11337 35947 11371 35981
rect 11371 35947 11405 35981
rect 11405 35947 11439 35981
rect 11439 35947 11473 35981
rect 11473 35947 11507 35981
rect 11507 35947 11541 35981
rect 11541 35947 11575 35981
rect 11575 35947 11609 35981
rect 11609 35947 11643 35981
rect 11643 35947 11677 35981
rect 11677 35947 11711 35981
rect 11711 35947 11745 35981
rect 11745 35947 11779 35981
rect 11779 35947 11813 35981
rect 11813 35947 11847 35981
rect 11847 35947 11881 35981
rect 11881 35947 11915 35981
rect 11915 35947 11949 35981
rect 11949 35947 11983 35981
rect 11983 35947 12017 35981
rect 12017 35947 12051 35981
rect 12051 35947 12085 35981
rect 12085 35947 12119 35981
rect 12119 35947 12153 35981
rect 12153 35947 12187 35981
rect 12187 35947 12221 35981
rect 12221 35947 12255 35981
rect 12255 35947 12289 35981
rect 12289 35947 12323 35981
rect 12323 35947 12357 35981
rect 12357 35947 12391 35981
rect 12391 35947 12425 35981
rect 12425 35947 12459 35981
rect 12459 35947 12493 35981
rect 12493 35947 12527 35981
rect 12527 35947 12561 35981
rect 12561 35947 12595 35981
rect 12595 35947 12629 35981
rect 12629 35947 12663 35981
rect 12663 35947 12697 35981
rect 12697 35947 12731 35981
rect 12731 35947 12765 35981
rect 12765 35947 12799 35981
rect 12799 35947 12833 35981
rect 12833 35947 12867 35981
rect 12867 35947 12901 35981
rect 12901 35947 12935 35981
rect 12935 35947 12969 35981
rect 12969 35947 13003 35981
rect 13003 35947 13037 35981
rect 13037 35947 13071 35981
rect 13071 35947 13105 35981
rect 13105 35947 13139 35981
rect 13139 35947 13173 35981
rect 13173 35947 13207 35981
rect 13207 35947 13241 35981
rect 13241 35947 13275 35981
rect 13275 35947 13309 35981
rect 13309 35947 13343 35981
rect 13343 35947 13377 35981
rect 13377 35947 13411 35981
rect 13411 35947 13445 35981
rect 13445 35947 13479 35981
rect 13479 35947 13513 35981
rect 13513 35947 13547 35981
rect 13547 35947 13581 35981
rect 13581 35947 13615 35981
rect 13615 35947 13649 35981
rect 13649 35947 13683 35981
rect 13683 35947 13717 35981
rect 13717 35947 13751 35981
rect 13751 35947 13785 35981
rect 13785 35947 13925 35981
rect 13925 35947 13959 35981
rect 13959 35947 13996 35981
rect 13996 35947 14030 35981
rect 14030 35947 14067 35981
rect 14067 35947 14101 35981
rect 14101 35947 14138 35981
rect 14138 35947 14172 35981
rect 14172 35947 14209 35981
rect 14209 35947 14243 35981
rect 14243 35947 14280 35981
rect 14280 35947 14314 35981
rect 14314 35947 14351 35981
rect 14351 35947 14385 35981
rect 14385 35947 14422 35981
rect 14422 35947 14456 35981
rect 14456 35947 14493 35981
rect 14493 35947 14527 35981
rect 14527 35947 14563 35981
rect 14563 35947 14597 35981
rect 14597 35947 14633 35981
rect 14633 35947 14667 35981
rect 14667 35947 14703 35981
rect 14703 35947 14737 35981
rect 14737 35947 14773 35981
rect 14773 35947 14807 35981
rect 14807 35947 14843 35981
rect 14843 35947 14877 35981
rect 14877 35947 14913 35981
rect 14913 35947 14947 35981
rect 14947 35947 14983 35981
rect 14983 35947 15017 35981
rect 15017 35947 15053 35981
rect 15053 35947 15087 35981
rect 15087 35947 15123 35981
rect 15123 35947 15157 35981
rect 15157 35947 15193 35981
rect 15193 35947 15227 35981
rect 15227 35947 15263 35981
rect 15263 35947 15297 35981
rect 15297 35947 15333 35981
rect 15333 35947 15367 35981
rect 15367 35947 15403 35981
rect 15403 35947 15437 35981
rect 15437 35947 15473 35981
rect 15473 35947 15507 35981
rect 15507 35947 15529 35981
rect 3157 35890 3191 35924
rect 3230 35890 3264 35924
rect 3303 35890 3337 35924
rect 3376 35890 3410 35924
rect 3449 35890 3483 35924
rect 3522 35890 3556 35924
rect 3595 35890 3629 35924
rect 3668 35890 3702 35924
rect 3741 35890 3775 35924
rect 3814 35890 3848 35924
rect 3887 35890 3921 35924
rect 3960 35890 3994 35924
rect 4033 35890 4067 35924
rect 4106 35890 4140 35924
rect 4179 35890 4213 35924
rect 4252 35890 4286 35924
rect 4325 35890 4359 35924
rect 4398 35890 4432 35924
rect 4471 35890 4505 35924
rect 4544 35890 4578 35924
rect 4617 35890 4651 35924
rect 4690 35890 4724 35924
rect 4763 35890 4797 35924
rect 4836 35890 4870 35924
rect 4909 35890 4943 35924
rect 4982 35890 5016 35924
rect 5055 35890 15529 35947
rect 463 35645 929 35648
rect 463 35637 843 35645
rect 463 35603 487 35637
rect 487 35603 521 35637
rect 521 35603 559 35637
rect 559 35603 593 35637
rect 593 35603 631 35637
rect 631 35603 665 35637
rect 665 35603 703 35637
rect 703 35603 737 35637
rect 737 35603 775 35637
rect 775 35603 809 35637
rect 809 35611 843 35637
rect 843 35611 877 35645
rect 877 35611 915 35645
rect 915 35611 929 35645
rect 809 35603 929 35611
rect 463 35569 929 35603
rect 463 35535 487 35569
rect 487 35535 521 35569
rect 521 35535 559 35569
rect 559 35535 593 35569
rect 593 35535 631 35569
rect 631 35535 665 35569
rect 665 35535 703 35569
rect 703 35535 737 35569
rect 737 35535 775 35569
rect 775 35535 809 35569
rect 809 35561 929 35569
rect 809 35535 843 35561
rect 463 35527 843 35535
rect 843 35527 877 35561
rect 877 35527 915 35561
rect 915 35527 929 35561
rect 463 35501 929 35527
rect 463 35467 487 35501
rect 487 35467 521 35501
rect 521 35467 559 35501
rect 559 35467 593 35501
rect 593 35467 631 35501
rect 631 35467 665 35501
rect 665 35467 703 35501
rect 703 35467 737 35501
rect 737 35467 775 35501
rect 775 35467 809 35501
rect 809 35477 929 35501
rect 809 35467 843 35477
rect 463 35443 843 35467
rect 843 35443 877 35477
rect 877 35443 915 35477
rect 915 35443 929 35477
rect 463 35433 929 35443
rect 463 35399 487 35433
rect 487 35399 521 35433
rect 521 35399 559 35433
rect 559 35399 593 35433
rect 593 35399 631 35433
rect 631 35399 665 35433
rect 665 35399 703 35433
rect 703 35399 737 35433
rect 737 35399 775 35433
rect 775 35399 809 35433
rect 809 35399 929 35433
rect 463 35393 929 35399
rect 463 35365 843 35393
rect 463 35331 487 35365
rect 487 35331 521 35365
rect 521 35331 559 35365
rect 559 35331 593 35365
rect 593 35331 631 35365
rect 631 35331 665 35365
rect 665 35331 703 35365
rect 703 35331 737 35365
rect 737 35331 775 35365
rect 775 35331 809 35365
rect 809 35359 843 35365
rect 843 35359 877 35393
rect 877 35359 915 35393
rect 915 35359 929 35393
rect 809 35331 929 35359
rect 463 35309 929 35331
rect 463 35297 843 35309
rect 463 35263 487 35297
rect 487 35263 521 35297
rect 521 35263 559 35297
rect 559 35263 593 35297
rect 593 35263 631 35297
rect 631 35263 665 35297
rect 665 35263 703 35297
rect 703 35263 737 35297
rect 737 35263 775 35297
rect 775 35263 809 35297
rect 809 35275 843 35297
rect 843 35275 877 35309
rect 877 35275 915 35309
rect 915 35275 929 35309
rect 809 35263 929 35275
rect 463 35229 929 35263
rect 463 35195 487 35229
rect 487 35195 521 35229
rect 521 35195 559 35229
rect 559 35195 593 35229
rect 593 35195 631 35229
rect 631 35195 665 35229
rect 665 35195 703 35229
rect 703 35195 737 35229
rect 737 35195 775 35229
rect 775 35195 809 35229
rect 809 35225 929 35229
rect 809 35195 843 35225
rect 463 35191 843 35195
rect 843 35191 877 35225
rect 877 35191 915 35225
rect 915 35191 929 35225
rect 463 35161 929 35191
rect 463 35127 487 35161
rect 487 35127 521 35161
rect 521 35127 559 35161
rect 559 35127 593 35161
rect 593 35127 631 35161
rect 631 35127 665 35161
rect 665 35127 703 35161
rect 703 35127 737 35161
rect 737 35127 775 35161
rect 775 35127 809 35161
rect 809 35141 929 35161
rect 809 35127 843 35141
rect 463 35107 843 35127
rect 843 35107 877 35141
rect 877 35107 915 35141
rect 915 35107 929 35141
rect 463 35093 929 35107
rect 463 35059 487 35093
rect 487 35059 521 35093
rect 521 35059 559 35093
rect 559 35059 593 35093
rect 593 35059 631 35093
rect 631 35059 665 35093
rect 665 35059 703 35093
rect 703 35059 737 35093
rect 737 35059 775 35093
rect 775 35059 809 35093
rect 809 35059 929 35093
rect 463 35057 929 35059
rect 463 35025 843 35057
rect 463 34991 487 35025
rect 487 34991 521 35025
rect 521 34991 559 35025
rect 559 34991 593 35025
rect 593 34991 631 35025
rect 631 34991 665 35025
rect 665 34991 703 35025
rect 703 34991 737 35025
rect 737 34991 775 35025
rect 775 34991 809 35025
rect 809 35023 843 35025
rect 843 35023 877 35057
rect 877 35023 915 35057
rect 915 35023 929 35057
rect 809 34991 929 35023
rect 463 34973 929 34991
rect 463 34957 843 34973
rect 463 34923 487 34957
rect 487 34923 521 34957
rect 521 34923 559 34957
rect 559 34923 593 34957
rect 593 34923 631 34957
rect 631 34923 665 34957
rect 665 34923 703 34957
rect 703 34923 737 34957
rect 737 34923 775 34957
rect 775 34923 809 34957
rect 809 34939 843 34957
rect 843 34939 877 34973
rect 877 34939 915 34973
rect 915 34939 929 34973
rect 809 34923 929 34939
rect 463 34889 929 34923
rect 463 34855 487 34889
rect 487 34855 521 34889
rect 521 34855 559 34889
rect 559 34855 593 34889
rect 593 34855 631 34889
rect 631 34855 665 34889
rect 665 34855 703 34889
rect 703 34855 737 34889
rect 737 34855 775 34889
rect 775 34855 809 34889
rect 809 34855 843 34889
rect 843 34855 877 34889
rect 877 34855 915 34889
rect 915 34855 929 34889
rect 463 34821 929 34855
rect 463 34787 487 34821
rect 487 34787 521 34821
rect 521 34787 559 34821
rect 559 34787 593 34821
rect 593 34787 631 34821
rect 631 34787 665 34821
rect 665 34787 703 34821
rect 703 34787 737 34821
rect 737 34787 775 34821
rect 775 34787 809 34821
rect 809 34805 929 34821
rect 809 34787 843 34805
rect 463 34771 843 34787
rect 843 34771 877 34805
rect 877 34771 915 34805
rect 915 34771 929 34805
rect 463 34753 929 34771
rect 463 34719 487 34753
rect 487 34719 521 34753
rect 521 34719 559 34753
rect 559 34719 593 34753
rect 593 34719 631 34753
rect 631 34719 665 34753
rect 665 34719 703 34753
rect 703 34719 737 34753
rect 737 34719 775 34753
rect 775 34719 809 34753
rect 809 34721 929 34753
rect 809 34719 843 34721
rect 463 34687 843 34719
rect 843 34687 877 34721
rect 877 34687 915 34721
rect 915 34687 929 34721
rect 463 34685 929 34687
rect 463 34651 487 34685
rect 487 34651 521 34685
rect 521 34651 559 34685
rect 559 34651 593 34685
rect 593 34651 631 34685
rect 631 34651 665 34685
rect 665 34651 703 34685
rect 703 34651 737 34685
rect 737 34651 775 34685
rect 775 34651 809 34685
rect 809 34651 929 34685
rect 463 34637 929 34651
rect 463 34617 843 34637
rect 463 34583 487 34617
rect 487 34583 521 34617
rect 521 34583 559 34617
rect 559 34583 593 34617
rect 593 34583 631 34617
rect 631 34583 665 34617
rect 665 34583 703 34617
rect 703 34583 737 34617
rect 737 34583 775 34617
rect 775 34583 809 34617
rect 809 34603 843 34617
rect 843 34603 877 34637
rect 877 34603 915 34637
rect 915 34603 929 34637
rect 809 34583 929 34603
rect 463 34553 929 34583
rect 463 34549 843 34553
rect 463 34515 487 34549
rect 487 34515 521 34549
rect 521 34515 559 34549
rect 559 34515 593 34549
rect 593 34515 631 34549
rect 631 34515 665 34549
rect 665 34515 703 34549
rect 703 34515 737 34549
rect 737 34515 775 34549
rect 775 34515 809 34549
rect 809 34519 843 34549
rect 843 34519 877 34553
rect 877 34519 915 34553
rect 915 34519 929 34553
rect 809 34515 929 34519
rect 463 34481 929 34515
rect 463 34447 487 34481
rect 487 34447 521 34481
rect 521 34447 559 34481
rect 559 34447 593 34481
rect 593 34447 631 34481
rect 631 34447 665 34481
rect 665 34447 703 34481
rect 703 34447 737 34481
rect 737 34447 775 34481
rect 775 34447 809 34481
rect 809 34469 929 34481
rect 809 34447 843 34469
rect 463 34435 843 34447
rect 843 34435 877 34469
rect 877 34435 915 34469
rect 915 34435 929 34469
rect 463 34413 929 34435
rect 463 34379 487 34413
rect 487 34379 521 34413
rect 521 34379 559 34413
rect 559 34379 593 34413
rect 593 34379 631 34413
rect 631 34379 665 34413
rect 665 34379 703 34413
rect 703 34379 737 34413
rect 737 34379 775 34413
rect 775 34379 809 34413
rect 809 34385 929 34413
rect 809 34379 843 34385
rect 463 34351 843 34379
rect 843 34351 877 34385
rect 877 34351 915 34385
rect 915 34351 929 34385
rect 463 34345 929 34351
rect 463 34311 487 34345
rect 487 34311 521 34345
rect 521 34311 559 34345
rect 559 34311 593 34345
rect 593 34311 631 34345
rect 631 34311 665 34345
rect 665 34311 703 34345
rect 703 34311 737 34345
rect 737 34311 775 34345
rect 775 34311 809 34345
rect 809 34311 929 34345
rect 463 34301 929 34311
rect 463 34277 843 34301
rect 463 34246 487 34277
rect 487 34246 521 34277
rect 521 34246 559 34277
rect 559 34246 593 34277
rect 593 34246 631 34277
rect 631 34246 665 34277
rect 665 34246 703 34277
rect 703 34246 737 34277
rect 737 34246 775 34277
rect 775 34246 809 34277
rect 809 34267 843 34277
rect 843 34267 877 34301
rect 877 34267 915 34301
rect 915 34267 929 34301
rect 809 34246 929 34267
rect 463 34175 487 34207
rect 487 34175 497 34207
rect 535 34175 559 34207
rect 559 34175 569 34207
rect 607 34175 631 34207
rect 631 34175 641 34207
rect 679 34175 703 34207
rect 703 34175 713 34207
rect 751 34175 775 34207
rect 775 34175 785 34207
rect 823 34183 843 34207
rect 843 34183 857 34207
rect 895 34183 915 34207
rect 915 34183 929 34207
rect 463 34173 497 34175
rect 535 34173 569 34175
rect 607 34173 641 34175
rect 679 34173 713 34175
rect 751 34173 785 34175
rect 823 34173 857 34183
rect 895 34173 929 34183
rect 463 34107 487 34134
rect 487 34107 497 34134
rect 535 34107 559 34134
rect 559 34107 569 34134
rect 607 34107 631 34134
rect 631 34107 641 34134
rect 679 34107 703 34134
rect 703 34107 713 34134
rect 751 34107 775 34134
rect 775 34107 785 34134
rect 823 34133 857 34134
rect 895 34133 929 34134
rect 463 34100 497 34107
rect 535 34100 569 34107
rect 607 34100 641 34107
rect 679 34100 713 34107
rect 751 34100 785 34107
rect 823 34100 843 34133
rect 843 34100 857 34133
rect 895 34100 915 34133
rect 915 34100 929 34133
rect 463 34039 487 34061
rect 487 34039 497 34061
rect 535 34039 559 34061
rect 559 34039 569 34061
rect 607 34039 631 34061
rect 631 34039 641 34061
rect 679 34039 703 34061
rect 703 34039 713 34061
rect 751 34039 775 34061
rect 775 34039 785 34061
rect 823 34049 857 34061
rect 895 34049 929 34061
rect 463 34027 497 34039
rect 535 34027 569 34039
rect 607 34027 641 34039
rect 679 34027 713 34039
rect 751 34027 785 34039
rect 823 34027 843 34049
rect 843 34027 857 34049
rect 895 34027 915 34049
rect 915 34027 929 34049
rect -17 33971 17 33986
rect 75 33971 89 33986
rect 89 33971 109 33986
rect 167 33971 199 33986
rect 199 33971 201 33986
rect 259 33971 271 33986
rect 271 33971 293 33986
rect 463 33971 487 33988
rect 487 33971 497 33988
rect 535 33971 559 33988
rect 559 33971 569 33988
rect 607 33971 631 33988
rect 631 33971 641 33988
rect 679 33971 703 33988
rect 703 33971 713 33988
rect 751 33971 775 33988
rect 775 33971 785 33988
rect -17 33952 17 33971
rect 75 33952 109 33971
rect 167 33952 201 33971
rect 259 33952 293 33971
rect 463 33954 497 33971
rect 535 33954 569 33971
rect 607 33954 641 33971
rect 679 33954 713 33971
rect 751 33954 785 33971
rect 823 33965 857 33988
rect 895 33965 929 33988
rect 823 33954 843 33965
rect 843 33954 857 33965
rect 895 33954 915 33965
rect 915 33954 929 33965
rect -17 33903 17 33914
rect 75 33903 89 33914
rect 89 33903 109 33914
rect 167 33903 199 33914
rect 199 33903 201 33914
rect 259 33903 271 33914
rect 271 33903 293 33914
rect 463 33903 487 33915
rect 487 33903 497 33915
rect 535 33903 559 33915
rect 559 33903 569 33915
rect 607 33903 631 33915
rect 631 33903 641 33915
rect 679 33903 703 33915
rect 703 33903 713 33915
rect 751 33903 775 33915
rect 775 33903 785 33915
rect -17 33880 17 33903
rect 75 33880 109 33903
rect 167 33880 201 33903
rect 259 33880 293 33903
rect 463 33881 497 33903
rect 535 33881 569 33903
rect 607 33881 641 33903
rect 679 33881 713 33903
rect 751 33881 785 33903
rect 823 33881 857 33915
rect 895 33881 929 33915
rect -17 33835 17 33842
rect 75 33835 89 33842
rect 89 33835 109 33842
rect 167 33835 199 33842
rect 199 33835 201 33842
rect 259 33835 271 33842
rect 271 33835 293 33842
rect 463 33835 487 33842
rect 487 33835 497 33842
rect 535 33835 559 33842
rect 559 33835 569 33842
rect 607 33835 631 33842
rect 631 33835 641 33842
rect 679 33835 703 33842
rect 703 33835 713 33842
rect 751 33835 775 33842
rect 775 33835 785 33842
rect -17 33808 17 33835
rect 75 33808 109 33835
rect 167 33808 201 33835
rect 259 33808 293 33835
rect 463 33808 497 33835
rect 535 33808 569 33835
rect 607 33808 641 33835
rect 679 33808 713 33835
rect 751 33808 785 33835
rect 823 33808 857 33842
rect 895 33808 929 33842
rect -17 33767 17 33769
rect 75 33767 89 33769
rect 89 33767 109 33769
rect 167 33767 199 33769
rect 199 33767 201 33769
rect 259 33767 271 33769
rect 271 33767 293 33769
rect 463 33767 487 33769
rect 487 33767 497 33769
rect 535 33767 559 33769
rect 559 33767 569 33769
rect 607 33767 631 33769
rect 631 33767 641 33769
rect 679 33767 703 33769
rect 703 33767 713 33769
rect 751 33767 775 33769
rect 775 33767 785 33769
rect -17 33735 17 33767
rect 75 33735 109 33767
rect 167 33735 201 33767
rect 259 33735 293 33767
rect 463 33735 497 33767
rect 535 33735 569 33767
rect 607 33735 641 33767
rect 679 33735 713 33767
rect 751 33735 785 33767
rect 823 33763 843 33769
rect 843 33763 857 33769
rect 895 33763 915 33769
rect 915 33763 929 33769
rect 823 33735 857 33763
rect 895 33735 929 33763
rect -17 33665 17 33696
rect 75 33665 109 33696
rect 167 33665 201 33696
rect 259 33665 293 33696
rect 463 33665 497 33696
rect 535 33665 569 33696
rect 607 33665 641 33696
rect 679 33665 713 33696
rect 751 33665 785 33696
rect 823 33679 843 33696
rect 843 33679 857 33696
rect 895 33679 915 33696
rect 915 33679 929 33696
rect -17 33662 17 33665
rect 75 33662 89 33665
rect 89 33662 109 33665
rect 167 33662 199 33665
rect 199 33662 201 33665
rect 259 33662 271 33665
rect 271 33662 293 33665
rect 463 33662 487 33665
rect 487 33662 497 33665
rect 535 33662 559 33665
rect 559 33662 569 33665
rect 607 33662 631 33665
rect 631 33662 641 33665
rect 679 33662 703 33665
rect 703 33662 713 33665
rect 751 33662 775 33665
rect 775 33662 785 33665
rect 823 33662 857 33679
rect 895 33662 929 33679
rect -17 33597 17 33623
rect 75 33597 109 33623
rect 167 33597 201 33623
rect 259 33597 293 33623
rect 463 33597 497 33623
rect 535 33597 569 33623
rect 607 33597 641 33623
rect 679 33597 713 33623
rect 751 33597 785 33623
rect -17 33589 17 33597
rect 75 33589 89 33597
rect 89 33589 109 33597
rect 167 33589 199 33597
rect 199 33589 201 33597
rect 259 33589 271 33597
rect 271 33589 293 33597
rect 463 33589 487 33597
rect 487 33589 497 33597
rect 535 33589 559 33597
rect 559 33589 569 33597
rect 607 33589 631 33597
rect 631 33589 641 33597
rect 679 33589 703 33597
rect 703 33589 713 33597
rect 751 33589 775 33597
rect 775 33589 785 33597
rect 823 33595 843 33623
rect 843 33595 857 33623
rect 895 33595 915 33623
rect 915 33595 929 33623
rect 823 33589 857 33595
rect 895 33589 929 33595
rect -17 33529 17 33550
rect 75 33529 109 33550
rect 167 33529 201 33550
rect 259 33529 293 33550
rect 463 33529 497 33550
rect 535 33529 569 33550
rect 607 33529 641 33550
rect 679 33529 713 33550
rect 751 33529 785 33550
rect 823 33545 857 33550
rect 895 33545 929 33550
rect -17 33516 17 33529
rect 75 33516 89 33529
rect 89 33516 109 33529
rect 167 33516 199 33529
rect 199 33516 201 33529
rect 259 33516 271 33529
rect 271 33516 293 33529
rect 463 33516 487 33529
rect 487 33516 497 33529
rect 535 33516 559 33529
rect 559 33516 569 33529
rect 607 33516 631 33529
rect 631 33516 641 33529
rect 679 33516 703 33529
rect 703 33516 713 33529
rect 751 33516 775 33529
rect 775 33516 785 33529
rect 823 33516 843 33545
rect 843 33516 857 33545
rect 895 33516 915 33545
rect 915 33516 929 33545
rect -17 33461 17 33477
rect 75 33461 109 33477
rect 167 33461 201 33477
rect 259 33461 293 33477
rect 463 33461 497 33477
rect 535 33461 569 33477
rect 607 33461 641 33477
rect 679 33461 713 33477
rect 751 33461 785 33477
rect 823 33461 857 33477
rect 895 33461 929 33477
rect -17 33443 17 33461
rect 75 33443 89 33461
rect 89 33443 109 33461
rect 167 33443 199 33461
rect 199 33443 201 33461
rect 259 33443 271 33461
rect 271 33443 293 33461
rect 463 33443 487 33461
rect 487 33443 497 33461
rect 535 33443 559 33461
rect 559 33443 569 33461
rect 607 33443 631 33461
rect 631 33443 641 33461
rect 679 33443 703 33461
rect 703 33443 713 33461
rect 751 33443 775 33461
rect 775 33443 785 33461
rect 823 33443 843 33461
rect 843 33443 857 33461
rect 895 33443 915 33461
rect 915 33443 929 33461
rect -17 33393 17 33404
rect 75 33393 109 33404
rect 167 33393 201 33404
rect 259 33393 293 33404
rect 463 33393 497 33404
rect 535 33393 569 33404
rect 607 33393 641 33404
rect 679 33393 713 33404
rect 751 33393 785 33404
rect -17 33370 17 33393
rect 75 33370 89 33393
rect 89 33370 109 33393
rect 167 33370 199 33393
rect 199 33370 201 33393
rect 259 33370 271 33393
rect 271 33370 293 33393
rect 463 33370 487 33393
rect 487 33370 497 33393
rect 535 33370 559 33393
rect 559 33370 569 33393
rect 607 33370 631 33393
rect 631 33370 641 33393
rect 679 33370 703 33393
rect 703 33370 713 33393
rect 751 33370 775 33393
rect 775 33370 785 33393
rect 823 33377 857 33404
rect 895 33377 929 33404
rect 823 33370 843 33377
rect 843 33370 857 33377
rect 895 33370 915 33377
rect 915 33370 929 33377
rect -17 33325 17 33331
rect 75 33325 109 33331
rect 167 33325 201 33331
rect 259 33325 293 33331
rect 463 33325 497 33331
rect 535 33325 569 33331
rect 607 33325 641 33331
rect 679 33325 713 33331
rect 751 33325 785 33331
rect -17 33297 17 33325
rect 75 33297 89 33325
rect 89 33297 109 33325
rect 167 33297 199 33325
rect 199 33297 201 33325
rect 259 33297 271 33325
rect 271 33297 293 33325
rect 463 33297 487 33325
rect 487 33297 497 33325
rect 535 33297 559 33325
rect 559 33297 569 33325
rect 607 33297 631 33325
rect 631 33297 641 33325
rect 679 33297 703 33325
rect 703 33297 713 33325
rect 751 33297 775 33325
rect 775 33297 785 33325
rect 823 33297 857 33331
rect 895 33297 929 33331
rect -17 33257 17 33258
rect 75 33257 109 33258
rect 167 33257 201 33258
rect 259 33257 293 33258
rect 463 33257 497 33258
rect 535 33257 569 33258
rect 607 33257 641 33258
rect 679 33257 713 33258
rect 751 33257 785 33258
rect -17 33224 17 33257
rect 75 33224 89 33257
rect 89 33224 109 33257
rect 167 33224 199 33257
rect 199 33224 201 33257
rect 259 33224 271 33257
rect 271 33224 293 33257
rect 463 33224 487 33257
rect 487 33224 497 33257
rect 535 33224 559 33257
rect 559 33224 569 33257
rect 607 33224 631 33257
rect 631 33224 641 33257
rect 679 33224 703 33257
rect 703 33224 713 33257
rect 751 33224 775 33257
rect 775 33224 785 33257
rect 823 33224 857 33258
rect 895 33224 929 33258
rect -17 33155 17 33185
rect 75 33155 89 33185
rect 89 33155 109 33185
rect 167 33155 199 33185
rect 199 33155 201 33185
rect 259 33155 271 33185
rect 271 33155 293 33185
rect 463 33155 487 33185
rect 487 33155 497 33185
rect 535 33155 559 33185
rect 559 33155 569 33185
rect 607 33155 631 33185
rect 631 33155 641 33185
rect 679 33155 703 33185
rect 703 33155 713 33185
rect 751 33155 775 33185
rect 775 33155 785 33185
rect 823 33175 843 33185
rect 843 33175 857 33185
rect 895 33175 915 33185
rect 915 33175 929 33185
rect -17 33151 17 33155
rect 75 33151 109 33155
rect 167 33151 201 33155
rect 259 33151 293 33155
rect 463 33151 497 33155
rect 535 33151 569 33155
rect 607 33151 641 33155
rect 679 33151 713 33155
rect 751 33151 785 33155
rect 823 33151 857 33175
rect 895 33151 929 33175
rect -17 33087 17 33112
rect 75 33087 89 33112
rect 89 33087 109 33112
rect 167 33087 199 33112
rect 199 33087 201 33112
rect 259 33087 271 33112
rect 271 33087 293 33112
rect 463 33087 487 33112
rect 487 33087 497 33112
rect 535 33087 559 33112
rect 559 33087 569 33112
rect 607 33087 631 33112
rect 631 33087 641 33112
rect 679 33087 703 33112
rect 703 33087 713 33112
rect 751 33087 775 33112
rect 775 33087 785 33112
rect 823 33091 843 33112
rect 843 33091 857 33112
rect 895 33091 915 33112
rect 915 33091 929 33112
rect -17 33078 17 33087
rect 75 33078 109 33087
rect 167 33078 201 33087
rect 259 33078 293 33087
rect 463 33078 497 33087
rect 535 33078 569 33087
rect 607 33078 641 33087
rect 679 33078 713 33087
rect 751 33078 785 33087
rect 823 33078 857 33091
rect 895 33078 929 33091
rect -17 33019 17 33039
rect 75 33019 89 33039
rect 89 33019 109 33039
rect 167 33019 199 33039
rect 199 33019 201 33039
rect 259 33019 271 33039
rect 271 33019 293 33039
rect 463 33019 487 33039
rect 487 33019 497 33039
rect 535 33019 559 33039
rect 559 33019 569 33039
rect 607 33019 631 33039
rect 631 33019 641 33039
rect 679 33019 703 33039
rect 703 33019 713 33039
rect 751 33019 775 33039
rect 775 33019 785 33039
rect -17 33005 17 33019
rect 75 33005 109 33019
rect 167 33005 201 33019
rect 259 33005 293 33019
rect 463 33005 497 33019
rect 535 33005 569 33019
rect 607 33005 641 33019
rect 679 33005 713 33019
rect 751 33005 785 33019
rect 823 33007 843 33039
rect 843 33007 857 33039
rect 895 33007 915 33039
rect 915 33007 929 33039
rect 823 33005 857 33007
rect 895 33005 929 33007
rect -17 32951 17 32966
rect 75 32951 89 32966
rect 89 32951 109 32966
rect 167 32951 199 32966
rect 199 32951 201 32966
rect 259 32951 271 32966
rect 271 32951 293 32966
rect 463 32951 487 32966
rect 487 32951 497 32966
rect 535 32951 559 32966
rect 559 32951 569 32966
rect 607 32951 631 32966
rect 631 32951 641 32966
rect 679 32951 703 32966
rect 703 32951 713 32966
rect 751 32951 775 32966
rect 775 32951 785 32966
rect 823 32957 857 32966
rect 895 32957 929 32966
rect -17 32932 17 32951
rect 75 32932 109 32951
rect 167 32932 201 32951
rect 259 32932 293 32951
rect 463 32932 497 32951
rect 535 32932 569 32951
rect 607 32932 641 32951
rect 679 32932 713 32951
rect 751 32932 785 32951
rect 823 32932 843 32957
rect 843 32932 857 32957
rect 895 32932 915 32957
rect 915 32932 929 32957
rect -17 32883 17 32893
rect 75 32883 89 32893
rect 89 32883 109 32893
rect 167 32883 199 32893
rect 199 32883 201 32893
rect 259 32883 271 32893
rect 271 32883 293 32893
rect 463 32883 487 32893
rect 487 32883 497 32893
rect 535 32883 559 32893
rect 559 32883 569 32893
rect 607 32883 631 32893
rect 631 32883 641 32893
rect 679 32883 703 32893
rect 703 32883 713 32893
rect 751 32883 775 32893
rect 775 32883 785 32893
rect -17 32859 17 32883
rect 75 32859 109 32883
rect 167 32859 201 32883
rect 259 32859 293 32883
rect 463 32859 497 32883
rect 535 32859 569 32883
rect 607 32859 641 32883
rect 679 32859 713 32883
rect 751 32859 785 32883
rect 823 32873 857 32893
rect 895 32873 929 32893
rect 823 32859 843 32873
rect 843 32859 857 32873
rect 895 32859 915 32873
rect 915 32859 929 32873
rect -17 32815 17 32820
rect 75 32815 89 32820
rect 89 32815 109 32820
rect 167 32815 199 32820
rect 199 32815 201 32820
rect 259 32815 271 32820
rect 271 32815 293 32820
rect 463 32815 487 32820
rect 487 32815 497 32820
rect 535 32815 559 32820
rect 559 32815 569 32820
rect 607 32815 631 32820
rect 631 32815 641 32820
rect 679 32815 703 32820
rect 703 32815 713 32820
rect 751 32815 775 32820
rect 775 32815 785 32820
rect -17 32786 17 32815
rect 75 32786 109 32815
rect 167 32786 201 32815
rect 259 32786 293 32815
rect 463 32786 497 32815
rect 535 32786 569 32815
rect 607 32786 641 32815
rect 679 32786 713 32815
rect 751 32786 785 32815
rect 823 32789 857 32820
rect 895 32789 929 32820
rect 823 32786 843 32789
rect 843 32786 857 32789
rect 895 32786 915 32789
rect 915 32786 929 32789
rect -17 32713 17 32747
rect 75 32713 109 32747
rect 167 32713 201 32747
rect 259 32713 293 32747
rect 463 32713 497 32747
rect 535 32713 569 32747
rect 607 32713 641 32747
rect 679 32713 713 32747
rect 751 32713 785 32747
rect 823 32713 857 32747
rect 895 32713 929 32747
rect -17 32645 17 32674
rect 75 32645 109 32674
rect 167 32645 201 32674
rect 259 32645 293 32674
rect 463 32645 497 32674
rect 535 32645 569 32674
rect 607 32645 641 32674
rect 679 32645 713 32674
rect 751 32645 785 32674
rect 823 32671 843 32674
rect 843 32671 857 32674
rect 895 32671 915 32674
rect 915 32671 929 32674
rect -17 32640 17 32645
rect 75 32640 89 32645
rect 89 32640 109 32645
rect 167 32640 199 32645
rect 199 32640 201 32645
rect 259 32640 271 32645
rect 271 32640 293 32645
rect 463 32640 487 32645
rect 487 32640 497 32645
rect 535 32640 559 32645
rect 559 32640 569 32645
rect 607 32640 631 32645
rect 631 32640 641 32645
rect 679 32640 703 32645
rect 703 32640 713 32645
rect 751 32640 775 32645
rect 775 32640 785 32645
rect 823 32640 857 32671
rect 895 32640 929 32671
rect -17 32577 17 32601
rect 75 32577 109 32601
rect 167 32577 201 32601
rect 259 32577 293 32601
rect 463 32577 497 32601
rect 535 32577 569 32601
rect 607 32577 641 32601
rect 679 32577 713 32601
rect 751 32577 785 32601
rect 823 32587 843 32601
rect 843 32587 857 32601
rect 895 32587 915 32601
rect 915 32587 929 32601
rect -17 32567 17 32577
rect 75 32567 89 32577
rect 89 32567 109 32577
rect 167 32567 199 32577
rect 199 32567 201 32577
rect 259 32567 271 32577
rect 271 32567 293 32577
rect 463 32567 487 32577
rect 487 32567 497 32577
rect 535 32567 559 32577
rect 559 32567 569 32577
rect 607 32567 631 32577
rect 631 32567 641 32577
rect 679 32567 703 32577
rect 703 32567 713 32577
rect 751 32567 775 32577
rect 775 32567 785 32577
rect 823 32567 857 32587
rect 895 32567 929 32587
rect -17 32509 17 32528
rect 75 32509 109 32528
rect 167 32509 201 32528
rect 259 32509 293 32528
rect 463 32509 497 32528
rect 535 32509 569 32528
rect 607 32509 641 32528
rect 679 32509 713 32528
rect 751 32509 785 32528
rect -17 32494 17 32509
rect 75 32494 89 32509
rect 89 32494 109 32509
rect 167 32494 199 32509
rect 199 32494 201 32509
rect 259 32494 271 32509
rect 271 32494 293 32509
rect 463 32494 487 32509
rect 487 32494 497 32509
rect 535 32494 559 32509
rect 559 32494 569 32509
rect 607 32494 631 32509
rect 631 32494 641 32509
rect 679 32494 703 32509
rect 703 32494 713 32509
rect 751 32494 775 32509
rect 775 32494 785 32509
rect 823 32503 843 32528
rect 843 32503 857 32528
rect 895 32503 915 32528
rect 915 32503 929 32528
rect 823 32494 857 32503
rect 895 32494 929 32503
rect -17 32441 17 32455
rect 75 32441 109 32455
rect 167 32441 201 32455
rect 259 32441 293 32455
rect 463 32441 497 32455
rect 535 32441 569 32455
rect 607 32441 641 32455
rect 679 32441 713 32455
rect 751 32441 785 32455
rect 823 32453 857 32455
rect 895 32453 929 32455
rect -17 32421 17 32441
rect 75 32421 89 32441
rect 89 32421 109 32441
rect 167 32421 199 32441
rect 199 32421 201 32441
rect 259 32421 271 32441
rect 271 32421 293 32441
rect 463 32421 487 32441
rect 487 32421 497 32441
rect 535 32421 559 32441
rect 559 32421 569 32441
rect 607 32421 631 32441
rect 631 32421 641 32441
rect 679 32421 703 32441
rect 703 32421 713 32441
rect 751 32421 775 32441
rect 775 32421 785 32441
rect 823 32421 843 32453
rect 843 32421 857 32453
rect 895 32421 915 32453
rect 915 32421 929 32453
rect -17 32373 17 32382
rect 75 32373 109 32382
rect 167 32373 201 32382
rect 259 32373 293 32382
rect 463 32373 497 32382
rect 535 32373 569 32382
rect 607 32373 641 32382
rect 679 32373 713 32382
rect 751 32373 785 32382
rect -17 32348 17 32373
rect 75 32348 89 32373
rect 89 32348 109 32373
rect 167 32348 199 32373
rect 199 32348 201 32373
rect 259 32348 271 32373
rect 271 32348 293 32373
rect 463 32348 487 32373
rect 487 32348 497 32373
rect 535 32348 559 32373
rect 559 32348 569 32373
rect 607 32348 631 32373
rect 631 32348 641 32373
rect 679 32348 703 32373
rect 703 32348 713 32373
rect 751 32348 775 32373
rect 775 32348 785 32373
rect 823 32369 857 32382
rect 895 32369 929 32382
rect 823 32348 843 32369
rect 843 32348 857 32369
rect 895 32348 915 32369
rect 915 32348 929 32369
rect -17 32305 17 32309
rect 75 32305 109 32309
rect 167 32305 201 32309
rect 259 32305 293 32309
rect 463 32305 497 32309
rect 535 32305 569 32309
rect 607 32305 641 32309
rect 679 32305 713 32309
rect 751 32305 785 32309
rect -17 32275 17 32305
rect 75 32275 89 32305
rect 89 32275 109 32305
rect 167 32275 199 32305
rect 199 32275 201 32305
rect 259 32275 271 32305
rect 271 32275 293 32305
rect 463 32275 487 32305
rect 487 32275 497 32305
rect 535 32275 559 32305
rect 559 32275 569 32305
rect 607 32275 631 32305
rect 631 32275 641 32305
rect 679 32275 703 32305
rect 703 32275 713 32305
rect 751 32275 775 32305
rect 775 32275 785 32305
rect 823 32285 857 32309
rect 895 32285 929 32309
rect 823 32275 843 32285
rect 843 32275 857 32285
rect 895 32275 915 32285
rect 915 32275 929 32285
rect -17 32203 17 32236
rect 75 32203 89 32236
rect 89 32203 109 32236
rect 167 32203 199 32236
rect 199 32203 201 32236
rect 259 32203 271 32236
rect 271 32203 293 32236
rect 463 32203 487 32236
rect 487 32203 497 32236
rect 535 32203 559 32236
rect 559 32203 569 32236
rect 607 32203 631 32236
rect 631 32203 641 32236
rect 679 32203 703 32236
rect 703 32203 713 32236
rect 751 32203 775 32236
rect 775 32203 785 32236
rect -17 32202 17 32203
rect 75 32202 109 32203
rect 167 32202 201 32203
rect 259 32202 293 32203
rect 463 32202 497 32203
rect 535 32202 569 32203
rect 607 32202 641 32203
rect 679 32202 713 32203
rect 751 32202 785 32203
rect 823 32202 857 32236
rect 895 32202 929 32236
rect -17 32135 17 32163
rect 75 32135 89 32163
rect 89 32135 109 32163
rect 167 32135 199 32163
rect 199 32135 201 32163
rect 259 32135 271 32163
rect 271 32135 293 32163
rect 463 32135 487 32163
rect 487 32135 497 32163
rect 535 32135 559 32163
rect 559 32135 569 32163
rect 607 32135 631 32163
rect 631 32135 641 32163
rect 679 32135 703 32163
rect 703 32135 713 32163
rect 751 32135 775 32163
rect 775 32135 785 32163
rect -17 32129 17 32135
rect 75 32129 109 32135
rect 167 32129 201 32135
rect 259 32129 293 32135
rect 463 32129 497 32135
rect 535 32129 569 32135
rect 607 32129 641 32135
rect 679 32129 713 32135
rect 751 32129 785 32135
rect 823 32129 857 32163
rect 895 32129 929 32163
rect -17 32067 17 32090
rect 75 32067 89 32090
rect 89 32067 109 32090
rect 167 32067 199 32090
rect 199 32067 201 32090
rect 259 32067 271 32090
rect 271 32067 293 32090
rect 463 32067 487 32090
rect 487 32067 497 32090
rect 535 32067 559 32090
rect 559 32067 569 32090
rect 607 32067 631 32090
rect 631 32067 641 32090
rect 679 32067 703 32090
rect 703 32067 713 32090
rect 751 32067 775 32090
rect 775 32067 785 32090
rect 823 32083 843 32090
rect 843 32083 857 32090
rect 895 32083 915 32090
rect 915 32083 929 32090
rect -17 32056 17 32067
rect 75 32056 109 32067
rect 167 32056 201 32067
rect 259 32056 293 32067
rect 463 32056 497 32067
rect 535 32056 569 32067
rect 607 32056 641 32067
rect 679 32056 713 32067
rect 751 32056 785 32067
rect 823 32056 857 32083
rect 895 32056 929 32083
rect -17 31999 17 32017
rect 75 31999 89 32017
rect 89 31999 109 32017
rect 167 31999 199 32017
rect 199 31999 201 32017
rect 259 31999 271 32017
rect 271 31999 293 32017
rect 463 31999 487 32017
rect 487 31999 497 32017
rect 535 31999 559 32017
rect 559 31999 569 32017
rect 607 31999 631 32017
rect 631 31999 641 32017
rect 679 31999 703 32017
rect 703 31999 713 32017
rect 751 31999 775 32017
rect 775 31999 785 32017
rect 823 31999 843 32017
rect 843 31999 857 32017
rect 895 31999 915 32017
rect 915 31999 929 32017
rect -17 31983 17 31999
rect 75 31983 109 31999
rect 167 31983 201 31999
rect 259 31983 293 31999
rect 463 31983 497 31999
rect 535 31983 569 31999
rect 607 31983 641 31999
rect 679 31983 713 31999
rect 751 31983 785 31999
rect 823 31983 857 31999
rect 895 31983 929 31999
rect -17 31931 17 31944
rect 75 31931 89 31944
rect 89 31931 109 31944
rect 167 31931 199 31944
rect 199 31931 201 31944
rect 259 31931 271 31944
rect 271 31931 293 31944
rect 463 31931 487 31944
rect 487 31931 497 31944
rect 535 31931 559 31944
rect 559 31931 569 31944
rect 607 31931 631 31944
rect 631 31931 641 31944
rect 679 31931 703 31944
rect 703 31931 713 31944
rect 751 31931 775 31944
rect 775 31931 785 31944
rect -17 31910 17 31931
rect 75 31910 109 31931
rect 167 31910 201 31931
rect 259 31910 293 31931
rect 463 31910 497 31931
rect 535 31910 569 31931
rect 607 31910 641 31931
rect 679 31910 713 31931
rect 751 31910 785 31931
rect 823 31915 843 31944
rect 843 31915 857 31944
rect 895 31915 915 31944
rect 915 31915 929 31944
rect 823 31910 857 31915
rect 895 31910 929 31915
rect -17 31863 17 31871
rect 75 31863 89 31871
rect 89 31863 109 31871
rect 167 31863 199 31871
rect 199 31863 201 31871
rect 259 31863 271 31871
rect 271 31863 293 31871
rect 463 31863 487 31871
rect 487 31863 497 31871
rect 535 31863 559 31871
rect 559 31863 569 31871
rect 607 31863 631 31871
rect 631 31863 641 31871
rect 679 31863 703 31871
rect 703 31863 713 31871
rect 751 31863 775 31871
rect 775 31863 785 31871
rect 823 31865 857 31871
rect 895 31865 929 31871
rect -17 31837 17 31863
rect 75 31837 109 31863
rect 167 31837 201 31863
rect 259 31837 293 31863
rect 463 31837 497 31863
rect 535 31837 569 31863
rect 607 31837 641 31863
rect 679 31837 713 31863
rect 751 31837 785 31863
rect 823 31837 843 31865
rect 843 31837 857 31865
rect 895 31837 915 31865
rect 915 31837 929 31865
rect -17 31795 17 31798
rect 75 31795 89 31798
rect 89 31795 109 31798
rect 167 31795 199 31798
rect 199 31795 201 31798
rect 259 31795 271 31798
rect 271 31795 293 31798
rect 463 31795 487 31798
rect 487 31795 497 31798
rect 535 31795 559 31798
rect 559 31795 569 31798
rect 607 31795 631 31798
rect 631 31795 641 31798
rect 679 31795 703 31798
rect 703 31795 713 31798
rect 751 31795 775 31798
rect 775 31795 785 31798
rect -17 31764 17 31795
rect 75 31764 109 31795
rect 167 31764 201 31795
rect 259 31764 293 31795
rect 463 31764 497 31795
rect 535 31764 569 31795
rect 607 31764 641 31795
rect 679 31764 713 31795
rect 751 31764 785 31795
rect 823 31781 857 31798
rect 895 31781 929 31798
rect 823 31764 843 31781
rect 843 31764 857 31781
rect 895 31764 915 31781
rect 915 31764 929 31781
rect -17 31693 17 31725
rect 75 31693 109 31725
rect 167 31693 201 31725
rect 259 31693 293 31725
rect 463 31693 497 31725
rect 535 31693 569 31725
rect 607 31693 641 31725
rect 679 31693 713 31725
rect 751 31693 785 31725
rect 823 31697 857 31725
rect 895 31697 929 31725
rect -17 31691 17 31693
rect 75 31691 89 31693
rect 89 31691 109 31693
rect 167 31691 199 31693
rect 199 31691 201 31693
rect 259 31691 271 31693
rect 271 31691 293 31693
rect 463 31691 487 31693
rect 487 31691 497 31693
rect 535 31691 559 31693
rect 559 31691 569 31693
rect 607 31691 631 31693
rect 631 31691 641 31693
rect 679 31691 703 31693
rect 703 31691 713 31693
rect 751 31691 775 31693
rect 775 31691 785 31693
rect 823 31691 843 31697
rect 843 31691 857 31697
rect 895 31691 915 31697
rect 915 31691 929 31697
rect -17 31625 17 31652
rect 75 31625 109 31652
rect 167 31625 201 31652
rect 259 31625 293 31652
rect 463 31625 497 31652
rect 535 31625 569 31652
rect 607 31625 641 31652
rect 679 31625 713 31652
rect 751 31625 785 31652
rect -17 31618 17 31625
rect 75 31618 89 31625
rect 89 31618 109 31625
rect 167 31618 199 31625
rect 199 31618 201 31625
rect 259 31618 271 31625
rect 271 31618 293 31625
rect 463 31618 487 31625
rect 487 31618 497 31625
rect 535 31618 559 31625
rect 559 31618 569 31625
rect 607 31618 631 31625
rect 631 31618 641 31625
rect 679 31618 703 31625
rect 703 31618 713 31625
rect 751 31618 775 31625
rect 775 31618 785 31625
rect 823 31618 857 31652
rect 895 31618 929 31652
rect -17 31557 17 31579
rect 75 31557 109 31579
rect 167 31557 201 31579
rect 259 31557 293 31579
rect 463 31557 497 31579
rect 535 31557 569 31579
rect 607 31557 641 31579
rect 679 31557 713 31579
rect 751 31557 785 31579
rect -17 31545 17 31557
rect 75 31545 89 31557
rect 89 31545 109 31557
rect 167 31545 199 31557
rect 199 31545 201 31557
rect 259 31545 271 31557
rect 271 31545 293 31557
rect 463 31545 487 31557
rect 487 31545 497 31557
rect 535 31545 559 31557
rect 559 31545 569 31557
rect 607 31545 631 31557
rect 631 31545 641 31557
rect 679 31545 703 31557
rect 703 31545 713 31557
rect 751 31545 775 31557
rect 775 31545 785 31557
rect 823 31545 857 31579
rect 895 31545 929 31579
rect -17 31489 17 31506
rect 75 31489 109 31506
rect 167 31489 201 31506
rect 259 31489 293 31506
rect 463 31489 497 31506
rect 535 31489 569 31506
rect 607 31489 641 31506
rect 679 31489 713 31506
rect 751 31489 785 31506
rect 823 31495 843 31506
rect 843 31495 857 31506
rect 895 31495 915 31506
rect 915 31495 929 31506
rect -17 31472 17 31489
rect 75 31472 89 31489
rect 89 31472 109 31489
rect 167 31472 199 31489
rect 199 31472 201 31489
rect 259 31472 271 31489
rect 271 31472 293 31489
rect 463 31472 487 31489
rect 487 31472 497 31489
rect 535 31472 559 31489
rect 559 31472 569 31489
rect 607 31472 631 31489
rect 631 31472 641 31489
rect 679 31472 703 31489
rect 703 31472 713 31489
rect 751 31472 775 31489
rect 775 31472 785 31489
rect 823 31472 857 31495
rect 895 31472 929 31495
rect -17 31421 17 31433
rect 75 31421 109 31433
rect 167 31421 201 31433
rect 259 31421 293 31433
rect 463 31421 497 31433
rect 535 31421 569 31433
rect 607 31421 641 31433
rect 679 31421 713 31433
rect 751 31421 785 31433
rect -17 31399 17 31421
rect 75 31399 89 31421
rect 89 31399 109 31421
rect 167 31399 199 31421
rect 199 31399 201 31421
rect 259 31399 271 31421
rect 271 31399 293 31421
rect 463 31399 487 31421
rect 487 31399 497 31421
rect 535 31399 559 31421
rect 559 31399 569 31421
rect 607 31399 631 31421
rect 631 31399 641 31421
rect 679 31399 703 31421
rect 703 31399 713 31421
rect 751 31399 775 31421
rect 775 31399 785 31421
rect 823 31411 843 31433
rect 843 31411 857 31433
rect 895 31411 915 31433
rect 915 31411 929 31433
rect 823 31399 857 31411
rect 895 31399 929 31411
rect -17 31353 17 31360
rect 75 31353 109 31360
rect 167 31353 201 31360
rect 259 31353 293 31360
rect 463 31353 497 31360
rect 535 31353 569 31360
rect 607 31353 641 31360
rect 679 31353 713 31360
rect 751 31353 785 31360
rect -17 31326 17 31353
rect 75 31326 89 31353
rect 89 31326 109 31353
rect 167 31326 199 31353
rect 199 31326 201 31353
rect 259 31326 271 31353
rect 271 31326 293 31353
rect 463 31326 487 31353
rect 487 31326 497 31353
rect 535 31326 559 31353
rect 559 31326 569 31353
rect 607 31326 631 31353
rect 631 31326 641 31353
rect 679 31326 703 31353
rect 703 31326 713 31353
rect 751 31326 775 31353
rect 775 31326 785 31353
rect 823 31327 843 31360
rect 843 31327 857 31360
rect 895 31327 915 31360
rect 915 31327 929 31360
rect 823 31326 857 31327
rect 895 31326 929 31327
rect -17 31285 17 31287
rect 75 31285 109 31287
rect 167 31285 201 31287
rect 259 31285 293 31287
rect 463 31285 497 31287
rect 535 31285 569 31287
rect 607 31285 641 31287
rect 679 31285 713 31287
rect 751 31285 785 31287
rect -17 31253 17 31285
rect 75 31253 89 31285
rect 89 31253 109 31285
rect 167 31253 199 31285
rect 199 31253 201 31285
rect 259 31253 271 31285
rect 271 31253 293 31285
rect 463 31253 487 31285
rect 487 31253 497 31285
rect 535 31253 559 31285
rect 559 31253 569 31285
rect 607 31253 631 31285
rect 631 31253 641 31285
rect 679 31253 703 31285
rect 703 31253 713 31285
rect 751 31253 775 31285
rect 775 31253 785 31285
rect 823 31277 857 31287
rect 895 31277 929 31287
rect 823 31253 843 31277
rect 843 31253 857 31277
rect 895 31253 915 31277
rect 915 31253 929 31277
rect -17 31183 17 31214
rect 75 31183 89 31214
rect 89 31183 109 31214
rect 167 31183 199 31214
rect 199 31183 201 31214
rect 259 31183 271 31214
rect 271 31183 293 31214
rect 463 31183 487 31214
rect 487 31183 497 31214
rect 535 31183 559 31214
rect 559 31183 569 31214
rect 607 31183 631 31214
rect 631 31183 641 31214
rect 679 31183 703 31214
rect 703 31183 713 31214
rect 751 31183 775 31214
rect 775 31183 785 31214
rect 823 31193 857 31214
rect 895 31193 929 31214
rect -17 31180 17 31183
rect 75 31180 109 31183
rect 167 31180 201 31183
rect 259 31180 293 31183
rect 463 31180 497 31183
rect 535 31180 569 31183
rect 607 31180 641 31183
rect 679 31180 713 31183
rect 751 31180 785 31183
rect 823 31180 843 31193
rect 843 31180 857 31193
rect 895 31180 915 31193
rect 915 31180 929 31193
rect -17 31115 17 31141
rect 75 31115 89 31141
rect 89 31115 109 31141
rect 167 31115 199 31141
rect 199 31115 201 31141
rect 259 31115 271 31141
rect 271 31115 293 31141
rect 463 31115 487 31141
rect 487 31115 497 31141
rect 535 31115 559 31141
rect 559 31115 569 31141
rect 607 31115 631 31141
rect 631 31115 641 31141
rect 679 31115 703 31141
rect 703 31115 713 31141
rect 751 31115 775 31141
rect 775 31115 785 31141
rect -17 31107 17 31115
rect 75 31107 109 31115
rect 167 31107 201 31115
rect 259 31107 293 31115
rect 463 31107 497 31115
rect 535 31107 569 31115
rect 607 31107 641 31115
rect 679 31107 713 31115
rect 751 31107 785 31115
rect 823 31109 857 31141
rect 895 31109 929 31141
rect 823 31107 843 31109
rect 843 31107 857 31109
rect 895 31107 915 31109
rect 915 31107 929 31109
rect -17 31047 17 31068
rect 75 31047 89 31068
rect 89 31047 109 31068
rect 167 31047 199 31068
rect 199 31047 201 31068
rect 259 31047 271 31068
rect 271 31047 293 31068
rect 463 31047 487 31068
rect 487 31047 497 31068
rect 535 31047 559 31068
rect 559 31047 569 31068
rect 607 31047 631 31068
rect 631 31047 641 31068
rect 679 31047 703 31068
rect 703 31047 713 31068
rect 751 31047 775 31068
rect 775 31047 785 31068
rect -17 31034 17 31047
rect 75 31034 109 31047
rect 167 31034 201 31047
rect 259 31034 293 31047
rect 463 31034 497 31047
rect 535 31034 569 31047
rect 607 31034 641 31047
rect 679 31034 713 31047
rect 751 31034 785 31047
rect 823 31034 857 31068
rect 895 31034 929 31068
rect -17 30979 17 30995
rect 75 30979 89 30995
rect 89 30979 109 30995
rect 167 30979 199 30995
rect 199 30979 201 30995
rect 259 30979 271 30995
rect 271 30979 293 30995
rect 463 30979 487 30995
rect 487 30979 497 30995
rect 535 30979 559 30995
rect 559 30979 569 30995
rect 607 30979 631 30995
rect 631 30979 641 30995
rect 679 30979 703 30995
rect 703 30979 713 30995
rect 751 30979 775 30995
rect 775 30979 785 30995
rect 823 30991 843 30995
rect 843 30991 857 30995
rect 895 30991 915 30995
rect 915 30991 929 30995
rect -17 30961 17 30979
rect 75 30961 109 30979
rect 167 30961 201 30979
rect 259 30961 293 30979
rect 463 30961 497 30979
rect 535 30961 569 30979
rect 607 30961 641 30979
rect 679 30961 713 30979
rect 751 30961 785 30979
rect 823 30961 857 30991
rect 895 30961 929 30991
rect -17 30911 17 30922
rect 75 30911 89 30922
rect 89 30911 109 30922
rect 167 30911 199 30922
rect 199 30911 201 30922
rect 259 30911 271 30922
rect 271 30911 293 30922
rect 463 30911 487 30922
rect 487 30911 497 30922
rect 535 30911 559 30922
rect 559 30911 569 30922
rect 607 30911 631 30922
rect 631 30911 641 30922
rect 679 30911 703 30922
rect 703 30911 713 30922
rect 751 30911 775 30922
rect 775 30911 785 30922
rect -17 30888 17 30911
rect 75 30888 109 30911
rect 167 30888 201 30911
rect 259 30888 293 30911
rect 463 30888 497 30911
rect 535 30888 569 30911
rect 607 30888 641 30911
rect 679 30888 713 30911
rect 751 30888 785 30911
rect 823 30907 843 30922
rect 843 30907 857 30922
rect 895 30907 915 30922
rect 915 30907 929 30922
rect 823 30888 857 30907
rect 895 30888 929 30907
rect -17 30843 17 30849
rect 75 30843 89 30849
rect 89 30843 109 30849
rect 167 30843 199 30849
rect 199 30843 201 30849
rect 259 30843 271 30849
rect 271 30843 293 30849
rect 463 30843 487 30849
rect 487 30843 497 30849
rect 535 30843 559 30849
rect 559 30843 569 30849
rect 607 30843 631 30849
rect 631 30843 641 30849
rect 679 30843 703 30849
rect 703 30843 713 30849
rect 751 30843 775 30849
rect 775 30843 785 30849
rect -17 30815 17 30843
rect 75 30815 109 30843
rect 167 30815 201 30843
rect 259 30815 293 30843
rect 463 30815 497 30843
rect 535 30815 569 30843
rect 607 30815 641 30843
rect 679 30815 713 30843
rect 751 30815 785 30843
rect 823 30823 843 30849
rect 843 30823 857 30849
rect 895 30823 915 30849
rect 915 30823 929 30849
rect 823 30815 857 30823
rect 895 30815 929 30823
rect -17 30775 17 30776
rect 75 30775 89 30776
rect 89 30775 109 30776
rect 167 30775 199 30776
rect 199 30775 201 30776
rect 259 30775 271 30776
rect 271 30775 293 30776
rect 463 30775 487 30776
rect 487 30775 497 30776
rect 535 30775 559 30776
rect 559 30775 569 30776
rect 607 30775 631 30776
rect 631 30775 641 30776
rect 679 30775 703 30776
rect 703 30775 713 30776
rect 751 30775 775 30776
rect 775 30775 785 30776
rect -17 30742 17 30775
rect 75 30742 109 30775
rect 167 30742 201 30775
rect 259 30742 293 30775
rect 463 30742 497 30775
rect 535 30742 569 30775
rect 607 30742 641 30775
rect 679 30742 713 30775
rect 751 30742 785 30775
rect 823 30773 857 30776
rect 895 30773 929 30776
rect 823 30742 843 30773
rect 843 30742 857 30773
rect 895 30742 915 30773
rect 915 30742 929 30773
rect -17 30673 17 30703
rect 75 30673 109 30703
rect 167 30673 201 30703
rect 259 30673 293 30703
rect 463 30673 497 30703
rect 535 30673 569 30703
rect 607 30673 641 30703
rect 679 30673 713 30703
rect 751 30673 785 30703
rect 823 30689 857 30703
rect 895 30689 929 30703
rect -17 30669 17 30673
rect 75 30669 89 30673
rect 89 30669 109 30673
rect 167 30669 199 30673
rect 199 30669 201 30673
rect 259 30669 271 30673
rect 271 30669 293 30673
rect 463 30669 487 30673
rect 487 30669 497 30673
rect 535 30669 559 30673
rect 559 30669 569 30673
rect 607 30669 631 30673
rect 631 30669 641 30673
rect 679 30669 703 30673
rect 703 30669 713 30673
rect 751 30669 775 30673
rect 775 30669 785 30673
rect 823 30669 843 30689
rect 843 30669 857 30689
rect 895 30669 915 30689
rect 915 30669 929 30689
rect -17 30605 17 30630
rect 75 30605 109 30630
rect 167 30605 201 30630
rect 259 30605 293 30630
rect 463 30605 497 30630
rect 535 30605 569 30630
rect 607 30605 641 30630
rect 679 30605 713 30630
rect 751 30605 785 30630
rect 823 30605 857 30630
rect 895 30605 929 30630
rect -17 30596 17 30605
rect 75 30596 89 30605
rect 89 30596 109 30605
rect 167 30596 199 30605
rect 199 30596 201 30605
rect 259 30596 271 30605
rect 271 30596 293 30605
rect 463 30596 487 30605
rect 487 30596 497 30605
rect 535 30596 559 30605
rect 559 30596 569 30605
rect 607 30596 631 30605
rect 631 30596 641 30605
rect 679 30596 703 30605
rect 703 30596 713 30605
rect 751 30596 775 30605
rect 775 30596 785 30605
rect 823 30596 843 30605
rect 843 30596 857 30605
rect 895 30596 915 30605
rect 915 30596 929 30605
rect -17 30537 17 30557
rect 75 30537 109 30557
rect 167 30537 201 30557
rect 259 30537 293 30557
rect 463 30537 497 30557
rect 535 30537 569 30557
rect 607 30537 641 30557
rect 679 30537 713 30557
rect 751 30537 785 30557
rect -17 30523 17 30537
rect 75 30523 89 30537
rect 89 30523 109 30537
rect 167 30523 199 30537
rect 199 30523 201 30537
rect 259 30523 271 30537
rect 271 30523 293 30537
rect 463 30523 487 30537
rect 487 30523 497 30537
rect 535 30523 559 30537
rect 559 30523 569 30537
rect 607 30523 631 30537
rect 631 30523 641 30537
rect 679 30523 703 30537
rect 703 30523 713 30537
rect 751 30523 775 30537
rect 775 30523 785 30537
rect 823 30523 857 30557
rect 895 30523 929 30557
rect -17 30469 17 30484
rect 75 30469 109 30484
rect 167 30469 201 30484
rect 259 30469 293 30484
rect 463 30469 497 30484
rect 535 30469 569 30484
rect 607 30469 641 30484
rect 679 30469 713 30484
rect 751 30469 785 30484
rect -17 30450 17 30469
rect 75 30450 89 30469
rect 89 30450 109 30469
rect 167 30450 199 30469
rect 199 30450 201 30469
rect 259 30450 271 30469
rect 271 30450 293 30469
rect 463 30450 487 30469
rect 487 30450 497 30469
rect 535 30450 559 30469
rect 559 30450 569 30469
rect 607 30450 631 30469
rect 631 30450 641 30469
rect 679 30450 703 30469
rect 703 30450 713 30469
rect 751 30450 775 30469
rect 775 30450 785 30469
rect 823 30450 857 30484
rect 895 30450 929 30484
rect -17 30401 17 30411
rect 75 30401 109 30411
rect 167 30401 201 30411
rect 259 30401 293 30411
rect 463 30401 497 30411
rect 535 30401 569 30411
rect 607 30401 641 30411
rect 679 30401 713 30411
rect 751 30401 785 30411
rect 823 30402 843 30411
rect 843 30402 857 30411
rect 895 30402 915 30411
rect 915 30402 929 30411
rect -17 30377 17 30401
rect 75 30377 89 30401
rect 89 30377 109 30401
rect 167 30377 199 30401
rect 199 30377 201 30401
rect 259 30377 271 30401
rect 271 30377 293 30401
rect 463 30377 487 30401
rect 487 30377 497 30401
rect 535 30377 559 30401
rect 559 30377 569 30401
rect 607 30377 631 30401
rect 631 30377 641 30401
rect 679 30377 703 30401
rect 703 30377 713 30401
rect 751 30377 775 30401
rect 775 30377 785 30401
rect 823 30377 857 30402
rect 895 30377 929 30402
rect -17 30333 17 30338
rect 75 30333 109 30338
rect 167 30333 201 30338
rect 259 30333 293 30338
rect 463 30333 497 30338
rect 535 30333 569 30338
rect 607 30333 641 30338
rect 679 30333 713 30338
rect 751 30333 785 30338
rect -17 30304 17 30333
rect 75 30304 89 30333
rect 89 30304 109 30333
rect 167 30304 199 30333
rect 199 30304 201 30333
rect 259 30304 271 30333
rect 271 30304 293 30333
rect 463 30304 487 30333
rect 487 30304 497 30333
rect 535 30304 559 30333
rect 559 30304 569 30333
rect 607 30304 631 30333
rect 631 30304 641 30333
rect 679 30304 703 30333
rect 703 30304 713 30333
rect 751 30304 775 30333
rect 775 30304 785 30333
rect 823 30317 843 30338
rect 843 30317 857 30338
rect 895 30317 915 30338
rect 915 30317 929 30338
rect 823 30304 857 30317
rect 895 30304 929 30317
rect -17 30231 17 30265
rect 75 30231 89 30265
rect 89 30231 109 30265
rect 167 30231 199 30265
rect 199 30231 201 30265
rect 259 30231 271 30265
rect 271 30231 293 30265
rect 463 30231 487 30265
rect 487 30231 497 30265
rect 535 30231 559 30265
rect 559 30231 569 30265
rect 607 30231 631 30265
rect 631 30231 641 30265
rect 679 30231 703 30265
rect 703 30231 713 30265
rect 751 30231 775 30265
rect 775 30231 785 30265
rect 823 30232 843 30265
rect 843 30232 857 30265
rect 895 30232 915 30265
rect 915 30232 929 30265
rect 823 30231 857 30232
rect 895 30231 929 30232
rect -17 30163 17 30192
rect 75 30163 89 30192
rect 89 30163 109 30192
rect 167 30163 199 30192
rect 199 30163 201 30192
rect 259 30163 271 30192
rect 271 30163 293 30192
rect 463 30163 487 30192
rect 487 30163 497 30192
rect 535 30163 559 30192
rect 559 30163 569 30192
rect 607 30163 631 30192
rect 631 30163 641 30192
rect 679 30163 703 30192
rect 703 30163 713 30192
rect 751 30163 775 30192
rect 775 30163 785 30192
rect 823 30181 857 30192
rect 895 30181 929 30192
rect -17 30158 17 30163
rect 75 30158 109 30163
rect 167 30158 201 30163
rect 259 30158 293 30163
rect 463 30158 497 30163
rect 535 30158 569 30163
rect 607 30158 641 30163
rect 679 30158 713 30163
rect 751 30158 785 30163
rect 823 30158 843 30181
rect 843 30158 857 30181
rect 895 30158 915 30181
rect 915 30158 929 30181
rect -17 30095 17 30119
rect 75 30095 89 30119
rect 89 30095 109 30119
rect 167 30095 199 30119
rect 199 30095 201 30119
rect 259 30095 271 30119
rect 271 30095 293 30119
rect 463 30095 487 30119
rect 487 30095 497 30119
rect 535 30095 559 30119
rect 559 30095 569 30119
rect 607 30095 631 30119
rect 631 30095 641 30119
rect 679 30095 703 30119
rect 703 30095 713 30119
rect 751 30095 775 30119
rect 775 30095 785 30119
rect 823 30096 857 30119
rect 895 30096 929 30119
rect -17 30085 17 30095
rect 75 30085 109 30095
rect 167 30085 201 30095
rect 259 30085 293 30095
rect 463 30085 497 30095
rect 535 30085 569 30095
rect 607 30085 641 30095
rect 679 30085 713 30095
rect 751 30085 785 30095
rect 823 30085 843 30096
rect 843 30085 857 30096
rect 895 30085 915 30096
rect 915 30085 929 30096
rect -17 30027 17 30046
rect 75 30027 89 30046
rect 89 30027 109 30046
rect 167 30027 199 30046
rect 199 30027 201 30046
rect 259 30027 271 30046
rect 271 30027 293 30046
rect 463 30027 487 30046
rect 487 30027 497 30046
rect 535 30027 559 30046
rect 559 30027 569 30046
rect 607 30027 631 30046
rect 631 30027 641 30046
rect 679 30027 703 30046
rect 703 30027 713 30046
rect 751 30027 775 30046
rect 775 30027 785 30046
rect -17 30012 17 30027
rect 75 30012 109 30027
rect 167 30012 201 30027
rect 259 30012 293 30027
rect 463 30012 497 30027
rect 535 30012 569 30027
rect 607 30012 641 30027
rect 679 30012 713 30027
rect 751 30012 785 30027
rect 823 30012 857 30046
rect 895 30012 929 30046
rect -17 29959 17 29973
rect 75 29959 89 29973
rect 89 29959 109 29973
rect 167 29959 199 29973
rect 199 29959 201 29973
rect 259 29959 271 29973
rect 271 29959 293 29973
rect 463 29959 487 29973
rect 487 29959 497 29973
rect 535 29959 559 29973
rect 559 29959 569 29973
rect 607 29959 631 29973
rect 631 29959 641 29973
rect 679 29959 703 29973
rect 703 29959 713 29973
rect 751 29959 775 29973
rect 775 29959 785 29973
rect -17 29939 17 29959
rect 75 29939 109 29959
rect 167 29939 201 29959
rect 259 29939 293 29959
rect 463 29939 497 29959
rect 535 29939 569 29959
rect 607 29939 641 29959
rect 679 29939 713 29959
rect 751 29939 785 29959
rect 823 29939 857 29973
rect 895 29939 929 29973
rect -17 29891 17 29900
rect 75 29891 89 29900
rect 89 29891 109 29900
rect 167 29891 199 29900
rect 199 29891 201 29900
rect 259 29891 271 29900
rect 271 29891 293 29900
rect 463 29891 487 29900
rect 487 29891 497 29900
rect 535 29891 559 29900
rect 559 29891 569 29900
rect 607 29891 631 29900
rect 631 29891 641 29900
rect 679 29891 703 29900
rect 703 29891 713 29900
rect 751 29891 775 29900
rect 775 29891 785 29900
rect 823 29892 843 29900
rect 843 29892 857 29900
rect 895 29892 915 29900
rect 915 29892 929 29900
rect -17 29866 17 29891
rect 75 29866 109 29891
rect 167 29866 201 29891
rect 259 29866 293 29891
rect 463 29866 497 29891
rect 535 29866 569 29891
rect 607 29866 641 29891
rect 679 29866 713 29891
rect 751 29866 785 29891
rect 823 29866 857 29892
rect 895 29866 929 29892
rect -17 29823 17 29827
rect 75 29823 89 29827
rect 89 29823 109 29827
rect 167 29823 199 29827
rect 199 29823 201 29827
rect 259 29823 271 29827
rect 271 29823 293 29827
rect 463 29823 487 29827
rect 487 29823 497 29827
rect 535 29823 559 29827
rect 559 29823 569 29827
rect 607 29823 631 29827
rect 631 29823 641 29827
rect 679 29823 703 29827
rect 703 29823 713 29827
rect 751 29823 775 29827
rect 775 29823 785 29827
rect -17 29793 17 29823
rect 75 29793 109 29823
rect 167 29793 201 29823
rect 259 29793 293 29823
rect 463 29793 497 29823
rect 535 29793 569 29823
rect 607 29793 641 29823
rect 679 29793 713 29823
rect 751 29793 785 29823
rect 823 29807 843 29827
rect 843 29807 857 29827
rect 895 29807 915 29827
rect 915 29807 929 29827
rect 823 29793 857 29807
rect 895 29793 929 29807
rect -17 29721 17 29754
rect 75 29721 109 29754
rect 167 29721 201 29754
rect 259 29721 293 29754
rect 463 29721 497 29754
rect 535 29721 569 29754
rect 607 29721 641 29754
rect 679 29721 713 29754
rect 751 29721 785 29754
rect 823 29722 843 29754
rect 843 29722 857 29754
rect 895 29722 915 29754
rect 915 29722 929 29754
rect -17 29720 17 29721
rect 75 29720 89 29721
rect 89 29720 109 29721
rect 167 29720 199 29721
rect 199 29720 201 29721
rect 259 29720 271 29721
rect 271 29720 293 29721
rect 463 29720 487 29721
rect 487 29720 497 29721
rect 535 29720 559 29721
rect 559 29720 569 29721
rect 607 29720 631 29721
rect 631 29720 641 29721
rect 679 29720 703 29721
rect 703 29720 713 29721
rect 751 29720 775 29721
rect 775 29720 785 29721
rect 823 29720 857 29722
rect 895 29720 929 29722
rect -17 29652 17 29681
rect 75 29652 109 29681
rect 167 29652 201 29681
rect 259 29652 293 29681
rect 463 29652 497 29681
rect 535 29652 569 29681
rect 607 29652 641 29681
rect 679 29652 713 29681
rect 751 29652 785 29681
rect 823 29671 857 29681
rect 895 29671 929 29681
rect -17 29647 17 29652
rect 75 29647 89 29652
rect 89 29647 109 29652
rect 167 29647 199 29652
rect 199 29647 201 29652
rect 259 29647 271 29652
rect 271 29647 293 29652
rect 463 29647 487 29652
rect 487 29647 497 29652
rect 535 29647 559 29652
rect 559 29647 569 29652
rect 607 29647 631 29652
rect 631 29647 641 29652
rect 679 29647 703 29652
rect 703 29647 713 29652
rect 751 29647 775 29652
rect 775 29647 785 29652
rect 823 29647 843 29671
rect 843 29647 857 29671
rect 895 29647 915 29671
rect 915 29647 929 29671
rect -17 29583 17 29608
rect 75 29583 109 29608
rect 167 29583 201 29608
rect 259 29583 293 29608
rect 463 29583 497 29608
rect 535 29583 569 29608
rect 607 29583 641 29608
rect 679 29583 713 29608
rect 751 29583 785 29608
rect 823 29586 857 29608
rect 895 29586 929 29608
rect -17 29574 17 29583
rect 75 29574 89 29583
rect 89 29574 109 29583
rect 167 29574 199 29583
rect 199 29574 201 29583
rect 259 29574 271 29583
rect 271 29574 293 29583
rect 463 29574 487 29583
rect 487 29574 497 29583
rect 535 29574 559 29583
rect 559 29574 569 29583
rect 607 29574 631 29583
rect 631 29574 641 29583
rect 679 29574 703 29583
rect 703 29574 713 29583
rect 751 29574 775 29583
rect 775 29574 785 29583
rect 823 29574 843 29586
rect 843 29574 857 29586
rect 895 29574 915 29586
rect 915 29574 929 29586
rect -17 29514 17 29535
rect 75 29514 109 29535
rect 167 29514 201 29535
rect 259 29514 293 29535
rect 463 29514 497 29535
rect 535 29514 569 29535
rect 607 29514 641 29535
rect 679 29514 713 29535
rect 751 29514 785 29535
rect -17 29501 17 29514
rect 75 29501 89 29514
rect 89 29501 109 29514
rect 167 29501 199 29514
rect 199 29501 201 29514
rect 259 29501 271 29514
rect 271 29501 293 29514
rect 463 29501 487 29514
rect 487 29501 497 29514
rect 535 29501 559 29514
rect 559 29501 569 29514
rect 607 29501 631 29514
rect 631 29501 641 29514
rect 679 29501 703 29514
rect 703 29501 713 29514
rect 751 29501 775 29514
rect 775 29501 785 29514
rect 823 29501 857 29535
rect 895 29501 929 29535
rect -17 29445 17 29462
rect 75 29445 109 29462
rect 167 29445 201 29462
rect 259 29445 293 29462
rect 463 29445 497 29462
rect 535 29445 569 29462
rect 607 29445 641 29462
rect 679 29445 713 29462
rect 751 29445 785 29462
rect -17 29428 17 29445
rect 75 29428 89 29445
rect 89 29428 109 29445
rect 167 29428 199 29445
rect 199 29428 201 29445
rect 259 29428 271 29445
rect 271 29428 293 29445
rect 463 29428 487 29445
rect 487 29428 497 29445
rect 535 29428 559 29445
rect 559 29428 569 29445
rect 607 29428 631 29445
rect 631 29428 641 29445
rect 679 29428 703 29445
rect 703 29428 713 29445
rect 751 29428 775 29445
rect 775 29428 785 29445
rect 823 29428 857 29462
rect 895 29428 929 29462
rect -17 29376 17 29389
rect 75 29376 109 29389
rect 167 29376 201 29389
rect 259 29376 293 29389
rect 463 29376 497 29389
rect 535 29376 569 29389
rect 607 29376 641 29389
rect 679 29376 713 29389
rect 751 29376 785 29389
rect 823 29382 843 29389
rect 843 29382 857 29389
rect 895 29382 915 29389
rect 915 29382 929 29389
rect -17 29355 17 29376
rect 75 29355 89 29376
rect 89 29355 109 29376
rect 167 29355 199 29376
rect 199 29355 201 29376
rect 259 29355 271 29376
rect 271 29355 293 29376
rect 463 29355 487 29376
rect 487 29355 497 29376
rect 535 29355 559 29376
rect 559 29355 569 29376
rect 607 29355 631 29376
rect 631 29355 641 29376
rect 679 29355 703 29376
rect 703 29355 713 29376
rect 751 29355 775 29376
rect 775 29355 785 29376
rect 823 29355 857 29382
rect 895 29355 929 29382
rect -17 29307 17 29316
rect 75 29307 109 29316
rect 167 29307 201 29316
rect 259 29307 293 29316
rect 463 29307 497 29316
rect 535 29307 569 29316
rect 607 29307 641 29316
rect 679 29307 713 29316
rect 751 29307 785 29316
rect -17 29282 17 29307
rect 75 29282 89 29307
rect 89 29282 109 29307
rect 167 29282 199 29307
rect 199 29282 201 29307
rect 259 29282 271 29307
rect 271 29282 293 29307
rect 463 29282 487 29307
rect 487 29282 497 29307
rect 535 29282 559 29307
rect 559 29282 569 29307
rect 607 29282 631 29307
rect 631 29282 641 29307
rect 679 29282 703 29307
rect 703 29282 713 29307
rect 751 29282 775 29307
rect 775 29282 785 29307
rect 823 29297 843 29316
rect 843 29297 857 29316
rect 895 29297 915 29316
rect 915 29297 929 29316
rect 823 29282 857 29297
rect 895 29282 929 29297
rect -17 29238 17 29243
rect 75 29238 109 29243
rect 167 29238 201 29243
rect 259 29238 293 29243
rect 463 29238 497 29243
rect 535 29238 569 29243
rect 607 29238 641 29243
rect 679 29238 713 29243
rect 751 29238 785 29243
rect -17 29209 17 29238
rect 75 29209 89 29238
rect 89 29209 109 29238
rect 167 29209 199 29238
rect 199 29209 201 29238
rect 259 29209 271 29238
rect 271 29209 293 29238
rect 463 29209 487 29238
rect 487 29209 497 29238
rect 535 29209 559 29238
rect 559 29209 569 29238
rect 607 29209 631 29238
rect 631 29209 641 29238
rect 679 29209 703 29238
rect 703 29209 713 29238
rect 751 29209 775 29238
rect 775 29209 785 29238
rect 823 29212 843 29243
rect 843 29212 857 29243
rect 895 29212 915 29243
rect 915 29212 929 29243
rect 823 29209 857 29212
rect 895 29209 929 29212
rect -17 29169 17 29170
rect 75 29169 109 29170
rect 167 29169 201 29170
rect 259 29169 293 29170
rect 463 29169 497 29170
rect 535 29169 569 29170
rect 607 29169 641 29170
rect 679 29169 713 29170
rect 751 29169 785 29170
rect -17 29136 17 29169
rect 75 29136 89 29169
rect 89 29136 109 29169
rect 167 29136 199 29169
rect 199 29136 201 29169
rect 259 29136 271 29169
rect 271 29136 293 29169
rect 463 29136 487 29169
rect 487 29136 497 29169
rect 535 29136 559 29169
rect 559 29136 569 29169
rect 607 29136 631 29169
rect 631 29136 641 29169
rect 679 29136 703 29169
rect 703 29136 713 29169
rect 751 29136 775 29169
rect 775 29136 785 29169
rect 823 29161 857 29170
rect 895 29161 929 29170
rect 823 29136 843 29161
rect 843 29136 857 29161
rect 895 29136 915 29161
rect 915 29136 929 29161
rect -17 29066 17 29097
rect 75 29066 89 29097
rect 89 29066 109 29097
rect 167 29066 199 29097
rect 199 29066 201 29097
rect 259 29066 271 29097
rect 271 29066 293 29097
rect 463 29066 487 29097
rect 487 29066 497 29097
rect 535 29066 559 29097
rect 559 29066 569 29097
rect 607 29066 631 29097
rect 631 29066 641 29097
rect 679 29066 703 29097
rect 703 29066 713 29097
rect 751 29066 775 29097
rect 775 29066 785 29097
rect 823 29076 857 29097
rect 895 29076 929 29097
rect -17 29063 17 29066
rect 75 29063 109 29066
rect 167 29063 201 29066
rect 259 29063 293 29066
rect 463 29063 497 29066
rect 535 29063 569 29066
rect 607 29063 641 29066
rect 679 29063 713 29066
rect 751 29063 785 29066
rect 823 29063 843 29076
rect 843 29063 857 29076
rect 895 29063 915 29076
rect 915 29063 929 29076
rect -17 27986 17 27998
rect 75 27986 109 27998
rect 167 27986 201 27998
rect 259 27986 293 27998
rect -17 27964 17 27986
rect 75 27964 89 27986
rect 89 27964 109 27986
rect 167 27964 199 27986
rect 199 27964 201 27986
rect 259 27964 271 27986
rect 271 27964 293 27986
rect 463 27952 487 27978
rect 487 27952 497 27978
rect 535 27952 559 27978
rect 559 27952 569 27978
rect 607 27952 631 27978
rect 631 27952 641 27978
rect 679 27952 703 27978
rect 703 27952 713 27978
rect 751 27952 775 27978
rect 775 27952 785 27978
rect 823 27976 843 27978
rect 843 27976 857 27978
rect 895 27976 915 27978
rect 915 27976 929 27978
rect 463 27944 497 27952
rect 535 27944 569 27952
rect 607 27944 641 27952
rect 679 27944 713 27952
rect 751 27944 785 27952
rect 823 27944 857 27976
rect 895 27944 929 27976
rect -17 27917 17 27925
rect 75 27917 109 27925
rect 167 27917 201 27925
rect 259 27917 293 27925
rect -17 27891 17 27917
rect 75 27891 89 27917
rect 89 27891 109 27917
rect 167 27891 199 27917
rect 199 27891 201 27917
rect 259 27891 271 27917
rect 271 27891 293 27917
rect 463 27883 487 27903
rect 487 27883 497 27903
rect 535 27883 559 27903
rect 559 27883 569 27903
rect 607 27883 631 27903
rect 631 27883 641 27903
rect 679 27883 703 27903
rect 703 27883 713 27903
rect 751 27883 775 27903
rect 775 27883 785 27903
rect 463 27869 497 27883
rect 535 27869 569 27883
rect 607 27869 641 27883
rect 679 27869 713 27883
rect 751 27869 785 27883
rect 823 27874 857 27903
rect 895 27874 929 27903
rect 823 27869 843 27874
rect 843 27869 857 27874
rect 895 27869 915 27874
rect 915 27869 929 27874
rect -17 27848 17 27852
rect 75 27848 109 27852
rect 167 27848 201 27852
rect 259 27848 293 27852
rect -17 27818 17 27848
rect 75 27818 89 27848
rect 89 27818 109 27848
rect 167 27818 199 27848
rect 199 27818 201 27848
rect 259 27818 271 27848
rect 271 27818 293 27848
rect 463 27814 487 27828
rect 487 27814 497 27828
rect 535 27814 559 27828
rect 559 27814 569 27828
rect 607 27814 631 27828
rect 631 27814 641 27828
rect 679 27814 703 27828
rect 703 27814 713 27828
rect 751 27814 775 27828
rect 775 27814 785 27828
rect 463 27794 497 27814
rect 535 27794 569 27814
rect 607 27794 641 27814
rect 679 27794 713 27814
rect 751 27794 785 27814
rect 823 27806 857 27828
rect 895 27806 929 27828
rect 823 27794 843 27806
rect 843 27794 857 27806
rect 895 27794 915 27806
rect 915 27794 929 27806
rect -17 27745 17 27779
rect 75 27745 89 27779
rect 89 27745 109 27779
rect 167 27745 199 27779
rect 199 27745 201 27779
rect 259 27745 271 27779
rect 271 27745 293 27779
rect 463 27745 487 27753
rect 487 27745 497 27753
rect 535 27745 559 27753
rect 559 27745 569 27753
rect 607 27745 631 27753
rect 631 27745 641 27753
rect 679 27745 703 27753
rect 703 27745 713 27753
rect 751 27745 775 27753
rect 775 27745 785 27753
rect 463 27719 497 27745
rect 535 27719 569 27745
rect 607 27719 641 27745
rect 679 27719 713 27745
rect 751 27719 785 27745
rect 823 27738 857 27753
rect 895 27738 929 27753
rect 823 27719 843 27738
rect 843 27719 857 27738
rect 895 27719 915 27738
rect 915 27719 929 27738
rect -17 27676 17 27706
rect 75 27676 89 27706
rect 89 27676 109 27706
rect 167 27676 199 27706
rect 199 27676 201 27706
rect 259 27676 271 27706
rect 271 27676 293 27706
rect 463 27676 487 27678
rect 487 27676 497 27678
rect 535 27676 559 27678
rect 559 27676 569 27678
rect 607 27676 631 27678
rect 631 27676 641 27678
rect 679 27676 703 27678
rect 703 27676 713 27678
rect 751 27676 775 27678
rect 775 27676 785 27678
rect -17 27672 17 27676
rect 75 27672 109 27676
rect 167 27672 201 27676
rect 259 27672 293 27676
rect 463 27644 497 27676
rect 535 27644 569 27676
rect 607 27644 641 27676
rect 679 27644 713 27676
rect 751 27644 785 27676
rect 823 27670 857 27678
rect 895 27670 929 27678
rect 823 27644 843 27670
rect 843 27644 857 27670
rect 895 27644 915 27670
rect 915 27644 929 27670
rect -17 27607 17 27633
rect 75 27607 89 27633
rect 89 27607 109 27633
rect 167 27607 199 27633
rect 199 27607 201 27633
rect 259 27607 271 27633
rect 271 27607 293 27633
rect -17 27599 17 27607
rect 75 27599 109 27607
rect 167 27599 201 27607
rect 259 27599 293 27607
rect 463 27572 497 27603
rect 535 27572 569 27603
rect 607 27572 641 27603
rect 679 27572 713 27603
rect 751 27572 785 27603
rect 823 27602 857 27603
rect 895 27602 929 27603
rect -17 27538 17 27560
rect 75 27538 89 27560
rect 89 27538 109 27560
rect 167 27538 199 27560
rect 199 27538 201 27560
rect 259 27538 271 27560
rect 271 27538 293 27560
rect 463 27569 487 27572
rect 487 27569 497 27572
rect 535 27569 559 27572
rect 559 27569 569 27572
rect 607 27569 631 27572
rect 631 27569 641 27572
rect 679 27569 703 27572
rect 703 27569 713 27572
rect 751 27569 775 27572
rect 775 27569 785 27572
rect 823 27569 843 27602
rect 843 27569 857 27602
rect 895 27569 915 27602
rect 915 27569 929 27602
rect -17 27526 17 27538
rect 75 27526 109 27538
rect 167 27526 201 27538
rect 259 27526 293 27538
rect 463 27503 497 27528
rect 535 27503 569 27528
rect 607 27503 641 27528
rect 679 27503 713 27528
rect 751 27503 785 27528
rect -17 27469 17 27487
rect 75 27469 89 27487
rect 89 27469 109 27487
rect 167 27469 199 27487
rect 199 27469 201 27487
rect 259 27469 271 27487
rect 271 27469 293 27487
rect 463 27494 487 27503
rect 487 27494 497 27503
rect 535 27494 559 27503
rect 559 27494 569 27503
rect 607 27494 631 27503
rect 631 27494 641 27503
rect 679 27494 703 27503
rect 703 27494 713 27503
rect 751 27494 775 27503
rect 775 27494 785 27503
rect 823 27500 843 27528
rect 843 27500 857 27528
rect 895 27500 915 27528
rect 915 27500 929 27528
rect 823 27494 857 27500
rect 895 27494 929 27500
rect -17 27453 17 27469
rect 75 27453 109 27469
rect 167 27453 201 27469
rect 259 27453 293 27469
rect 463 27434 497 27453
rect 535 27434 569 27453
rect 607 27434 641 27453
rect 679 27434 713 27453
rect 751 27434 785 27453
rect -17 27400 17 27414
rect 75 27400 89 27414
rect 89 27400 109 27414
rect 167 27400 199 27414
rect 199 27400 201 27414
rect 259 27400 271 27414
rect 271 27400 293 27414
rect 463 27419 487 27434
rect 487 27419 497 27434
rect 535 27419 559 27434
rect 559 27419 569 27434
rect 607 27419 631 27434
rect 631 27419 641 27434
rect 679 27419 703 27434
rect 703 27419 713 27434
rect 751 27419 775 27434
rect 775 27419 785 27434
rect 823 27432 843 27453
rect 843 27432 857 27453
rect 895 27432 915 27453
rect 915 27432 929 27453
rect 823 27419 857 27432
rect 895 27419 929 27432
rect -17 27380 17 27400
rect 75 27380 109 27400
rect 167 27380 201 27400
rect 259 27380 293 27400
rect 463 27365 497 27378
rect 535 27365 569 27378
rect 607 27365 641 27378
rect 679 27365 713 27378
rect 751 27365 785 27378
rect -17 27331 17 27341
rect 75 27331 89 27341
rect 89 27331 109 27341
rect 167 27331 199 27341
rect 199 27331 201 27341
rect 259 27331 271 27341
rect 271 27331 293 27341
rect 463 27344 487 27365
rect 487 27344 497 27365
rect 535 27344 559 27365
rect 559 27344 569 27365
rect 607 27344 631 27365
rect 631 27344 641 27365
rect 679 27344 703 27365
rect 703 27344 713 27365
rect 751 27344 775 27365
rect 775 27344 785 27365
rect 823 27364 843 27378
rect 843 27364 857 27378
rect 895 27364 915 27378
rect 915 27364 929 27378
rect 823 27344 857 27364
rect 895 27344 929 27364
rect -17 27307 17 27331
rect 75 27307 109 27331
rect 167 27307 201 27331
rect 259 27307 293 27331
rect 463 27296 497 27303
rect 535 27296 569 27303
rect 607 27296 641 27303
rect 679 27296 713 27303
rect 751 27296 785 27303
rect 823 27296 843 27303
rect 843 27296 857 27303
rect 895 27296 915 27303
rect 915 27296 929 27303
rect -17 27262 17 27268
rect 75 27262 89 27268
rect 89 27262 109 27268
rect 167 27262 199 27268
rect 199 27262 201 27268
rect 259 27262 271 27268
rect 271 27262 293 27268
rect 463 27269 487 27296
rect 487 27269 497 27296
rect 535 27269 559 27296
rect 559 27269 569 27296
rect 607 27269 631 27296
rect 631 27269 641 27296
rect 679 27269 703 27296
rect 703 27269 713 27296
rect 751 27269 775 27296
rect 775 27269 785 27296
rect 823 27269 857 27296
rect 895 27269 929 27296
rect -17 27234 17 27262
rect 75 27234 109 27262
rect 167 27234 201 27262
rect 259 27234 293 27262
rect 463 27227 497 27228
rect 535 27227 569 27228
rect 607 27227 641 27228
rect 679 27227 713 27228
rect 751 27227 785 27228
rect -17 27193 17 27195
rect 75 27193 89 27195
rect 89 27193 109 27195
rect 167 27193 199 27195
rect 199 27193 201 27195
rect 259 27193 271 27195
rect 271 27193 293 27195
rect 463 27194 487 27227
rect 487 27194 497 27227
rect 535 27194 559 27227
rect 559 27194 569 27227
rect 607 27194 631 27227
rect 631 27194 641 27227
rect 679 27194 703 27227
rect 703 27194 713 27227
rect 751 27194 775 27227
rect 775 27194 785 27227
rect 823 27194 857 27228
rect 895 27194 929 27228
rect -17 27161 17 27193
rect 75 27161 109 27193
rect 167 27161 201 27193
rect 259 27161 293 27193
rect 463 27124 487 27153
rect 487 27124 497 27153
rect 535 27124 559 27153
rect 559 27124 569 27153
rect 607 27124 631 27153
rect 631 27124 641 27153
rect 679 27124 703 27153
rect 703 27124 713 27153
rect 751 27124 775 27153
rect 775 27124 785 27153
rect 823 27126 857 27153
rect 895 27126 929 27153
rect -17 27089 17 27122
rect 75 27089 109 27122
rect 167 27089 201 27122
rect 259 27089 293 27122
rect 463 27119 497 27124
rect 535 27119 569 27124
rect 607 27119 641 27124
rect 679 27119 713 27124
rect 751 27119 785 27124
rect 823 27119 843 27126
rect 843 27119 857 27126
rect 895 27119 915 27126
rect 915 27119 929 27126
rect -17 27088 17 27089
rect 75 27088 89 27089
rect 89 27088 109 27089
rect 167 27088 199 27089
rect 199 27088 201 27089
rect 259 27088 271 27089
rect 271 27088 293 27089
rect 463 27055 487 27079
rect 487 27055 497 27079
rect 535 27055 559 27079
rect 559 27055 569 27079
rect 607 27055 631 27079
rect 631 27055 641 27079
rect 679 27055 703 27079
rect 703 27055 713 27079
rect 751 27055 775 27079
rect 775 27055 785 27079
rect 823 27058 857 27079
rect 895 27058 929 27079
rect -17 27020 17 27049
rect 75 27020 109 27049
rect 167 27020 201 27049
rect 259 27020 293 27049
rect 463 27045 497 27055
rect 535 27045 569 27055
rect 607 27045 641 27055
rect 679 27045 713 27055
rect 751 27045 785 27055
rect 823 27045 843 27058
rect 843 27045 857 27058
rect 895 27045 915 27058
rect 915 27045 929 27058
rect -17 27015 17 27020
rect 75 27015 89 27020
rect 89 27015 109 27020
rect 167 27015 199 27020
rect 199 27015 201 27020
rect 259 27015 271 27020
rect 271 27015 293 27020
rect 463 26986 487 27005
rect 487 26986 497 27005
rect 535 26986 559 27005
rect 559 26986 569 27005
rect 607 26986 631 27005
rect 631 26986 641 27005
rect 679 26986 703 27005
rect 703 26986 713 27005
rect 751 26986 775 27005
rect 775 26986 785 27005
rect 823 26990 857 27005
rect 895 26990 929 27005
rect -17 26951 17 26976
rect 75 26951 109 26976
rect 167 26951 201 26976
rect 259 26951 293 26976
rect 463 26971 497 26986
rect 535 26971 569 26986
rect 607 26971 641 26986
rect 679 26971 713 26986
rect 751 26971 785 26986
rect 823 26971 843 26990
rect 843 26971 857 26990
rect 895 26971 915 26990
rect 915 26971 929 26990
rect -17 26942 17 26951
rect 75 26942 89 26951
rect 89 26942 109 26951
rect 167 26942 199 26951
rect 199 26942 201 26951
rect 259 26942 271 26951
rect 271 26942 293 26951
rect 463 26917 487 26931
rect 487 26917 497 26931
rect 535 26917 559 26931
rect 559 26917 569 26931
rect 607 26917 631 26931
rect 631 26917 641 26931
rect 679 26917 703 26931
rect 703 26917 713 26931
rect 751 26917 775 26931
rect 775 26917 785 26931
rect 823 26922 857 26931
rect 895 26922 929 26931
rect -17 26882 17 26903
rect 75 26882 109 26903
rect 167 26882 201 26903
rect 259 26882 293 26903
rect 463 26897 497 26917
rect 535 26897 569 26917
rect 607 26897 641 26917
rect 679 26897 713 26917
rect 751 26897 785 26917
rect 823 26897 843 26922
rect 843 26897 857 26922
rect 895 26897 915 26922
rect 915 26897 929 26922
rect -17 26869 17 26882
rect 75 26869 89 26882
rect 89 26869 109 26882
rect 167 26869 199 26882
rect 199 26869 201 26882
rect 259 26869 271 26882
rect 271 26869 293 26882
rect 463 26848 487 26857
rect 487 26848 497 26857
rect 535 26848 559 26857
rect 559 26848 569 26857
rect 607 26848 631 26857
rect 631 26848 641 26857
rect 679 26848 703 26857
rect 703 26848 713 26857
rect 751 26848 775 26857
rect 775 26848 785 26857
rect 823 26854 857 26857
rect 895 26854 929 26857
rect -17 26813 17 26830
rect 75 26813 109 26830
rect 167 26813 201 26830
rect 259 26813 293 26830
rect 463 26823 497 26848
rect 535 26823 569 26848
rect 607 26823 641 26848
rect 679 26823 713 26848
rect 751 26823 785 26848
rect 823 26823 843 26854
rect 843 26823 857 26854
rect 895 26823 915 26854
rect 915 26823 929 26854
rect -17 26796 17 26813
rect 75 26796 89 26813
rect 89 26796 109 26813
rect 167 26796 199 26813
rect 199 26796 201 26813
rect 259 26796 271 26813
rect 271 26796 293 26813
rect 463 26779 487 26783
rect 487 26779 497 26783
rect 535 26779 559 26783
rect 559 26779 569 26783
rect 607 26779 631 26783
rect 631 26779 641 26783
rect 679 26779 703 26783
rect 703 26779 713 26783
rect 751 26779 775 26783
rect 775 26779 785 26783
rect -17 26744 17 26757
rect 75 26744 109 26757
rect 167 26744 201 26757
rect 259 26744 293 26757
rect 463 26749 497 26779
rect 535 26749 569 26779
rect 607 26749 641 26779
rect 679 26749 713 26779
rect 751 26749 785 26779
rect 823 26751 843 26783
rect 843 26751 857 26783
rect 895 26751 915 26783
rect 915 26751 929 26783
rect 823 26749 857 26751
rect 895 26749 929 26751
rect -17 26723 17 26744
rect 75 26723 89 26744
rect 89 26723 109 26744
rect 167 26723 199 26744
rect 199 26723 201 26744
rect 259 26723 271 26744
rect 271 26723 293 26744
rect -17 26675 17 26684
rect 75 26675 109 26684
rect 167 26675 201 26684
rect 259 26675 293 26684
rect 463 26675 497 26709
rect 535 26675 569 26709
rect 607 26675 641 26709
rect 679 26675 713 26709
rect 751 26675 785 26709
rect 823 26682 843 26709
rect 843 26682 857 26709
rect 895 26682 915 26709
rect 915 26682 929 26709
rect 823 26675 857 26682
rect 895 26675 929 26682
rect -17 26650 17 26675
rect 75 26650 89 26675
rect 89 26650 109 26675
rect 167 26650 199 26675
rect 199 26650 201 26675
rect 259 26650 271 26675
rect 271 26650 293 26675
rect -17 26606 17 26611
rect 75 26606 109 26611
rect 167 26606 201 26611
rect 259 26606 293 26611
rect 463 26606 497 26635
rect 535 26606 569 26635
rect 607 26606 641 26635
rect 679 26606 713 26635
rect 751 26606 785 26635
rect 823 26613 843 26635
rect 843 26613 857 26635
rect 895 26613 915 26635
rect 915 26613 929 26635
rect -17 26577 17 26606
rect 75 26577 89 26606
rect 89 26577 109 26606
rect 167 26577 199 26606
rect 199 26577 201 26606
rect 259 26577 271 26606
rect 271 26577 293 26606
rect 463 26601 487 26606
rect 487 26601 497 26606
rect 535 26601 559 26606
rect 559 26601 569 26606
rect 607 26601 631 26606
rect 631 26601 641 26606
rect 679 26601 703 26606
rect 703 26601 713 26606
rect 751 26601 775 26606
rect 775 26601 785 26606
rect 823 26601 857 26613
rect 895 26601 929 26613
rect -17 26537 17 26538
rect 75 26537 109 26538
rect 167 26537 201 26538
rect 259 26537 293 26538
rect 463 26537 497 26561
rect 535 26537 569 26561
rect 607 26537 641 26561
rect 679 26537 713 26561
rect 751 26537 785 26561
rect 823 26544 843 26561
rect 843 26544 857 26561
rect 895 26544 915 26561
rect 915 26544 929 26561
rect -17 26504 17 26537
rect 75 26504 89 26537
rect 89 26504 109 26537
rect 167 26504 199 26537
rect 199 26504 201 26537
rect 259 26504 271 26537
rect 271 26504 293 26537
rect 463 26527 487 26537
rect 487 26527 497 26537
rect 535 26527 559 26537
rect 559 26527 569 26537
rect 607 26527 631 26537
rect 631 26527 641 26537
rect 679 26527 703 26537
rect 703 26527 713 26537
rect 751 26527 775 26537
rect 775 26527 785 26537
rect 823 26527 857 26544
rect 895 26527 929 26544
rect 463 26467 497 26487
rect 535 26467 569 26487
rect 607 26467 641 26487
rect 679 26467 713 26487
rect 751 26467 785 26487
rect 823 26475 843 26487
rect 843 26475 857 26487
rect 895 26475 915 26487
rect 915 26475 929 26487
rect -17 26433 17 26465
rect 75 26433 89 26465
rect 89 26433 109 26465
rect 167 26433 199 26465
rect 199 26433 201 26465
rect 259 26433 271 26465
rect 271 26433 293 26465
rect 463 26453 487 26467
rect 487 26453 497 26467
rect 535 26453 559 26467
rect 559 26453 569 26467
rect 607 26453 631 26467
rect 631 26453 641 26467
rect 679 26453 703 26467
rect 703 26453 713 26467
rect 751 26453 775 26467
rect 775 26453 785 26467
rect 823 26453 857 26475
rect 895 26453 929 26475
rect -17 26431 17 26433
rect 75 26431 109 26433
rect 167 26431 201 26433
rect 259 26431 293 26433
rect 463 26397 497 26413
rect 535 26397 569 26413
rect 607 26397 641 26413
rect 679 26397 713 26413
rect 751 26397 785 26413
rect 823 26406 843 26413
rect 843 26406 857 26413
rect 895 26406 915 26413
rect 915 26406 929 26413
rect -17 26363 17 26393
rect 75 26363 89 26393
rect 89 26363 109 26393
rect 167 26363 199 26393
rect 199 26363 201 26393
rect 259 26363 271 26393
rect 271 26363 293 26393
rect 463 26379 487 26397
rect 487 26379 497 26397
rect 535 26379 559 26397
rect 559 26379 569 26397
rect 607 26379 631 26397
rect 631 26379 641 26397
rect 679 26379 703 26397
rect 703 26379 713 26397
rect 751 26379 775 26397
rect 775 26379 785 26397
rect 823 26379 857 26406
rect 895 26379 929 26406
rect -17 26359 17 26363
rect 75 26359 109 26363
rect 167 26359 201 26363
rect 259 26359 293 26363
rect 463 26327 497 26339
rect 535 26327 569 26339
rect 607 26327 641 26339
rect 679 26327 713 26339
rect 751 26327 785 26339
rect 823 26337 843 26339
rect 843 26337 857 26339
rect 895 26337 915 26339
rect 915 26337 929 26339
rect -17 26293 17 26321
rect 75 26293 89 26321
rect 89 26293 109 26321
rect 167 26293 199 26321
rect 199 26293 201 26321
rect 259 26293 271 26321
rect 271 26293 293 26321
rect 463 26305 487 26327
rect 487 26305 497 26327
rect 535 26305 559 26327
rect 559 26305 569 26327
rect 607 26305 631 26327
rect 631 26305 641 26327
rect 679 26305 703 26327
rect 703 26305 713 26327
rect 751 26305 775 26327
rect 775 26305 785 26327
rect 823 26305 857 26337
rect 895 26305 929 26337
rect -17 26287 17 26293
rect 75 26287 109 26293
rect 167 26287 201 26293
rect 259 26287 293 26293
rect 463 26257 497 26265
rect 535 26257 569 26265
rect 607 26257 641 26265
rect 679 26257 713 26265
rect 751 26257 785 26265
rect 463 26231 487 26257
rect 487 26231 497 26257
rect 535 26231 559 26257
rect 559 26231 569 26257
rect 607 26231 631 26257
rect 631 26231 641 26257
rect 679 26231 703 26257
rect 703 26231 713 26257
rect 751 26231 775 26257
rect 775 26231 785 26257
rect 823 26233 857 26265
rect 895 26233 929 26265
rect 823 26231 843 26233
rect 843 26231 857 26233
rect 895 26231 915 26233
rect 915 26231 929 26233
rect -17 25987 17 26012
rect 75 25987 89 26012
rect 89 25987 109 26012
rect 167 25987 199 26012
rect 199 25987 201 26012
rect 259 25987 271 26012
rect 271 25987 293 26012
rect 459 25987 487 26012
rect 487 25987 493 26012
rect 537 25987 559 26012
rect 559 25987 571 26012
rect 615 25987 631 26012
rect 631 25987 649 26012
rect 693 25987 703 26012
rect 703 25987 727 26012
rect 771 25987 775 26012
rect 775 25987 805 26012
rect -17 25978 17 25987
rect 75 25978 109 25987
rect 167 25978 201 25987
rect 259 25978 293 25987
rect 459 25978 493 25987
rect 537 25978 571 25987
rect 615 25978 649 25987
rect 693 25978 727 25987
rect 771 25978 805 25987
rect 863 25972 897 25988
rect 863 25954 877 25972
rect 877 25954 897 25972
rect -17 25918 17 25940
rect 75 25918 89 25940
rect 89 25918 109 25940
rect 167 25918 199 25940
rect 199 25918 201 25940
rect 259 25918 271 25940
rect 271 25918 293 25940
rect 459 25918 487 25940
rect 487 25918 493 25940
rect 537 25918 559 25940
rect 559 25918 571 25940
rect 615 25918 631 25940
rect 631 25918 649 25940
rect 693 25918 703 25940
rect 703 25918 727 25940
rect 771 25918 775 25940
rect 775 25918 805 25940
rect -17 25906 17 25918
rect 75 25906 109 25918
rect 167 25906 201 25918
rect 259 25906 293 25918
rect 459 25906 493 25918
rect 537 25906 571 25918
rect 615 25906 649 25918
rect 693 25906 727 25918
rect 771 25906 805 25918
rect 863 25899 897 25915
rect -17 25849 17 25868
rect 75 25849 89 25868
rect 89 25849 109 25868
rect 167 25849 199 25868
rect 199 25849 201 25868
rect 259 25849 271 25868
rect 271 25849 293 25868
rect 459 25849 487 25868
rect 487 25849 493 25868
rect 537 25849 559 25868
rect 559 25849 571 25868
rect 615 25849 631 25868
rect 631 25849 649 25868
rect 693 25849 703 25868
rect 703 25849 727 25868
rect 771 25849 775 25868
rect 775 25849 805 25868
rect 863 25881 877 25899
rect 877 25881 897 25899
rect -17 25834 17 25849
rect 75 25834 109 25849
rect 167 25834 201 25849
rect 259 25834 293 25849
rect 459 25834 493 25849
rect 537 25834 571 25849
rect 615 25834 649 25849
rect 693 25834 727 25849
rect 771 25834 805 25849
rect 863 25826 897 25842
rect -17 25780 17 25796
rect 75 25780 89 25796
rect 89 25780 109 25796
rect 167 25780 199 25796
rect 199 25780 201 25796
rect 259 25780 271 25796
rect 271 25780 293 25796
rect 459 25780 487 25796
rect 487 25780 493 25796
rect 537 25780 559 25796
rect 559 25780 571 25796
rect 615 25780 631 25796
rect 631 25780 649 25796
rect 693 25780 703 25796
rect 703 25780 727 25796
rect 771 25780 775 25796
rect 775 25780 805 25796
rect 863 25808 877 25826
rect 877 25808 897 25826
rect -17 25762 17 25780
rect 75 25762 109 25780
rect 167 25762 201 25780
rect 259 25762 293 25780
rect 459 25762 493 25780
rect 537 25762 571 25780
rect 615 25762 649 25780
rect 693 25762 727 25780
rect 771 25762 805 25780
rect 863 25753 897 25769
rect -17 25711 17 25724
rect 75 25711 89 25724
rect 89 25711 109 25724
rect 167 25711 199 25724
rect 199 25711 201 25724
rect 259 25711 271 25724
rect 271 25711 293 25724
rect 459 25711 487 25724
rect 487 25711 493 25724
rect 537 25711 559 25724
rect 559 25711 571 25724
rect 615 25711 631 25724
rect 631 25711 649 25724
rect 693 25711 703 25724
rect 703 25711 727 25724
rect 771 25711 775 25724
rect 775 25711 805 25724
rect 863 25735 877 25753
rect 877 25735 897 25753
rect -17 25690 17 25711
rect 75 25690 109 25711
rect 167 25690 201 25711
rect 259 25690 293 25711
rect 459 25690 493 25711
rect 537 25690 571 25711
rect 615 25690 649 25711
rect 693 25690 727 25711
rect 771 25690 805 25711
rect 863 25680 897 25696
rect 13833 25987 13867 26021
rect 13906 25987 13940 26021
rect 13979 25987 14013 26021
rect 14052 25987 14086 26021
rect 14125 25987 14159 26021
rect 14198 25987 14232 26021
rect 14271 25987 14305 26021
rect 14344 25987 14378 26021
rect 14417 25987 14451 26021
rect 14490 25987 14524 26021
rect 14563 25987 14597 26021
rect 14636 25987 14670 26021
rect 14709 25987 14743 26021
rect 14782 25987 14816 26021
rect 14855 25987 14889 26021
rect 14928 25987 14962 26021
rect 15001 25987 15035 26021
rect 15074 25987 15108 26021
rect 15147 25987 15181 26021
rect 15220 25987 15254 26021
rect 15293 25987 15327 26021
rect 15366 25987 15400 26021
rect 15439 25987 15473 26021
rect 15513 25987 15547 26021
rect 15587 25987 15621 26021
rect 15661 25987 15695 26021
rect 15735 25987 15769 26021
rect 15809 25987 15843 26021
rect 15883 25987 15917 26021
rect 13833 25913 13867 25947
rect 13906 25913 13940 25947
rect 13979 25913 14013 25947
rect 14052 25913 14086 25947
rect 14125 25913 14159 25947
rect 14198 25913 14232 25947
rect 14271 25913 14305 25947
rect 14344 25913 14378 25947
rect 14417 25913 14451 25947
rect 14490 25913 14524 25947
rect 14563 25913 14597 25947
rect 14636 25913 14670 25947
rect 14709 25913 14743 25947
rect 14782 25913 14816 25947
rect 14855 25913 14889 25947
rect 14928 25913 14962 25947
rect 15001 25913 15035 25947
rect 15074 25913 15108 25947
rect 15147 25913 15181 25947
rect 15220 25913 15254 25947
rect 15293 25913 15327 25947
rect 15366 25913 15400 25947
rect 15439 25913 15473 25947
rect 15513 25913 15547 25947
rect 15587 25913 15621 25947
rect 15661 25913 15695 25947
rect 15735 25913 15769 25947
rect 15809 25913 15843 25947
rect 15883 25913 15917 25947
rect 13833 25839 13867 25873
rect 13906 25839 13940 25873
rect 13979 25839 14013 25873
rect 14052 25839 14086 25873
rect 14125 25839 14159 25873
rect 14198 25839 14232 25873
rect 14271 25839 14305 25873
rect 14344 25839 14378 25873
rect 14417 25839 14451 25873
rect 14490 25839 14524 25873
rect 14563 25839 14597 25873
rect 14636 25839 14670 25873
rect 14709 25839 14743 25873
rect 14782 25839 14816 25873
rect 14855 25839 14889 25873
rect 14928 25839 14962 25873
rect 15001 25839 15035 25873
rect 15074 25839 15108 25873
rect 15147 25839 15181 25873
rect 15220 25839 15254 25873
rect 15293 25839 15327 25873
rect 15366 25839 15400 25873
rect 15439 25839 15473 25873
rect 15513 25839 15547 25873
rect 15587 25839 15621 25873
rect 15661 25839 15695 25873
rect 15735 25839 15769 25873
rect 15809 25839 15843 25873
rect 15883 25839 15917 25873
rect 13833 25765 13867 25799
rect 13906 25765 13940 25799
rect 13979 25765 14013 25799
rect 14052 25765 14086 25799
rect 14125 25765 14159 25799
rect 14198 25765 14232 25799
rect 14271 25765 14305 25799
rect 14344 25765 14378 25799
rect 14417 25765 14451 25799
rect 14490 25765 14524 25799
rect 14563 25765 14597 25799
rect 14636 25765 14670 25799
rect 14709 25765 14743 25799
rect 14782 25765 14816 25799
rect 14855 25765 14889 25799
rect 14928 25765 14962 25799
rect 15001 25765 15035 25799
rect 15074 25765 15108 25799
rect 15147 25765 15181 25799
rect 15220 25765 15254 25799
rect 15293 25765 15327 25799
rect 15366 25765 15400 25799
rect 15439 25765 15473 25799
rect 15513 25765 15547 25799
rect 15587 25765 15621 25799
rect 15661 25765 15695 25799
rect 15735 25765 15769 25799
rect 15809 25765 15843 25799
rect 15883 25765 15917 25799
rect 13833 25691 13867 25725
rect 13906 25691 13940 25725
rect 13979 25691 14013 25725
rect 14052 25691 14086 25725
rect 14125 25691 14159 25725
rect 14198 25691 14232 25725
rect 14271 25691 14305 25725
rect 14344 25691 14378 25725
rect 14417 25691 14451 25725
rect 14490 25691 14524 25725
rect 14563 25691 14597 25725
rect 14636 25691 14670 25725
rect 14709 25691 14743 25725
rect 14782 25691 14816 25725
rect 14855 25691 14889 25725
rect 14928 25691 14962 25725
rect 15001 25691 15035 25725
rect 15074 25691 15108 25725
rect 15147 25691 15181 25725
rect 15220 25691 15254 25725
rect 15293 25691 15327 25725
rect 15366 25691 15400 25725
rect 15439 25691 15473 25725
rect 15513 25691 15547 25725
rect 15587 25691 15621 25725
rect 15661 25691 15695 25725
rect 15735 25691 15769 25725
rect 15809 25691 15843 25725
rect 15883 25691 15917 25725
rect -17 25642 17 25652
rect 75 25642 89 25652
rect 89 25642 109 25652
rect 167 25642 199 25652
rect 199 25642 201 25652
rect 259 25642 271 25652
rect 271 25642 293 25652
rect 459 25642 487 25652
rect 487 25642 493 25652
rect 537 25642 559 25652
rect 559 25642 571 25652
rect 615 25642 631 25652
rect 631 25642 649 25652
rect 693 25642 703 25652
rect 703 25642 727 25652
rect 771 25642 775 25652
rect 775 25642 805 25652
rect 863 25662 877 25680
rect 877 25662 897 25680
rect -17 25618 17 25642
rect 75 25618 109 25642
rect 167 25618 201 25642
rect 259 25618 293 25642
rect 459 25618 493 25642
rect 537 25618 571 25642
rect 615 25618 649 25642
rect 693 25618 727 25642
rect 771 25618 805 25642
rect 863 25607 897 25623
rect -17 25573 17 25580
rect 75 25573 89 25580
rect 89 25573 109 25580
rect 167 25573 199 25580
rect 199 25573 201 25580
rect 259 25573 271 25580
rect 271 25573 293 25580
rect 459 25573 487 25580
rect 487 25573 493 25580
rect 537 25573 559 25580
rect 559 25573 571 25580
rect 615 25573 631 25580
rect 631 25573 649 25580
rect 693 25573 703 25580
rect 703 25573 727 25580
rect 771 25573 775 25580
rect 775 25573 805 25580
rect 863 25589 877 25607
rect 877 25589 897 25607
rect -17 25546 17 25573
rect 75 25546 109 25573
rect 167 25546 201 25573
rect 259 25546 293 25573
rect 459 25546 493 25573
rect 537 25546 571 25573
rect 615 25546 649 25573
rect 693 25546 727 25573
rect 771 25546 805 25573
rect -17 25505 17 25508
rect 75 25505 89 25508
rect 89 25505 109 25508
rect 167 25505 199 25508
rect 199 25505 201 25508
rect 259 25505 271 25508
rect 271 25505 293 25508
rect 863 25534 897 25550
rect 459 25505 487 25508
rect 487 25505 493 25508
rect 537 25505 559 25508
rect 559 25505 571 25508
rect 615 25505 631 25508
rect 631 25505 649 25508
rect 693 25505 703 25508
rect 703 25505 727 25508
rect 771 25505 775 25508
rect 775 25505 805 25508
rect 863 25516 877 25534
rect 877 25516 897 25534
rect -17 25474 17 25505
rect 75 25474 109 25505
rect 167 25474 201 25505
rect 259 25474 293 25505
rect 459 25474 493 25505
rect 537 25474 571 25505
rect 615 25474 649 25505
rect 693 25474 727 25505
rect 771 25474 805 25505
rect 863 25461 897 25476
rect 863 25442 877 25461
rect 877 25442 897 25461
rect -17 25403 17 25436
rect 75 25403 109 25436
rect 167 25403 201 25436
rect 259 25403 293 25436
rect 459 25403 493 25436
rect 537 25403 571 25436
rect 615 25403 649 25436
rect 693 25403 727 25436
rect 771 25403 805 25436
rect -17 25402 17 25403
rect 75 25402 89 25403
rect 89 25402 109 25403
rect 167 25402 199 25403
rect 199 25402 201 25403
rect 259 25402 271 25403
rect 271 25402 293 25403
rect 459 25402 487 25403
rect 487 25402 493 25403
rect 537 25402 559 25403
rect 559 25402 571 25403
rect 615 25402 631 25403
rect 631 25402 649 25403
rect 693 25402 703 25403
rect 703 25402 727 25403
rect 771 25402 775 25403
rect 775 25402 805 25403
rect 863 25388 897 25402
rect 863 25368 877 25388
rect 877 25368 897 25388
rect -17 25335 17 25364
rect 75 25335 109 25364
rect 167 25335 201 25364
rect 259 25335 293 25364
rect 459 25335 493 25364
rect 537 25335 571 25364
rect 615 25335 649 25364
rect 693 25335 727 25364
rect 771 25335 805 25364
rect -17 25330 17 25335
rect 75 25330 89 25335
rect 89 25330 109 25335
rect 167 25330 199 25335
rect 199 25330 201 25335
rect 259 25330 271 25335
rect 271 25330 293 25335
rect 459 25330 487 25335
rect 487 25330 493 25335
rect 537 25330 559 25335
rect 559 25330 571 25335
rect 615 25330 631 25335
rect 631 25330 649 25335
rect 693 25330 703 25335
rect 703 25330 727 25335
rect 771 25330 775 25335
rect 775 25330 805 25335
rect 863 25316 897 25328
rect 863 25294 877 25316
rect 877 25294 897 25316
rect -17 25267 17 25292
rect 75 25267 109 25292
rect 167 25267 201 25292
rect 259 25267 293 25292
rect 459 25267 493 25292
rect 537 25267 571 25292
rect 615 25267 649 25292
rect 693 25267 727 25292
rect 771 25267 805 25292
rect -17 25258 17 25267
rect 75 25258 89 25267
rect 89 25258 109 25267
rect 167 25258 199 25267
rect 199 25258 201 25267
rect 259 25258 271 25267
rect 271 25258 293 25267
rect 459 25258 487 25267
rect 487 25258 493 25267
rect 537 25258 559 25267
rect 559 25258 571 25267
rect 615 25258 631 25267
rect 631 25258 649 25267
rect 693 25258 703 25267
rect 703 25258 727 25267
rect 771 25258 775 25267
rect 775 25258 805 25267
rect -17 25199 17 25220
rect 75 25199 109 25220
rect 167 25199 201 25220
rect 259 25199 293 25220
rect 459 25199 493 25220
rect 537 25199 571 25220
rect 615 25199 649 25220
rect 693 25199 727 25220
rect 771 25199 805 25220
rect -17 25186 17 25199
rect 75 25186 89 25199
rect 89 25186 109 25199
rect 167 25186 199 25199
rect 199 25186 201 25199
rect 259 25186 271 25199
rect 271 25186 293 25199
rect 459 25186 487 25199
rect 487 25186 493 25199
rect 537 25186 559 25199
rect 559 25186 571 25199
rect 615 25186 631 25199
rect 631 25186 649 25199
rect 693 25186 703 25199
rect 703 25186 727 25199
rect 771 25186 775 25199
rect 775 25186 805 25199
rect -17 25131 17 25148
rect 75 25131 109 25148
rect 167 25131 201 25148
rect 259 25131 293 25148
rect 459 25131 493 25148
rect 537 25131 571 25148
rect 615 25131 649 25148
rect 693 25131 727 25148
rect 771 25131 805 25148
rect -17 25114 17 25131
rect 75 25114 89 25131
rect 89 25114 109 25131
rect 167 25114 199 25131
rect 199 25114 201 25131
rect 259 25114 271 25131
rect 271 25114 293 25131
rect 459 25114 487 25131
rect 487 25114 493 25131
rect 537 25114 559 25131
rect 559 25114 571 25131
rect 615 25114 631 25131
rect 631 25114 649 25131
rect 693 25114 703 25131
rect 703 25114 727 25131
rect 771 25114 775 25131
rect 775 25114 805 25131
rect -17 25063 17 25076
rect 75 25063 109 25076
rect 167 25063 201 25076
rect 259 25063 293 25076
rect 459 25063 493 25076
rect 537 25063 571 25076
rect 615 25063 649 25076
rect 693 25063 727 25076
rect 771 25063 805 25076
rect -17 25042 17 25063
rect 75 25042 89 25063
rect 89 25042 109 25063
rect 167 25042 199 25063
rect 199 25042 201 25063
rect 259 25042 271 25063
rect 271 25042 293 25063
rect 459 25042 487 25063
rect 487 25042 493 25063
rect 537 25042 559 25063
rect 559 25042 571 25063
rect 615 25042 631 25063
rect 631 25042 649 25063
rect 693 25042 703 25063
rect 703 25042 727 25063
rect 771 25042 775 25063
rect 775 25042 805 25063
rect -17 24995 17 25004
rect 75 24995 109 25004
rect 167 24995 201 25004
rect 259 24995 293 25004
rect 459 24995 493 25004
rect 537 24995 571 25004
rect 615 24995 649 25004
rect 693 24995 727 25004
rect 771 24995 805 25004
rect -17 24970 17 24995
rect 75 24970 89 24995
rect 89 24970 109 24995
rect 167 24970 199 24995
rect 199 24970 201 24995
rect 259 24970 271 24995
rect 271 24970 293 24995
rect 459 24970 487 24995
rect 487 24970 493 24995
rect 537 24970 559 24995
rect 559 24970 571 24995
rect 615 24970 631 24995
rect 631 24970 649 24995
rect 693 24970 703 24995
rect 703 24970 727 24995
rect 771 24970 775 24995
rect 775 24970 805 24995
rect -17 24927 17 24932
rect 75 24927 109 24932
rect 167 24927 201 24932
rect 259 24927 293 24932
rect 459 24927 493 24932
rect 537 24927 571 24932
rect 615 24927 649 24932
rect 693 24927 727 24932
rect 771 24927 805 24932
rect -17 24898 17 24927
rect 75 24898 89 24927
rect 89 24898 109 24927
rect 167 24898 199 24927
rect 199 24898 201 24927
rect 259 24898 271 24927
rect 271 24898 293 24927
rect 459 24898 487 24927
rect 487 24898 493 24927
rect 537 24898 559 24927
rect 559 24898 571 24927
rect 615 24898 631 24927
rect 631 24898 649 24927
rect 693 24898 703 24927
rect 703 24898 727 24927
rect 771 24898 775 24927
rect 775 24898 805 24927
rect -17 24859 17 24860
rect 75 24859 109 24860
rect 167 24859 201 24860
rect 259 24859 293 24860
rect 459 24859 493 24860
rect 537 24859 571 24860
rect 615 24859 649 24860
rect 693 24859 727 24860
rect 771 24859 805 24860
rect -17 24826 17 24859
rect 75 24826 89 24859
rect 89 24826 109 24859
rect 167 24826 199 24859
rect 199 24826 201 24859
rect 259 24826 271 24859
rect 271 24826 293 24859
rect 459 24826 487 24859
rect 487 24826 493 24859
rect 537 24826 559 24859
rect 559 24826 571 24859
rect 615 24826 631 24859
rect 631 24826 649 24859
rect 693 24826 703 24859
rect 703 24826 727 24859
rect 771 24826 775 24859
rect 775 24826 805 24859
rect -17 24757 17 24788
rect 75 24757 89 24788
rect 89 24757 109 24788
rect 167 24757 199 24788
rect 199 24757 201 24788
rect 259 24757 271 24788
rect 271 24757 293 24788
rect 459 24757 487 24788
rect 487 24757 493 24788
rect 537 24757 559 24788
rect 559 24757 571 24788
rect 615 24757 631 24788
rect 631 24757 649 24788
rect 693 24757 703 24788
rect 703 24757 727 24788
rect 771 24757 775 24788
rect 775 24757 805 24788
rect -17 24754 17 24757
rect 75 24754 109 24757
rect 167 24754 201 24757
rect 259 24754 293 24757
rect 459 24754 493 24757
rect 537 24754 571 24757
rect 615 24754 649 24757
rect 693 24754 727 24757
rect 771 24754 805 24757
rect -17 24689 17 24716
rect 75 24689 89 24716
rect 89 24689 109 24716
rect 167 24689 199 24716
rect 199 24689 201 24716
rect 259 24689 271 24716
rect 271 24689 293 24716
rect 459 24689 487 24716
rect 487 24689 493 24716
rect 537 24689 559 24716
rect 559 24689 571 24716
rect 615 24689 631 24716
rect 631 24689 649 24716
rect 693 24689 703 24716
rect 703 24689 727 24716
rect 771 24689 775 24716
rect 775 24689 805 24716
rect -17 24682 17 24689
rect 75 24682 109 24689
rect 167 24682 201 24689
rect 259 24682 293 24689
rect 459 24682 493 24689
rect 537 24682 571 24689
rect 615 24682 649 24689
rect 693 24682 727 24689
rect 771 24682 805 24689
rect -17 24621 17 24644
rect 75 24621 89 24644
rect 89 24621 109 24644
rect 167 24621 199 24644
rect 199 24621 201 24644
rect 259 24621 271 24644
rect 271 24621 293 24644
rect 459 24621 487 24644
rect 487 24621 493 24644
rect 537 24621 559 24644
rect 559 24621 571 24644
rect 615 24621 631 24644
rect 631 24621 649 24644
rect 693 24621 703 24644
rect 703 24621 727 24644
rect 771 24621 775 24644
rect 775 24621 805 24644
rect -17 24610 17 24621
rect 75 24610 109 24621
rect 167 24610 201 24621
rect 259 24610 293 24621
rect 459 24610 493 24621
rect 537 24610 571 24621
rect 615 24610 649 24621
rect 693 24610 727 24621
rect 771 24610 805 24621
rect -17 24553 17 24572
rect 75 24553 89 24572
rect 89 24553 109 24572
rect 167 24553 199 24572
rect 199 24553 201 24572
rect 259 24553 271 24572
rect 271 24553 293 24572
rect 459 24553 487 24572
rect 487 24553 493 24572
rect 537 24553 559 24572
rect 559 24553 571 24572
rect 615 24553 631 24572
rect 631 24553 649 24572
rect 693 24553 703 24572
rect 703 24553 727 24572
rect 771 24553 775 24572
rect 775 24553 805 24572
rect -17 24538 17 24553
rect 75 24538 109 24553
rect 167 24538 201 24553
rect 259 24538 293 24553
rect 459 24538 493 24553
rect 537 24538 571 24553
rect 615 24538 649 24553
rect 693 24538 727 24553
rect 771 24538 805 24553
rect -17 24485 17 24500
rect 75 24485 89 24500
rect 89 24485 109 24500
rect 167 24485 199 24500
rect 199 24485 201 24500
rect 259 24485 271 24500
rect 271 24485 293 24500
rect 459 24485 487 24500
rect 487 24485 493 24500
rect 537 24485 559 24500
rect 559 24485 571 24500
rect 615 24485 631 24500
rect 631 24485 649 24500
rect 693 24485 703 24500
rect 703 24485 727 24500
rect 771 24485 775 24500
rect 775 24485 805 24500
rect -17 24466 17 24485
rect 75 24466 109 24485
rect 167 24466 201 24485
rect 259 24466 293 24485
rect 459 24466 493 24485
rect 537 24466 571 24485
rect 615 24466 649 24485
rect 693 24466 727 24485
rect 771 24466 805 24485
rect -17 24417 17 24428
rect 75 24417 89 24428
rect 89 24417 109 24428
rect 167 24417 199 24428
rect 199 24417 201 24428
rect 259 24417 271 24428
rect 271 24417 293 24428
rect 459 24417 487 24428
rect 487 24417 493 24428
rect 537 24417 559 24428
rect 559 24417 571 24428
rect 615 24417 631 24428
rect 631 24417 649 24428
rect 693 24417 703 24428
rect 703 24417 727 24428
rect 771 24417 775 24428
rect 775 24417 805 24428
rect -17 24394 17 24417
rect 75 24394 109 24417
rect 167 24394 201 24417
rect 259 24394 293 24417
rect 459 24394 493 24417
rect 537 24394 571 24417
rect 615 24394 649 24417
rect 693 24394 727 24417
rect 771 24394 805 24417
rect -17 24349 17 24355
rect 75 24349 89 24355
rect 89 24349 109 24355
rect 167 24349 199 24355
rect 199 24349 201 24355
rect 259 24349 271 24355
rect 271 24349 293 24355
rect 459 24349 487 24355
rect 487 24349 493 24355
rect 537 24349 559 24355
rect 559 24349 571 24355
rect 615 24349 631 24355
rect 631 24349 649 24355
rect 693 24349 703 24355
rect 703 24349 727 24355
rect 771 24349 775 24355
rect 775 24349 805 24355
rect -17 24321 17 24349
rect 75 24321 109 24349
rect 167 24321 201 24349
rect 259 24321 293 24349
rect 459 24321 493 24349
rect 537 24321 571 24349
rect 615 24321 649 24349
rect 693 24321 727 24349
rect 771 24321 805 24349
rect -17 24281 17 24282
rect 75 24281 89 24282
rect 89 24281 109 24282
rect 167 24281 199 24282
rect 199 24281 201 24282
rect 259 24281 271 24282
rect 271 24281 293 24282
rect 459 24281 487 24282
rect 487 24281 493 24282
rect 537 24281 559 24282
rect 559 24281 571 24282
rect 615 24281 631 24282
rect 631 24281 649 24282
rect 693 24281 703 24282
rect 703 24281 727 24282
rect 771 24281 775 24282
rect 775 24281 805 24282
rect -17 24248 17 24281
rect 75 24248 109 24281
rect 167 24248 201 24281
rect 259 24248 293 24281
rect 459 24248 493 24281
rect 537 24248 571 24281
rect 615 24248 649 24281
rect 693 24248 727 24281
rect 771 24248 805 24281
rect -17 24179 17 24209
rect 75 24179 109 24209
rect 167 24179 201 24209
rect 259 24179 293 24209
rect 459 24179 493 24209
rect 537 24179 571 24209
rect 615 24179 649 24209
rect 693 24179 727 24209
rect 771 24179 805 24209
rect -17 24175 17 24179
rect 75 24175 89 24179
rect 89 24175 109 24179
rect 167 24175 199 24179
rect 199 24175 201 24179
rect 259 24175 271 24179
rect 271 24175 293 24179
rect 459 24175 487 24179
rect 487 24175 493 24179
rect 537 24175 559 24179
rect 559 24175 571 24179
rect 615 24175 631 24179
rect 631 24175 649 24179
rect 693 24175 703 24179
rect 703 24175 727 24179
rect 771 24175 775 24179
rect 775 24175 805 24179
rect -17 24111 17 24136
rect 75 24111 109 24136
rect 167 24111 201 24136
rect 259 24111 293 24136
rect 459 24111 493 24136
rect 537 24111 571 24136
rect 615 24111 649 24136
rect 693 24111 727 24136
rect 771 24111 805 24136
rect -17 24102 17 24111
rect 75 24102 89 24111
rect 89 24102 109 24111
rect 167 24102 199 24111
rect 199 24102 201 24111
rect 259 24102 271 24111
rect 271 24102 293 24111
rect 459 24102 487 24111
rect 487 24102 493 24111
rect 537 24102 559 24111
rect 559 24102 571 24111
rect 615 24102 631 24111
rect 631 24102 649 24111
rect 693 24102 703 24111
rect 703 24102 727 24111
rect 771 24102 775 24111
rect 775 24102 805 24111
rect -17 24043 17 24063
rect 75 24043 109 24063
rect 167 24043 201 24063
rect 259 24043 293 24063
rect 459 24043 493 24063
rect 537 24043 571 24063
rect 615 24043 649 24063
rect 693 24043 727 24063
rect 771 24043 805 24063
rect -17 24029 17 24043
rect 75 24029 89 24043
rect 89 24029 109 24043
rect 167 24029 199 24043
rect 199 24029 201 24043
rect 259 24029 271 24043
rect 271 24029 293 24043
rect 459 24029 487 24043
rect 487 24029 493 24043
rect 537 24029 559 24043
rect 559 24029 571 24043
rect 615 24029 631 24043
rect 631 24029 649 24043
rect 693 24029 703 24043
rect 703 24029 727 24043
rect 771 24029 775 24043
rect 775 24029 805 24043
rect -17 23975 17 23990
rect 75 23975 109 23990
rect 167 23975 201 23990
rect 259 23975 293 23990
rect 459 23975 493 23990
rect 537 23975 571 23990
rect 615 23975 649 23990
rect 693 23975 727 23990
rect 771 23975 805 23990
rect -17 23956 17 23975
rect 75 23956 89 23975
rect 89 23956 109 23975
rect 167 23956 199 23975
rect 199 23956 201 23975
rect 259 23956 271 23975
rect 271 23956 293 23975
rect 459 23956 487 23975
rect 487 23956 493 23975
rect 537 23956 559 23975
rect 559 23956 571 23975
rect 615 23956 631 23975
rect 631 23956 649 23975
rect 693 23956 703 23975
rect 703 23956 727 23975
rect 771 23956 775 23975
rect 775 23956 805 23975
rect -17 23907 17 23917
rect 75 23907 109 23917
rect 167 23907 201 23917
rect 259 23907 293 23917
rect 459 23907 493 23917
rect 537 23907 571 23917
rect 615 23907 649 23917
rect 693 23907 727 23917
rect 771 23907 805 23917
rect -17 23883 17 23907
rect 75 23883 89 23907
rect 89 23883 109 23907
rect 167 23883 199 23907
rect 199 23883 201 23907
rect 259 23883 271 23907
rect 271 23883 293 23907
rect 459 23883 487 23907
rect 487 23883 493 23907
rect 537 23883 559 23907
rect 559 23883 571 23907
rect 615 23883 631 23907
rect 631 23883 649 23907
rect 693 23883 703 23907
rect 703 23883 727 23907
rect 771 23883 775 23907
rect 775 23883 805 23907
rect -17 23839 17 23844
rect 75 23839 109 23844
rect 167 23839 201 23844
rect 259 23839 293 23844
rect 459 23839 493 23844
rect 537 23839 571 23844
rect 615 23839 649 23844
rect 693 23839 727 23844
rect 771 23839 805 23844
rect -17 23810 17 23839
rect 75 23810 89 23839
rect 89 23810 109 23839
rect 167 23810 199 23839
rect 199 23810 201 23839
rect 259 23810 271 23839
rect 271 23810 293 23839
rect 459 23810 487 23839
rect 487 23810 493 23839
rect 537 23810 559 23839
rect 559 23810 571 23839
rect 615 23810 631 23839
rect 631 23810 649 23839
rect 693 23810 703 23839
rect 703 23810 727 23839
rect 771 23810 775 23839
rect 775 23810 805 23839
rect -17 23737 17 23771
rect 75 23737 89 23771
rect 89 23737 109 23771
rect 167 23737 199 23771
rect 199 23737 201 23771
rect 259 23737 271 23771
rect 271 23737 293 23771
rect 459 23737 487 23771
rect 487 23737 493 23771
rect 537 23737 559 23771
rect 559 23737 571 23771
rect 615 23737 631 23771
rect 631 23737 649 23771
rect 693 23737 703 23771
rect 703 23737 727 23771
rect 771 23737 775 23771
rect 775 23737 805 23771
rect -17 23669 17 23698
rect 75 23669 89 23698
rect 89 23669 109 23698
rect 167 23669 199 23698
rect 199 23669 201 23698
rect 259 23669 271 23698
rect 271 23669 293 23698
rect 459 23669 487 23698
rect 487 23669 493 23698
rect 537 23669 559 23698
rect 559 23669 571 23698
rect 615 23669 631 23698
rect 631 23669 649 23698
rect 693 23669 703 23698
rect 703 23669 727 23698
rect 771 23669 775 23698
rect 775 23669 805 23698
rect -17 23664 17 23669
rect 75 23664 109 23669
rect 167 23664 201 23669
rect 259 23664 293 23669
rect 459 23664 493 23669
rect 537 23664 571 23669
rect 615 23664 649 23669
rect 693 23664 727 23669
rect 771 23664 805 23669
rect -17 23601 17 23625
rect 75 23601 89 23625
rect 89 23601 109 23625
rect 167 23601 199 23625
rect 199 23601 201 23625
rect 259 23601 271 23625
rect 271 23601 293 23625
rect 459 23601 487 23625
rect 487 23601 493 23625
rect 537 23601 559 23625
rect 559 23601 571 23625
rect 615 23601 631 23625
rect 631 23601 649 23625
rect 693 23601 703 23625
rect 703 23601 727 23625
rect 771 23601 775 23625
rect 775 23601 805 23625
rect -17 23591 17 23601
rect 75 23591 109 23601
rect 167 23591 201 23601
rect 259 23591 293 23601
rect 459 23591 493 23601
rect 537 23591 571 23601
rect 615 23591 649 23601
rect 693 23591 727 23601
rect 771 23591 805 23601
rect -17 23533 17 23552
rect 75 23533 89 23552
rect 89 23533 109 23552
rect 167 23533 199 23552
rect 199 23533 201 23552
rect 259 23533 271 23552
rect 271 23533 293 23552
rect 459 23533 487 23552
rect 487 23533 493 23552
rect 537 23533 559 23552
rect 559 23533 571 23552
rect 615 23533 631 23552
rect 631 23533 649 23552
rect 693 23533 703 23552
rect 703 23533 727 23552
rect 771 23533 775 23552
rect 775 23533 805 23552
rect -17 23518 17 23533
rect 75 23518 109 23533
rect 167 23518 201 23533
rect 259 23518 293 23533
rect 459 23518 493 23533
rect 537 23518 571 23533
rect 615 23518 649 23533
rect 693 23518 727 23533
rect 771 23518 805 23533
rect -17 23465 17 23479
rect 75 23465 89 23479
rect 89 23465 109 23479
rect 167 23465 199 23479
rect 199 23465 201 23479
rect 259 23465 271 23479
rect 271 23465 293 23479
rect 459 23465 487 23479
rect 487 23465 493 23479
rect 537 23465 559 23479
rect 559 23465 571 23479
rect 615 23465 631 23479
rect 631 23465 649 23479
rect 693 23465 703 23479
rect 703 23465 727 23479
rect 771 23465 775 23479
rect 775 23465 805 23479
rect -17 23445 17 23465
rect 75 23445 109 23465
rect 167 23445 201 23465
rect 259 23445 293 23465
rect 459 23445 493 23465
rect 537 23445 571 23465
rect 615 23445 649 23465
rect 693 23445 727 23465
rect 771 23445 805 23465
rect -17 23397 17 23406
rect 75 23397 89 23406
rect 89 23397 109 23406
rect 167 23397 199 23406
rect 199 23397 201 23406
rect 259 23397 271 23406
rect 271 23397 293 23406
rect 459 23397 487 23406
rect 487 23397 493 23406
rect 537 23397 559 23406
rect 559 23397 571 23406
rect 615 23397 631 23406
rect 631 23397 649 23406
rect 693 23397 703 23406
rect 703 23397 727 23406
rect 771 23397 775 23406
rect 775 23397 805 23406
rect -17 23372 17 23397
rect 75 23372 109 23397
rect 167 23372 201 23397
rect 259 23372 293 23397
rect 459 23372 493 23397
rect 537 23372 571 23397
rect 615 23372 649 23397
rect 693 23372 727 23397
rect 771 23372 805 23397
rect -17 23329 17 23333
rect 75 23329 89 23333
rect 89 23329 109 23333
rect 167 23329 199 23333
rect 199 23329 201 23333
rect 259 23329 271 23333
rect 271 23329 293 23333
rect 459 23329 487 23333
rect 487 23329 493 23333
rect 537 23329 559 23333
rect 559 23329 571 23333
rect 615 23329 631 23333
rect 631 23329 649 23333
rect 693 23329 703 23333
rect 703 23329 727 23333
rect 771 23329 775 23333
rect 775 23329 805 23333
rect -17 23299 17 23329
rect 75 23299 109 23329
rect 167 23299 201 23329
rect 259 23299 293 23329
rect 459 23299 493 23329
rect 537 23299 571 23329
rect 615 23299 649 23329
rect 693 23299 727 23329
rect 771 23299 805 23329
rect -17 23227 17 23260
rect 75 23227 109 23260
rect 167 23227 201 23260
rect 259 23227 293 23260
rect 459 23227 493 23260
rect 537 23227 571 23260
rect 615 23227 649 23260
rect 693 23227 727 23260
rect 771 23227 805 23260
rect -17 23226 17 23227
rect 75 23226 89 23227
rect 89 23226 109 23227
rect 167 23226 199 23227
rect 199 23226 201 23227
rect 259 23226 271 23227
rect 271 23226 293 23227
rect 459 23226 487 23227
rect 487 23226 493 23227
rect 537 23226 559 23227
rect 559 23226 571 23227
rect 615 23226 631 23227
rect 631 23226 649 23227
rect 693 23226 703 23227
rect 703 23226 727 23227
rect 771 23226 775 23227
rect 775 23226 805 23227
rect -17 23159 17 23187
rect 75 23159 109 23187
rect 167 23159 201 23187
rect 259 23159 293 23187
rect 459 23159 493 23187
rect 537 23159 571 23187
rect 615 23159 649 23187
rect 693 23159 727 23187
rect 771 23159 805 23187
rect -17 23153 17 23159
rect 75 23153 89 23159
rect 89 23153 109 23159
rect 167 23153 199 23159
rect 199 23153 201 23159
rect 259 23153 271 23159
rect 271 23153 293 23159
rect 459 23153 487 23159
rect 487 23153 493 23159
rect 537 23153 559 23159
rect 559 23153 571 23159
rect 615 23153 631 23159
rect 631 23153 649 23159
rect 693 23153 703 23159
rect 703 23153 727 23159
rect 771 23153 775 23159
rect 775 23153 805 23159
rect -17 23091 17 23114
rect 75 23091 109 23114
rect 167 23091 201 23114
rect 259 23091 293 23114
rect 459 23091 493 23114
rect 537 23091 571 23114
rect 615 23091 649 23114
rect 693 23091 727 23114
rect 771 23091 805 23114
rect -17 23080 17 23091
rect 75 23080 89 23091
rect 89 23080 109 23091
rect 167 23080 199 23091
rect 199 23080 201 23091
rect 259 23080 271 23091
rect 271 23080 293 23091
rect 459 23080 487 23091
rect 487 23080 493 23091
rect 537 23080 559 23091
rect 559 23080 571 23091
rect 615 23080 631 23091
rect 631 23080 649 23091
rect 693 23080 703 23091
rect 703 23080 727 23091
rect 771 23080 775 23091
rect 775 23080 805 23091
rect -17 23023 17 23041
rect 75 23023 109 23041
rect 167 23023 201 23041
rect 259 23023 293 23041
rect 459 23023 493 23041
rect 537 23023 571 23041
rect 615 23023 649 23041
rect 693 23023 727 23041
rect 771 23023 805 23041
rect -17 23007 17 23023
rect 75 23007 89 23023
rect 89 23007 109 23023
rect 167 23007 199 23023
rect 199 23007 201 23023
rect 259 23007 271 23023
rect 271 23007 293 23023
rect 459 23007 487 23023
rect 487 23007 493 23023
rect 537 23007 559 23023
rect 559 23007 571 23023
rect 615 23007 631 23023
rect 631 23007 649 23023
rect 693 23007 703 23023
rect 703 23007 727 23023
rect 771 23007 775 23023
rect 775 23007 805 23023
rect -17 22955 17 22968
rect 75 22955 109 22968
rect 167 22955 201 22968
rect 259 22955 293 22968
rect 459 22955 493 22968
rect 537 22955 571 22968
rect 615 22955 649 22968
rect 693 22955 727 22968
rect 771 22955 805 22968
rect -17 22934 17 22955
rect 75 22934 89 22955
rect 89 22934 109 22955
rect 167 22934 199 22955
rect 199 22934 201 22955
rect 259 22934 271 22955
rect 271 22934 293 22955
rect 459 22934 487 22955
rect 487 22934 493 22955
rect 537 22934 559 22955
rect 559 22934 571 22955
rect 615 22934 631 22955
rect 631 22934 649 22955
rect 693 22934 703 22955
rect 703 22934 727 22955
rect 771 22934 775 22955
rect 775 22934 805 22955
rect -17 22887 17 22895
rect 75 22887 109 22895
rect 167 22887 201 22895
rect 259 22887 293 22895
rect 459 22887 493 22895
rect 537 22887 571 22895
rect 615 22887 649 22895
rect 693 22887 727 22895
rect 771 22887 805 22895
rect -17 22861 17 22887
rect 75 22861 89 22887
rect 89 22861 109 22887
rect 167 22861 199 22887
rect 199 22861 201 22887
rect 259 22861 271 22887
rect 271 22861 293 22887
rect 459 22861 487 22887
rect 487 22861 493 22887
rect 537 22861 559 22887
rect 559 22861 571 22887
rect 615 22861 631 22887
rect 631 22861 649 22887
rect 693 22861 703 22887
rect 703 22861 727 22887
rect 771 22861 775 22887
rect 775 22861 805 22887
rect -17 22819 17 22822
rect 75 22819 109 22822
rect 167 22819 201 22822
rect 259 22819 293 22822
rect 459 22819 493 22822
rect 537 22819 571 22822
rect 615 22819 649 22822
rect 693 22819 727 22822
rect 771 22819 805 22822
rect -17 22788 17 22819
rect 75 22788 89 22819
rect 89 22788 109 22819
rect 167 22788 199 22819
rect 199 22788 201 22819
rect 259 22788 271 22819
rect 271 22788 293 22819
rect 459 22788 487 22819
rect 487 22788 493 22819
rect 537 22788 559 22819
rect 559 22788 571 22819
rect 615 22788 631 22819
rect 631 22788 649 22819
rect 693 22788 703 22819
rect 703 22788 727 22819
rect 771 22788 775 22819
rect 775 22788 805 22819
rect -17 22717 17 22749
rect 75 22717 89 22749
rect 89 22717 109 22749
rect 167 22717 199 22749
rect 199 22717 201 22749
rect 259 22717 271 22749
rect 271 22717 293 22749
rect 459 22717 487 22749
rect 487 22717 493 22749
rect 537 22717 559 22749
rect 559 22717 571 22749
rect 615 22717 631 22749
rect 631 22717 649 22749
rect 693 22717 703 22749
rect 703 22717 727 22749
rect 771 22717 775 22749
rect 775 22717 805 22749
rect -17 22715 17 22717
rect 75 22715 109 22717
rect 167 22715 201 22717
rect 259 22715 293 22717
rect 459 22715 493 22717
rect 537 22715 571 22717
rect 615 22715 649 22717
rect 693 22715 727 22717
rect 771 22715 805 22717
rect -17 22649 17 22676
rect 75 22649 89 22676
rect 89 22649 109 22676
rect 167 22649 199 22676
rect 199 22649 201 22676
rect 259 22649 271 22676
rect 271 22649 293 22676
rect 459 22649 487 22676
rect 487 22649 493 22676
rect 537 22649 559 22676
rect 559 22649 571 22676
rect 615 22649 631 22676
rect 631 22649 649 22676
rect 693 22649 703 22676
rect 703 22649 727 22676
rect 771 22649 775 22676
rect 775 22649 805 22676
rect -17 22642 17 22649
rect 75 22642 109 22649
rect 167 22642 201 22649
rect 259 22642 293 22649
rect 459 22642 493 22649
rect 537 22642 571 22649
rect 615 22642 649 22649
rect 693 22642 727 22649
rect 771 22642 805 22649
rect -17 22581 17 22603
rect 75 22581 89 22603
rect 89 22581 109 22603
rect 167 22581 199 22603
rect 199 22581 201 22603
rect 259 22581 271 22603
rect 271 22581 293 22603
rect 459 22581 487 22603
rect 487 22581 493 22603
rect 537 22581 559 22603
rect 559 22581 571 22603
rect 615 22581 631 22603
rect 631 22581 649 22603
rect 693 22581 703 22603
rect 703 22581 727 22603
rect 771 22581 775 22603
rect 775 22581 805 22603
rect -17 22569 17 22581
rect 75 22569 109 22581
rect 167 22569 201 22581
rect 259 22569 293 22581
rect 459 22569 493 22581
rect 537 22569 571 22581
rect 615 22569 649 22581
rect 693 22569 727 22581
rect 771 22569 805 22581
rect -17 22513 17 22530
rect 75 22513 89 22530
rect 89 22513 109 22530
rect 167 22513 199 22530
rect 199 22513 201 22530
rect 259 22513 271 22530
rect 271 22513 293 22530
rect 459 22513 487 22530
rect 487 22513 493 22530
rect 537 22513 559 22530
rect 559 22513 571 22530
rect 615 22513 631 22530
rect 631 22513 649 22530
rect 693 22513 703 22530
rect 703 22513 727 22530
rect 771 22513 775 22530
rect 775 22513 805 22530
rect -17 22496 17 22513
rect 75 22496 109 22513
rect 167 22496 201 22513
rect 259 22496 293 22513
rect 459 22496 493 22513
rect 537 22496 571 22513
rect 615 22496 649 22513
rect 693 22496 727 22513
rect 771 22496 805 22513
rect -17 22445 17 22457
rect 75 22445 89 22457
rect 89 22445 109 22457
rect 167 22445 199 22457
rect 199 22445 201 22457
rect 259 22445 271 22457
rect 271 22445 293 22457
rect 459 22445 487 22457
rect 487 22445 493 22457
rect 537 22445 559 22457
rect 559 22445 571 22457
rect 615 22445 631 22457
rect 631 22445 649 22457
rect 693 22445 703 22457
rect 703 22445 727 22457
rect 771 22445 775 22457
rect 775 22445 805 22457
rect -17 22423 17 22445
rect 75 22423 109 22445
rect 167 22423 201 22445
rect 259 22423 293 22445
rect 459 22423 493 22445
rect 537 22423 571 22445
rect 615 22423 649 22445
rect 693 22423 727 22445
rect 771 22423 805 22445
rect -17 22377 17 22384
rect 75 22377 89 22384
rect 89 22377 109 22384
rect 167 22377 199 22384
rect 199 22377 201 22384
rect 259 22377 271 22384
rect 271 22377 293 22384
rect 459 22377 487 22384
rect 487 22377 493 22384
rect 537 22377 559 22384
rect 559 22377 571 22384
rect 615 22377 631 22384
rect 631 22377 649 22384
rect 693 22377 703 22384
rect 703 22377 727 22384
rect 771 22377 775 22384
rect 775 22377 805 22384
rect -17 22350 17 22377
rect 75 22350 109 22377
rect 167 22350 201 22377
rect 259 22350 293 22377
rect 459 22350 493 22377
rect 537 22350 571 22377
rect 615 22350 649 22377
rect 693 22350 727 22377
rect 771 22350 805 22377
rect -17 22309 17 22311
rect 75 22309 89 22311
rect 89 22309 109 22311
rect 167 22309 199 22311
rect 199 22309 201 22311
rect 259 22309 271 22311
rect 271 22309 293 22311
rect 459 22309 487 22311
rect 487 22309 493 22311
rect 537 22309 559 22311
rect 559 22309 571 22311
rect 615 22309 631 22311
rect 631 22309 649 22311
rect 693 22309 703 22311
rect 703 22309 727 22311
rect 771 22309 775 22311
rect 775 22309 805 22311
rect -17 22277 17 22309
rect 75 22277 109 22309
rect 167 22277 201 22309
rect 259 22277 293 22309
rect 459 22277 493 22309
rect 537 22277 571 22309
rect 615 22277 649 22309
rect 693 22277 727 22309
rect 771 22277 805 22309
rect -17 22207 17 22238
rect 75 22207 109 22238
rect 167 22207 201 22238
rect 259 22207 293 22238
rect 459 22207 493 22238
rect 537 22207 571 22238
rect 615 22207 649 22238
rect 693 22207 727 22238
rect 771 22207 805 22238
rect -17 22204 17 22207
rect 75 22204 89 22207
rect 89 22204 109 22207
rect 167 22204 199 22207
rect 199 22204 201 22207
rect 259 22204 271 22207
rect 271 22204 293 22207
rect 459 22204 487 22207
rect 487 22204 493 22207
rect 537 22204 559 22207
rect 559 22204 571 22207
rect 615 22204 631 22207
rect 631 22204 649 22207
rect 693 22204 703 22207
rect 703 22204 727 22207
rect 771 22204 775 22207
rect 775 22204 805 22207
rect -17 22139 17 22165
rect 75 22139 109 22165
rect 167 22139 201 22165
rect 259 22139 293 22165
rect 459 22139 493 22165
rect 537 22139 571 22165
rect 615 22139 649 22165
rect 693 22139 727 22165
rect 771 22139 805 22165
rect -17 22131 17 22139
rect 75 22131 89 22139
rect 89 22131 109 22139
rect 167 22131 199 22139
rect 199 22131 201 22139
rect 259 22131 271 22139
rect 271 22131 293 22139
rect 459 22131 487 22139
rect 487 22131 493 22139
rect 537 22131 559 22139
rect 559 22131 571 22139
rect 615 22131 631 22139
rect 631 22131 649 22139
rect 693 22131 703 22139
rect 703 22131 727 22139
rect 771 22131 775 22139
rect 775 22131 805 22139
rect -17 22071 17 22092
rect 75 22071 109 22092
rect 167 22071 201 22092
rect 259 22071 293 22092
rect 459 22071 493 22092
rect 537 22071 571 22092
rect 615 22071 649 22092
rect 693 22071 727 22092
rect 771 22071 805 22092
rect -17 22058 17 22071
rect 75 22058 89 22071
rect 89 22058 109 22071
rect 167 22058 199 22071
rect 199 22058 201 22071
rect 259 22058 271 22071
rect 271 22058 293 22071
rect 459 22058 487 22071
rect 487 22058 493 22071
rect 537 22058 559 22071
rect 559 22058 571 22071
rect 615 22058 631 22071
rect 631 22058 649 22071
rect 693 22058 703 22071
rect 703 22058 727 22071
rect 771 22058 775 22071
rect 775 22058 805 22071
rect -17 22003 17 22019
rect 75 22003 109 22019
rect 167 22003 201 22019
rect 259 22003 293 22019
rect 459 22003 493 22019
rect 537 22003 571 22019
rect 615 22003 649 22019
rect 693 22003 727 22019
rect 771 22003 805 22019
rect -17 21985 17 22003
rect 75 21985 89 22003
rect 89 21985 109 22003
rect 167 21985 199 22003
rect 199 21985 201 22003
rect 259 21985 271 22003
rect 271 21985 293 22003
rect 459 21985 487 22003
rect 487 21985 493 22003
rect 537 21985 559 22003
rect 559 21985 571 22003
rect 615 21985 631 22003
rect 631 21985 649 22003
rect 693 21985 703 22003
rect 703 21985 727 22003
rect 771 21985 775 22003
rect 775 21985 805 22003
rect -17 21935 17 21946
rect 75 21935 109 21946
rect 167 21935 201 21946
rect 259 21935 293 21946
rect 459 21935 493 21946
rect 537 21935 571 21946
rect 615 21935 649 21946
rect 693 21935 727 21946
rect 771 21935 805 21946
rect -17 21912 17 21935
rect 75 21912 89 21935
rect 89 21912 109 21935
rect 167 21912 199 21935
rect 199 21912 201 21935
rect 259 21912 271 21935
rect 271 21912 293 21935
rect 459 21912 487 21935
rect 487 21912 493 21935
rect 537 21912 559 21935
rect 559 21912 571 21935
rect 615 21912 631 21935
rect 631 21912 649 21935
rect 693 21912 703 21935
rect 703 21912 727 21935
rect 771 21912 775 21935
rect 775 21912 805 21935
rect -17 21867 17 21873
rect 75 21867 109 21873
rect 167 21867 201 21873
rect 259 21867 293 21873
rect 459 21867 493 21873
rect 537 21867 571 21873
rect 615 21867 649 21873
rect 693 21867 727 21873
rect 771 21867 805 21873
rect -17 21839 17 21867
rect 75 21839 89 21867
rect 89 21839 109 21867
rect 167 21839 199 21867
rect 199 21839 201 21867
rect 259 21839 271 21867
rect 271 21839 293 21867
rect 459 21839 487 21867
rect 487 21839 493 21867
rect 537 21839 559 21867
rect 559 21839 571 21867
rect 615 21839 631 21867
rect 631 21839 649 21867
rect 693 21839 703 21867
rect 703 21839 727 21867
rect 771 21839 775 21867
rect 775 21839 805 21867
rect -17 21799 17 21800
rect 75 21799 109 21800
rect 167 21799 201 21800
rect 259 21799 293 21800
rect 459 21799 493 21800
rect 537 21799 571 21800
rect 615 21799 649 21800
rect 693 21799 727 21800
rect 771 21799 805 21800
rect -17 21766 17 21799
rect 75 21766 89 21799
rect 89 21766 109 21799
rect 167 21766 199 21799
rect 199 21766 201 21799
rect 259 21766 271 21799
rect 271 21766 293 21799
rect 459 21766 487 21799
rect 487 21766 493 21799
rect 537 21766 559 21799
rect 559 21766 571 21799
rect 615 21766 631 21799
rect 631 21766 649 21799
rect 693 21766 703 21799
rect 703 21766 727 21799
rect 771 21766 775 21799
rect 775 21766 805 21799
rect -17 21697 17 21727
rect 75 21697 89 21727
rect 89 21697 109 21727
rect 167 21697 199 21727
rect 199 21697 201 21727
rect 259 21697 271 21727
rect 271 21697 293 21727
rect 459 21697 487 21727
rect 487 21697 493 21727
rect 537 21697 559 21727
rect 559 21697 571 21727
rect 615 21697 631 21727
rect 631 21697 649 21727
rect 693 21697 703 21727
rect 703 21697 727 21727
rect 771 21697 775 21727
rect 775 21697 805 21727
rect -17 21693 17 21697
rect 75 21693 109 21697
rect 167 21693 201 21697
rect 259 21693 293 21697
rect 459 21693 493 21697
rect 537 21693 571 21697
rect 615 21693 649 21697
rect 693 21693 727 21697
rect 771 21693 805 21697
rect -17 21629 17 21654
rect 75 21629 89 21654
rect 89 21629 109 21654
rect 167 21629 199 21654
rect 199 21629 201 21654
rect 259 21629 271 21654
rect 271 21629 293 21654
rect 459 21629 487 21654
rect 487 21629 493 21654
rect 537 21629 559 21654
rect 559 21629 571 21654
rect 615 21629 631 21654
rect 631 21629 649 21654
rect 693 21629 703 21654
rect 703 21629 727 21654
rect 771 21629 775 21654
rect 775 21629 805 21654
rect -17 21620 17 21629
rect 75 21620 109 21629
rect 167 21620 201 21629
rect 259 21620 293 21629
rect 459 21620 493 21629
rect 537 21620 571 21629
rect 615 21620 649 21629
rect 693 21620 727 21629
rect 771 21620 805 21629
rect -17 21561 17 21581
rect 75 21561 89 21581
rect 89 21561 109 21581
rect 167 21561 199 21581
rect 199 21561 201 21581
rect 259 21561 271 21581
rect 271 21561 293 21581
rect 459 21561 487 21581
rect 487 21561 493 21581
rect 537 21561 559 21581
rect 559 21561 571 21581
rect 615 21561 631 21581
rect 631 21561 649 21581
rect 693 21561 703 21581
rect 703 21561 727 21581
rect 771 21561 775 21581
rect 775 21561 805 21581
rect -17 21547 17 21561
rect 75 21547 109 21561
rect 167 21547 201 21561
rect 259 21547 293 21561
rect 459 21547 493 21561
rect 537 21547 571 21561
rect 615 21547 649 21561
rect 693 21547 727 21561
rect 771 21547 805 21561
rect -17 21493 17 21508
rect 75 21493 89 21508
rect 89 21493 109 21508
rect 167 21493 199 21508
rect 199 21493 201 21508
rect 259 21493 271 21508
rect 271 21493 293 21508
rect 459 21493 487 21508
rect 487 21493 493 21508
rect 537 21493 559 21508
rect 559 21493 571 21508
rect 615 21493 631 21508
rect 631 21493 649 21508
rect 693 21493 703 21508
rect 703 21493 727 21508
rect 771 21493 775 21508
rect 775 21493 805 21508
rect -17 21474 17 21493
rect 75 21474 109 21493
rect 167 21474 201 21493
rect 259 21474 293 21493
rect 459 21474 493 21493
rect 537 21474 571 21493
rect 615 21474 649 21493
rect 693 21474 727 21493
rect 771 21474 805 21493
rect -17 21425 17 21435
rect 75 21425 89 21435
rect 89 21425 109 21435
rect 167 21425 199 21435
rect 199 21425 201 21435
rect 259 21425 271 21435
rect 271 21425 293 21435
rect 459 21425 487 21435
rect 487 21425 493 21435
rect 537 21425 559 21435
rect 559 21425 571 21435
rect 615 21425 631 21435
rect 631 21425 649 21435
rect 693 21425 703 21435
rect 703 21425 727 21435
rect 771 21425 775 21435
rect 775 21425 805 21435
rect -17 21401 17 21425
rect 75 21401 109 21425
rect 167 21401 201 21425
rect 259 21401 293 21425
rect 459 21401 493 21425
rect 537 21401 571 21425
rect 615 21401 649 21425
rect 693 21401 727 21425
rect 771 21401 805 21425
rect -17 21357 17 21362
rect 75 21357 89 21362
rect 89 21357 109 21362
rect 167 21357 199 21362
rect 199 21357 201 21362
rect 259 21357 271 21362
rect 271 21357 293 21362
rect 459 21357 487 21362
rect 487 21357 493 21362
rect 537 21357 559 21362
rect 559 21357 571 21362
rect 615 21357 631 21362
rect 631 21357 649 21362
rect 693 21357 703 21362
rect 703 21357 727 21362
rect 771 21357 775 21362
rect 775 21357 805 21362
rect -17 21328 17 21357
rect 75 21328 109 21357
rect 167 21328 201 21357
rect 259 21328 293 21357
rect 459 21328 493 21357
rect 537 21328 571 21357
rect 615 21328 649 21357
rect 693 21328 727 21357
rect 771 21328 805 21357
rect -17 21255 17 21289
rect 75 21255 109 21289
rect 167 21255 201 21289
rect 259 21255 293 21289
rect 459 21255 493 21289
rect 537 21255 571 21289
rect 615 21255 649 21289
rect 693 21255 727 21289
rect 771 21255 805 21289
rect -17 21187 17 21216
rect 75 21187 109 21216
rect 167 21187 201 21216
rect 259 21187 293 21216
rect 459 21187 493 21216
rect 537 21187 571 21216
rect 615 21187 649 21216
rect 693 21187 727 21216
rect 771 21187 805 21216
rect -17 21182 17 21187
rect 75 21182 89 21187
rect 89 21182 109 21187
rect 167 21182 199 21187
rect 199 21182 201 21187
rect 259 21182 271 21187
rect 271 21182 293 21187
rect 459 21182 487 21187
rect 487 21182 493 21187
rect 537 21182 559 21187
rect 559 21182 571 21187
rect 615 21182 631 21187
rect 631 21182 649 21187
rect 693 21182 703 21187
rect 703 21182 727 21187
rect 771 21182 775 21187
rect 775 21182 805 21187
rect -17 21119 17 21143
rect 75 21119 109 21143
rect 167 21119 201 21143
rect 259 21119 293 21143
rect 459 21119 493 21143
rect 537 21119 571 21143
rect 615 21119 649 21143
rect 693 21119 727 21143
rect 771 21119 805 21143
rect -17 21109 17 21119
rect 75 21109 89 21119
rect 89 21109 109 21119
rect 167 21109 199 21119
rect 199 21109 201 21119
rect 259 21109 271 21119
rect 271 21109 293 21119
rect 459 21109 487 21119
rect 487 21109 493 21119
rect 537 21109 559 21119
rect 559 21109 571 21119
rect 615 21109 631 21119
rect 631 21109 649 21119
rect 693 21109 703 21119
rect 703 21109 727 21119
rect 771 21109 775 21119
rect 775 21109 805 21119
rect -17 21051 17 21070
rect 75 21051 109 21070
rect 167 21051 201 21070
rect 259 21051 293 21070
rect 459 21051 493 21070
rect 537 21051 571 21070
rect 615 21051 649 21070
rect 693 21051 727 21070
rect 771 21051 805 21070
rect -17 21036 17 21051
rect 75 21036 89 21051
rect 89 21036 109 21051
rect 167 21036 199 21051
rect 199 21036 201 21051
rect 259 21036 271 21051
rect 271 21036 293 21051
rect 459 21036 487 21051
rect 487 21036 493 21051
rect 537 21036 559 21051
rect 559 21036 571 21051
rect 615 21036 631 21051
rect 631 21036 649 21051
rect 693 21036 703 21051
rect 703 21036 727 21051
rect 771 21036 775 21051
rect 775 21036 805 21051
rect -17 20983 17 20997
rect 75 20983 109 20997
rect 167 20983 201 20997
rect 259 20983 293 20997
rect 459 20983 493 20997
rect 537 20983 571 20997
rect 615 20983 649 20997
rect 693 20983 727 20997
rect 771 20983 805 20997
rect -17 20963 17 20983
rect 75 20963 89 20983
rect 89 20963 109 20983
rect 167 20963 199 20983
rect 199 20963 201 20983
rect 259 20963 271 20983
rect 271 20963 293 20983
rect 459 20963 487 20983
rect 487 20963 493 20983
rect 537 20963 559 20983
rect 559 20963 571 20983
rect 615 20963 631 20983
rect 631 20963 649 20983
rect 693 20963 703 20983
rect 703 20963 727 20983
rect 771 20963 775 20983
rect 775 20963 805 20983
rect -17 20915 17 20924
rect 75 20915 109 20924
rect 167 20915 201 20924
rect 259 20915 293 20924
rect 459 20915 493 20924
rect 537 20915 571 20924
rect 615 20915 649 20924
rect 693 20915 727 20924
rect 771 20915 805 20924
rect -17 20890 17 20915
rect 75 20890 89 20915
rect 89 20890 109 20915
rect 167 20890 199 20915
rect 199 20890 201 20915
rect 259 20890 271 20915
rect 271 20890 293 20915
rect 459 20890 487 20915
rect 487 20890 493 20915
rect 537 20890 559 20915
rect 559 20890 571 20915
rect 615 20890 631 20915
rect 631 20890 649 20915
rect 693 20890 703 20915
rect 703 20890 727 20915
rect 771 20890 775 20915
rect 775 20890 805 20915
rect -17 20847 17 20851
rect 75 20847 109 20851
rect 167 20847 201 20851
rect 259 20847 293 20851
rect 459 20847 493 20851
rect 537 20847 571 20851
rect 615 20847 649 20851
rect 693 20847 727 20851
rect 771 20847 805 20851
rect -17 20817 17 20847
rect 75 20817 89 20847
rect 89 20817 109 20847
rect 167 20817 199 20847
rect 199 20817 201 20847
rect 259 20817 271 20847
rect 271 20817 293 20847
rect 459 20817 487 20847
rect 487 20817 493 20847
rect 537 20817 559 20847
rect 559 20817 571 20847
rect 615 20817 631 20847
rect 631 20817 649 20847
rect 693 20817 703 20847
rect 703 20817 727 20847
rect 771 20817 775 20847
rect 775 20817 805 20847
rect -17 20745 17 20778
rect 75 20745 89 20778
rect 89 20745 109 20778
rect 167 20745 199 20778
rect 199 20745 201 20778
rect 259 20745 271 20778
rect 271 20745 293 20778
rect 459 20745 487 20778
rect 487 20745 493 20778
rect 537 20745 559 20778
rect 559 20745 571 20778
rect 615 20745 631 20778
rect 631 20745 649 20778
rect 693 20745 703 20778
rect 703 20745 727 20778
rect 771 20745 775 20778
rect 775 20745 805 20778
rect -17 20744 17 20745
rect 75 20744 109 20745
rect 167 20744 201 20745
rect 259 20744 293 20745
rect 459 20744 493 20745
rect 537 20744 571 20745
rect 615 20744 649 20745
rect 693 20744 727 20745
rect 771 20744 805 20745
rect -17 20677 17 20705
rect 75 20677 89 20705
rect 89 20677 109 20705
rect 167 20677 199 20705
rect 199 20677 201 20705
rect 259 20677 271 20705
rect 271 20677 293 20705
rect 459 20677 487 20705
rect 487 20677 493 20705
rect 537 20677 559 20705
rect 559 20677 571 20705
rect 615 20677 631 20705
rect 631 20677 649 20705
rect 693 20677 703 20705
rect 703 20677 727 20705
rect 771 20677 775 20705
rect 775 20677 805 20705
rect -17 20671 17 20677
rect 75 20671 109 20677
rect 167 20671 201 20677
rect 259 20671 293 20677
rect 459 20671 493 20677
rect 537 20671 571 20677
rect 615 20671 649 20677
rect 693 20671 727 20677
rect 771 20671 805 20677
rect -17 20609 17 20632
rect 75 20609 89 20632
rect 89 20609 109 20632
rect 167 20609 199 20632
rect 199 20609 201 20632
rect 259 20609 271 20632
rect 271 20609 293 20632
rect 459 20609 487 20632
rect 487 20609 493 20632
rect 537 20609 559 20632
rect 559 20609 571 20632
rect 615 20609 631 20632
rect 631 20609 649 20632
rect 693 20609 703 20632
rect 703 20609 727 20632
rect 771 20609 775 20632
rect 775 20609 805 20632
rect -17 20598 17 20609
rect 75 20598 109 20609
rect 167 20598 201 20609
rect 259 20598 293 20609
rect 459 20598 493 20609
rect 537 20598 571 20609
rect 615 20598 649 20609
rect 693 20598 727 20609
rect 771 20598 805 20609
rect -17 20541 17 20559
rect 75 20541 89 20559
rect 89 20541 109 20559
rect 167 20541 199 20559
rect 199 20541 201 20559
rect 259 20541 271 20559
rect 271 20541 293 20559
rect 459 20541 487 20559
rect 487 20541 493 20559
rect 537 20541 559 20559
rect 559 20541 571 20559
rect 615 20541 631 20559
rect 631 20541 649 20559
rect 693 20541 703 20559
rect 703 20541 727 20559
rect 771 20541 775 20559
rect 775 20541 805 20559
rect -17 20525 17 20541
rect 75 20525 109 20541
rect 167 20525 201 20541
rect 259 20525 293 20541
rect 459 20525 493 20541
rect 537 20525 571 20541
rect 615 20525 649 20541
rect 693 20525 727 20541
rect 771 20525 805 20541
rect -17 20473 17 20486
rect 75 20473 89 20486
rect 89 20473 109 20486
rect 167 20473 199 20486
rect 199 20473 201 20486
rect 259 20473 271 20486
rect 271 20473 293 20486
rect 459 20473 487 20486
rect 487 20473 493 20486
rect 537 20473 559 20486
rect 559 20473 571 20486
rect 615 20473 631 20486
rect 631 20473 649 20486
rect 693 20473 703 20486
rect 703 20473 727 20486
rect 771 20473 775 20486
rect 775 20473 805 20486
rect -17 20452 17 20473
rect 75 20452 109 20473
rect 167 20452 201 20473
rect 259 20452 293 20473
rect 459 20452 493 20473
rect 537 20452 571 20473
rect 615 20452 649 20473
rect 693 20452 727 20473
rect 771 20452 805 20473
rect -17 20405 17 20413
rect 75 20405 89 20413
rect 89 20405 109 20413
rect 167 20405 199 20413
rect 199 20405 201 20413
rect 259 20405 271 20413
rect 271 20405 293 20413
rect 868 20415 902 20418
rect 459 20405 487 20413
rect 487 20405 493 20413
rect 537 20405 559 20413
rect 559 20405 571 20413
rect 615 20405 631 20413
rect 631 20405 649 20413
rect 693 20405 703 20413
rect 703 20405 727 20413
rect -17 20379 17 20405
rect 75 20379 109 20405
rect 167 20379 201 20405
rect 259 20379 293 20405
rect 459 20379 493 20405
rect 537 20379 571 20405
rect 615 20379 649 20405
rect 693 20379 727 20405
rect 771 20379 775 20413
rect 775 20379 805 20413
rect 868 20384 877 20415
rect 877 20384 902 20415
rect -17 20337 17 20340
rect 75 20337 89 20340
rect 89 20337 109 20340
rect 167 20337 199 20340
rect 199 20337 201 20340
rect 259 20337 271 20340
rect 271 20337 293 20340
rect 459 20337 487 20340
rect 487 20337 493 20340
rect 537 20337 559 20340
rect 559 20337 571 20340
rect 615 20337 631 20340
rect 631 20337 649 20340
rect 693 20337 703 20340
rect 703 20337 727 20340
rect -17 20306 17 20337
rect 75 20306 109 20337
rect 167 20306 201 20337
rect 259 20306 293 20337
rect 459 20306 493 20337
rect 537 20306 571 20337
rect 615 20306 649 20337
rect 693 20306 727 20337
rect 771 20306 775 20340
rect 775 20306 805 20340
rect 868 20309 877 20343
rect 877 20309 902 20343
rect -17 20235 17 20267
rect 75 20235 109 20267
rect 167 20235 201 20267
rect 259 20235 293 20267
rect 459 20235 493 20267
rect 537 20235 571 20267
rect 615 20235 649 20267
rect 693 20235 727 20267
rect -17 20233 17 20235
rect 75 20233 89 20235
rect 89 20233 109 20235
rect 167 20233 199 20235
rect 199 20233 201 20235
rect 259 20233 271 20235
rect 271 20233 293 20235
rect 459 20233 487 20235
rect 487 20233 493 20235
rect 537 20233 559 20235
rect 559 20233 571 20235
rect 615 20233 631 20235
rect 631 20233 649 20235
rect 693 20233 703 20235
rect 703 20233 727 20235
rect 771 20233 775 20267
rect 775 20233 805 20267
rect 868 20234 877 20268
rect 877 20234 902 20268
rect -17 20167 17 20194
rect 75 20167 109 20194
rect 167 20167 201 20194
rect 259 20167 293 20194
rect 459 20167 493 20194
rect 537 20167 571 20194
rect 615 20167 649 20194
rect 693 20167 727 20194
rect -17 20160 17 20167
rect 75 20160 89 20167
rect 89 20160 109 20167
rect 167 20160 199 20167
rect 199 20160 201 20167
rect 259 20160 271 20167
rect 271 20160 293 20167
rect 459 20160 487 20167
rect 487 20160 493 20167
rect 537 20160 559 20167
rect 559 20160 571 20167
rect 615 20160 631 20167
rect 631 20160 649 20167
rect 693 20160 703 20167
rect 703 20160 727 20167
rect 771 20160 775 20194
rect 775 20160 805 20194
rect 868 20159 877 20193
rect 877 20159 902 20193
rect -17 20099 17 20121
rect 75 20099 109 20121
rect 167 20099 201 20121
rect 259 20099 293 20121
rect 459 20099 493 20121
rect 537 20099 571 20121
rect 615 20099 649 20121
rect 693 20099 727 20121
rect -17 20087 17 20099
rect 75 20087 89 20099
rect 89 20087 109 20099
rect 167 20087 199 20099
rect 199 20087 201 20099
rect 259 20087 271 20099
rect 271 20087 293 20099
rect 459 20087 487 20099
rect 487 20087 493 20099
rect 537 20087 559 20099
rect 559 20087 571 20099
rect 615 20087 631 20099
rect 631 20087 649 20099
rect 693 20087 703 20099
rect 703 20087 727 20099
rect 771 20087 775 20121
rect 775 20087 805 20121
rect 868 20083 877 20117
rect 877 20083 902 20117
rect -17 20031 17 20048
rect 75 20031 109 20048
rect 167 20031 201 20048
rect 259 20031 293 20048
rect 459 20031 493 20048
rect 537 20031 571 20048
rect 615 20031 649 20048
rect 693 20031 727 20048
rect -17 20014 17 20031
rect 75 20014 89 20031
rect 89 20014 109 20031
rect 167 20014 199 20031
rect 199 20014 201 20031
rect 259 20014 271 20031
rect 271 20014 293 20031
rect 459 20014 487 20031
rect 487 20014 493 20031
rect 537 20014 559 20031
rect 559 20014 571 20031
rect 615 20014 631 20031
rect 631 20014 649 20031
rect 693 20014 703 20031
rect 703 20014 727 20031
rect 771 20014 775 20048
rect 775 20014 805 20048
rect 868 20007 877 20041
rect 877 20007 902 20041
rect -17 19963 17 19975
rect 75 19963 109 19975
rect 167 19963 201 19975
rect 259 19963 293 19975
rect 459 19963 493 19975
rect 537 19963 571 19975
rect 615 19963 649 19975
rect 693 19963 727 19975
rect -17 19941 17 19963
rect 75 19941 89 19963
rect 89 19941 109 19963
rect 167 19941 199 19963
rect 199 19941 201 19963
rect 259 19941 271 19963
rect 271 19941 293 19963
rect 459 19941 487 19963
rect 487 19941 493 19963
rect 537 19941 559 19963
rect 559 19941 571 19963
rect 615 19941 631 19963
rect 631 19941 649 19963
rect 693 19941 703 19963
rect 703 19941 727 19963
rect 771 19941 775 19975
rect 775 19941 805 19975
rect 868 19931 877 19965
rect 877 19931 902 19965
rect -17 19895 17 19902
rect 75 19895 109 19902
rect 167 19895 201 19902
rect 259 19895 293 19902
rect 459 19895 493 19902
rect 537 19895 571 19902
rect 615 19895 649 19902
rect 693 19895 727 19902
rect -17 19868 17 19895
rect 75 19868 89 19895
rect 89 19868 109 19895
rect 167 19868 199 19895
rect 199 19868 201 19895
rect 259 19868 271 19895
rect 271 19868 293 19895
rect 459 19868 487 19895
rect 487 19868 493 19895
rect 537 19868 559 19895
rect 559 19868 571 19895
rect 615 19868 631 19895
rect 631 19868 649 19895
rect 693 19868 703 19895
rect 703 19868 727 19895
rect 771 19868 775 19902
rect 775 19868 805 19902
rect 868 19855 877 19889
rect 877 19855 902 19889
rect -17 19827 17 19829
rect 75 19827 109 19829
rect 167 19827 201 19829
rect 259 19827 293 19829
rect 459 19827 493 19829
rect 537 19827 571 19829
rect 615 19827 649 19829
rect 693 19827 727 19829
rect -17 19795 17 19827
rect 75 19795 89 19827
rect 89 19795 109 19827
rect 167 19795 199 19827
rect 199 19795 201 19827
rect 259 19795 271 19827
rect 271 19795 293 19827
rect 459 19795 487 19827
rect 487 19795 493 19827
rect 537 19795 559 19827
rect 559 19795 571 19827
rect 615 19795 631 19827
rect 631 19795 649 19827
rect 693 19795 703 19827
rect 703 19795 727 19827
rect 771 19795 775 19829
rect 775 19795 805 19829
rect 868 19779 877 19813
rect 877 19779 902 19813
rect -17 19725 17 19756
rect 75 19725 89 19756
rect 89 19725 109 19756
rect 167 19725 199 19756
rect 199 19725 201 19756
rect 259 19725 271 19756
rect 271 19725 293 19756
rect 459 19725 487 19756
rect 487 19725 493 19756
rect 537 19725 559 19756
rect 559 19725 571 19756
rect 615 19725 631 19756
rect 631 19725 649 19756
rect 693 19725 703 19756
rect 703 19725 727 19756
rect -17 19722 17 19725
rect 75 19722 109 19725
rect 167 19722 201 19725
rect 259 19722 293 19725
rect 459 19722 493 19725
rect 537 19722 571 19725
rect 615 19722 649 19725
rect 693 19722 727 19725
rect 771 19722 775 19756
rect 775 19722 805 19756
rect 868 19703 877 19737
rect 877 19703 902 19737
rect -17 19657 17 19683
rect 75 19657 89 19683
rect 89 19657 109 19683
rect 167 19657 199 19683
rect 199 19657 201 19683
rect 259 19657 271 19683
rect 271 19657 293 19683
rect 459 19657 487 19683
rect 487 19657 493 19683
rect 537 19657 559 19683
rect 559 19657 571 19683
rect 615 19657 631 19683
rect 631 19657 649 19683
rect 693 19657 703 19683
rect 703 19657 727 19683
rect -17 19649 17 19657
rect 75 19649 109 19657
rect 167 19649 201 19657
rect 259 19649 293 19657
rect 459 19649 493 19657
rect 537 19649 571 19657
rect 615 19649 649 19657
rect 693 19649 727 19657
rect 771 19649 775 19683
rect 775 19649 805 19683
rect 868 19627 877 19661
rect 877 19627 902 19661
rect -17 19589 17 19610
rect 75 19589 89 19610
rect 89 19589 109 19610
rect 167 19589 199 19610
rect 199 19589 201 19610
rect 259 19589 271 19610
rect 271 19589 293 19610
rect 459 19589 487 19610
rect 487 19589 493 19610
rect 537 19589 559 19610
rect 559 19589 571 19610
rect 615 19589 631 19610
rect 631 19589 649 19610
rect 693 19589 703 19610
rect 703 19589 727 19610
rect -17 19576 17 19589
rect 75 19576 109 19589
rect 167 19576 201 19589
rect 259 19576 293 19589
rect 459 19576 493 19589
rect 537 19576 571 19589
rect 615 19576 649 19589
rect 693 19576 727 19589
rect 771 19576 775 19610
rect 775 19576 805 19610
rect -17 19521 17 19537
rect 75 19521 89 19537
rect 89 19521 109 19537
rect 167 19521 199 19537
rect 199 19521 201 19537
rect 259 19521 271 19537
rect 271 19521 293 19537
rect 868 19551 877 19585
rect 877 19551 902 19585
rect 459 19521 487 19537
rect 487 19521 493 19537
rect 537 19521 559 19537
rect 559 19521 571 19537
rect 615 19521 631 19537
rect 631 19521 649 19537
rect 693 19521 703 19537
rect 703 19521 727 19537
rect -17 19503 17 19521
rect 75 19503 109 19521
rect 167 19503 201 19521
rect 259 19503 293 19521
rect 459 19503 493 19521
rect 537 19503 571 19521
rect 615 19503 649 19521
rect 693 19503 727 19521
rect 771 19503 775 19537
rect 775 19503 805 19537
rect -17 19453 17 19464
rect 75 19453 89 19464
rect 89 19453 109 19464
rect 167 19453 199 19464
rect 199 19453 201 19464
rect 259 19453 271 19464
rect 271 19453 293 19464
rect 868 19475 877 19509
rect 877 19475 902 19509
rect 459 19453 487 19464
rect 487 19453 493 19464
rect 537 19453 559 19464
rect 559 19453 571 19464
rect 615 19453 631 19464
rect 631 19453 649 19464
rect 693 19453 703 19464
rect 703 19453 727 19464
rect -17 19430 17 19453
rect 75 19430 109 19453
rect 167 19430 201 19453
rect 259 19430 293 19453
rect 459 19430 493 19453
rect 537 19430 571 19453
rect 615 19430 649 19453
rect 693 19430 727 19453
rect 771 19430 775 19464
rect 775 19430 805 19464
rect -17 19385 17 19391
rect 75 19385 89 19391
rect 89 19385 109 19391
rect 167 19385 199 19391
rect 199 19385 201 19391
rect 259 19385 271 19391
rect 271 19385 293 19391
rect 868 19399 877 19433
rect 877 19399 902 19433
rect 459 19385 487 19391
rect 487 19385 493 19391
rect 537 19385 559 19391
rect 559 19385 571 19391
rect 615 19385 631 19391
rect 631 19385 649 19391
rect 693 19385 703 19391
rect 703 19385 727 19391
rect -17 19357 17 19385
rect 75 19357 109 19385
rect 167 19357 201 19385
rect 259 19357 293 19385
rect 459 19357 493 19385
rect 537 19357 571 19385
rect 615 19357 649 19385
rect 693 19357 727 19385
rect 771 19357 775 19391
rect 775 19357 805 19391
rect -17 19317 17 19318
rect 75 19317 89 19318
rect 89 19317 109 19318
rect 167 19317 199 19318
rect 199 19317 201 19318
rect 259 19317 271 19318
rect 271 19317 293 19318
rect 868 19323 877 19357
rect 877 19323 902 19357
rect 459 19317 487 19318
rect 487 19317 493 19318
rect 537 19317 559 19318
rect 559 19317 571 19318
rect 615 19317 631 19318
rect 631 19317 649 19318
rect 693 19317 703 19318
rect 703 19317 727 19318
rect -17 19284 17 19317
rect 75 19284 109 19317
rect 167 19284 201 19317
rect 259 19284 293 19317
rect 459 19284 493 19317
rect 537 19284 571 19317
rect 615 19284 649 19317
rect 693 19284 727 19317
rect 771 19284 775 19318
rect 775 19284 805 19318
rect 868 19247 877 19281
rect 877 19247 902 19281
rect -17 19215 17 19245
rect 75 19215 109 19245
rect 167 19215 201 19245
rect 259 19215 293 19245
rect 459 19215 493 19245
rect 537 19215 571 19245
rect 615 19215 649 19245
rect 693 19215 727 19245
rect -17 19211 17 19215
rect 75 19211 89 19215
rect 89 19211 109 19215
rect 167 19211 199 19215
rect 199 19211 201 19215
rect 259 19211 271 19215
rect 271 19211 293 19215
rect 459 19211 487 19215
rect 487 19211 493 19215
rect 537 19211 559 19215
rect 559 19211 571 19215
rect 615 19211 631 19215
rect 631 19211 649 19215
rect 693 19211 703 19215
rect 703 19211 727 19215
rect 771 19211 775 19245
rect 775 19211 805 19245
rect 472 19147 506 19153
rect 545 19147 579 19153
rect 618 19147 652 19153
rect 691 19147 725 19153
rect 472 19119 487 19147
rect 487 19119 506 19147
rect 545 19119 559 19147
rect 559 19119 579 19147
rect 618 19119 631 19147
rect 631 19119 652 19147
rect 691 19119 703 19147
rect 703 19119 725 19147
rect 764 19119 775 19153
rect 775 19119 798 19153
rect 837 19119 871 19153
rect 910 19119 915 19153
rect 915 19119 944 19153
rect 983 19119 1017 19153
rect 1056 19123 1058 19153
rect 1058 19123 1090 19153
rect 1129 19123 1133 19153
rect 1133 19123 1163 19153
rect 1202 19123 1208 19153
rect 1208 19123 1236 19153
rect 1275 19123 1283 19153
rect 1283 19123 1309 19153
rect 1348 19123 1358 19153
rect 1358 19123 1382 19153
rect 1420 19123 1433 19153
rect 1433 19123 1454 19153
rect 1492 19123 1508 19153
rect 1508 19123 1526 19153
rect 1564 19123 1583 19153
rect 1583 19123 1598 19153
rect 1636 19123 1658 19153
rect 1658 19123 1670 19153
rect 1056 19119 1090 19123
rect 1129 19119 1163 19123
rect 1202 19119 1236 19123
rect 1275 19119 1309 19123
rect 1348 19119 1382 19123
rect 1420 19119 1454 19123
rect 1492 19119 1526 19123
rect 1564 19119 1598 19123
rect 1636 19119 1670 19123
rect 1708 19119 1729 19153
rect 1729 19119 1742 19153
rect 472 19045 487 19063
rect 487 19045 506 19063
rect 545 19045 559 19063
rect 559 19045 579 19063
rect 618 19045 631 19063
rect 631 19045 652 19063
rect 691 19045 703 19063
rect 703 19045 725 19063
rect 472 19029 506 19045
rect 545 19029 579 19045
rect 618 19029 652 19045
rect 691 19029 725 19045
rect 764 19029 775 19063
rect 775 19029 798 19063
rect 837 19029 871 19063
rect 910 19029 915 19063
rect 915 19029 944 19063
rect 983 19029 1017 19063
rect 1056 19055 1058 19063
rect 1058 19055 1090 19063
rect 1129 19055 1133 19063
rect 1133 19055 1163 19063
rect 1202 19055 1208 19063
rect 1208 19055 1236 19063
rect 1275 19055 1283 19063
rect 1283 19055 1309 19063
rect 1348 19055 1358 19063
rect 1358 19055 1382 19063
rect 1420 19055 1433 19063
rect 1433 19055 1454 19063
rect 1492 19055 1508 19063
rect 1508 19055 1526 19063
rect 1564 19055 1583 19063
rect 1583 19055 1598 19063
rect 1636 19055 1658 19063
rect 1658 19055 1670 19063
rect 1056 19029 1090 19055
rect 1129 19029 1163 19055
rect 1202 19029 1236 19055
rect 1275 19029 1309 19055
rect 1348 19029 1382 19055
rect 1420 19029 1454 19055
rect 1492 19029 1526 19055
rect 1564 19029 1598 19055
rect 1636 19029 1670 19055
rect 1708 19047 1729 19063
rect 1729 19047 1742 19063
rect 1708 19029 1742 19047
rect 1584 18135 1606 18158
rect 1606 18135 1652 18158
rect 1652 18135 1686 18158
rect 1686 18135 1732 18158
rect 1732 18135 1762 18158
rect 1584 18100 1762 18135
rect 1584 18066 1606 18100
rect 1606 18066 1652 18100
rect 1652 18066 1686 18100
rect 1686 18066 1732 18100
rect 1732 18066 1762 18100
rect 1584 18031 1762 18066
rect 1584 17997 1606 18031
rect 1606 17997 1652 18031
rect 1652 17997 1686 18031
rect 1686 17997 1732 18031
rect 1732 17997 1762 18031
rect 1584 17962 1762 17997
rect 1584 17928 1606 17962
rect 1606 17928 1652 17962
rect 1652 17928 1686 17962
rect 1686 17928 1732 17962
rect 1732 17928 1762 17962
rect 1584 17908 1762 17928
rect 1584 17859 1606 17869
rect 1606 17859 1618 17869
rect 1656 17859 1686 17869
rect 1686 17859 1690 17869
rect 1584 17835 1618 17859
rect 1656 17835 1690 17859
rect 1728 17859 1732 17869
rect 1732 17859 1762 17869
rect 1728 17835 1762 17859
rect 5535 13855 5569 13889
rect 5608 13855 5642 13889
rect 5681 13855 5715 13889
rect 5754 13855 5788 13889
rect 5827 13855 5861 13889
rect 5900 13855 5934 13889
rect 5535 13747 5569 13781
rect 5608 13747 5642 13781
rect 5681 13747 5715 13781
rect 5754 13747 5788 13781
rect 5827 13747 5861 13781
rect 5900 13747 5934 13781
rect 5305 13529 5339 13563
rect 5380 13529 5414 13563
rect 5455 13529 5489 13563
rect 5530 13529 5564 13563
rect 5604 13529 5638 13563
rect 5678 13529 5712 13563
rect 5752 13529 5786 13563
rect 5826 13529 5860 13563
rect 5900 13529 5934 13563
rect 5305 13421 5339 13455
rect 5380 13421 5414 13455
rect 5455 13421 5489 13455
rect 5530 13421 5564 13455
rect 5604 13421 5638 13455
rect 5678 13421 5712 13455
rect 5752 13421 5786 13455
rect 5826 13421 5860 13455
rect 5900 13421 5934 13455
rect 5498 12876 5532 12910
rect 5581 12876 5615 12910
rect 5664 12876 5698 12910
rect 5747 12876 5781 12910
rect 5829 12876 5863 12910
rect 5498 12794 5532 12828
rect 5581 12794 5615 12828
rect 5664 12794 5698 12828
rect 5747 12794 5781 12828
rect 5829 12794 5863 12828
rect 5186 11991 5220 12025
rect 5266 11991 5300 12025
rect 5346 11991 5380 12025
rect 5426 11991 5460 12025
rect 5506 11991 5540 12025
rect 5586 11991 5620 12025
rect 5186 11905 5220 11939
rect 5266 11905 5300 11939
rect 5346 11905 5380 11939
rect 5426 11905 5460 11939
rect 5506 11905 5540 11939
rect 5586 11905 5620 11939
rect 5186 11819 5220 11853
rect 5266 11819 5300 11853
rect 5346 11819 5380 11853
rect 5426 11819 5460 11853
rect 5506 11819 5540 11853
rect 5586 11819 5620 11853
rect 5668 11908 5702 11942
rect 5668 11836 5702 11870
rect 5187 11739 5221 11773
rect 5260 11739 5294 11773
rect 5333 11739 5367 11773
rect 5406 11739 5440 11773
rect 5479 11739 5513 11773
rect 5552 11739 5586 11773
rect 5624 11739 5658 11773
rect 5696 11739 5730 11773
rect 5768 11739 5802 11773
rect 5840 11739 5874 11773
rect 5187 11665 5221 11699
rect 5260 11665 5294 11699
rect 5333 11665 5367 11699
rect 5406 11665 5440 11699
rect 5479 11665 5513 11699
rect 5552 11665 5586 11699
rect 5624 11665 5658 11699
rect 5696 11665 5730 11699
rect 5768 11665 5802 11699
rect 5840 11665 5874 11699
rect 5187 11591 5221 11625
rect 5260 11591 5294 11625
rect 5333 11591 5367 11625
rect 5406 11591 5440 11625
rect 5479 11591 5513 11625
rect 5552 11591 5586 11625
rect 5624 11591 5658 11625
rect 5696 11591 5730 11625
rect 5768 11591 5802 11625
rect 5840 11591 5874 11625
rect 5187 11517 5221 11551
rect 5260 11517 5294 11551
rect 5333 11517 5367 11551
rect 5406 11517 5440 11551
rect 5479 11517 5513 11551
rect 5552 11517 5586 11551
rect 5624 11517 5658 11551
rect 5696 11517 5730 11551
rect 5768 11517 5802 11551
rect 5840 11517 5874 11551
rect 5807 11351 5913 11457
rect 359 9109 362 9143
rect 362 9109 393 9143
rect 443 9109 467 9143
rect 467 9109 477 9143
rect 527 9109 538 9143
rect 538 9109 561 9143
rect 611 9109 645 9143
rect 694 9109 717 9143
rect 717 9109 728 9143
rect 777 9109 788 9143
rect 788 9109 811 9143
rect 860 9109 893 9143
rect 893 9109 894 9143
rect 15983 7121 16017 7133
rect 15983 7099 16017 7121
rect 15983 7052 16017 7061
rect 15983 7027 16017 7052
rect 15983 6983 16017 6989
rect 15983 6955 16017 6983
rect 15983 6914 16017 6917
rect 15983 6883 16017 6914
rect 15983 6811 16017 6845
rect 15983 6742 16017 6773
rect 15983 6739 16017 6742
rect 15983 6673 16017 6701
rect 15983 6667 16017 6673
rect 15983 6604 16017 6629
rect 15983 6595 16017 6604
rect 15983 6535 16017 6557
rect 15983 6523 16017 6535
rect 15983 6466 16017 6485
rect 15983 6451 16017 6466
rect 15983 6397 16017 6413
rect 15983 6379 16017 6397
rect 15983 6327 16017 6341
rect 15983 6307 16017 6327
rect 15983 6257 16017 6269
rect 15983 6235 16017 6257
rect 15983 6187 16017 6197
rect 15983 6163 16017 6187
rect 15983 6117 16017 6125
rect 15983 6091 16017 6117
rect 15983 4979 16017 4991
rect 15983 4957 16017 4979
rect 15983 4911 16017 4919
rect 15983 4885 16017 4911
rect 15983 4843 16017 4847
rect 15983 4813 16017 4843
rect 15983 4741 16017 4775
rect 15983 4673 16017 4703
rect 15983 4669 16017 4673
rect 15983 4605 16017 4631
rect 15983 4597 16017 4605
rect 15983 4537 16017 4559
rect 15983 4525 16017 4537
rect 15983 4469 16017 4487
rect 15983 4453 16017 4469
rect 15983 4401 16017 4415
rect 15983 4381 16017 4401
rect 15983 4333 16017 4343
rect 15983 4309 16017 4333
rect 15983 4265 16017 4271
rect 15983 4237 16017 4265
rect 15983 4197 16017 4199
rect 15983 4165 16017 4197
rect 15983 4093 16017 4127
rect 15983 4024 16017 4055
rect 15983 4021 16017 4024
rect 15983 3955 16017 3983
rect 15983 3949 16017 3955
rect 13949 2061 13967 2068
rect 13967 2061 13983 2068
rect 14031 2061 14040 2068
rect 14040 2061 14065 2068
rect 13949 2034 13983 2061
rect 14031 2034 14065 2061
rect 14113 2034 14147 2068
rect 14195 2061 14224 2068
rect 14224 2061 14229 2068
rect 14277 2061 14296 2068
rect 14296 2061 14311 2068
rect 14195 2034 14229 2061
rect 14277 2034 14311 2061
rect 13782 2003 13796 2024
rect 13796 2003 13816 2024
rect 13854 2003 13865 2024
rect 13865 2003 13888 2024
rect 13782 1990 13816 2003
rect 13854 1990 13888 2003
rect 13451 1915 13485 1949
rect 13529 1915 13554 1949
rect 13554 1915 13563 1949
rect 13607 1915 13623 1949
rect 13623 1915 13641 1949
rect 13685 1915 13692 1949
rect 13692 1915 13719 1949
rect 13762 1915 13796 1949
rect 13839 1915 13865 1949
rect 13865 1915 13873 1949
rect 13379 1846 13385 1873
rect 13385 1846 13413 1873
rect 13379 1839 13413 1846
rect 13379 1776 13385 1797
rect 13385 1776 13413 1797
rect 13379 1763 13413 1776
rect 13379 1706 13385 1721
rect 13385 1706 13413 1721
rect 13379 1687 13413 1706
rect 12312 1050 12346 1069
rect 12387 1050 12421 1069
rect 12462 1050 12496 1069
rect 12536 1050 12570 1069
rect 12610 1050 12644 1069
rect 12684 1050 12718 1069
rect 12312 1035 12332 1050
rect 12332 1035 12346 1050
rect 12387 1035 12403 1050
rect 12403 1035 12421 1050
rect 12462 1035 12474 1050
rect 12474 1035 12496 1050
rect 12536 1035 12545 1050
rect 12545 1035 12570 1050
rect 12610 1035 12616 1050
rect 12616 1035 12644 1050
rect 12684 1035 12687 1050
rect 12687 1035 12718 1050
rect 12758 1035 12792 1069
rect 12832 1035 12866 1069
rect 12906 1050 12940 1069
rect 12980 1050 13014 1069
rect 13054 1050 13088 1069
rect 13128 1050 13162 1069
rect 13202 1050 13236 1069
rect 13276 1050 13310 1069
rect 13350 1050 13384 1069
rect 12906 1035 12937 1050
rect 12937 1035 12940 1050
rect 12980 1035 13008 1050
rect 13008 1035 13014 1050
rect 13054 1035 13079 1050
rect 13079 1035 13088 1050
rect 13128 1035 13150 1050
rect 13150 1035 13162 1050
rect 13202 1035 13221 1050
rect 13221 1035 13236 1050
rect 13276 1035 13292 1050
rect 13292 1035 13310 1050
rect 13350 1035 13362 1050
rect 13362 1035 13384 1050
rect 13424 1035 13458 1069
rect 12312 953 12346 987
rect 12387 953 12421 987
rect 12462 953 12496 987
rect 12536 953 12570 987
rect 12610 953 12644 987
rect 12684 953 12718 987
rect 12758 953 12792 987
rect 12832 953 12866 987
rect 12906 953 12940 987
rect 12980 953 13014 987
rect 13054 953 13088 987
rect 13128 953 13162 987
rect 13202 953 13236 987
rect 13276 953 13310 987
rect 13350 953 13384 987
rect 13424 953 13458 987
rect 15439 1000 15473 1034
rect 15521 1000 15555 1034
rect 15439 914 15473 948
rect 15521 914 15555 948
rect 11899 524 11933 558
rect 11899 452 11933 486
rect 13664 606 13770 784
rect 13664 533 13698 567
rect 13736 533 13770 567
rect 13664 460 13698 494
rect 13736 460 13770 494
rect 15439 828 15473 862
rect 15521 828 15555 862
rect 15439 741 15473 775
rect 15521 741 15555 775
rect 12887 142 12909 171
rect 12909 142 12921 171
rect 12887 137 12921 142
rect 12960 142 12977 171
rect 12977 142 12994 171
rect 12960 137 12994 142
rect 13033 137 13067 171
rect 13105 142 13113 171
rect 13113 142 13139 171
rect 13105 137 13139 142
rect 13177 142 13181 171
rect 13181 142 13211 171
rect 13177 137 13211 142
rect 12887 74 12909 93
rect 12909 74 12921 93
rect 12887 59 12921 74
rect 12960 74 12977 93
rect 12977 74 12994 93
rect 12960 59 12994 74
rect 13033 59 13067 93
rect 13105 74 13113 93
rect 13113 74 13139 93
rect 13105 59 13139 74
rect 13177 74 13181 93
rect 13181 74 13211 93
rect 13177 59 13211 74
<< metal1 >>
rect 14399 39998 15371 40000
rect 3154 39994 11343 39995
rect 3154 39942 3160 39994
rect 3212 39942 3225 39994
rect 3277 39942 3290 39994
rect 3342 39942 3355 39994
rect 3407 39942 3420 39994
rect 3472 39942 3485 39994
rect 3537 39942 3550 39994
rect 3602 39942 3615 39994
rect 3667 39942 3680 39994
rect 3732 39942 3745 39994
rect 3797 39942 3810 39994
rect 3862 39942 3875 39994
rect 3927 39942 3940 39994
rect 3992 39942 4005 39994
rect 4057 39942 4070 39994
rect 4122 39942 4135 39994
rect 4187 39942 4200 39994
rect 4252 39942 4265 39994
rect 4317 39942 4330 39994
rect 4382 39942 4395 39994
rect 4447 39942 4460 39994
rect 4512 39942 4525 39994
rect 4577 39942 4590 39994
rect 4642 39942 4655 39994
rect 4707 39942 4720 39994
rect 4772 39942 4785 39994
rect 4837 39942 4850 39994
rect 4902 39942 4915 39994
rect 4967 39942 4980 39994
rect 5032 39942 5045 39994
rect 5097 39942 5110 39994
rect 5162 39942 5175 39994
rect 5227 39942 5240 39994
rect 5292 39942 5305 39994
rect 5357 39942 5370 39994
rect 5422 39942 5435 39994
rect 5487 39942 5500 39994
rect 5552 39942 5565 39994
rect 5617 39942 5630 39994
rect 5682 39942 5695 39994
rect 5747 39942 5760 39994
rect 5812 39942 5825 39994
rect 5877 39942 5890 39994
rect 5942 39942 5955 39994
rect 6007 39942 6020 39994
rect 6072 39942 6085 39994
rect 6137 39942 6150 39994
rect 6202 39942 6215 39994
rect 6267 39942 6280 39994
rect 6332 39942 6345 39994
rect 6397 39942 6410 39994
rect 6462 39942 6475 39994
rect 6527 39942 6540 39994
rect 6592 39942 6605 39994
rect 6657 39942 6670 39994
rect 6722 39942 6735 39994
rect 6787 39942 6800 39994
rect 6852 39942 6865 39994
rect 6917 39942 6930 39994
rect 6982 39942 6995 39994
rect 7047 39942 7060 39994
rect 7112 39942 7125 39994
rect 7177 39942 7189 39994
rect 7241 39942 7253 39994
rect 7305 39942 7317 39994
rect 7369 39942 7381 39994
rect 7433 39942 7445 39994
rect 7497 39942 7509 39994
rect 7561 39942 7573 39994
rect 7625 39942 7637 39994
rect 7689 39942 7701 39994
rect 7753 39942 7765 39994
rect 7817 39942 7829 39994
rect 7881 39942 7893 39994
rect 7945 39942 7957 39994
rect 8009 39942 8021 39994
rect 8073 39942 8085 39994
rect 8137 39942 8149 39994
rect 8201 39942 8213 39994
rect 8265 39942 8277 39994
rect 8329 39942 8341 39994
rect 8393 39942 8405 39994
rect 8457 39942 8469 39994
rect 8521 39942 8533 39994
rect 8585 39942 8597 39994
rect 8649 39942 8661 39994
rect 8713 39942 8725 39994
rect 8777 39942 8789 39994
rect 8841 39942 8853 39994
rect 8905 39942 8917 39994
rect 8969 39942 8981 39994
rect 9033 39942 9045 39994
rect 9097 39942 9109 39994
rect 9161 39942 9173 39994
rect 9225 39942 9237 39994
rect 9289 39942 9301 39994
rect 9353 39942 9365 39994
rect 9417 39942 9429 39994
rect 9481 39942 9493 39994
rect 9545 39942 9557 39994
rect 9609 39942 9621 39994
rect 9673 39942 9685 39994
rect 9737 39942 9749 39994
rect 9801 39942 9813 39994
rect 9865 39942 9877 39994
rect 9929 39942 9941 39994
rect 9993 39942 10005 39994
rect 10057 39942 10069 39994
rect 10121 39942 10133 39994
rect 10185 39942 10197 39994
rect 10249 39942 10261 39994
rect 10313 39942 10325 39994
rect 10377 39942 10389 39994
rect 10441 39942 10453 39994
rect 10505 39942 10517 39994
rect 10569 39942 10581 39994
rect 10633 39942 10645 39994
rect 10697 39942 10709 39994
rect 10761 39942 10773 39994
rect 10825 39942 10837 39994
rect 10889 39942 10901 39994
rect 10953 39942 10965 39994
rect 11017 39942 11029 39994
rect 11081 39942 11093 39994
rect 11145 39942 11157 39994
rect 11209 39942 11221 39994
rect 11273 39942 11285 39994
rect 11337 39942 11343 39994
rect 3154 39926 11343 39942
rect 3154 39874 3160 39926
rect 3212 39874 3225 39926
rect 3277 39874 3290 39926
rect 3342 39874 3355 39926
rect 3407 39874 3420 39926
rect 3472 39874 3485 39926
rect 3537 39874 3550 39926
rect 3602 39874 3615 39926
rect 3667 39874 3680 39926
rect 3732 39874 3745 39926
rect 3797 39874 3810 39926
rect 3862 39874 3875 39926
rect 3927 39874 3940 39926
rect 3992 39874 4005 39926
rect 4057 39874 4070 39926
rect 4122 39874 4135 39926
rect 4187 39874 4200 39926
rect 4252 39874 4265 39926
rect 4317 39874 4330 39926
rect 4382 39874 4395 39926
rect 4447 39874 4460 39926
rect 4512 39874 4525 39926
rect 4577 39874 4590 39926
rect 4642 39874 4655 39926
rect 4707 39874 4720 39926
rect 4772 39874 4785 39926
rect 4837 39874 4850 39926
rect 4902 39874 4915 39926
rect 4967 39874 4980 39926
rect 5032 39874 5045 39926
rect 5097 39874 5110 39926
rect 5162 39874 5175 39926
rect 5227 39874 5240 39926
rect 5292 39874 5305 39926
rect 5357 39874 5370 39926
rect 5422 39874 5435 39926
rect 5487 39874 5500 39926
rect 5552 39874 5565 39926
rect 5617 39874 5630 39926
rect 5682 39874 5695 39926
rect 5747 39874 5760 39926
rect 5812 39874 5825 39926
rect 5877 39874 5890 39926
rect 5942 39874 5955 39926
rect 6007 39874 6020 39926
rect 6072 39874 6085 39926
rect 6137 39874 6150 39926
rect 6202 39874 6215 39926
rect 6267 39874 6280 39926
rect 6332 39874 6345 39926
rect 6397 39874 6410 39926
rect 6462 39874 6475 39926
rect 6527 39874 6540 39926
rect 6592 39874 6605 39926
rect 6657 39874 6670 39926
rect 6722 39874 6735 39926
rect 6787 39874 6800 39926
rect 6852 39874 6865 39926
rect 6917 39874 6930 39926
rect 6982 39874 6995 39926
rect 7047 39874 7060 39926
rect 7112 39874 7125 39926
rect 7177 39874 7189 39926
rect 7241 39874 7253 39926
rect 7305 39874 7317 39926
rect 7369 39874 7381 39926
rect 7433 39874 7445 39926
rect 7497 39874 7509 39926
rect 7561 39874 7573 39926
rect 7625 39874 7637 39926
rect 7689 39874 7701 39926
rect 7753 39874 7765 39926
rect 7817 39874 7829 39926
rect 7881 39874 7893 39926
rect 7945 39874 7957 39926
rect 8009 39874 8021 39926
rect 8073 39874 8085 39926
rect 8137 39874 8149 39926
rect 8201 39874 8213 39926
rect 8265 39874 8277 39926
rect 8329 39874 8341 39926
rect 8393 39874 8405 39926
rect 8457 39874 8469 39926
rect 8521 39874 8533 39926
rect 8585 39874 8597 39926
rect 8649 39874 8661 39926
rect 8713 39874 8725 39926
rect 8777 39874 8789 39926
rect 8841 39874 8853 39926
rect 8905 39874 8917 39926
rect 8969 39874 8981 39926
rect 9033 39874 9045 39926
rect 9097 39874 9109 39926
rect 9161 39874 9173 39926
rect 9225 39874 9237 39926
rect 9289 39874 9301 39926
rect 9353 39874 9365 39926
rect 9417 39874 9429 39926
rect 9481 39874 9493 39926
rect 9545 39874 9557 39926
rect 9609 39874 9621 39926
rect 9673 39874 9685 39926
rect 9737 39874 9749 39926
rect 9801 39874 9813 39926
rect 9865 39874 9877 39926
rect 9929 39874 9941 39926
rect 9993 39874 10005 39926
rect 10057 39874 10069 39926
rect 10121 39874 10133 39926
rect 10185 39874 10197 39926
rect 10249 39874 10261 39926
rect 10313 39874 10325 39926
rect 10377 39874 10389 39926
rect 10441 39874 10453 39926
rect 10505 39874 10517 39926
rect 10569 39874 10581 39926
rect 10633 39874 10645 39926
rect 10697 39874 10709 39926
rect 10761 39874 10773 39926
rect 10825 39874 10837 39926
rect 10889 39874 10901 39926
rect 10953 39874 10965 39926
rect 11017 39874 11029 39926
rect 11081 39874 11093 39926
rect 11145 39874 11157 39926
rect 11209 39874 11221 39926
rect 11273 39874 11285 39926
rect 11337 39874 11343 39926
rect 3154 39858 11343 39874
rect 3154 39806 3160 39858
rect 3212 39806 3225 39858
rect 3277 39806 3290 39858
rect 3342 39806 3355 39858
rect 3407 39806 3420 39858
rect 3472 39806 3485 39858
rect 3537 39806 3550 39858
rect 3602 39806 3615 39858
rect 3667 39806 3680 39858
rect 3732 39806 3745 39858
rect 3797 39806 3810 39858
rect 3862 39806 3875 39858
rect 3927 39806 3940 39858
rect 3992 39806 4005 39858
rect 4057 39806 4070 39858
rect 4122 39806 4135 39858
rect 4187 39806 4200 39858
rect 4252 39806 4265 39858
rect 4317 39806 4330 39858
rect 4382 39806 4395 39858
rect 4447 39806 4460 39858
rect 4512 39806 4525 39858
rect 4577 39806 4590 39858
rect 4642 39806 4655 39858
rect 4707 39806 4720 39858
rect 4772 39806 4785 39858
rect 4837 39806 4850 39858
rect 4902 39806 4915 39858
rect 4967 39806 4980 39858
rect 5032 39806 5045 39858
rect 5097 39806 5110 39858
rect 5162 39806 5175 39858
rect 5227 39806 5240 39858
rect 5292 39806 5305 39858
rect 5357 39806 5370 39858
rect 5422 39806 5435 39858
rect 5487 39806 5500 39858
rect 5552 39806 5565 39858
rect 5617 39806 5630 39858
rect 5682 39806 5695 39858
rect 5747 39806 5760 39858
rect 5812 39806 5825 39858
rect 5877 39806 5890 39858
rect 5942 39806 5955 39858
rect 6007 39806 6020 39858
rect 6072 39806 6085 39858
rect 6137 39806 6150 39858
rect 6202 39806 6215 39858
rect 6267 39806 6280 39858
rect 6332 39806 6345 39858
rect 6397 39806 6410 39858
rect 6462 39806 6475 39858
rect 6527 39806 6540 39858
rect 6592 39806 6605 39858
rect 6657 39806 6670 39858
rect 6722 39806 6735 39858
rect 6787 39806 6800 39858
rect 6852 39806 6865 39858
rect 6917 39806 6930 39858
rect 6982 39806 6995 39858
rect 7047 39806 7060 39858
rect 7112 39806 7125 39858
rect 7177 39806 7189 39858
rect 7241 39806 7253 39858
rect 7305 39806 7317 39858
rect 7369 39806 7381 39858
rect 7433 39806 7445 39858
rect 7497 39806 7509 39858
rect 7561 39806 7573 39858
rect 7625 39806 7637 39858
rect 7689 39806 7701 39858
rect 7753 39806 7765 39858
rect 7817 39806 7829 39858
rect 7881 39806 7893 39858
rect 7945 39806 7957 39858
rect 8009 39806 8021 39858
rect 8073 39806 8085 39858
rect 8137 39806 8149 39858
rect 8201 39806 8213 39858
rect 8265 39806 8277 39858
rect 8329 39806 8341 39858
rect 8393 39806 8405 39858
rect 8457 39806 8469 39858
rect 8521 39806 8533 39858
rect 8585 39806 8597 39858
rect 8649 39806 8661 39858
rect 8713 39806 8725 39858
rect 8777 39806 8789 39858
rect 8841 39806 8853 39858
rect 8905 39806 8917 39858
rect 8969 39806 8981 39858
rect 9033 39806 9045 39858
rect 9097 39806 9109 39858
rect 9161 39806 9173 39858
rect 9225 39806 9237 39858
rect 9289 39806 9301 39858
rect 9353 39806 9365 39858
rect 9417 39806 9429 39858
rect 9481 39806 9493 39858
rect 9545 39806 9557 39858
rect 9609 39806 9621 39858
rect 9673 39806 9685 39858
rect 9737 39806 9749 39858
rect 9801 39806 9813 39858
rect 9865 39806 9877 39858
rect 9929 39806 9941 39858
rect 9993 39806 10005 39858
rect 10057 39806 10069 39858
rect 10121 39806 10133 39858
rect 10185 39806 10197 39858
rect 10249 39806 10261 39858
rect 10313 39806 10325 39858
rect 10377 39806 10389 39858
rect 10441 39806 10453 39858
rect 10505 39806 10517 39858
rect 10569 39806 10581 39858
rect 10633 39806 10645 39858
rect 10697 39806 10709 39858
rect 10761 39806 10773 39858
rect 10825 39806 10837 39858
rect 10889 39806 10901 39858
rect 10953 39806 10965 39858
rect 11017 39806 11029 39858
rect 11081 39806 11093 39858
rect 11145 39806 11157 39858
rect 11209 39806 11221 39858
rect 11273 39806 11285 39858
rect 11337 39806 11343 39858
rect 3154 39790 11343 39806
rect 3154 39738 3160 39790
rect 3212 39738 3225 39790
rect 3277 39738 3290 39790
rect 3342 39738 3355 39790
rect 3407 39738 3420 39790
rect 3472 39738 3485 39790
rect 3537 39738 3550 39790
rect 3602 39738 3615 39790
rect 3667 39738 3680 39790
rect 3732 39738 3745 39790
rect 3797 39738 3810 39790
rect 3862 39738 3875 39790
rect 3927 39738 3940 39790
rect 3992 39738 4005 39790
rect 4057 39738 4070 39790
rect 4122 39738 4135 39790
rect 4187 39738 4200 39790
rect 4252 39738 4265 39790
rect 4317 39738 4330 39790
rect 4382 39738 4395 39790
rect 4447 39738 4460 39790
rect 4512 39738 4525 39790
rect 4577 39738 4590 39790
rect 4642 39738 4655 39790
rect 4707 39738 4720 39790
rect 4772 39738 4785 39790
rect 4837 39738 4850 39790
rect 4902 39738 4915 39790
rect 4967 39738 4980 39790
rect 5032 39738 5045 39790
rect 5097 39738 5110 39790
rect 5162 39738 5175 39790
rect 5227 39738 5240 39790
rect 5292 39738 5305 39790
rect 5357 39738 5370 39790
rect 5422 39738 5435 39790
rect 5487 39738 5500 39790
rect 5552 39738 5565 39790
rect 5617 39738 5630 39790
rect 5682 39738 5695 39790
rect 5747 39738 5760 39790
rect 5812 39738 5825 39790
rect 5877 39738 5890 39790
rect 5942 39738 5955 39790
rect 6007 39738 6020 39790
rect 6072 39738 6085 39790
rect 6137 39738 6150 39790
rect 6202 39738 6215 39790
rect 6267 39738 6280 39790
rect 6332 39738 6345 39790
rect 6397 39738 6410 39790
rect 6462 39738 6475 39790
rect 6527 39738 6540 39790
rect 6592 39738 6605 39790
rect 6657 39738 6670 39790
rect 6722 39738 6735 39790
rect 6787 39738 6800 39790
rect 6852 39738 6865 39790
rect 6917 39738 6930 39790
rect 6982 39738 6995 39790
rect 7047 39738 7060 39790
rect 7112 39738 7125 39790
rect 7177 39738 7189 39790
rect 7241 39738 7253 39790
rect 7305 39738 7317 39790
rect 7369 39738 7381 39790
rect 7433 39738 7445 39790
rect 7497 39738 7509 39790
rect 7561 39738 7573 39790
rect 7625 39738 7637 39790
rect 7689 39738 7701 39790
rect 7753 39738 7765 39790
rect 7817 39738 7829 39790
rect 7881 39738 7893 39790
rect 7945 39738 7957 39790
rect 8009 39738 8021 39790
rect 8073 39738 8085 39790
rect 8137 39738 8149 39790
rect 8201 39738 8213 39790
rect 8265 39738 8277 39790
rect 8329 39738 8341 39790
rect 8393 39738 8405 39790
rect 8457 39738 8469 39790
rect 8521 39738 8533 39790
rect 8585 39738 8597 39790
rect 8649 39738 8661 39790
rect 8713 39738 8725 39790
rect 8777 39738 8789 39790
rect 8841 39738 8853 39790
rect 8905 39738 8917 39790
rect 8969 39738 8981 39790
rect 9033 39738 9045 39790
rect 9097 39738 9109 39790
rect 9161 39738 9173 39790
rect 9225 39738 9237 39790
rect 9289 39738 9301 39790
rect 9353 39738 9365 39790
rect 9417 39738 9429 39790
rect 9481 39738 9493 39790
rect 9545 39738 9557 39790
rect 9609 39738 9621 39790
rect 9673 39738 9685 39790
rect 9737 39738 9749 39790
rect 9801 39738 9813 39790
rect 9865 39738 9877 39790
rect 9929 39738 9941 39790
rect 9993 39738 10005 39790
rect 10057 39738 10069 39790
rect 10121 39738 10133 39790
rect 10185 39738 10197 39790
rect 10249 39738 10261 39790
rect 10313 39738 10325 39790
rect 10377 39738 10389 39790
rect 10441 39738 10453 39790
rect 10505 39738 10517 39790
rect 10569 39738 10581 39790
rect 10633 39738 10645 39790
rect 10697 39738 10709 39790
rect 10761 39738 10773 39790
rect 10825 39738 10837 39790
rect 10889 39738 10901 39790
rect 10953 39738 10965 39790
rect 11017 39738 11029 39790
rect 11081 39738 11093 39790
rect 11145 39738 11157 39790
rect 11209 39738 11221 39790
rect 11273 39738 11285 39790
rect 11337 39738 11343 39790
rect 14399 39946 14405 39998
rect 14457 39946 14470 39998
rect 14522 39946 14535 39998
rect 14587 39946 14600 39998
rect 14652 39946 14665 39998
rect 14717 39946 14730 39998
rect 14782 39946 14795 39998
rect 14847 39946 14860 39998
rect 14912 39946 14925 39998
rect 14977 39946 14990 39998
rect 15042 39946 15055 39998
rect 15107 39946 15120 39998
rect 15172 39946 15185 39998
rect 15237 39946 15249 39998
rect 15301 39946 15313 39998
rect 15365 39946 15371 39998
rect 14399 39930 15371 39946
rect 14399 39878 14405 39930
rect 14457 39878 14470 39930
rect 14522 39878 14535 39930
rect 14587 39878 14600 39930
rect 14652 39878 14665 39930
rect 14717 39878 14730 39930
rect 14782 39878 14795 39930
rect 14847 39878 14860 39930
rect 14912 39878 14925 39930
rect 14977 39878 14990 39930
rect 15042 39878 15055 39930
rect 15107 39878 15120 39930
rect 15172 39878 15185 39930
rect 15237 39878 15249 39930
rect 15301 39878 15313 39930
rect 15365 39878 15371 39930
rect 14399 39862 15371 39878
rect 14399 39810 14405 39862
rect 14457 39810 14470 39862
rect 14522 39810 14535 39862
rect 14587 39810 14600 39862
rect 14652 39810 14665 39862
rect 14717 39810 14730 39862
rect 14782 39810 14795 39862
rect 14847 39810 14860 39862
rect 14912 39810 14925 39862
rect 14977 39810 14990 39862
rect 15042 39810 15055 39862
rect 15107 39810 15120 39862
rect 15172 39810 15185 39862
rect 15237 39810 15249 39862
rect 15301 39810 15313 39862
rect 15365 39810 15371 39862
rect 14399 39794 15371 39810
rect 14399 39742 14405 39794
rect 14457 39742 14470 39794
rect 14522 39742 14535 39794
rect 14587 39742 14600 39794
rect 14652 39742 14665 39794
rect 14717 39742 14730 39794
rect 14782 39742 14795 39794
rect 14847 39742 14860 39794
rect 14912 39742 14925 39794
rect 14977 39742 14990 39794
rect 15042 39742 15055 39794
rect 15107 39742 15120 39794
rect 15172 39742 15185 39794
rect 15237 39742 15249 39794
rect 15301 39742 15313 39794
rect 15365 39742 15371 39794
rect 14399 39740 15371 39742
rect 3154 39737 11343 39738
tri 8054 36568 8055 36569 sw
rect 2786 36079 3773 36080
rect 2786 36027 2792 36079
rect 2844 36027 2858 36079
rect 2910 36027 2924 36079
rect 2976 36027 2990 36079
rect 3042 36027 3056 36079
rect 3108 36027 3122 36079
rect 3174 36027 3188 36079
rect 3240 36027 3254 36079
rect 3306 36027 3320 36079
rect 3372 36027 3386 36079
rect 3438 36027 3452 36079
rect 3504 36027 3518 36079
rect 3570 36027 3584 36079
rect 3636 36027 3650 36079
rect 3702 36027 3715 36079
rect 3767 36027 3773 36079
rect 2786 36002 3773 36027
rect 2786 36001 15541 36002
rect 2786 35949 2792 36001
rect 2844 35949 2858 36001
rect 2910 35949 2924 36001
rect 2976 35949 2990 36001
rect 3042 35949 3056 36001
rect 3108 35949 3122 36001
rect 3174 35996 3188 36001
rect 3240 35996 3254 36001
rect 3306 35996 3320 36001
rect 3372 35996 3386 36001
rect 3438 35996 3452 36001
rect 3372 35962 3376 35996
rect 3438 35962 3449 35996
rect 3174 35949 3188 35962
rect 3240 35949 3254 35962
rect 3306 35949 3320 35962
rect 3372 35949 3386 35962
rect 3438 35949 3452 35962
rect 3504 35949 3518 36001
rect 3570 35949 3584 36001
rect 3636 35949 3650 36001
rect 3702 35949 3715 36001
rect 3767 35996 15541 36001
rect 3775 35962 3814 35996
rect 3848 35962 3887 35996
rect 3921 35962 3960 35996
rect 3994 35962 4033 35996
rect 4067 35962 4106 35996
rect 4140 35962 4179 35996
rect 4213 35962 4252 35996
rect 4286 35962 4325 35996
rect 4359 35962 4398 35996
rect 4432 35962 4471 35996
rect 4505 35962 4544 35996
rect 4578 35962 4617 35996
rect 4651 35962 4690 35996
rect 4724 35962 4763 35996
rect 4797 35962 4836 35996
rect 4870 35962 4909 35996
rect 4943 35962 4982 35996
rect 5016 35962 5055 35996
rect 3767 35949 5055 35962
rect 2786 35924 5055 35949
rect 2786 35923 3157 35924
rect 3191 35923 3230 35924
rect 3264 35923 3303 35924
rect 3337 35923 3376 35924
rect 3410 35923 3449 35924
rect 3483 35923 3522 35924
rect 3556 35923 3595 35924
rect 3629 35923 3668 35924
rect 3702 35923 3741 35924
rect 2786 35871 2792 35923
rect 2844 35871 2858 35923
rect 2910 35871 2924 35923
rect 2976 35871 2990 35923
rect 3042 35871 3056 35923
rect 3108 35871 3122 35923
rect 3372 35890 3376 35923
rect 3438 35890 3449 35923
rect 3174 35871 3188 35890
rect 3240 35871 3254 35890
rect 3306 35871 3320 35890
rect 3372 35871 3386 35890
rect 3438 35871 3452 35890
rect 3504 35871 3518 35923
rect 3570 35871 3584 35923
rect 3636 35871 3650 35923
rect 3702 35871 3715 35923
rect 3775 35890 3814 35924
rect 3848 35890 3887 35924
rect 3921 35890 3960 35924
rect 3994 35890 4033 35924
rect 4067 35890 4106 35924
rect 4140 35890 4179 35924
rect 4213 35890 4252 35924
rect 4286 35890 4325 35924
rect 4359 35890 4398 35924
rect 4432 35890 4471 35924
rect 4505 35890 4544 35924
rect 4578 35890 4617 35924
rect 4651 35890 4690 35924
rect 4724 35890 4763 35924
rect 4797 35890 4836 35924
rect 4870 35890 4909 35924
rect 4943 35890 4982 35924
rect 5016 35890 5055 35924
rect 15529 35890 15541 35996
rect 3767 35884 15541 35890
rect 3767 35871 3773 35884
rect 2786 35845 3773 35871
rect 2786 35793 2792 35845
rect 2844 35793 2858 35845
rect 2910 35793 2924 35845
rect 2976 35793 2990 35845
rect 3042 35793 3056 35845
rect 3108 35793 3122 35845
rect 3174 35793 3188 35845
rect 3240 35793 3254 35845
rect 3306 35793 3320 35845
rect 3372 35793 3386 35845
rect 3438 35793 3452 35845
rect 3504 35793 3518 35845
rect 3570 35793 3584 35845
rect 3636 35793 3650 35845
rect 3702 35793 3715 35845
rect 3767 35793 3773 35845
rect 2786 35792 3773 35793
rect 452 35674 972 35680
rect 452 35622 454 35674
rect 506 35648 528 35674
rect 580 35648 602 35674
rect 654 35648 972 35674
rect 1487 35655 1880 35701
rect 452 35610 463 35622
rect 452 35558 454 35610
rect 452 35546 463 35558
rect 452 35494 454 35546
rect 452 35482 463 35494
rect 452 35430 454 35482
rect 452 35418 463 35430
rect 452 35366 454 35418
rect 452 35354 463 35366
rect 452 35302 454 35354
rect 452 35290 463 35302
rect 452 35238 454 35290
rect 452 35226 463 35238
rect 452 35174 454 35226
rect 452 35162 463 35174
rect 452 35110 454 35162
rect 452 35098 463 35110
rect 452 35046 454 35098
rect 452 35034 463 35046
rect 452 34982 454 35034
rect 452 34970 463 34982
rect 452 34918 454 34970
rect 929 34927 972 35648
tri 972 34927 1194 35149 sw
rect 452 34906 463 34918
rect 452 34854 454 34906
rect 452 34842 463 34854
rect 452 34790 454 34842
rect 452 34778 463 34790
rect 452 34726 454 34778
rect 452 34714 463 34726
rect 452 34662 454 34714
rect 452 34650 463 34662
rect 452 34598 454 34650
rect 452 34586 463 34598
rect 452 34534 454 34586
rect 452 34522 463 34534
rect 452 34470 454 34522
rect 452 34458 463 34470
rect 452 34406 454 34458
rect 452 34394 463 34406
rect 452 34342 454 34394
rect 452 34330 463 34342
rect 452 34278 454 34330
rect 452 34266 463 34278
rect 452 34214 454 34266
rect 929 34246 1296 34927
rect 506 34214 528 34246
rect 580 34214 602 34246
rect 654 34214 1296 34246
rect 452 34207 1296 34214
rect 452 34202 463 34207
rect 497 34202 535 34207
rect 569 34202 607 34207
rect 641 34202 679 34207
rect 452 34150 454 34202
rect 506 34150 528 34202
rect 580 34150 602 34202
rect 654 34173 679 34202
rect 713 34173 751 34207
rect 785 34173 823 34207
rect 857 34173 895 34207
rect 929 34173 1296 34207
rect 654 34150 1296 34173
rect 452 34138 1296 34150
rect 452 34086 454 34138
rect 506 34086 528 34138
rect 580 34086 602 34138
rect 654 34134 1296 34138
rect 654 34100 679 34134
rect 713 34100 751 34134
rect 785 34100 823 34134
rect 857 34100 895 34134
rect 929 34100 1296 34134
rect 654 34086 1296 34100
rect 452 34074 1296 34086
rect 452 34022 454 34074
rect 506 34022 528 34074
rect 580 34022 602 34074
rect 654 34061 1296 34074
rect 654 34027 679 34061
rect 713 34027 751 34061
rect 785 34027 823 34061
rect 857 34027 895 34061
rect 929 34027 1296 34061
rect 654 34022 1296 34027
rect -23 34012 299 34018
rect -23 33986 149 34012
rect -23 33952 -17 33986
rect 17 33952 75 33986
rect 109 33960 149 33986
rect 201 33960 247 34012
rect 109 33952 167 33960
rect 201 33952 259 33960
rect 293 33952 299 33960
rect -23 33948 299 33952
rect -23 33914 149 33948
rect -23 33880 -17 33914
rect 17 33880 75 33914
rect 109 33896 149 33914
rect 201 33896 247 33948
rect 109 33884 167 33896
rect 201 33884 259 33896
rect 293 33884 299 33896
rect 109 33880 149 33884
rect -23 33842 149 33880
rect -23 33808 -17 33842
rect 17 33808 75 33842
rect 109 33832 149 33842
rect 201 33832 247 33884
rect 109 33820 167 33832
rect 201 33820 259 33832
rect 293 33820 299 33832
rect 109 33808 149 33820
rect -23 33769 149 33808
rect -23 33735 -17 33769
rect 17 33735 75 33769
rect 109 33768 149 33769
rect 201 33768 247 33820
rect 109 33756 167 33768
rect 201 33756 259 33768
rect 293 33756 299 33768
rect 109 33735 149 33756
rect -23 33704 149 33735
rect 201 33704 247 33756
rect -23 33696 299 33704
rect -23 33662 -17 33696
rect 17 33662 75 33696
rect 109 33692 167 33696
rect 201 33692 259 33696
rect 293 33692 299 33696
rect 109 33662 149 33692
rect -23 33640 149 33662
rect 201 33640 247 33692
rect -23 33628 299 33640
rect -23 33623 149 33628
rect -23 33589 -17 33623
rect 17 33589 75 33623
rect 109 33589 149 33623
rect -23 33576 149 33589
rect 201 33576 247 33628
rect -23 33564 299 33576
rect -23 33550 149 33564
rect -23 33516 -17 33550
rect 17 33516 75 33550
rect 109 33516 149 33550
rect -23 33512 149 33516
rect 201 33512 247 33564
rect -23 33500 299 33512
rect -23 33477 149 33500
rect -23 33443 -17 33477
rect 17 33443 75 33477
rect 109 33448 149 33477
rect 201 33448 247 33500
rect 109 33443 167 33448
rect 201 33443 259 33448
rect 293 33443 299 33448
rect -23 33436 299 33443
rect -23 33404 149 33436
rect -23 33370 -17 33404
rect 17 33370 75 33404
rect 109 33384 149 33404
rect 201 33384 247 33436
rect 109 33372 167 33384
rect 201 33372 259 33384
rect 293 33372 299 33384
rect 109 33370 149 33372
rect -23 33331 149 33370
rect -23 33297 -17 33331
rect 17 33297 75 33331
rect 109 33320 149 33331
rect 201 33320 247 33372
rect 109 33308 167 33320
rect 201 33308 259 33320
rect 293 33308 299 33320
rect 109 33297 149 33308
rect -23 33258 149 33297
rect -23 33224 -17 33258
rect 17 33224 75 33258
rect 109 33256 149 33258
rect 201 33256 247 33308
rect 109 33244 167 33256
rect 201 33244 259 33256
rect 293 33244 299 33256
rect 109 33224 149 33244
rect -23 33192 149 33224
rect 201 33192 247 33244
rect -23 33185 299 33192
rect -23 33151 -17 33185
rect 17 33151 75 33185
rect 109 33180 167 33185
rect 201 33180 259 33185
rect 293 33180 299 33185
rect 109 33151 149 33180
rect -23 33128 149 33151
rect 201 33128 247 33180
rect -23 33116 299 33128
rect -23 33112 149 33116
rect -23 33078 -17 33112
rect 17 33078 75 33112
rect 109 33078 149 33112
rect -23 33064 149 33078
rect 201 33064 247 33116
rect -23 33052 299 33064
rect -23 33039 149 33052
rect -23 33005 -17 33039
rect 17 33005 75 33039
rect 109 33005 149 33039
rect -23 33000 149 33005
rect 201 33000 247 33052
rect -23 32988 299 33000
rect -23 32966 149 32988
rect -23 32932 -17 32966
rect 17 32932 75 32966
rect 109 32936 149 32966
rect 201 32936 247 32988
rect 109 32932 167 32936
rect 201 32932 259 32936
rect 293 32932 299 32936
rect -23 32924 299 32932
rect -23 32893 149 32924
rect -23 32859 -17 32893
rect 17 32859 75 32893
rect 109 32872 149 32893
rect 201 32872 247 32924
rect 109 32859 167 32872
rect 201 32859 259 32872
rect 293 32859 299 32872
rect -23 32820 149 32859
rect -23 32786 -17 32820
rect 17 32786 75 32820
rect 109 32807 149 32820
rect 201 32807 247 32859
rect 109 32794 167 32807
rect 201 32794 259 32807
rect 293 32794 299 32807
rect 109 32786 149 32794
rect -23 32747 149 32786
rect -23 32713 -17 32747
rect 17 32713 75 32747
rect 109 32742 149 32747
rect 201 32742 247 32794
rect 109 32729 167 32742
rect 201 32729 259 32742
rect 293 32729 299 32742
rect 109 32713 149 32729
rect -23 32677 149 32713
rect 201 32677 247 32729
rect -23 32674 299 32677
rect -23 32640 -17 32674
rect 17 32640 75 32674
rect 109 32664 167 32674
rect 201 32664 259 32674
rect 293 32664 299 32674
rect 109 32640 149 32664
rect -23 32612 149 32640
rect 201 32612 247 32664
rect -23 32601 299 32612
rect -23 32567 -17 32601
rect 17 32567 75 32601
rect 109 32599 167 32601
rect 201 32599 259 32601
rect 293 32599 299 32601
rect 109 32567 149 32599
rect -23 32547 149 32567
rect 201 32547 247 32599
rect -23 32534 299 32547
rect -23 32528 149 32534
rect -23 32494 -17 32528
rect 17 32494 75 32528
rect 109 32494 149 32528
rect -23 32482 149 32494
rect 201 32482 247 32534
rect -23 32469 299 32482
rect -23 32455 149 32469
rect -23 32421 -17 32455
rect 17 32421 75 32455
rect 109 32421 149 32455
rect -23 32417 149 32421
rect 201 32417 247 32469
rect -23 32404 299 32417
rect -23 32382 149 32404
rect -23 32348 -17 32382
rect 17 32348 75 32382
rect 109 32352 149 32382
rect 201 32352 247 32404
rect 109 32348 167 32352
rect 201 32348 259 32352
rect 293 32348 299 32352
rect -23 32339 299 32348
rect -23 32309 149 32339
rect -23 32275 -17 32309
rect 17 32275 75 32309
rect 109 32287 149 32309
rect 201 32287 247 32339
rect 109 32275 167 32287
rect 201 32275 259 32287
rect 293 32275 299 32287
rect -23 32274 299 32275
rect -23 32236 149 32274
rect -23 32202 -17 32236
rect 17 32202 75 32236
rect 109 32222 149 32236
rect 201 32222 247 32274
rect 109 32209 167 32222
rect 201 32209 259 32222
rect 293 32209 299 32222
rect 109 32202 149 32209
rect -23 32163 149 32202
rect -23 32129 -17 32163
rect 17 32129 75 32163
rect 109 32157 149 32163
rect 201 32157 247 32209
rect 109 32144 167 32157
rect 201 32144 259 32157
rect 293 32144 299 32157
rect 109 32129 149 32144
rect -23 32092 149 32129
rect 201 32092 247 32144
rect -23 32090 299 32092
rect -23 32056 -17 32090
rect 17 32056 75 32090
rect 109 32079 167 32090
rect 201 32079 259 32090
rect 293 32079 299 32090
rect 109 32056 149 32079
rect -23 32027 149 32056
rect 201 32027 247 32079
rect -23 32017 299 32027
rect -23 31983 -17 32017
rect 17 31983 75 32017
rect 109 32014 167 32017
rect 201 32014 259 32017
rect 293 32014 299 32017
rect 109 31983 149 32014
rect -23 31962 149 31983
rect 201 31962 247 32014
rect -23 31949 299 31962
rect -23 31944 149 31949
rect -23 31910 -17 31944
rect 17 31910 75 31944
rect 109 31910 149 31944
rect -23 31897 149 31910
rect 201 31897 247 31949
rect -23 31884 299 31897
rect -23 31871 149 31884
rect -23 31837 -17 31871
rect 17 31837 75 31871
rect 109 31837 149 31871
rect -23 31832 149 31837
rect 201 31832 247 31884
rect -23 31819 299 31832
rect -23 31798 149 31819
rect -23 31764 -17 31798
rect 17 31764 75 31798
rect 109 31767 149 31798
rect 201 31767 247 31819
rect 109 31764 167 31767
rect 201 31764 259 31767
rect 293 31764 299 31767
rect -23 31754 299 31764
rect -23 31725 149 31754
rect -23 31691 -17 31725
rect 17 31691 75 31725
rect 109 31702 149 31725
rect 201 31702 247 31754
rect 109 31691 167 31702
rect 201 31691 259 31702
rect 293 31691 299 31702
rect -23 31689 299 31691
rect -23 31652 149 31689
rect -23 31618 -17 31652
rect 17 31618 75 31652
rect 109 31637 149 31652
rect 201 31637 247 31689
rect 109 31624 167 31637
rect 201 31624 259 31637
rect 293 31624 299 31637
rect 109 31618 149 31624
rect -23 31579 149 31618
rect -23 31545 -17 31579
rect 17 31545 75 31579
rect 109 31572 149 31579
rect 201 31572 247 31624
rect 109 31559 167 31572
rect 201 31559 259 31572
rect 293 31559 299 31572
rect 109 31545 149 31559
rect -23 31507 149 31545
rect 201 31507 247 31559
rect -23 31506 299 31507
rect -23 31472 -17 31506
rect 17 31472 75 31506
rect 109 31494 167 31506
rect 201 31494 259 31506
rect 293 31494 299 31506
rect 109 31472 149 31494
rect -23 31442 149 31472
rect 201 31442 247 31494
rect -23 31433 299 31442
rect -23 31399 -17 31433
rect 17 31399 75 31433
rect 109 31429 167 31433
rect 201 31429 259 31433
rect 293 31429 299 31433
rect 109 31399 149 31429
rect -23 31377 149 31399
rect 201 31377 247 31429
rect -23 31364 299 31377
rect -23 31360 149 31364
rect -23 31326 -17 31360
rect 17 31326 75 31360
rect 109 31326 149 31360
rect -23 31312 149 31326
rect 201 31312 247 31364
rect -23 31299 299 31312
rect -23 31287 149 31299
rect -23 31253 -17 31287
rect 17 31253 75 31287
rect 109 31253 149 31287
rect -23 31247 149 31253
rect 201 31247 247 31299
rect -23 31234 299 31247
rect -23 31214 149 31234
rect -23 31180 -17 31214
rect 17 31180 75 31214
rect 109 31182 149 31214
rect 201 31182 247 31234
rect 109 31180 167 31182
rect 201 31180 259 31182
rect 293 31180 299 31182
rect -23 31169 299 31180
rect -23 31141 149 31169
rect -23 31107 -17 31141
rect 17 31107 75 31141
rect 109 31117 149 31141
rect 201 31117 247 31169
rect 109 31107 167 31117
rect 201 31107 259 31117
rect 293 31107 299 31117
rect -23 31104 299 31107
rect -23 31068 149 31104
rect -23 31034 -17 31068
rect 17 31034 75 31068
rect 109 31052 149 31068
rect 201 31052 247 31104
rect 109 31039 167 31052
rect 201 31039 259 31052
rect 293 31039 299 31052
rect 109 31034 149 31039
rect -23 30995 149 31034
rect -23 30961 -17 30995
rect 17 30961 75 30995
rect 109 30987 149 30995
rect 201 30987 247 31039
rect 109 30974 167 30987
rect 201 30974 259 30987
rect 293 30974 299 30987
rect 109 30961 149 30974
rect -23 30922 149 30961
rect 201 30922 247 30974
rect -23 30888 -17 30922
rect 17 30888 75 30922
rect 109 30909 167 30922
rect 201 30909 259 30922
rect 293 30909 299 30922
rect 109 30888 149 30909
rect -23 30857 149 30888
rect 201 30857 247 30909
rect -23 30849 299 30857
rect -23 30815 -17 30849
rect 17 30815 75 30849
rect 109 30844 167 30849
rect 201 30844 259 30849
rect 293 30844 299 30849
rect 109 30815 149 30844
rect -23 30792 149 30815
rect 201 30792 247 30844
rect -23 30779 299 30792
rect -23 30776 149 30779
rect -23 30742 -17 30776
rect 17 30742 75 30776
rect 109 30742 149 30776
rect -23 30727 149 30742
rect 201 30727 247 30779
rect -23 30714 299 30727
rect -23 30703 149 30714
rect -23 30669 -17 30703
rect 17 30669 75 30703
rect 109 30669 149 30703
rect -23 30662 149 30669
rect 201 30662 247 30714
rect -23 30649 299 30662
rect -23 30630 149 30649
rect -23 30596 -17 30630
rect 17 30596 75 30630
rect 109 30597 149 30630
rect 201 30597 247 30649
rect 109 30596 167 30597
rect 201 30596 259 30597
rect 293 30596 299 30597
rect -23 30584 299 30596
rect -23 30557 149 30584
rect -23 30523 -17 30557
rect 17 30523 75 30557
rect 109 30532 149 30557
rect 201 30532 247 30584
rect 109 30523 167 30532
rect 201 30523 259 30532
rect 293 30523 299 30532
rect -23 30519 299 30523
rect -23 30484 149 30519
rect -23 30450 -17 30484
rect 17 30450 75 30484
rect 109 30467 149 30484
rect 201 30467 247 30519
rect 109 30454 167 30467
rect 201 30454 259 30467
rect 293 30454 299 30467
rect 109 30450 149 30454
rect -23 30411 149 30450
rect -23 30377 -17 30411
rect 17 30377 75 30411
rect 109 30402 149 30411
rect 201 30402 247 30454
rect 109 30389 167 30402
rect 201 30389 259 30402
rect 293 30389 299 30402
rect 109 30377 149 30389
rect -23 30338 149 30377
rect -23 30304 -17 30338
rect 17 30304 75 30338
rect 109 30337 149 30338
rect 201 30337 247 30389
rect 109 30324 167 30337
rect 201 30324 259 30337
rect 293 30324 299 30337
rect 109 30304 149 30324
rect -23 30272 149 30304
rect 201 30272 247 30324
rect -23 30265 299 30272
rect -23 30231 -17 30265
rect 17 30231 75 30265
rect 109 30259 167 30265
rect 201 30259 259 30265
rect 293 30259 299 30265
rect 109 30231 149 30259
rect -23 30207 149 30231
rect 201 30207 247 30259
rect -23 30194 299 30207
rect -23 30192 149 30194
rect -23 30158 -17 30192
rect 17 30158 75 30192
rect 109 30158 149 30192
rect -23 30142 149 30158
rect 201 30142 247 30194
rect -23 30129 299 30142
rect -23 30119 149 30129
rect -23 30085 -17 30119
rect 17 30085 75 30119
rect 109 30085 149 30119
rect -23 30077 149 30085
rect 201 30077 247 30129
rect -23 30064 299 30077
rect -23 30046 149 30064
rect -23 30012 -17 30046
rect 17 30012 75 30046
rect 109 30012 149 30046
rect 201 30012 247 30064
rect -23 29999 299 30012
rect -23 29973 149 29999
rect -23 29939 -17 29973
rect 17 29939 75 29973
rect 109 29947 149 29973
rect 201 29947 247 29999
rect 109 29939 167 29947
rect 201 29939 259 29947
rect 293 29939 299 29947
rect -23 29934 299 29939
rect -23 29900 149 29934
rect -23 29866 -17 29900
rect 17 29866 75 29900
rect 109 29882 149 29900
rect 201 29882 247 29934
rect 109 29869 167 29882
rect 201 29869 259 29882
rect 293 29869 299 29882
rect 109 29866 149 29869
rect -23 29827 149 29866
rect -23 29793 -17 29827
rect 17 29793 75 29827
rect 109 29817 149 29827
rect 201 29817 247 29869
rect 109 29804 167 29817
rect 201 29804 259 29817
rect 293 29804 299 29817
rect 109 29793 149 29804
rect -23 29754 149 29793
rect -23 29720 -17 29754
rect 17 29720 75 29754
rect 109 29752 149 29754
rect 201 29752 247 29804
rect 109 29739 167 29752
rect 201 29739 259 29752
rect 293 29739 299 29752
rect 109 29720 149 29739
rect -23 29687 149 29720
rect 201 29687 247 29739
rect -23 29681 299 29687
rect -23 29647 -17 29681
rect 17 29647 75 29681
rect 109 29674 167 29681
rect 201 29674 259 29681
rect 293 29674 299 29681
rect 109 29647 149 29674
rect -23 29622 149 29647
rect 201 29622 247 29674
rect -23 29609 299 29622
rect -23 29608 149 29609
rect -23 29574 -17 29608
rect 17 29574 75 29608
rect 109 29574 149 29608
rect -23 29557 149 29574
rect 201 29557 247 29609
rect -23 29544 299 29557
rect -23 29535 149 29544
rect -23 29501 -17 29535
rect 17 29501 75 29535
rect 109 29501 149 29535
rect -23 29492 149 29501
rect 201 29492 247 29544
rect -23 29479 299 29492
rect -23 29462 149 29479
rect -23 29428 -17 29462
rect 17 29428 75 29462
rect 109 29428 149 29462
rect -23 29427 149 29428
rect 201 29427 247 29479
rect -23 29414 299 29427
rect -23 29389 149 29414
rect -23 29355 -17 29389
rect 17 29355 75 29389
rect 109 29362 149 29389
rect 201 29362 247 29414
rect 109 29355 167 29362
rect 201 29355 259 29362
rect 293 29355 299 29362
rect -23 29349 299 29355
rect -23 29316 149 29349
rect -23 29282 -17 29316
rect 17 29282 75 29316
rect 109 29297 149 29316
rect 201 29297 247 29349
rect 109 29284 167 29297
rect 201 29284 259 29297
rect 293 29284 299 29297
rect 109 29282 149 29284
rect -23 29243 149 29282
rect -23 29209 -17 29243
rect 17 29209 75 29243
rect 109 29232 149 29243
rect 201 29232 247 29284
rect 109 29219 167 29232
rect 201 29219 259 29232
rect 293 29219 299 29232
rect 109 29209 149 29219
rect -23 29170 149 29209
rect -23 29136 -17 29170
rect 17 29136 75 29170
rect 109 29167 149 29170
rect 201 29167 247 29219
rect 109 29154 167 29167
rect 201 29154 259 29167
rect 293 29154 299 29167
rect 109 29136 149 29154
rect -23 29102 149 29136
rect 201 29102 247 29154
rect -23 29097 299 29102
rect -23 29063 -17 29097
rect 17 29063 75 29097
rect 109 29089 167 29097
rect 201 29089 259 29097
rect 293 29089 299 29097
rect 109 29063 149 29089
rect -23 29037 149 29063
rect 201 29037 247 29089
rect -23 28024 299 29037
rect 452 34010 1296 34022
rect 452 33958 454 34010
rect 506 33958 528 34010
rect 580 33958 602 34010
rect 654 33991 1296 34010
rect 13523 33991 16029 34018
rect 654 33988 972 33991
rect 654 33958 679 33988
rect 452 33954 463 33958
rect 497 33954 535 33958
rect 569 33954 607 33958
rect 641 33954 679 33958
rect 713 33954 751 33988
rect 785 33954 823 33988
rect 857 33954 895 33988
rect 929 33954 972 33988
rect 452 33946 972 33954
rect 452 33894 454 33946
rect 506 33894 528 33946
rect 580 33894 602 33946
rect 654 33915 972 33946
rect 654 33894 679 33915
rect 452 33882 463 33894
rect 497 33882 535 33894
rect 569 33882 607 33894
rect 641 33882 679 33894
rect 452 33830 454 33882
rect 506 33830 528 33882
rect 580 33830 602 33882
rect 654 33881 679 33882
rect 713 33881 751 33915
rect 785 33881 823 33915
rect 857 33881 895 33915
rect 929 33881 972 33915
rect 654 33842 972 33881
rect 654 33830 679 33842
rect 452 33818 463 33830
rect 497 33818 535 33830
rect 569 33818 607 33830
rect 641 33818 679 33830
rect 452 33766 454 33818
rect 506 33766 528 33818
rect 580 33766 602 33818
rect 654 33808 679 33818
rect 713 33808 751 33842
rect 785 33808 823 33842
rect 857 33808 895 33842
rect 929 33808 972 33842
rect 654 33769 972 33808
rect 654 33766 679 33769
rect 452 33754 463 33766
rect 497 33754 535 33766
rect 569 33754 607 33766
rect 641 33754 679 33766
rect 452 33702 454 33754
rect 506 33702 528 33754
rect 580 33702 602 33754
rect 654 33735 679 33754
rect 713 33735 751 33769
rect 785 33735 823 33769
rect 857 33735 895 33769
rect 929 33735 972 33769
rect 654 33702 972 33735
rect 452 33696 972 33702
rect 452 33690 463 33696
rect 497 33690 535 33696
rect 569 33690 607 33696
rect 641 33690 679 33696
rect 452 33638 454 33690
rect 506 33638 528 33690
rect 580 33638 602 33690
rect 654 33662 679 33690
rect 713 33662 751 33696
rect 785 33662 823 33696
rect 857 33662 895 33696
rect 929 33662 972 33696
rect 654 33638 972 33662
rect 452 33626 972 33638
rect 452 33574 454 33626
rect 506 33574 528 33626
rect 580 33574 602 33626
rect 654 33623 972 33626
rect 654 33589 679 33623
rect 713 33589 751 33623
rect 785 33589 823 33623
rect 857 33589 895 33623
rect 929 33589 972 33623
rect 654 33574 972 33589
rect 452 33562 972 33574
rect 452 33510 454 33562
rect 506 33510 528 33562
rect 580 33510 602 33562
rect 654 33550 972 33562
rect 654 33516 679 33550
rect 713 33516 751 33550
rect 785 33516 823 33550
rect 857 33516 895 33550
rect 929 33516 972 33550
rect 654 33510 972 33516
rect 452 33498 972 33510
rect 452 33446 454 33498
rect 506 33446 528 33498
rect 580 33446 602 33498
rect 654 33477 972 33498
rect 654 33446 679 33477
rect 452 33443 463 33446
rect 497 33443 535 33446
rect 569 33443 607 33446
rect 641 33443 679 33446
rect 713 33443 751 33477
rect 785 33443 823 33477
rect 857 33443 895 33477
rect 929 33443 972 33477
rect 452 33434 972 33443
rect 452 33382 454 33434
rect 506 33382 528 33434
rect 580 33382 602 33434
rect 654 33404 972 33434
rect 654 33382 679 33404
rect 452 33370 463 33382
rect 497 33370 535 33382
rect 569 33370 607 33382
rect 641 33370 679 33382
rect 713 33370 751 33404
rect 785 33370 823 33404
rect 857 33370 895 33404
rect 929 33370 972 33404
rect 452 33318 454 33370
rect 506 33318 528 33370
rect 580 33318 602 33370
rect 654 33331 972 33370
rect 654 33318 679 33331
rect 452 33306 463 33318
rect 497 33306 535 33318
rect 569 33306 607 33318
rect 641 33306 679 33318
rect 452 33254 454 33306
rect 506 33254 528 33306
rect 580 33254 602 33306
rect 654 33297 679 33306
rect 713 33297 751 33331
rect 785 33297 823 33331
rect 857 33297 895 33331
rect 929 33297 972 33331
rect 654 33258 972 33297
rect 654 33254 679 33258
rect 452 33242 463 33254
rect 497 33242 535 33254
rect 569 33242 607 33254
rect 641 33242 679 33254
rect 452 33190 454 33242
rect 506 33190 528 33242
rect 580 33190 602 33242
rect 654 33224 679 33242
rect 713 33224 751 33258
rect 785 33224 823 33258
rect 857 33224 895 33258
rect 929 33224 972 33258
rect 654 33190 972 33224
rect 452 33185 972 33190
rect 452 33178 463 33185
rect 497 33178 535 33185
rect 569 33178 607 33185
rect 641 33178 679 33185
rect 452 33126 454 33178
rect 506 33126 528 33178
rect 580 33126 602 33178
rect 654 33151 679 33178
rect 713 33151 751 33185
rect 785 33151 823 33185
rect 857 33151 895 33185
rect 929 33151 972 33185
rect 654 33126 972 33151
rect 452 33114 972 33126
rect 452 33062 454 33114
rect 506 33062 528 33114
rect 580 33062 602 33114
rect 654 33112 972 33114
rect 654 33078 679 33112
rect 713 33078 751 33112
rect 785 33078 823 33112
rect 857 33078 895 33112
rect 929 33078 972 33112
rect 654 33062 972 33078
rect 452 33050 972 33062
rect 452 32998 454 33050
rect 506 32998 528 33050
rect 580 32998 602 33050
rect 654 33039 972 33050
rect 654 33005 679 33039
rect 713 33005 751 33039
rect 785 33005 823 33039
rect 857 33005 895 33039
rect 929 33005 972 33039
rect 654 32998 972 33005
rect 452 32986 972 32998
rect 452 32934 454 32986
rect 506 32934 528 32986
rect 580 32934 602 32986
rect 654 32966 972 32986
rect 654 32934 679 32966
rect 452 32932 463 32934
rect 497 32932 535 32934
rect 569 32932 607 32934
rect 641 32932 679 32934
rect 713 32932 751 32966
rect 785 32932 823 32966
rect 857 32932 895 32966
rect 929 32932 972 32966
rect 452 32922 972 32932
rect 452 32870 454 32922
rect 506 32870 528 32922
rect 580 32870 602 32922
rect 654 32893 972 32922
rect 654 32870 679 32893
rect 452 32859 463 32870
rect 497 32859 535 32870
rect 569 32859 607 32870
rect 641 32859 679 32870
rect 713 32859 751 32893
rect 785 32859 823 32893
rect 857 32859 895 32893
rect 929 32859 972 32893
rect 452 32858 972 32859
rect 452 32806 454 32858
rect 506 32806 528 32858
rect 580 32806 602 32858
rect 654 32820 972 32858
rect 654 32806 679 32820
rect 452 32794 463 32806
rect 497 32794 535 32806
rect 569 32794 607 32806
rect 641 32794 679 32806
rect 452 32742 454 32794
rect 506 32742 528 32794
rect 580 32742 602 32794
rect 654 32786 679 32794
rect 713 32786 751 32820
rect 785 32786 823 32820
rect 857 32786 895 32820
rect 929 32786 972 32820
rect 654 32747 972 32786
rect 654 32742 679 32747
rect 452 32729 463 32742
rect 497 32729 535 32742
rect 569 32729 607 32742
rect 641 32729 679 32742
rect 452 32677 454 32729
rect 506 32677 528 32729
rect 580 32677 602 32729
rect 654 32713 679 32729
rect 713 32713 751 32747
rect 785 32713 823 32747
rect 857 32713 895 32747
rect 929 32713 972 32747
rect 654 32677 972 32713
rect 452 32674 972 32677
rect 452 32664 463 32674
rect 497 32664 535 32674
rect 569 32664 607 32674
rect 641 32664 679 32674
rect 452 32612 454 32664
rect 506 32612 528 32664
rect 580 32612 602 32664
rect 654 32640 679 32664
rect 713 32640 751 32674
rect 785 32640 823 32674
rect 857 32640 895 32674
rect 929 32640 972 32674
rect 654 32612 972 32640
rect 452 32601 972 32612
rect 452 32599 463 32601
rect 497 32599 535 32601
rect 569 32599 607 32601
rect 641 32599 679 32601
rect 452 32547 454 32599
rect 506 32547 528 32599
rect 580 32547 602 32599
rect 654 32567 679 32599
rect 713 32567 751 32601
rect 785 32567 823 32601
rect 857 32567 895 32601
rect 929 32567 972 32601
rect 654 32547 972 32567
rect 452 32534 972 32547
rect 452 32482 454 32534
rect 506 32482 528 32534
rect 580 32482 602 32534
rect 654 32528 972 32534
rect 654 32494 679 32528
rect 713 32494 751 32528
rect 785 32494 823 32528
rect 857 32494 895 32528
rect 929 32494 972 32528
rect 654 32482 972 32494
rect 452 32469 972 32482
rect 452 32417 454 32469
rect 506 32417 528 32469
rect 580 32417 602 32469
rect 654 32455 972 32469
rect 654 32421 679 32455
rect 713 32421 751 32455
rect 785 32421 823 32455
rect 857 32421 895 32455
rect 929 32421 972 32455
rect 654 32417 972 32421
rect 452 32404 972 32417
rect 452 32352 454 32404
rect 506 32352 528 32404
rect 580 32352 602 32404
rect 654 32382 972 32404
rect 654 32352 679 32382
rect 452 32348 463 32352
rect 497 32348 535 32352
rect 569 32348 607 32352
rect 641 32348 679 32352
rect 713 32348 751 32382
rect 785 32348 823 32382
rect 857 32348 895 32382
rect 929 32348 972 32382
rect 452 32339 972 32348
rect 452 32287 454 32339
rect 506 32287 528 32339
rect 580 32287 602 32339
rect 654 32309 972 32339
rect 654 32287 679 32309
rect 452 32275 463 32287
rect 497 32275 535 32287
rect 569 32275 607 32287
rect 641 32275 679 32287
rect 713 32275 751 32309
rect 785 32275 823 32309
rect 857 32275 895 32309
rect 929 32275 972 32309
rect 452 32274 972 32275
rect 452 32222 454 32274
rect 506 32222 528 32274
rect 580 32222 602 32274
rect 654 32236 972 32274
rect 654 32222 679 32236
rect 452 32209 463 32222
rect 497 32209 535 32222
rect 569 32209 607 32222
rect 641 32209 679 32222
rect 452 32157 454 32209
rect 506 32157 528 32209
rect 580 32157 602 32209
rect 654 32202 679 32209
rect 713 32202 751 32236
rect 785 32202 823 32236
rect 857 32202 895 32236
rect 929 32202 972 32236
rect 654 32163 972 32202
rect 654 32157 679 32163
rect 452 32144 463 32157
rect 497 32144 535 32157
rect 569 32144 607 32157
rect 641 32144 679 32157
rect 452 32092 454 32144
rect 506 32092 528 32144
rect 580 32092 602 32144
rect 654 32129 679 32144
rect 713 32129 751 32163
rect 785 32129 823 32163
rect 857 32129 895 32163
rect 929 32129 972 32163
rect 654 32092 972 32129
rect 452 32090 972 32092
rect 452 32079 463 32090
rect 497 32079 535 32090
rect 569 32079 607 32090
rect 641 32079 679 32090
rect 452 32027 454 32079
rect 506 32027 528 32079
rect 580 32027 602 32079
rect 654 32056 679 32079
rect 713 32056 751 32090
rect 785 32056 823 32090
rect 857 32056 895 32090
rect 929 32056 972 32090
rect 654 32027 972 32056
rect 452 32017 972 32027
rect 452 32014 463 32017
rect 497 32014 535 32017
rect 569 32014 607 32017
rect 641 32014 679 32017
rect 452 31962 454 32014
rect 506 31962 528 32014
rect 580 31962 602 32014
rect 654 31983 679 32014
rect 713 31983 751 32017
rect 785 31983 823 32017
rect 857 31983 895 32017
rect 929 31983 972 32017
rect 654 31962 972 31983
rect 452 31949 972 31962
rect 452 31897 454 31949
rect 506 31897 528 31949
rect 580 31897 602 31949
rect 654 31944 972 31949
rect 654 31910 679 31944
rect 713 31910 751 31944
rect 785 31910 823 31944
rect 857 31910 895 31944
rect 929 31910 972 31944
rect 654 31897 972 31910
rect 452 31884 972 31897
rect 452 31832 454 31884
rect 506 31832 528 31884
rect 580 31832 602 31884
rect 654 31871 972 31884
rect 654 31837 679 31871
rect 713 31837 751 31871
rect 785 31837 823 31871
rect 857 31837 895 31871
rect 929 31837 972 31871
rect 654 31832 972 31837
rect 452 31819 972 31832
rect 452 31767 454 31819
rect 506 31767 528 31819
rect 580 31767 602 31819
rect 654 31798 972 31819
rect 654 31767 679 31798
rect 452 31764 463 31767
rect 497 31764 535 31767
rect 569 31764 607 31767
rect 641 31764 679 31767
rect 713 31764 751 31798
rect 785 31764 823 31798
rect 857 31764 895 31798
rect 929 31764 972 31798
rect 452 31754 972 31764
rect 452 31702 454 31754
rect 506 31702 528 31754
rect 580 31702 602 31754
rect 654 31725 972 31754
rect 654 31702 679 31725
rect 452 31691 463 31702
rect 497 31691 535 31702
rect 569 31691 607 31702
rect 641 31691 679 31702
rect 713 31691 751 31725
rect 785 31691 823 31725
rect 857 31691 895 31725
rect 929 31691 972 31725
rect 452 31689 972 31691
rect 452 31637 454 31689
rect 506 31637 528 31689
rect 580 31637 602 31689
rect 654 31652 972 31689
rect 654 31637 679 31652
rect 452 31624 463 31637
rect 497 31624 535 31637
rect 569 31624 607 31637
rect 641 31624 679 31637
rect 452 31572 454 31624
rect 506 31572 528 31624
rect 580 31572 602 31624
rect 654 31618 679 31624
rect 713 31618 751 31652
rect 785 31618 823 31652
rect 857 31618 895 31652
rect 929 31618 972 31652
rect 654 31579 972 31618
rect 654 31572 679 31579
rect 452 31559 463 31572
rect 497 31559 535 31572
rect 569 31559 607 31572
rect 641 31559 679 31572
rect 452 31507 454 31559
rect 506 31507 528 31559
rect 580 31507 602 31559
rect 654 31545 679 31559
rect 713 31545 751 31579
rect 785 31545 823 31579
rect 857 31545 895 31579
rect 929 31545 972 31579
rect 654 31507 972 31545
rect 452 31506 972 31507
rect 452 31494 463 31506
rect 497 31494 535 31506
rect 569 31494 607 31506
rect 641 31494 679 31506
rect 452 31442 454 31494
rect 506 31442 528 31494
rect 580 31442 602 31494
rect 654 31472 679 31494
rect 713 31472 751 31506
rect 785 31472 823 31506
rect 857 31472 895 31506
rect 929 31472 972 31506
rect 654 31442 972 31472
rect 452 31433 972 31442
rect 452 31429 463 31433
rect 497 31429 535 31433
rect 569 31429 607 31433
rect 641 31429 679 31433
rect 452 31377 454 31429
rect 506 31377 528 31429
rect 580 31377 602 31429
rect 654 31399 679 31429
rect 713 31399 751 31433
rect 785 31399 823 31433
rect 857 31399 895 31433
rect 929 31399 972 31433
rect 654 31377 972 31399
rect 452 31364 972 31377
rect 452 31312 454 31364
rect 506 31312 528 31364
rect 580 31312 602 31364
rect 654 31360 972 31364
rect 654 31326 679 31360
rect 713 31326 751 31360
rect 785 31326 823 31360
rect 857 31326 895 31360
rect 929 31326 972 31360
rect 654 31312 972 31326
rect 452 31299 972 31312
rect 452 31247 454 31299
rect 506 31247 528 31299
rect 580 31247 602 31299
rect 654 31287 972 31299
rect 654 31253 679 31287
rect 713 31253 751 31287
rect 785 31253 823 31287
rect 857 31253 895 31287
rect 929 31253 972 31287
rect 654 31247 972 31253
rect 452 31234 972 31247
rect 452 31182 454 31234
rect 506 31182 528 31234
rect 580 31182 602 31234
rect 654 31214 972 31234
rect 654 31182 679 31214
rect 452 31180 463 31182
rect 497 31180 535 31182
rect 569 31180 607 31182
rect 641 31180 679 31182
rect 713 31180 751 31214
rect 785 31180 823 31214
rect 857 31180 895 31214
rect 929 31180 972 31214
rect 452 31169 972 31180
rect 452 31117 454 31169
rect 506 31117 528 31169
rect 580 31117 602 31169
rect 654 31141 972 31169
rect 654 31117 679 31141
rect 452 31107 463 31117
rect 497 31107 535 31117
rect 569 31107 607 31117
rect 641 31107 679 31117
rect 713 31107 751 31141
rect 785 31107 823 31141
rect 857 31107 895 31141
rect 929 31107 972 31141
rect 452 31104 972 31107
rect 452 31052 454 31104
rect 506 31052 528 31104
rect 580 31052 602 31104
rect 654 31068 972 31104
rect 654 31052 679 31068
rect 452 31039 463 31052
rect 497 31039 535 31052
rect 569 31039 607 31052
rect 641 31039 679 31052
rect 452 30987 454 31039
rect 506 30987 528 31039
rect 580 30987 602 31039
rect 654 31034 679 31039
rect 713 31034 751 31068
rect 785 31034 823 31068
rect 857 31034 895 31068
rect 929 31034 972 31068
rect 654 30995 972 31034
rect 654 30987 679 30995
rect 452 30974 463 30987
rect 497 30974 535 30987
rect 569 30974 607 30987
rect 641 30974 679 30987
rect 452 30922 454 30974
rect 506 30922 528 30974
rect 580 30922 602 30974
rect 654 30961 679 30974
rect 713 30961 751 30995
rect 785 30961 823 30995
rect 857 30961 895 30995
rect 929 30961 972 30995
rect 654 30922 972 30961
rect 452 30909 463 30922
rect 497 30909 535 30922
rect 569 30909 607 30922
rect 641 30909 679 30922
rect 452 30857 454 30909
rect 506 30857 528 30909
rect 580 30857 602 30909
rect 654 30888 679 30909
rect 713 30888 751 30922
rect 785 30888 823 30922
rect 857 30888 895 30922
rect 929 30888 972 30922
rect 654 30857 972 30888
rect 452 30849 972 30857
rect 452 30844 463 30849
rect 497 30844 535 30849
rect 569 30844 607 30849
rect 641 30844 679 30849
rect 452 30792 454 30844
rect 506 30792 528 30844
rect 580 30792 602 30844
rect 654 30815 679 30844
rect 713 30815 751 30849
rect 785 30815 823 30849
rect 857 30815 895 30849
rect 929 30815 972 30849
rect 654 30792 972 30815
rect 452 30779 972 30792
rect 452 30727 454 30779
rect 506 30727 528 30779
rect 580 30727 602 30779
rect 654 30776 972 30779
rect 654 30742 679 30776
rect 713 30742 751 30776
rect 785 30742 823 30776
rect 857 30742 895 30776
rect 929 30742 972 30776
rect 654 30727 972 30742
rect 452 30714 972 30727
rect 452 30662 454 30714
rect 506 30662 528 30714
rect 580 30662 602 30714
rect 654 30703 972 30714
rect 654 30669 679 30703
rect 713 30669 751 30703
rect 785 30669 823 30703
rect 857 30669 895 30703
rect 929 30669 972 30703
rect 654 30662 972 30669
rect 452 30649 972 30662
rect 452 30597 454 30649
rect 506 30597 528 30649
rect 580 30597 602 30649
rect 654 30630 972 30649
rect 654 30597 679 30630
rect 452 30596 463 30597
rect 497 30596 535 30597
rect 569 30596 607 30597
rect 641 30596 679 30597
rect 713 30596 751 30630
rect 785 30596 823 30630
rect 857 30596 895 30630
rect 929 30596 972 30630
rect 452 30584 972 30596
rect 452 30532 454 30584
rect 506 30532 528 30584
rect 580 30532 602 30584
rect 654 30557 972 30584
rect 654 30532 679 30557
rect 452 30523 463 30532
rect 497 30523 535 30532
rect 569 30523 607 30532
rect 641 30523 679 30532
rect 713 30523 751 30557
rect 785 30523 823 30557
rect 857 30523 895 30557
rect 929 30523 972 30557
rect 452 30519 972 30523
rect 452 30467 454 30519
rect 506 30467 528 30519
rect 580 30467 602 30519
rect 654 30484 972 30519
rect 654 30467 679 30484
rect 452 30454 463 30467
rect 497 30454 535 30467
rect 569 30454 607 30467
rect 641 30454 679 30467
rect 452 30402 454 30454
rect 506 30402 528 30454
rect 580 30402 602 30454
rect 654 30450 679 30454
rect 713 30450 751 30484
rect 785 30450 823 30484
rect 857 30450 895 30484
rect 929 30450 972 30484
rect 654 30411 972 30450
rect 654 30402 679 30411
rect 452 30389 463 30402
rect 497 30389 535 30402
rect 569 30389 607 30402
rect 641 30389 679 30402
rect 452 30337 454 30389
rect 506 30337 528 30389
rect 580 30337 602 30389
rect 654 30377 679 30389
rect 713 30377 751 30411
rect 785 30377 823 30411
rect 857 30377 895 30411
rect 929 30377 972 30411
rect 654 30338 972 30377
rect 654 30337 679 30338
rect 452 30324 463 30337
rect 497 30324 535 30337
rect 569 30324 607 30337
rect 641 30324 679 30337
rect 452 30272 454 30324
rect 506 30272 528 30324
rect 580 30272 602 30324
rect 654 30304 679 30324
rect 713 30304 751 30338
rect 785 30304 823 30338
rect 857 30304 895 30338
rect 929 30304 972 30338
rect 654 30272 972 30304
rect 452 30265 972 30272
rect 452 30259 463 30265
rect 497 30259 535 30265
rect 569 30259 607 30265
rect 641 30259 679 30265
rect 452 30207 454 30259
rect 506 30207 528 30259
rect 580 30207 602 30259
rect 654 30231 679 30259
rect 713 30231 751 30265
rect 785 30231 823 30265
rect 857 30231 895 30265
rect 929 30231 972 30265
rect 654 30207 972 30231
rect 452 30194 972 30207
rect 452 30142 454 30194
rect 506 30142 528 30194
rect 580 30142 602 30194
rect 654 30192 972 30194
rect 654 30158 679 30192
rect 713 30158 751 30192
rect 785 30158 823 30192
rect 857 30158 895 30192
rect 929 30158 972 30192
rect 654 30142 972 30158
rect 452 30129 972 30142
rect 452 30077 454 30129
rect 506 30077 528 30129
rect 580 30077 602 30129
rect 654 30119 972 30129
rect 654 30085 679 30119
rect 713 30085 751 30119
rect 785 30085 823 30119
rect 857 30085 895 30119
rect 929 30085 972 30119
rect 654 30077 972 30085
rect 452 30064 972 30077
rect 452 30012 454 30064
rect 506 30012 528 30064
rect 580 30012 602 30064
rect 654 30046 972 30064
rect 654 30012 679 30046
rect 713 30012 751 30046
rect 785 30012 823 30046
rect 857 30012 895 30046
rect 929 30012 972 30046
rect 452 29999 972 30012
rect 452 29947 454 29999
rect 506 29947 528 29999
rect 580 29947 602 29999
rect 654 29973 972 29999
rect 654 29947 679 29973
rect 452 29939 463 29947
rect 497 29939 535 29947
rect 569 29939 607 29947
rect 641 29939 679 29947
rect 713 29939 751 29973
rect 785 29939 823 29973
rect 857 29939 895 29973
rect 929 29939 972 29973
rect 452 29934 972 29939
rect 452 29882 454 29934
rect 506 29882 528 29934
rect 580 29882 602 29934
rect 654 29900 972 29934
rect 654 29882 679 29900
rect 452 29869 463 29882
rect 497 29869 535 29882
rect 569 29869 607 29882
rect 641 29869 679 29882
rect 452 29817 454 29869
rect 506 29817 528 29869
rect 580 29817 602 29869
rect 654 29866 679 29869
rect 713 29866 751 29900
rect 785 29866 823 29900
rect 857 29866 895 29900
rect 929 29866 972 29900
rect 654 29827 972 29866
rect 654 29817 679 29827
rect 452 29804 463 29817
rect 497 29804 535 29817
rect 569 29804 607 29817
rect 641 29804 679 29817
rect 452 29752 454 29804
rect 506 29752 528 29804
rect 580 29752 602 29804
rect 654 29793 679 29804
rect 713 29793 751 29827
rect 785 29793 823 29827
rect 857 29793 895 29827
rect 929 29793 972 29827
rect 654 29754 972 29793
rect 654 29752 679 29754
rect 452 29739 463 29752
rect 497 29739 535 29752
rect 569 29739 607 29752
rect 641 29739 679 29752
rect 452 29687 454 29739
rect 506 29687 528 29739
rect 580 29687 602 29739
rect 654 29720 679 29739
rect 713 29720 751 29754
rect 785 29720 823 29754
rect 857 29720 895 29754
rect 929 29720 972 29754
rect 654 29687 972 29720
rect 452 29681 972 29687
rect 452 29674 463 29681
rect 497 29674 535 29681
rect 569 29674 607 29681
rect 641 29674 679 29681
rect 452 29622 454 29674
rect 506 29622 528 29674
rect 580 29622 602 29674
rect 654 29647 679 29674
rect 713 29647 751 29681
rect 785 29647 823 29681
rect 857 29647 895 29681
rect 929 29647 972 29681
rect 654 29622 972 29647
rect 452 29609 972 29622
rect 452 29557 454 29609
rect 506 29557 528 29609
rect 580 29557 602 29609
rect 654 29608 972 29609
rect 654 29574 679 29608
rect 713 29574 751 29608
rect 785 29574 823 29608
rect 857 29574 895 29608
rect 929 29574 972 29608
rect 654 29557 972 29574
rect 452 29544 972 29557
rect 452 29492 454 29544
rect 506 29492 528 29544
rect 580 29492 602 29544
rect 654 29535 972 29544
rect 654 29501 679 29535
rect 713 29501 751 29535
rect 785 29501 823 29535
rect 857 29501 895 29535
rect 929 29501 972 29535
rect 654 29492 972 29501
rect 452 29479 972 29492
rect 452 29427 454 29479
rect 506 29427 528 29479
rect 580 29427 602 29479
rect 654 29462 972 29479
rect 654 29428 679 29462
rect 713 29428 751 29462
rect 785 29428 823 29462
rect 857 29428 895 29462
rect 929 29428 972 29462
rect 654 29427 972 29428
rect 452 29414 972 29427
rect 452 29362 454 29414
rect 506 29362 528 29414
rect 580 29362 602 29414
rect 654 29389 972 29414
rect 654 29362 679 29389
rect 452 29355 463 29362
rect 497 29355 535 29362
rect 569 29355 607 29362
rect 641 29355 679 29362
rect 713 29355 751 29389
rect 785 29355 823 29389
rect 857 29355 895 29389
rect 929 29355 972 29389
rect 452 29349 972 29355
rect 452 29297 454 29349
rect 506 29297 528 29349
rect 580 29297 602 29349
rect 654 29316 972 29349
rect 654 29297 679 29316
rect 452 29284 463 29297
rect 497 29284 535 29297
rect 569 29284 607 29297
rect 641 29284 679 29297
rect 452 29232 454 29284
rect 506 29232 528 29284
rect 580 29232 602 29284
rect 654 29282 679 29284
rect 713 29282 751 29316
rect 785 29282 823 29316
rect 857 29282 895 29316
rect 929 29282 972 29316
rect 654 29243 972 29282
rect 654 29232 679 29243
rect 452 29219 463 29232
rect 497 29219 535 29232
rect 569 29219 607 29232
rect 641 29219 679 29232
rect 452 29167 454 29219
rect 506 29167 528 29219
rect 580 29167 602 29219
rect 654 29209 679 29219
rect 713 29209 751 29243
rect 785 29209 823 29243
rect 857 29209 895 29243
rect 929 29209 972 29243
rect 654 29170 972 29209
rect 654 29167 679 29170
rect 452 29154 463 29167
rect 497 29154 535 29167
rect 569 29154 607 29167
rect 641 29154 679 29167
rect 452 29102 454 29154
rect 506 29102 528 29154
rect 580 29102 602 29154
rect 654 29136 679 29154
rect 713 29136 751 29170
rect 785 29136 823 29170
rect 857 29136 895 29170
rect 929 29136 972 29170
rect 654 29102 972 29136
rect 452 29097 972 29102
rect 452 29089 463 29097
rect 497 29089 535 29097
rect 569 29089 607 29097
rect 641 29089 679 29097
rect 452 29037 454 29089
rect 506 29037 528 29089
rect 580 29037 602 29089
rect 654 29063 679 29089
rect 713 29063 751 29097
rect 785 29063 823 29097
rect 857 29063 895 29097
rect 929 29063 972 29097
rect 654 29037 972 29063
rect 452 29031 972 29037
rect 2782 28561 3757 28562
rect 2782 28509 2788 28561
rect 2840 28509 2854 28561
rect 2906 28509 2919 28561
rect 2971 28509 2984 28561
rect 3036 28509 3049 28561
rect 3101 28509 3114 28561
rect 3166 28509 3179 28561
rect 3231 28509 3244 28561
rect 3296 28509 3309 28561
rect 3361 28509 3374 28561
rect 3426 28509 3439 28561
rect 3491 28509 3504 28561
rect 3556 28509 3569 28561
rect 3621 28509 3634 28561
rect 3686 28509 3699 28561
rect 3751 28509 3757 28561
rect 2782 28491 3757 28509
rect 2782 28439 2788 28491
rect 2840 28439 2854 28491
rect 2906 28439 2919 28491
rect 2971 28439 2984 28491
rect 3036 28439 3049 28491
rect 3101 28439 3114 28491
rect 3166 28439 3179 28491
rect 3231 28439 3244 28491
rect 3296 28439 3309 28491
rect 3361 28439 3374 28491
rect 3426 28439 3439 28491
rect 3491 28439 3504 28491
rect 3556 28439 3569 28491
rect 3621 28439 3634 28491
rect 3686 28439 3699 28491
rect 3751 28439 3757 28491
rect 2782 28421 3757 28439
rect 2782 28369 2788 28421
rect 2840 28369 2854 28421
rect 2906 28369 2919 28421
rect 2971 28369 2984 28421
rect 3036 28369 3049 28421
rect 3101 28369 3114 28421
rect 3166 28369 3179 28421
rect 3231 28369 3244 28421
rect 3296 28369 3309 28421
rect 3361 28369 3374 28421
rect 3426 28369 3439 28421
rect 3491 28369 3504 28421
rect 3556 28369 3569 28421
rect 3621 28369 3634 28421
rect 3686 28369 3699 28421
rect 3751 28369 3757 28421
rect 2782 28368 3757 28369
rect -23 27998 149 28024
rect -23 27964 -17 27998
rect 17 27964 75 27998
rect 109 27972 149 27998
rect 201 27972 247 28024
rect 109 27964 167 27972
rect 201 27964 259 27972
rect 293 27964 299 27972
rect -23 27958 299 27964
rect -23 27925 149 27958
rect -23 27891 -17 27925
rect 17 27891 75 27925
rect 109 27906 149 27925
rect 201 27906 247 27958
rect 109 27892 167 27906
rect 201 27892 259 27906
rect 293 27892 299 27906
rect 109 27891 149 27892
rect -23 27852 149 27891
rect -23 27818 -17 27852
rect 17 27818 75 27852
rect 109 27840 149 27852
rect 201 27840 247 27892
rect 109 27826 167 27840
rect 201 27826 259 27840
rect 293 27826 299 27840
rect 109 27818 149 27826
rect -23 27779 149 27818
rect -23 27745 -17 27779
rect 17 27745 75 27779
rect 109 27774 149 27779
rect 201 27774 247 27826
rect 109 27760 167 27774
rect 201 27760 259 27774
rect 293 27760 299 27774
rect 109 27745 149 27760
rect -23 27708 149 27745
rect 201 27708 247 27760
rect -23 27706 299 27708
rect -23 27672 -17 27706
rect 17 27672 75 27706
rect 109 27694 167 27706
rect 201 27694 259 27706
rect 293 27694 299 27706
rect 109 27672 149 27694
rect -23 27642 149 27672
rect 201 27642 247 27694
rect -23 27633 299 27642
rect -23 27599 -17 27633
rect 17 27599 75 27633
rect 109 27628 167 27633
rect 201 27628 259 27633
rect 293 27628 299 27633
rect 109 27599 149 27628
rect -23 27576 149 27599
rect 201 27576 247 27628
rect -23 27562 299 27576
rect -23 27560 149 27562
rect -23 27526 -17 27560
rect 17 27526 75 27560
rect 109 27526 149 27560
rect -23 27510 149 27526
rect 201 27510 247 27562
rect -23 27496 299 27510
rect -23 27487 149 27496
rect -23 27453 -17 27487
rect 17 27453 75 27487
rect 109 27453 149 27487
rect -23 27444 149 27453
rect 201 27444 247 27496
rect -23 27430 299 27444
rect -23 27414 149 27430
rect -23 27380 -17 27414
rect 17 27380 75 27414
rect 109 27380 149 27414
rect -23 27378 149 27380
rect 201 27378 247 27430
rect -23 27364 299 27378
rect -23 27341 149 27364
rect -23 27307 -17 27341
rect 17 27307 75 27341
rect 109 27312 149 27341
rect 201 27312 247 27364
rect 109 27307 167 27312
rect 201 27307 259 27312
rect 293 27307 299 27312
rect -23 27298 299 27307
rect -23 27268 149 27298
rect -23 27234 -17 27268
rect 17 27234 75 27268
rect 109 27246 149 27268
rect 201 27246 247 27298
rect 109 27234 167 27246
rect 201 27234 259 27246
rect 293 27234 299 27246
rect -23 27232 299 27234
rect -23 27195 149 27232
rect -23 27161 -17 27195
rect 17 27161 75 27195
rect 109 27180 149 27195
rect 201 27180 247 27232
rect 109 27166 167 27180
rect 201 27166 259 27180
rect 293 27166 299 27180
rect 109 27161 149 27166
rect -23 27122 149 27161
rect -23 27088 -17 27122
rect 17 27088 75 27122
rect 109 27114 149 27122
rect 201 27114 247 27166
rect 109 27100 167 27114
rect 201 27100 259 27114
rect 293 27100 299 27114
rect 109 27088 149 27100
rect -23 27049 149 27088
rect -23 27015 -17 27049
rect 17 27015 75 27049
rect 109 27048 149 27049
rect 201 27048 247 27100
rect 109 27034 167 27048
rect 201 27034 259 27048
rect 293 27034 299 27048
rect 109 27015 149 27034
rect -23 26982 149 27015
rect 201 26982 247 27034
rect -23 26976 299 26982
rect -23 26942 -17 26976
rect 17 26942 75 26976
rect 109 26968 167 26976
rect 201 26968 259 26976
rect 293 26968 299 26976
rect 109 26942 149 26968
rect -23 26916 149 26942
rect 201 26916 247 26968
rect -23 26903 299 26916
rect -23 26869 -17 26903
rect 17 26869 75 26903
rect 109 26902 167 26903
rect 201 26902 259 26903
rect 293 26902 299 26903
rect 109 26869 149 26902
rect -23 26850 149 26869
rect 201 26850 247 26902
rect -23 26836 299 26850
rect -23 26830 149 26836
rect -23 26796 -17 26830
rect 17 26796 75 26830
rect 109 26796 149 26830
rect -23 26784 149 26796
rect 201 26784 247 26836
rect -23 26770 299 26784
rect -23 26757 149 26770
rect -23 26723 -17 26757
rect 17 26723 75 26757
rect 109 26723 149 26757
rect -23 26718 149 26723
rect 201 26718 247 26770
rect -23 26704 299 26718
rect -23 26684 149 26704
rect -23 26650 -17 26684
rect 17 26650 75 26684
rect 109 26652 149 26684
rect 201 26652 247 26704
rect 109 26650 167 26652
rect 201 26650 259 26652
rect 293 26650 299 26652
rect -23 26638 299 26650
rect -23 26611 149 26638
rect -23 26577 -17 26611
rect 17 26577 75 26611
rect 109 26586 149 26611
rect 201 26586 247 26638
rect 109 26577 167 26586
rect 201 26577 259 26586
rect 293 26577 299 26586
rect -23 26573 299 26577
rect -23 26538 149 26573
rect -23 26504 -17 26538
rect 17 26504 75 26538
rect 109 26521 149 26538
rect 201 26521 247 26573
rect 109 26508 167 26521
rect 201 26508 259 26521
rect 293 26508 299 26521
rect 109 26504 149 26508
rect -23 26465 149 26504
rect -23 26431 -17 26465
rect 17 26431 75 26465
rect 109 26456 149 26465
rect 201 26456 247 26508
rect 109 26443 167 26456
rect 201 26443 259 26456
rect 293 26443 299 26456
rect 109 26431 149 26443
rect -23 26393 149 26431
rect -23 26359 -17 26393
rect 17 26359 75 26393
rect 109 26391 149 26393
rect 201 26391 247 26443
rect 109 26378 167 26391
rect 201 26378 259 26391
rect 293 26378 299 26391
rect 109 26359 149 26378
rect -23 26326 149 26359
rect 201 26326 247 26378
rect -23 26321 299 26326
rect -23 26287 -17 26321
rect 17 26287 75 26321
rect 109 26313 167 26321
rect 201 26313 259 26321
rect 293 26313 299 26321
rect 109 26287 149 26313
rect -23 26261 149 26287
rect 201 26261 247 26313
rect -23 26255 299 26261
rect 452 28024 971 28030
rect 452 27972 454 28024
rect 506 27972 528 28024
rect 580 27972 602 28024
rect 654 27978 971 28024
rect 654 27972 679 27978
rect 452 27958 463 27972
rect 497 27958 535 27972
rect 569 27958 607 27972
rect 641 27958 679 27972
rect 452 27906 454 27958
rect 506 27906 528 27958
rect 580 27906 602 27958
rect 654 27944 679 27958
rect 713 27944 751 27978
rect 785 27944 823 27978
rect 857 27944 895 27978
rect 929 27944 971 27978
rect 654 27906 971 27944
rect 452 27904 971 27906
rect 452 27903 1198 27904
rect 452 27892 463 27903
rect 497 27892 535 27903
rect 569 27892 607 27903
rect 641 27892 679 27903
rect 452 27840 454 27892
rect 506 27840 528 27892
rect 580 27840 602 27892
rect 654 27869 679 27892
rect 713 27869 751 27903
rect 785 27869 823 27903
rect 857 27869 895 27903
rect 929 27902 1198 27903
tri 1198 27902 1200 27904 nw
rect 929 27869 940 27902
rect 654 27840 940 27869
rect 452 27828 940 27840
rect 452 27826 463 27828
rect 497 27826 535 27828
rect 569 27826 607 27828
rect 641 27826 679 27828
rect 452 27774 454 27826
rect 506 27774 528 27826
rect 580 27774 602 27826
rect 654 27794 679 27826
rect 713 27794 751 27828
rect 785 27794 823 27828
rect 857 27794 895 27828
rect 929 27794 940 27828
rect 654 27774 940 27794
rect 452 27760 940 27774
rect 452 27708 454 27760
rect 506 27708 528 27760
rect 580 27708 602 27760
rect 654 27753 940 27760
rect 654 27719 679 27753
rect 713 27719 751 27753
rect 785 27719 823 27753
rect 857 27719 895 27753
rect 929 27719 940 27753
rect 654 27708 940 27719
rect 452 27694 940 27708
rect 452 27642 454 27694
rect 506 27642 528 27694
rect 580 27642 602 27694
rect 654 27678 940 27694
rect 654 27644 679 27678
rect 713 27644 751 27678
rect 785 27644 823 27678
rect 857 27644 895 27678
rect 929 27644 940 27678
tri 940 27644 1198 27902 nw
rect 654 27642 940 27644
rect 452 27628 940 27642
rect 452 27576 454 27628
rect 506 27576 528 27628
rect 580 27576 602 27628
rect 654 27603 940 27628
rect 654 27576 679 27603
rect 452 27569 463 27576
rect 497 27569 535 27576
rect 569 27569 607 27576
rect 641 27569 679 27576
rect 713 27569 751 27603
rect 785 27569 823 27603
rect 857 27569 895 27603
rect 929 27569 940 27603
rect 452 27562 940 27569
rect 452 27510 454 27562
rect 506 27510 528 27562
rect 580 27510 602 27562
rect 654 27528 940 27562
rect 654 27510 679 27528
rect 452 27496 463 27510
rect 497 27496 535 27510
rect 569 27496 607 27510
rect 641 27496 679 27510
rect 452 27444 454 27496
rect 506 27444 528 27496
rect 580 27444 602 27496
rect 654 27494 679 27496
rect 713 27494 751 27528
rect 785 27494 823 27528
rect 857 27494 895 27528
rect 929 27494 940 27528
rect 654 27453 940 27494
rect 654 27444 679 27453
rect 452 27430 463 27444
rect 497 27430 535 27444
rect 569 27430 607 27444
rect 641 27430 679 27444
rect 452 27378 454 27430
rect 506 27378 528 27430
rect 580 27378 602 27430
rect 654 27419 679 27430
rect 713 27419 751 27453
rect 785 27419 823 27453
rect 857 27419 895 27453
rect 929 27419 940 27453
rect 654 27378 940 27419
rect 452 27364 463 27378
rect 497 27364 535 27378
rect 569 27364 607 27378
rect 641 27364 679 27378
rect 452 27312 454 27364
rect 506 27312 528 27364
rect 580 27312 602 27364
rect 654 27344 679 27364
rect 713 27344 751 27378
rect 785 27344 823 27378
rect 857 27344 895 27378
rect 929 27344 940 27378
rect 654 27312 940 27344
rect 452 27303 940 27312
rect 452 27298 463 27303
rect 497 27298 535 27303
rect 569 27298 607 27303
rect 641 27298 679 27303
rect 452 27246 454 27298
rect 506 27246 528 27298
rect 580 27246 602 27298
rect 654 27269 679 27298
rect 713 27269 751 27303
rect 785 27269 823 27303
rect 857 27269 895 27303
rect 929 27269 940 27303
rect 654 27246 940 27269
rect 452 27232 940 27246
rect 452 27180 454 27232
rect 506 27180 528 27232
rect 580 27180 602 27232
rect 654 27228 940 27232
rect 654 27194 679 27228
rect 713 27194 751 27228
rect 785 27194 823 27228
rect 857 27194 895 27228
rect 929 27194 940 27228
rect 654 27180 940 27194
rect 452 27167 940 27180
rect 452 27115 454 27167
rect 506 27115 528 27167
rect 580 27115 602 27167
rect 654 27153 940 27167
rect 654 27119 679 27153
rect 713 27119 751 27153
rect 785 27119 823 27153
rect 857 27119 895 27153
rect 929 27119 940 27153
rect 654 27115 940 27119
rect 452 27102 940 27115
rect 452 27050 454 27102
rect 506 27050 528 27102
rect 580 27050 602 27102
rect 654 27079 940 27102
rect 14213 27483 14409 27489
rect 14265 27431 14285 27483
rect 14337 27431 14357 27483
rect 14213 27416 14409 27431
rect 14265 27364 14285 27416
rect 14337 27364 14357 27416
rect 14213 27349 14409 27364
rect 14265 27297 14285 27349
rect 14337 27297 14357 27349
rect 14213 27281 14409 27297
rect 14265 27229 14285 27281
rect 14337 27229 14357 27281
rect 14213 27213 14409 27229
rect 14265 27161 14285 27213
rect 14337 27161 14357 27213
rect 14213 27145 14409 27161
rect 14265 27093 14285 27145
rect 14337 27093 14357 27145
rect 14213 27087 14409 27093
rect 654 27050 679 27079
rect 452 27045 463 27050
rect 497 27045 535 27050
rect 569 27045 607 27050
rect 641 27045 679 27050
rect 713 27045 751 27079
rect 785 27045 823 27079
rect 857 27045 895 27079
rect 929 27045 940 27079
rect 452 27037 940 27045
rect 452 26985 454 27037
rect 506 26985 528 27037
rect 580 26985 602 27037
rect 654 27005 940 27037
rect 654 26985 679 27005
rect 452 26972 463 26985
rect 497 26972 535 26985
rect 569 26972 607 26985
rect 641 26972 679 26985
rect 452 26920 454 26972
rect 506 26920 528 26972
rect 580 26920 602 26972
rect 654 26971 679 26972
rect 713 26971 751 27005
rect 785 26971 823 27005
rect 857 26971 895 27005
rect 929 26971 940 27005
rect 654 26931 940 26971
rect 654 26920 679 26931
rect 452 26907 463 26920
rect 497 26907 535 26920
rect 569 26907 607 26920
rect 641 26907 679 26920
rect 452 26855 454 26907
rect 506 26855 528 26907
rect 580 26855 602 26907
rect 654 26897 679 26907
rect 713 26897 751 26931
rect 785 26897 823 26931
rect 857 26897 895 26931
rect 929 26897 940 26931
rect 654 26857 940 26897
rect 654 26855 679 26857
rect 452 26842 463 26855
rect 497 26842 535 26855
rect 569 26842 607 26855
rect 641 26842 679 26855
rect 452 26790 454 26842
rect 506 26790 528 26842
rect 580 26790 602 26842
rect 654 26823 679 26842
rect 713 26823 751 26857
rect 785 26823 823 26857
rect 857 26823 895 26857
rect 929 26823 940 26857
rect 654 26790 940 26823
rect 452 26783 940 26790
rect 452 26777 463 26783
rect 497 26777 535 26783
rect 569 26777 607 26783
rect 641 26777 679 26783
rect 452 26725 454 26777
rect 506 26725 528 26777
rect 580 26725 602 26777
rect 654 26749 679 26777
rect 713 26749 751 26783
rect 785 26749 823 26783
rect 857 26749 895 26783
rect 929 26749 940 26783
rect 654 26725 940 26749
rect 452 26712 940 26725
rect 452 26660 454 26712
rect 506 26660 528 26712
rect 580 26660 602 26712
rect 654 26709 940 26712
rect 654 26675 679 26709
rect 713 26675 751 26709
rect 785 26675 823 26709
rect 857 26675 895 26709
rect 929 26675 940 26709
rect 654 26660 940 26675
rect 452 26647 940 26660
rect 452 26595 454 26647
rect 506 26595 528 26647
rect 580 26595 602 26647
rect 654 26635 940 26647
rect 654 26601 679 26635
rect 713 26601 751 26635
rect 785 26601 823 26635
rect 857 26601 895 26635
rect 929 26601 940 26635
rect 654 26595 940 26601
rect 452 26582 940 26595
rect 452 26530 454 26582
rect 506 26530 528 26582
rect 580 26530 602 26582
rect 654 26561 940 26582
rect 654 26530 679 26561
rect 452 26527 463 26530
rect 497 26527 535 26530
rect 569 26527 607 26530
rect 641 26527 679 26530
rect 713 26527 751 26561
rect 785 26527 823 26561
rect 857 26527 895 26561
rect 929 26527 940 26561
rect 452 26517 940 26527
rect 452 26465 454 26517
rect 506 26465 528 26517
rect 580 26465 602 26517
rect 654 26487 940 26517
rect 654 26465 679 26487
rect 452 26453 463 26465
rect 497 26453 535 26465
rect 569 26453 607 26465
rect 641 26453 679 26465
rect 713 26453 751 26487
rect 785 26453 823 26487
rect 857 26453 895 26487
rect 929 26453 940 26487
rect 452 26452 940 26453
rect 452 26400 454 26452
rect 506 26400 528 26452
rect 580 26400 602 26452
rect 654 26413 940 26452
rect 654 26400 679 26413
rect 452 26387 463 26400
rect 497 26387 535 26400
rect 569 26387 607 26400
rect 641 26387 679 26400
rect 452 26335 454 26387
rect 506 26335 528 26387
rect 580 26335 602 26387
rect 654 26379 679 26387
rect 713 26379 751 26413
rect 785 26379 823 26413
rect 857 26379 895 26413
rect 929 26379 940 26413
rect 654 26339 940 26379
rect 654 26335 679 26339
rect 452 26322 463 26335
rect 497 26322 535 26335
rect 569 26322 607 26335
rect 641 26322 679 26335
rect 452 26270 454 26322
rect 506 26270 528 26322
rect 580 26270 602 26322
rect 654 26305 679 26322
rect 713 26305 751 26339
rect 785 26305 823 26339
rect 857 26305 895 26339
rect 929 26305 940 26339
rect 654 26270 940 26305
rect 452 26265 940 26270
rect 452 26257 463 26265
rect 497 26257 535 26265
rect 569 26257 607 26265
rect 641 26257 679 26265
rect 452 26205 454 26257
rect 506 26205 528 26257
rect 580 26205 602 26257
rect 654 26231 679 26257
rect 713 26231 751 26265
rect 785 26231 823 26265
rect 857 26231 895 26265
rect 929 26231 940 26265
rect 654 26205 940 26231
rect 452 26199 940 26205
tri 14158 26199 14596 26637 sw
rect 14158 26044 14596 26199
tri 14596 26044 14751 26199 sw
rect -23 26038 299 26044
rect -23 26012 149 26038
rect -23 25978 -17 26012
rect 17 25978 75 26012
rect 109 25986 149 26012
rect 201 25986 247 26038
rect 109 25978 167 25986
rect 201 25978 259 25986
rect 293 25978 299 25986
rect -23 25974 299 25978
rect -23 25940 149 25974
rect -23 25906 -17 25940
rect 17 25906 75 25940
rect 109 25922 149 25940
rect 201 25922 247 25974
rect 109 25910 167 25922
rect 201 25910 259 25922
rect 293 25910 299 25922
rect 109 25906 149 25910
rect -23 25868 149 25906
rect -23 25834 -17 25868
rect 17 25834 75 25868
rect 109 25858 149 25868
rect 201 25858 247 25910
rect 109 25846 167 25858
rect 201 25846 259 25858
rect 293 25846 299 25858
rect 109 25834 149 25846
rect -23 25796 149 25834
rect -23 25762 -17 25796
rect 17 25762 75 25796
rect 109 25794 149 25796
rect 201 25794 247 25846
rect 109 25782 167 25794
rect 201 25782 259 25794
rect 293 25782 299 25794
rect 109 25762 149 25782
rect -23 25730 149 25762
rect 201 25730 247 25782
rect -23 25724 299 25730
rect -23 25690 -17 25724
rect 17 25690 75 25724
rect 109 25718 167 25724
rect 201 25718 259 25724
rect 293 25718 299 25724
rect 109 25690 149 25718
rect -23 25666 149 25690
rect 201 25666 247 25718
rect -23 25654 299 25666
rect -23 25652 149 25654
rect -23 25618 -17 25652
rect 17 25618 75 25652
rect 109 25618 149 25652
rect -23 25602 149 25618
rect 201 25602 247 25654
rect -23 25590 299 25602
rect -23 25580 149 25590
rect -23 25546 -17 25580
rect 17 25546 75 25580
rect 109 25546 149 25580
rect -23 25538 149 25546
rect 201 25538 247 25590
rect -23 25526 299 25538
rect -23 25508 149 25526
rect -23 25474 -17 25508
rect 17 25474 75 25508
rect 109 25474 149 25508
rect 201 25474 247 25526
rect -23 25462 299 25474
rect -23 25436 149 25462
rect -23 25402 -17 25436
rect 17 25402 75 25436
rect 109 25410 149 25436
rect 201 25410 247 25462
rect 109 25402 167 25410
rect 201 25402 259 25410
rect 293 25402 299 25410
rect -23 25398 299 25402
rect -23 25364 149 25398
rect -23 25330 -17 25364
rect 17 25330 75 25364
rect 109 25346 149 25364
rect 201 25346 247 25398
rect 109 25334 167 25346
rect 201 25334 259 25346
rect 293 25334 299 25346
rect 109 25330 149 25334
rect -23 25292 149 25330
rect -23 25258 -17 25292
rect 17 25258 75 25292
rect 109 25282 149 25292
rect 201 25282 247 25334
rect 109 25270 167 25282
rect 201 25270 259 25282
rect 293 25270 299 25282
rect 109 25258 149 25270
rect -23 25220 149 25258
rect -23 25186 -17 25220
rect 17 25186 75 25220
rect 109 25218 149 25220
rect 201 25218 247 25270
rect 109 25206 167 25218
rect 201 25206 259 25218
rect 293 25206 299 25218
rect 109 25186 149 25206
rect -23 25154 149 25186
rect 201 25154 247 25206
rect -23 25148 299 25154
rect -23 25114 -17 25148
rect 17 25114 75 25148
rect 109 25142 167 25148
rect 201 25142 259 25148
rect 293 25142 299 25148
rect 109 25114 149 25142
rect -23 25090 149 25114
rect 201 25090 247 25142
rect -23 25078 299 25090
rect -23 25076 149 25078
rect -23 25042 -17 25076
rect 17 25042 75 25076
rect 109 25042 149 25076
rect -23 25026 149 25042
rect 201 25026 247 25078
rect -23 25014 299 25026
rect -23 25004 149 25014
rect -23 24970 -17 25004
rect 17 24970 75 25004
rect 109 24970 149 25004
rect -23 24962 149 24970
rect 201 24962 247 25014
rect -23 24950 299 24962
rect -23 24932 149 24950
rect -23 24898 -17 24932
rect 17 24898 75 24932
rect 109 24898 149 24932
rect 201 24898 247 24950
rect -23 24886 299 24898
rect -23 24860 149 24886
rect -23 24826 -17 24860
rect 17 24826 75 24860
rect 109 24834 149 24860
rect 201 24834 247 24886
rect 109 24826 167 24834
rect 201 24826 259 24834
rect 293 24826 299 24834
rect -23 24822 299 24826
rect -23 24788 149 24822
rect -23 24754 -17 24788
rect 17 24754 75 24788
rect 109 24770 149 24788
rect 201 24770 247 24822
rect 109 24758 167 24770
rect 201 24758 259 24770
rect 293 24758 299 24770
rect 109 24754 149 24758
rect -23 24716 149 24754
rect -23 24682 -17 24716
rect 17 24682 75 24716
rect 109 24706 149 24716
rect 201 24706 247 24758
rect 109 24694 167 24706
rect 201 24694 259 24706
rect 293 24694 299 24706
rect 109 24682 149 24694
rect -23 24644 149 24682
rect -23 24610 -17 24644
rect 17 24610 75 24644
rect 109 24642 149 24644
rect 201 24642 247 24694
rect 109 24630 167 24642
rect 201 24630 259 24642
rect 293 24630 299 24642
rect 109 24610 149 24630
rect -23 24578 149 24610
rect 201 24578 247 24630
rect -23 24572 299 24578
rect -23 24538 -17 24572
rect 17 24538 75 24572
rect 109 24566 167 24572
rect 201 24566 259 24572
rect 293 24566 299 24572
rect 109 24538 149 24566
rect -23 24514 149 24538
rect 201 24514 247 24566
rect -23 24502 299 24514
rect -23 24500 149 24502
rect -23 24466 -17 24500
rect 17 24466 75 24500
rect 109 24466 149 24500
rect -23 24450 149 24466
rect 201 24450 247 24502
rect -23 24438 299 24450
rect -23 24428 149 24438
rect -23 24394 -17 24428
rect 17 24394 75 24428
rect 109 24394 149 24428
rect -23 24386 149 24394
rect 201 24386 247 24438
rect -23 24374 299 24386
rect -23 24355 149 24374
rect -23 24321 -17 24355
rect 17 24321 75 24355
rect 109 24322 149 24355
rect 201 24322 247 24374
rect 109 24321 167 24322
rect 201 24321 259 24322
rect 293 24321 299 24322
rect -23 24310 299 24321
rect -23 24282 149 24310
rect -23 24248 -17 24282
rect 17 24248 75 24282
rect 109 24258 149 24282
rect 201 24258 247 24310
rect 109 24248 167 24258
rect 201 24248 259 24258
rect 293 24248 299 24258
rect -23 24246 299 24248
rect -23 24209 149 24246
rect -23 24175 -17 24209
rect 17 24175 75 24209
rect 109 24194 149 24209
rect 201 24194 247 24246
rect 109 24182 167 24194
rect 201 24182 259 24194
rect 293 24182 299 24194
rect 109 24175 149 24182
rect -23 24136 149 24175
rect -23 24102 -17 24136
rect 17 24102 75 24136
rect 109 24130 149 24136
rect 201 24130 247 24182
rect 109 24118 167 24130
rect 201 24118 259 24130
rect 293 24118 299 24130
rect 109 24102 149 24118
rect -23 24066 149 24102
rect 201 24066 247 24118
rect -23 24063 299 24066
rect -23 24029 -17 24063
rect 17 24029 75 24063
rect 109 24054 167 24063
rect 201 24054 259 24063
rect 293 24054 299 24063
rect 109 24029 149 24054
rect -23 24002 149 24029
rect 201 24002 247 24054
rect -23 23990 299 24002
rect -23 23956 -17 23990
rect 17 23956 75 23990
rect 109 23956 149 23990
rect -23 23938 149 23956
rect 201 23938 247 23990
rect -23 23926 299 23938
rect -23 23917 149 23926
rect -23 23883 -17 23917
rect 17 23883 75 23917
rect 109 23883 149 23917
rect -23 23874 149 23883
rect 201 23874 247 23926
rect -23 23862 299 23874
rect -23 23844 149 23862
rect -23 23810 -17 23844
rect 17 23810 75 23844
rect 109 23810 149 23844
rect 201 23810 247 23862
rect -23 23798 299 23810
rect -23 23771 149 23798
rect -23 23737 -17 23771
rect 17 23737 75 23771
rect 109 23746 149 23771
rect 201 23746 247 23798
rect 109 23737 167 23746
rect 201 23737 259 23746
rect 293 23737 299 23746
rect -23 23734 299 23737
rect -23 23698 149 23734
rect -23 23664 -17 23698
rect 17 23664 75 23698
rect 109 23682 149 23698
rect 201 23682 247 23734
rect 109 23670 167 23682
rect 201 23670 259 23682
rect 293 23670 299 23682
rect 109 23664 149 23670
rect -23 23625 149 23664
rect -23 23591 -17 23625
rect 17 23591 75 23625
rect 109 23618 149 23625
rect 201 23618 247 23670
rect 109 23606 167 23618
rect 201 23606 259 23618
rect 293 23606 299 23618
rect 109 23591 149 23606
rect -23 23554 149 23591
rect 201 23554 247 23606
rect -23 23552 299 23554
rect -23 23518 -17 23552
rect 17 23518 75 23552
rect 109 23542 167 23552
rect 201 23542 259 23552
rect 293 23542 299 23552
rect 109 23518 149 23542
rect -23 23490 149 23518
rect 201 23490 247 23542
rect -23 23479 299 23490
rect -23 23445 -17 23479
rect 17 23445 75 23479
rect 109 23478 167 23479
rect 201 23478 259 23479
rect 293 23478 299 23479
rect 109 23445 149 23478
rect -23 23426 149 23445
rect 201 23426 247 23478
rect -23 23414 299 23426
rect -23 23406 149 23414
rect -23 23372 -17 23406
rect 17 23372 75 23406
rect 109 23372 149 23406
rect -23 23362 149 23372
rect 201 23362 247 23414
rect -23 23350 299 23362
rect -23 23333 149 23350
rect -23 23299 -17 23333
rect 17 23299 75 23333
rect 109 23299 149 23333
rect -23 23298 149 23299
rect 201 23298 247 23350
rect -23 23286 299 23298
rect -23 23260 149 23286
rect -23 23226 -17 23260
rect 17 23226 75 23260
rect 109 23234 149 23260
rect 201 23234 247 23286
rect 109 23226 167 23234
rect 201 23226 259 23234
rect 293 23226 299 23234
rect -23 23222 299 23226
rect -23 23187 149 23222
rect -23 23153 -17 23187
rect 17 23153 75 23187
rect 109 23170 149 23187
rect 201 23170 247 23222
rect 109 23158 167 23170
rect 201 23158 259 23170
rect 293 23158 299 23170
rect 109 23153 149 23158
rect -23 23114 149 23153
rect -23 23080 -17 23114
rect 17 23080 75 23114
rect 109 23106 149 23114
rect 201 23106 247 23158
rect 109 23094 167 23106
rect 201 23094 259 23106
rect 293 23094 299 23106
rect 109 23080 149 23094
rect -23 23042 149 23080
rect 201 23042 247 23094
rect -23 23041 299 23042
rect -23 23007 -17 23041
rect 17 23007 75 23041
rect 109 23030 167 23041
rect 201 23030 259 23041
rect 293 23030 299 23041
rect 109 23007 149 23030
rect -23 22978 149 23007
rect 201 22978 247 23030
rect -23 22968 299 22978
rect -23 22934 -17 22968
rect 17 22934 75 22968
rect 109 22966 167 22968
rect 201 22966 259 22968
rect 293 22966 299 22968
rect 109 22934 149 22966
rect -23 22914 149 22934
rect 201 22914 247 22966
rect -23 22902 299 22914
rect -23 22895 149 22902
rect -23 22861 -17 22895
rect 17 22861 75 22895
rect 109 22861 149 22895
rect -23 22850 149 22861
rect 201 22850 247 22902
rect -23 22838 299 22850
rect -23 22822 149 22838
rect -23 22788 -17 22822
rect 17 22788 75 22822
rect 109 22788 149 22822
rect -23 22786 149 22788
rect 201 22786 247 22838
rect -23 22774 299 22786
rect -23 22749 149 22774
rect -23 22715 -17 22749
rect 17 22715 75 22749
rect 109 22722 149 22749
rect 201 22722 247 22774
rect 109 22715 167 22722
rect 201 22715 259 22722
rect 293 22715 299 22722
rect -23 22710 299 22715
rect -23 22676 149 22710
rect -23 22642 -17 22676
rect 17 22642 75 22676
rect 109 22658 149 22676
rect 201 22658 247 22710
rect 109 22646 167 22658
rect 201 22646 259 22658
rect 293 22646 299 22658
rect 109 22642 149 22646
rect -23 22603 149 22642
rect -23 22569 -17 22603
rect 17 22569 75 22603
rect 109 22594 149 22603
rect 201 22594 247 22646
rect 109 22582 167 22594
rect 201 22582 259 22594
rect 293 22582 299 22594
rect 109 22569 149 22582
rect -23 22530 149 22569
rect 201 22530 247 22582
rect -23 22496 -17 22530
rect 17 22496 75 22530
rect 109 22518 167 22530
rect 201 22518 259 22530
rect 293 22518 299 22530
rect 109 22496 149 22518
rect -23 22466 149 22496
rect 201 22466 247 22518
rect -23 22457 299 22466
rect -23 22423 -17 22457
rect 17 22423 75 22457
rect 109 22454 167 22457
rect 201 22454 259 22457
rect 293 22454 299 22457
rect 109 22423 149 22454
rect -23 22402 149 22423
rect 201 22402 247 22454
rect -23 22390 299 22402
rect -23 22384 149 22390
rect -23 22350 -17 22384
rect 17 22350 75 22384
rect 109 22350 149 22384
rect -23 22338 149 22350
rect 201 22338 247 22390
rect -23 22326 299 22338
rect -23 22311 149 22326
rect -23 22277 -17 22311
rect 17 22277 75 22311
rect 109 22277 149 22311
rect -23 22274 149 22277
rect 201 22274 247 22326
rect -23 22262 299 22274
rect -23 22238 149 22262
rect -23 22204 -17 22238
rect 17 22204 75 22238
rect 109 22210 149 22238
rect 201 22210 247 22262
rect 109 22204 167 22210
rect 201 22204 259 22210
rect 293 22204 299 22210
rect -23 22198 299 22204
rect -23 22165 149 22198
rect -23 22131 -17 22165
rect 17 22131 75 22165
rect 109 22146 149 22165
rect 201 22146 247 22198
rect 109 22134 167 22146
rect 201 22134 259 22146
rect 293 22134 299 22146
rect 109 22131 149 22134
rect -23 22092 149 22131
rect -23 22058 -17 22092
rect 17 22058 75 22092
rect 109 22082 149 22092
rect 201 22082 247 22134
rect 109 22070 167 22082
rect 201 22070 259 22082
rect 293 22070 299 22082
rect 109 22058 149 22070
rect -23 22019 149 22058
rect -23 21985 -17 22019
rect 17 21985 75 22019
rect 109 22018 149 22019
rect 201 22018 247 22070
rect 109 22006 167 22018
rect 201 22006 259 22018
rect 293 22006 299 22018
rect 109 21985 149 22006
rect -23 21954 149 21985
rect 201 21954 247 22006
rect -23 21946 299 21954
rect -23 21912 -17 21946
rect 17 21912 75 21946
rect 109 21942 167 21946
rect 201 21942 259 21946
rect 293 21942 299 21946
rect 109 21912 149 21942
rect -23 21890 149 21912
rect 201 21890 247 21942
rect -23 21878 299 21890
rect -23 21873 149 21878
rect -23 21839 -17 21873
rect 17 21839 75 21873
rect 109 21839 149 21873
rect -23 21826 149 21839
rect 201 21826 247 21878
rect -23 21814 299 21826
rect -23 21800 149 21814
rect -23 21766 -17 21800
rect 17 21766 75 21800
rect 109 21766 149 21800
rect -23 21762 149 21766
rect 201 21762 247 21814
rect -23 21750 299 21762
rect -23 21727 149 21750
rect -23 21693 -17 21727
rect 17 21693 75 21727
rect 109 21698 149 21727
rect 201 21698 247 21750
rect 109 21693 167 21698
rect 201 21693 259 21698
rect 293 21693 299 21698
rect -23 21686 299 21693
rect -23 21654 149 21686
rect -23 21620 -17 21654
rect 17 21620 75 21654
rect 109 21634 149 21654
rect 201 21634 247 21686
rect 109 21622 167 21634
rect 201 21622 259 21634
rect 293 21622 299 21634
rect 109 21620 149 21622
rect -23 21581 149 21620
rect -23 21547 -17 21581
rect 17 21547 75 21581
rect 109 21570 149 21581
rect 201 21570 247 21622
rect 109 21558 167 21570
rect 201 21558 259 21570
rect 293 21558 299 21570
rect 109 21547 149 21558
rect -23 21508 149 21547
rect -23 21474 -17 21508
rect 17 21474 75 21508
rect 109 21506 149 21508
rect 201 21506 247 21558
rect 109 21494 167 21506
rect 201 21494 259 21506
rect 293 21494 299 21506
rect 109 21474 149 21494
rect -23 21442 149 21474
rect 201 21442 247 21494
rect -23 21435 299 21442
rect -23 21401 -17 21435
rect 17 21401 75 21435
rect 109 21430 167 21435
rect 201 21430 259 21435
rect 293 21430 299 21435
rect 109 21401 149 21430
rect -23 21378 149 21401
rect 201 21378 247 21430
rect -23 21366 299 21378
rect -23 21362 149 21366
rect -23 21328 -17 21362
rect 17 21328 75 21362
rect 109 21328 149 21362
rect -23 21314 149 21328
rect 201 21314 247 21366
rect -23 21302 299 21314
rect -23 21289 149 21302
rect -23 21255 -17 21289
rect 17 21255 75 21289
rect 109 21255 149 21289
rect -23 21250 149 21255
rect 201 21250 247 21302
rect -23 21238 299 21250
rect -23 21216 149 21238
rect -23 21182 -17 21216
rect 17 21182 75 21216
rect 109 21186 149 21216
rect 201 21186 247 21238
rect 109 21182 167 21186
rect 201 21182 259 21186
rect 293 21182 299 21186
rect -23 21174 299 21182
rect -23 21143 149 21174
rect -23 21109 -17 21143
rect 17 21109 75 21143
rect 109 21122 149 21143
rect 201 21122 247 21174
rect 109 21110 167 21122
rect 201 21110 259 21122
rect 293 21110 299 21122
rect 109 21109 149 21110
rect -23 21070 149 21109
rect -23 21036 -17 21070
rect 17 21036 75 21070
rect 109 21058 149 21070
rect 201 21058 247 21110
rect 109 21046 167 21058
rect 201 21046 259 21058
rect 293 21046 299 21058
rect 109 21036 149 21046
rect -23 20997 149 21036
rect -23 20963 -17 20997
rect 17 20963 75 20997
rect 109 20994 149 20997
rect 201 20994 247 21046
rect 109 20982 167 20994
rect 201 20982 259 20994
rect 293 20982 299 20994
rect 109 20963 149 20982
rect -23 20930 149 20963
rect 201 20930 247 20982
rect -23 20924 299 20930
rect -23 20890 -17 20924
rect 17 20890 75 20924
rect 109 20918 167 20924
rect 201 20918 259 20924
rect 293 20918 299 20924
rect 109 20890 149 20918
rect -23 20866 149 20890
rect 201 20866 247 20918
rect -23 20854 299 20866
rect -23 20851 149 20854
rect -23 20817 -17 20851
rect 17 20817 75 20851
rect 109 20817 149 20851
rect -23 20802 149 20817
rect 201 20802 247 20854
rect -23 20790 299 20802
rect -23 20778 149 20790
rect -23 20744 -17 20778
rect 17 20744 75 20778
rect 109 20744 149 20778
rect -23 20738 149 20744
rect 201 20738 247 20790
rect -23 20726 299 20738
rect -23 20705 149 20726
rect -23 20671 -17 20705
rect 17 20671 75 20705
rect 109 20674 149 20705
rect 201 20674 247 20726
rect 109 20671 167 20674
rect 201 20671 259 20674
rect 293 20671 299 20674
rect -23 20662 299 20671
rect -23 20632 149 20662
rect -23 20598 -17 20632
rect 17 20598 75 20632
rect 109 20610 149 20632
rect 201 20610 247 20662
rect 109 20598 167 20610
rect 201 20598 259 20610
rect 293 20598 299 20610
rect -23 20559 149 20598
rect -23 20525 -17 20559
rect 17 20525 75 20559
rect 109 20546 149 20559
rect 201 20546 247 20598
rect 109 20534 167 20546
rect 201 20534 259 20546
rect 293 20534 299 20546
rect 109 20525 149 20534
rect -23 20486 149 20525
rect -23 20452 -17 20486
rect 17 20452 75 20486
rect 109 20482 149 20486
rect 201 20482 247 20534
rect 109 20470 167 20482
rect 201 20470 259 20482
rect 293 20470 299 20482
rect 109 20452 149 20470
rect -23 20418 149 20452
rect 201 20418 247 20470
rect -23 20413 299 20418
rect -23 20379 -17 20413
rect 17 20379 75 20413
rect 109 20406 167 20413
rect 201 20406 259 20413
rect 293 20406 299 20413
rect 109 20379 149 20406
rect -23 20354 149 20379
rect 201 20354 247 20406
rect -23 20342 299 20354
rect -23 20340 149 20342
rect -23 20306 -17 20340
rect 17 20306 75 20340
rect 109 20306 149 20340
rect -23 20290 149 20306
rect 201 20290 247 20342
rect -23 20277 299 20290
rect -23 20267 149 20277
rect -23 20233 -17 20267
rect 17 20233 75 20267
rect 109 20233 149 20267
rect -23 20225 149 20233
rect 201 20225 247 20277
rect -23 20212 299 20225
rect -23 20194 149 20212
rect -23 20160 -17 20194
rect 17 20160 75 20194
rect 109 20160 149 20194
rect 201 20160 247 20212
rect -23 20147 299 20160
rect -23 20121 149 20147
rect -23 20087 -17 20121
rect 17 20087 75 20121
rect 109 20095 149 20121
rect 201 20095 247 20147
rect 109 20087 167 20095
rect 201 20087 259 20095
rect 293 20087 299 20095
rect -23 20082 299 20087
rect -23 20048 149 20082
rect -23 20014 -17 20048
rect 17 20014 75 20048
rect 109 20030 149 20048
rect 201 20030 247 20082
rect 109 20017 167 20030
rect 201 20017 259 20030
rect 293 20017 299 20030
rect 109 20014 149 20017
rect -23 19975 149 20014
rect -23 19941 -17 19975
rect 17 19941 75 19975
rect 109 19965 149 19975
rect 201 19965 247 20017
rect 109 19952 167 19965
rect 201 19952 259 19965
rect 293 19952 299 19965
rect 109 19941 149 19952
rect -23 19902 149 19941
rect -23 19868 -17 19902
rect 17 19868 75 19902
rect 109 19900 149 19902
rect 201 19900 247 19952
rect 109 19887 167 19900
rect 201 19887 259 19900
rect 293 19887 299 19900
rect 109 19868 149 19887
rect -23 19835 149 19868
rect 201 19835 247 19887
rect -23 19829 299 19835
rect -23 19795 -17 19829
rect 17 19795 75 19829
rect 109 19822 167 19829
rect 201 19822 259 19829
rect 293 19822 299 19829
rect 109 19795 149 19822
rect -23 19770 149 19795
rect 201 19770 247 19822
rect -23 19757 299 19770
rect -23 19756 149 19757
rect -23 19722 -17 19756
rect 17 19722 75 19756
rect 109 19722 149 19756
rect -23 19705 149 19722
rect 201 19705 247 19757
rect -23 19692 299 19705
rect -23 19683 149 19692
rect -23 19649 -17 19683
rect 17 19649 75 19683
rect 109 19649 149 19683
rect -23 19640 149 19649
rect 201 19640 247 19692
rect -23 19627 299 19640
rect -23 19610 149 19627
rect -23 19576 -17 19610
rect 17 19576 75 19610
rect 109 19576 149 19610
rect -23 19575 149 19576
rect 201 19575 247 19627
rect -23 19562 299 19575
rect -23 19537 149 19562
rect -23 19503 -17 19537
rect 17 19503 75 19537
rect 109 19510 149 19537
rect 201 19510 247 19562
rect 109 19503 167 19510
rect 201 19503 259 19510
rect 293 19503 299 19510
rect -23 19497 299 19503
rect -23 19464 149 19497
rect -23 19430 -17 19464
rect 17 19430 75 19464
rect 109 19445 149 19464
rect 201 19445 247 19497
rect 109 19432 167 19445
rect 201 19432 259 19445
rect 293 19432 299 19445
rect 109 19430 149 19432
rect -23 19391 149 19430
rect -23 19357 -17 19391
rect 17 19357 75 19391
rect 109 19380 149 19391
rect 201 19380 247 19432
rect 109 19367 167 19380
rect 201 19367 259 19380
rect 293 19367 299 19380
rect 109 19357 149 19367
rect -23 19318 149 19357
rect -23 19284 -17 19318
rect 17 19284 75 19318
rect 109 19315 149 19318
rect 201 19315 247 19367
rect 109 19302 167 19315
rect 201 19302 259 19315
rect 293 19302 299 19315
rect 109 19284 149 19302
rect -23 19250 149 19284
rect 201 19250 247 19302
rect -23 19245 299 19250
rect -23 19211 -17 19245
rect 17 19211 75 19245
rect 109 19237 167 19245
rect 201 19237 259 19245
rect 293 19237 299 19245
rect 109 19211 149 19237
rect -23 19185 149 19211
rect 201 19185 247 19237
rect -23 19179 299 19185
rect 453 26038 973 26044
rect 453 25986 456 26038
rect 508 25986 524 26038
rect 576 25986 592 26038
rect 644 26012 660 26038
rect 712 26012 728 26038
rect 780 26012 796 26038
rect 848 26029 973 26038
tri 973 26029 988 26044 sw
rect 14076 26029 16029 26044
rect 848 26021 988 26029
tri 988 26021 996 26029 sw
rect 13821 26021 16029 26029
rect 649 25986 660 26012
rect 727 25986 728 26012
rect 848 25988 996 26021
rect 848 25986 863 25988
rect 453 25978 459 25986
rect 493 25978 537 25986
rect 571 25978 615 25986
rect 649 25978 693 25986
rect 727 25978 771 25986
rect 805 25978 863 25986
rect 453 25974 863 25978
rect 453 25922 456 25974
rect 508 25922 524 25974
rect 576 25922 592 25974
rect 644 25940 660 25974
rect 712 25940 728 25974
rect 780 25940 796 25974
rect 848 25954 863 25974
rect 897 25987 996 25988
tri 996 25987 1030 26021 sw
rect 13821 25987 13833 26021
rect 13867 25987 13906 26021
rect 13940 25987 13979 26021
rect 14013 25987 14052 26021
rect 14086 25987 14125 26021
rect 14159 25987 14198 26021
rect 14232 25987 14271 26021
rect 14305 25987 14344 26021
rect 14378 25987 14417 26021
rect 14451 25987 14490 26021
rect 14524 25987 14563 26021
rect 14597 25987 14636 26021
rect 14670 25987 14709 26021
rect 14743 25987 14782 26021
rect 14816 25987 14855 26021
rect 14889 25987 14928 26021
rect 14962 25987 15001 26021
rect 15035 25987 15074 26021
rect 15108 25987 15147 26021
rect 15181 25987 15220 26021
rect 15254 25987 15293 26021
rect 15327 25987 15366 26021
rect 15400 25987 15439 26021
rect 15473 25987 15513 26021
rect 15547 25987 15587 26021
rect 15621 25987 15661 26021
rect 15695 25987 15735 26021
rect 15769 25987 15809 26021
rect 15843 25987 15883 26021
rect 15917 25987 16029 26021
rect 897 25954 1030 25987
rect 848 25947 1030 25954
tri 1030 25947 1070 25987 sw
rect 13821 25947 16029 25987
rect 649 25922 660 25940
rect 727 25922 728 25940
rect 848 25922 1070 25947
rect 453 25910 459 25922
rect 493 25910 537 25922
rect 571 25910 615 25922
rect 649 25910 693 25922
rect 727 25910 771 25922
rect 805 25915 1070 25922
rect 805 25910 863 25915
rect 453 25858 456 25910
rect 508 25858 524 25910
rect 576 25858 592 25910
rect 649 25906 660 25910
rect 727 25906 728 25910
rect 644 25868 660 25906
rect 712 25868 728 25906
rect 780 25868 796 25906
rect 848 25881 863 25910
rect 897 25913 1070 25915
tri 1070 25913 1104 25947 sw
rect 13821 25913 13833 25947
rect 13867 25913 13906 25947
rect 13940 25913 13979 25947
rect 14013 25913 14052 25947
rect 14086 25913 14125 25947
rect 14159 25913 14198 25947
rect 14232 25913 14271 25947
rect 14305 25913 14344 25947
rect 14378 25913 14417 25947
rect 14451 25913 14490 25947
rect 14524 25913 14563 25947
rect 14597 25913 14636 25947
rect 14670 25913 14709 25947
rect 14743 25913 14782 25947
rect 14816 25913 14855 25947
rect 14889 25913 14928 25947
rect 14962 25913 15001 25947
rect 15035 25913 15074 25947
rect 15108 25913 15147 25947
rect 15181 25913 15220 25947
rect 15254 25913 15293 25947
rect 15327 25913 15366 25947
rect 15400 25913 15439 25947
rect 15473 25913 15513 25947
rect 15547 25913 15587 25947
rect 15621 25913 15661 25947
rect 15695 25913 15735 25947
rect 15769 25913 15809 25947
rect 15843 25913 15883 25947
rect 15917 25913 16029 25947
rect 897 25881 1104 25913
rect 848 25873 1104 25881
tri 1104 25873 1144 25913 sw
rect 13821 25873 16029 25913
rect 649 25858 660 25868
rect 727 25858 728 25868
rect 848 25858 1144 25873
rect 453 25846 459 25858
rect 493 25846 537 25858
rect 571 25846 615 25858
rect 649 25846 693 25858
rect 727 25846 771 25858
rect 805 25846 1144 25858
rect 453 25794 456 25846
rect 508 25794 524 25846
rect 576 25794 592 25846
rect 649 25834 660 25846
rect 727 25834 728 25846
rect 848 25842 1144 25846
rect 644 25796 660 25834
rect 712 25796 728 25834
rect 780 25796 796 25834
rect 848 25808 863 25842
rect 897 25839 1144 25842
tri 1144 25839 1178 25873 sw
rect 13821 25839 13833 25873
rect 13867 25839 13906 25873
rect 13940 25839 13979 25873
rect 14013 25839 14052 25873
rect 14086 25839 14125 25873
rect 14159 25839 14198 25873
rect 14232 25839 14271 25873
rect 14305 25839 14344 25873
rect 14378 25839 14417 25873
rect 14451 25839 14490 25873
rect 14524 25839 14563 25873
rect 14597 25839 14636 25873
rect 14670 25839 14709 25873
rect 14743 25839 14782 25873
rect 14816 25839 14855 25873
rect 14889 25839 14928 25873
rect 14962 25839 15001 25873
rect 15035 25839 15074 25873
rect 15108 25839 15147 25873
rect 15181 25839 15220 25873
rect 15254 25839 15293 25873
rect 15327 25839 15366 25873
rect 15400 25839 15439 25873
rect 15473 25839 15513 25873
rect 15547 25839 15587 25873
rect 15621 25839 15661 25873
rect 15695 25839 15735 25873
rect 15769 25839 15809 25873
rect 15843 25839 15883 25873
rect 15917 25839 16029 25873
rect 897 25808 1178 25839
rect 848 25799 1178 25808
tri 1178 25799 1218 25839 sw
rect 13821 25799 16029 25839
rect 649 25794 660 25796
rect 727 25794 728 25796
rect 848 25794 1218 25799
rect 453 25782 459 25794
rect 493 25782 537 25794
rect 571 25782 615 25794
rect 649 25782 693 25794
rect 727 25782 771 25794
rect 805 25782 1218 25794
rect 453 25730 456 25782
rect 508 25730 524 25782
rect 576 25730 592 25782
rect 649 25762 660 25782
rect 727 25762 728 25782
rect 848 25769 1218 25782
rect 644 25730 660 25762
rect 712 25730 728 25762
rect 780 25730 796 25762
rect 848 25735 863 25769
rect 897 25765 1218 25769
tri 1218 25765 1252 25799 sw
rect 13821 25765 13833 25799
rect 13867 25765 13906 25799
rect 13940 25765 13979 25799
rect 14013 25765 14052 25799
rect 14086 25765 14125 25799
rect 14159 25765 14198 25799
rect 14232 25765 14271 25799
rect 14305 25765 14344 25799
rect 14378 25765 14417 25799
rect 14451 25765 14490 25799
rect 14524 25765 14563 25799
rect 14597 25765 14636 25799
rect 14670 25765 14709 25799
rect 14743 25765 14782 25799
rect 14816 25765 14855 25799
rect 14889 25765 14928 25799
rect 14962 25765 15001 25799
rect 15035 25765 15074 25799
rect 15108 25765 15147 25799
rect 15181 25765 15220 25799
rect 15254 25765 15293 25799
rect 15327 25765 15366 25799
rect 15400 25765 15439 25799
rect 15473 25765 15513 25799
rect 15547 25765 15587 25799
rect 15621 25765 15661 25799
rect 15695 25765 15735 25799
rect 15769 25765 15809 25799
rect 15843 25765 15883 25799
rect 15917 25765 16029 25799
rect 897 25735 1252 25765
rect 848 25730 1252 25735
rect 453 25725 1252 25730
tri 1252 25725 1292 25765 sw
rect 13821 25725 16029 25765
rect 453 25724 1292 25725
rect 453 25718 459 25724
rect 493 25718 537 25724
rect 571 25718 615 25724
rect 649 25718 693 25724
rect 727 25718 771 25724
rect 805 25718 1292 25724
rect 453 25666 456 25718
rect 508 25666 524 25718
rect 576 25666 592 25718
rect 649 25690 660 25718
rect 727 25690 728 25718
rect 848 25696 1292 25718
rect 644 25666 660 25690
rect 712 25666 728 25690
rect 780 25666 796 25690
rect 848 25666 863 25696
rect 453 25662 863 25666
rect 897 25691 1292 25696
tri 1292 25691 1326 25725 sw
rect 13821 25691 13833 25725
rect 13867 25691 13906 25725
rect 13940 25691 13979 25725
rect 14013 25691 14052 25725
rect 14086 25691 14125 25725
rect 14159 25691 14198 25725
rect 14232 25691 14271 25725
rect 14305 25691 14344 25725
rect 14378 25691 14417 25725
rect 14451 25691 14490 25725
rect 14524 25691 14563 25725
rect 14597 25691 14636 25725
rect 14670 25691 14709 25725
rect 14743 25691 14782 25725
rect 14816 25691 14855 25725
rect 14889 25691 14928 25725
rect 14962 25691 15001 25725
rect 15035 25691 15074 25725
rect 15108 25691 15147 25725
rect 15181 25691 15220 25725
rect 15254 25691 15293 25725
rect 15327 25691 15366 25725
rect 15400 25691 15439 25725
rect 15473 25691 15513 25725
rect 15547 25691 15587 25725
rect 15621 25691 15661 25725
rect 15695 25691 15735 25725
rect 15769 25691 15809 25725
rect 15843 25691 15883 25725
rect 15917 25691 16029 25725
rect 897 25683 1326 25691
tri 1326 25683 1334 25691 sw
rect 13821 25683 16029 25691
rect 897 25662 1334 25683
rect 453 25654 1334 25662
rect 453 25602 456 25654
rect 508 25602 524 25654
rect 576 25602 592 25654
rect 644 25652 660 25654
rect 712 25652 728 25654
rect 780 25652 796 25654
rect 649 25618 660 25652
rect 727 25618 728 25652
rect 848 25646 1334 25654
tri 1334 25646 1371 25683 sw
rect 14076 25652 16029 25683
rect 848 25623 971 25646
rect 644 25602 660 25618
rect 712 25602 728 25618
rect 780 25602 796 25618
rect 848 25602 863 25623
rect 453 25590 863 25602
rect 453 25538 456 25590
rect 508 25538 524 25590
rect 576 25538 592 25590
rect 644 25580 660 25590
rect 712 25580 728 25590
rect 780 25580 796 25590
rect 848 25589 863 25590
rect 897 25589 971 25623
rect 649 25546 660 25580
rect 727 25546 728 25580
rect 848 25550 971 25589
rect 644 25538 660 25546
rect 712 25538 728 25546
rect 780 25538 796 25546
rect 848 25538 863 25550
rect 453 25526 863 25538
rect 453 25474 456 25526
rect 508 25474 524 25526
rect 576 25474 592 25526
rect 644 25508 660 25526
rect 712 25508 728 25526
rect 780 25508 796 25526
rect 848 25516 863 25526
rect 897 25516 971 25550
rect 649 25474 660 25508
rect 727 25474 728 25508
rect 848 25476 971 25516
rect 848 25474 863 25476
rect 453 25462 863 25474
rect 453 25410 456 25462
rect 508 25410 524 25462
rect 576 25410 592 25462
rect 644 25436 660 25462
rect 712 25436 728 25462
rect 780 25436 796 25462
rect 848 25442 863 25462
rect 897 25442 971 25476
rect 649 25410 660 25436
rect 727 25410 728 25436
rect 848 25410 971 25442
rect 453 25402 459 25410
rect 493 25402 537 25410
rect 571 25402 615 25410
rect 649 25402 693 25410
rect 727 25402 771 25410
rect 805 25402 971 25410
rect 453 25398 863 25402
rect 453 25346 456 25398
rect 508 25346 524 25398
rect 576 25346 592 25398
rect 644 25364 660 25398
rect 712 25364 728 25398
rect 780 25364 796 25398
rect 848 25368 863 25398
rect 897 25368 971 25402
rect 649 25346 660 25364
rect 727 25346 728 25364
rect 848 25346 971 25368
rect 453 25334 459 25346
rect 493 25334 537 25346
rect 571 25334 615 25346
rect 649 25334 693 25346
rect 727 25334 771 25346
rect 805 25334 971 25346
rect 453 25282 456 25334
rect 508 25282 524 25334
rect 576 25282 592 25334
rect 649 25330 660 25334
rect 727 25330 728 25334
rect 644 25292 660 25330
rect 712 25292 728 25330
rect 780 25292 796 25330
rect 848 25328 971 25334
rect 848 25294 863 25328
rect 897 25294 971 25328
rect 649 25282 660 25292
rect 727 25282 728 25292
rect 848 25282 971 25294
rect 453 25270 459 25282
rect 493 25270 537 25282
rect 571 25270 615 25282
rect 649 25270 693 25282
rect 727 25270 771 25282
rect 805 25270 971 25282
rect 453 25218 456 25270
rect 508 25218 524 25270
rect 576 25218 592 25270
rect 649 25258 660 25270
rect 727 25258 728 25270
rect 848 25263 971 25270
rect 644 25220 660 25258
rect 712 25220 728 25258
rect 780 25220 796 25258
rect 649 25218 660 25220
rect 727 25218 728 25220
rect 848 25218 850 25263
rect 453 25206 459 25218
rect 493 25206 537 25218
rect 571 25206 615 25218
rect 649 25206 693 25218
rect 727 25206 771 25218
rect 805 25206 850 25218
rect 453 25154 456 25206
rect 508 25154 524 25206
rect 576 25154 592 25206
rect 649 25186 660 25206
rect 727 25186 728 25206
rect 644 25154 660 25186
rect 712 25154 728 25186
rect 780 25154 796 25186
rect 848 25154 850 25206
rect 453 25148 850 25154
rect 453 25142 459 25148
rect 493 25142 537 25148
rect 571 25142 615 25148
rect 649 25142 693 25148
rect 727 25142 771 25148
rect 805 25142 850 25148
rect 453 25090 456 25142
rect 508 25090 524 25142
rect 576 25090 592 25142
rect 649 25114 660 25142
rect 727 25114 728 25142
rect 644 25090 660 25114
rect 712 25090 728 25114
rect 780 25090 796 25114
rect 848 25090 850 25142
rect 453 25078 850 25090
rect 453 25026 456 25078
rect 508 25026 524 25078
rect 576 25026 592 25078
rect 644 25076 660 25078
rect 712 25076 728 25078
rect 780 25076 796 25078
rect 649 25042 660 25076
rect 727 25042 728 25076
rect 644 25026 660 25042
rect 712 25026 728 25042
rect 780 25026 796 25042
rect 848 25026 850 25078
rect 453 25014 850 25026
rect 453 24962 456 25014
rect 508 24962 524 25014
rect 576 24962 592 25014
rect 644 25004 660 25014
rect 712 25004 728 25014
rect 780 25004 796 25014
rect 649 24970 660 25004
rect 727 24970 728 25004
rect 644 24962 660 24970
rect 712 24962 728 24970
rect 780 24962 796 24970
rect 848 24962 850 25014
rect 453 24950 850 24962
rect 453 24898 456 24950
rect 508 24898 524 24950
rect 576 24898 592 24950
rect 644 24932 660 24950
rect 712 24932 728 24950
rect 780 24932 796 24950
rect 649 24898 660 24932
rect 727 24898 728 24932
rect 848 24898 850 24950
rect 453 24886 850 24898
rect 453 24834 456 24886
rect 508 24834 524 24886
rect 576 24834 592 24886
rect 644 24860 660 24886
rect 712 24860 728 24886
rect 780 24860 796 24886
rect 649 24834 660 24860
rect 727 24834 728 24860
rect 848 24834 850 24886
rect 453 24826 459 24834
rect 493 24826 537 24834
rect 571 24826 615 24834
rect 649 24826 693 24834
rect 727 24826 771 24834
rect 805 24826 850 24834
rect 453 24822 850 24826
rect 453 24770 456 24822
rect 508 24770 524 24822
rect 576 24770 592 24822
rect 644 24788 660 24822
rect 712 24788 728 24822
rect 780 24788 796 24822
rect 649 24770 660 24788
rect 727 24770 728 24788
rect 848 24770 850 24822
rect 453 24758 459 24770
rect 493 24758 537 24770
rect 571 24758 615 24770
rect 649 24758 693 24770
rect 727 24758 771 24770
rect 805 24758 850 24770
rect 453 24706 456 24758
rect 508 24706 524 24758
rect 576 24706 592 24758
rect 649 24754 660 24758
rect 727 24754 728 24758
rect 644 24716 660 24754
rect 712 24716 728 24754
rect 780 24716 796 24754
rect 649 24706 660 24716
rect 727 24706 728 24716
rect 848 24706 850 24758
rect 453 24694 459 24706
rect 493 24694 537 24706
rect 571 24694 615 24706
rect 649 24694 693 24706
rect 727 24694 771 24706
rect 805 24694 850 24706
rect 453 24642 456 24694
rect 508 24642 524 24694
rect 576 24642 592 24694
rect 649 24682 660 24694
rect 727 24682 728 24694
rect 644 24644 660 24682
rect 712 24644 728 24682
rect 780 24644 796 24682
rect 649 24642 660 24644
rect 727 24642 728 24644
rect 848 24642 850 24694
rect 453 24630 459 24642
rect 493 24630 537 24642
rect 571 24630 615 24642
rect 649 24630 693 24642
rect 727 24630 771 24642
rect 805 24630 850 24642
rect 453 24578 456 24630
rect 508 24578 524 24630
rect 576 24578 592 24630
rect 649 24610 660 24630
rect 727 24610 728 24630
rect 644 24578 660 24610
rect 712 24578 728 24610
rect 780 24578 796 24610
rect 848 24578 850 24630
rect 453 24572 850 24578
rect 453 24566 459 24572
rect 493 24566 537 24572
rect 571 24566 615 24572
rect 649 24566 693 24572
rect 727 24566 771 24572
rect 805 24566 850 24572
rect 453 24514 456 24566
rect 508 24514 524 24566
rect 576 24514 592 24566
rect 649 24538 660 24566
rect 727 24538 728 24566
rect 644 24514 660 24538
rect 712 24514 728 24538
rect 780 24514 796 24538
rect 848 24514 850 24566
rect 453 24502 850 24514
rect 453 24450 456 24502
rect 508 24450 524 24502
rect 576 24450 592 24502
rect 644 24500 660 24502
rect 712 24500 728 24502
rect 780 24500 796 24502
rect 649 24466 660 24500
rect 727 24466 728 24500
rect 644 24450 660 24466
rect 712 24450 728 24466
rect 780 24450 796 24466
rect 848 24450 850 24502
rect 453 24438 850 24450
rect 453 24386 456 24438
rect 508 24386 524 24438
rect 576 24386 592 24438
rect 644 24428 660 24438
rect 712 24428 728 24438
rect 780 24428 796 24438
rect 649 24394 660 24428
rect 727 24394 728 24428
rect 644 24386 660 24394
rect 712 24386 728 24394
rect 780 24386 796 24394
rect 848 24386 850 24438
rect 453 24374 850 24386
rect 453 24322 456 24374
rect 508 24322 524 24374
rect 576 24322 592 24374
rect 644 24355 660 24374
rect 712 24355 728 24374
rect 780 24355 796 24374
rect 649 24322 660 24355
rect 727 24322 728 24355
rect 848 24322 850 24374
rect 453 24321 459 24322
rect 493 24321 537 24322
rect 571 24321 615 24322
rect 649 24321 693 24322
rect 727 24321 771 24322
rect 805 24321 850 24322
rect 453 24310 850 24321
rect 453 24258 456 24310
rect 508 24258 524 24310
rect 576 24258 592 24310
rect 644 24282 660 24310
rect 712 24282 728 24310
rect 780 24282 796 24310
rect 649 24258 660 24282
rect 727 24258 728 24282
rect 848 24258 850 24310
rect 453 24248 459 24258
rect 493 24248 537 24258
rect 571 24248 615 24258
rect 649 24248 693 24258
rect 727 24248 771 24258
rect 805 24248 850 24258
rect 453 24246 850 24248
rect 453 24194 456 24246
rect 508 24194 524 24246
rect 576 24194 592 24246
rect 644 24209 660 24246
rect 712 24209 728 24246
rect 780 24209 796 24246
rect 649 24194 660 24209
rect 727 24194 728 24209
rect 848 24194 850 24246
rect 453 24182 459 24194
rect 493 24182 537 24194
rect 571 24182 615 24194
rect 649 24182 693 24194
rect 727 24182 771 24194
rect 805 24182 850 24194
rect 453 24130 456 24182
rect 508 24130 524 24182
rect 576 24130 592 24182
rect 649 24175 660 24182
rect 727 24175 728 24182
rect 644 24136 660 24175
rect 712 24136 728 24175
rect 780 24136 796 24175
rect 649 24130 660 24136
rect 727 24130 728 24136
rect 848 24130 850 24182
rect 453 24118 459 24130
rect 493 24118 537 24130
rect 571 24118 615 24130
rect 649 24118 693 24130
rect 727 24118 771 24130
rect 805 24118 850 24130
rect 453 24066 456 24118
rect 508 24066 524 24118
rect 576 24066 592 24118
rect 649 24102 660 24118
rect 727 24102 728 24118
rect 644 24066 660 24102
rect 712 24066 728 24102
rect 780 24066 796 24102
rect 848 24066 850 24118
rect 453 24063 850 24066
rect 453 24054 459 24063
rect 493 24054 537 24063
rect 571 24054 615 24063
rect 649 24054 693 24063
rect 727 24054 771 24063
rect 805 24054 850 24063
rect 453 24002 456 24054
rect 508 24002 524 24054
rect 576 24002 592 24054
rect 649 24029 660 24054
rect 727 24029 728 24054
rect 644 24002 660 24029
rect 712 24002 728 24029
rect 780 24002 796 24029
rect 848 24002 850 24054
rect 453 23990 850 24002
rect 453 23938 456 23990
rect 508 23938 524 23990
rect 576 23938 592 23990
rect 649 23956 660 23990
rect 727 23956 728 23990
rect 644 23938 660 23956
rect 712 23938 728 23956
rect 780 23938 796 23956
rect 848 23938 850 23990
rect 453 23926 850 23938
rect 453 23874 456 23926
rect 508 23874 524 23926
rect 576 23874 592 23926
rect 644 23917 660 23926
rect 712 23917 728 23926
rect 780 23917 796 23926
rect 649 23883 660 23917
rect 727 23883 728 23917
rect 644 23874 660 23883
rect 712 23874 728 23883
rect 780 23874 796 23883
rect 848 23874 850 23926
rect 453 23862 850 23874
rect 453 23810 456 23862
rect 508 23810 524 23862
rect 576 23810 592 23862
rect 644 23844 660 23862
rect 712 23844 728 23862
rect 780 23844 796 23862
rect 649 23810 660 23844
rect 727 23810 728 23844
rect 848 23810 850 23862
rect 453 23798 850 23810
rect 453 23746 456 23798
rect 508 23746 524 23798
rect 576 23746 592 23798
rect 644 23771 660 23798
rect 712 23771 728 23798
rect 780 23771 796 23798
rect 649 23746 660 23771
rect 727 23746 728 23771
rect 848 23746 850 23798
rect 453 23737 459 23746
rect 493 23737 537 23746
rect 571 23737 615 23746
rect 649 23737 693 23746
rect 727 23737 771 23746
rect 805 23737 850 23746
rect 453 23734 850 23737
rect 453 23682 456 23734
rect 508 23682 524 23734
rect 576 23682 592 23734
rect 644 23698 660 23734
rect 712 23698 728 23734
rect 780 23698 796 23734
rect 649 23682 660 23698
rect 727 23682 728 23698
rect 848 23682 850 23734
rect 453 23670 459 23682
rect 493 23670 537 23682
rect 571 23670 615 23682
rect 649 23670 693 23682
rect 727 23670 771 23682
rect 805 23670 850 23682
rect 453 23618 456 23670
rect 508 23618 524 23670
rect 576 23618 592 23670
rect 649 23664 660 23670
rect 727 23664 728 23670
rect 644 23625 660 23664
rect 712 23625 728 23664
rect 780 23625 796 23664
rect 649 23618 660 23625
rect 727 23618 728 23625
rect 848 23618 850 23670
rect 453 23606 459 23618
rect 493 23606 537 23618
rect 571 23606 615 23618
rect 649 23606 693 23618
rect 727 23606 771 23618
rect 805 23606 850 23618
rect 453 23554 456 23606
rect 508 23554 524 23606
rect 576 23554 592 23606
rect 649 23591 660 23606
rect 727 23591 728 23606
rect 644 23554 660 23591
rect 712 23554 728 23591
rect 780 23554 796 23591
rect 848 23554 850 23606
rect 453 23552 850 23554
rect 453 23542 459 23552
rect 493 23542 537 23552
rect 571 23542 615 23552
rect 649 23542 693 23552
rect 727 23542 771 23552
rect 805 23542 850 23552
rect 453 23490 456 23542
rect 508 23490 524 23542
rect 576 23490 592 23542
rect 649 23518 660 23542
rect 727 23518 728 23542
rect 644 23490 660 23518
rect 712 23490 728 23518
rect 780 23490 796 23518
rect 848 23490 850 23542
rect 453 23479 850 23490
rect 453 23478 459 23479
rect 493 23478 537 23479
rect 571 23478 615 23479
rect 649 23478 693 23479
rect 727 23478 771 23479
rect 805 23478 850 23479
rect 453 23426 456 23478
rect 508 23426 524 23478
rect 576 23426 592 23478
rect 649 23445 660 23478
rect 727 23445 728 23478
rect 644 23426 660 23445
rect 712 23426 728 23445
rect 780 23426 796 23445
rect 848 23426 850 23478
rect 453 23414 850 23426
rect 453 23362 456 23414
rect 508 23362 524 23414
rect 576 23362 592 23414
rect 644 23406 660 23414
rect 712 23406 728 23414
rect 780 23406 796 23414
rect 649 23372 660 23406
rect 727 23372 728 23406
rect 644 23362 660 23372
rect 712 23362 728 23372
rect 780 23362 796 23372
rect 848 23362 850 23414
rect 453 23350 850 23362
rect 453 23298 456 23350
rect 508 23298 524 23350
rect 576 23298 592 23350
rect 644 23333 660 23350
rect 712 23333 728 23350
rect 780 23333 796 23350
rect 649 23299 660 23333
rect 727 23299 728 23333
rect 644 23298 660 23299
rect 712 23298 728 23299
rect 780 23298 796 23299
rect 848 23298 850 23350
rect 453 23286 850 23298
rect 453 23234 456 23286
rect 508 23234 524 23286
rect 576 23234 592 23286
rect 644 23260 660 23286
rect 712 23260 728 23286
rect 780 23260 796 23286
rect 649 23234 660 23260
rect 727 23234 728 23260
rect 848 23234 850 23286
rect 453 23226 459 23234
rect 493 23226 537 23234
rect 571 23226 615 23234
rect 649 23226 693 23234
rect 727 23226 771 23234
rect 805 23226 850 23234
rect 453 23222 850 23226
rect 453 23170 456 23222
rect 508 23170 524 23222
rect 576 23170 592 23222
rect 644 23187 660 23222
rect 712 23187 728 23222
rect 780 23187 796 23222
rect 649 23170 660 23187
rect 727 23170 728 23187
rect 848 23170 850 23222
rect 453 23158 459 23170
rect 493 23158 537 23170
rect 571 23158 615 23170
rect 649 23158 693 23170
rect 727 23158 771 23170
rect 805 23158 850 23170
rect 453 23106 456 23158
rect 508 23106 524 23158
rect 576 23106 592 23158
rect 649 23153 660 23158
rect 727 23153 728 23158
rect 644 23114 660 23153
rect 712 23114 728 23153
rect 780 23114 796 23153
rect 649 23106 660 23114
rect 727 23106 728 23114
rect 848 23106 850 23158
rect 453 23094 459 23106
rect 493 23094 537 23106
rect 571 23094 615 23106
rect 649 23094 693 23106
rect 727 23094 771 23106
rect 805 23094 850 23106
rect 453 23042 456 23094
rect 508 23042 524 23094
rect 576 23042 592 23094
rect 649 23080 660 23094
rect 727 23080 728 23094
rect 644 23042 660 23080
rect 712 23042 728 23080
rect 780 23042 796 23080
rect 848 23042 850 23094
rect 453 23041 850 23042
rect 453 23030 459 23041
rect 493 23030 537 23041
rect 571 23030 615 23041
rect 649 23030 693 23041
rect 727 23030 771 23041
rect 805 23030 850 23041
rect 453 22978 456 23030
rect 508 22978 524 23030
rect 576 22978 592 23030
rect 649 23007 660 23030
rect 727 23007 728 23030
rect 644 22978 660 23007
rect 712 22978 728 23007
rect 780 22978 796 23007
rect 848 22978 850 23030
rect 453 22968 850 22978
rect 453 22966 459 22968
rect 493 22966 537 22968
rect 571 22966 615 22968
rect 649 22966 693 22968
rect 727 22966 771 22968
rect 805 22966 850 22968
rect 453 22914 456 22966
rect 508 22914 524 22966
rect 576 22914 592 22966
rect 649 22934 660 22966
rect 727 22934 728 22966
rect 644 22914 660 22934
rect 712 22914 728 22934
rect 780 22914 796 22934
rect 848 22914 850 22966
rect 453 22902 850 22914
rect 453 22850 456 22902
rect 508 22850 524 22902
rect 576 22850 592 22902
rect 644 22895 660 22902
rect 712 22895 728 22902
rect 780 22895 796 22902
rect 649 22861 660 22895
rect 727 22861 728 22895
rect 644 22850 660 22861
rect 712 22850 728 22861
rect 780 22850 796 22861
rect 848 22850 850 22902
rect 453 22838 850 22850
rect 453 22786 456 22838
rect 508 22786 524 22838
rect 576 22786 592 22838
rect 644 22822 660 22838
rect 712 22822 728 22838
rect 780 22822 796 22838
rect 649 22788 660 22822
rect 727 22788 728 22822
rect 644 22786 660 22788
rect 712 22786 728 22788
rect 780 22786 796 22788
rect 848 22786 850 22838
rect 453 22774 850 22786
rect 453 22722 456 22774
rect 508 22722 524 22774
rect 576 22722 592 22774
rect 644 22749 660 22774
rect 712 22749 728 22774
rect 780 22749 796 22774
rect 649 22722 660 22749
rect 727 22722 728 22749
rect 848 22722 850 22774
rect 453 22715 459 22722
rect 493 22715 537 22722
rect 571 22715 615 22722
rect 649 22715 693 22722
rect 727 22715 771 22722
rect 805 22715 850 22722
rect 453 22710 850 22715
rect 453 22658 456 22710
rect 508 22658 524 22710
rect 576 22658 592 22710
rect 644 22676 660 22710
rect 712 22676 728 22710
rect 780 22676 796 22710
rect 649 22658 660 22676
rect 727 22658 728 22676
rect 848 22658 850 22710
rect 453 22646 459 22658
rect 493 22646 537 22658
rect 571 22646 615 22658
rect 649 22646 693 22658
rect 727 22646 771 22658
rect 805 22646 850 22658
rect 453 22594 456 22646
rect 508 22594 524 22646
rect 576 22594 592 22646
rect 649 22642 660 22646
rect 727 22642 728 22646
rect 644 22603 660 22642
rect 712 22603 728 22642
rect 780 22603 796 22642
rect 649 22594 660 22603
rect 727 22594 728 22603
rect 848 22594 850 22646
rect 453 22582 459 22594
rect 493 22582 537 22594
rect 571 22582 615 22594
rect 649 22582 693 22594
rect 727 22582 771 22594
rect 805 22582 850 22594
rect 453 22530 456 22582
rect 508 22530 524 22582
rect 576 22530 592 22582
rect 649 22569 660 22582
rect 727 22569 728 22582
rect 644 22530 660 22569
rect 712 22530 728 22569
rect 780 22530 796 22569
rect 848 22530 850 22582
rect 453 22518 459 22530
rect 493 22518 537 22530
rect 571 22518 615 22530
rect 649 22518 693 22530
rect 727 22518 771 22530
rect 805 22518 850 22530
rect 453 22466 456 22518
rect 508 22466 524 22518
rect 576 22466 592 22518
rect 649 22496 660 22518
rect 727 22496 728 22518
rect 644 22466 660 22496
rect 712 22466 728 22496
rect 780 22466 796 22496
rect 848 22466 850 22518
rect 453 22457 850 22466
rect 453 22454 459 22457
rect 493 22454 537 22457
rect 571 22454 615 22457
rect 649 22454 693 22457
rect 727 22454 771 22457
rect 805 22454 850 22457
rect 453 22402 456 22454
rect 508 22402 524 22454
rect 576 22402 592 22454
rect 649 22423 660 22454
rect 727 22423 728 22454
rect 644 22402 660 22423
rect 712 22402 728 22423
rect 780 22402 796 22423
rect 848 22402 850 22454
rect 453 22390 850 22402
rect 453 22338 456 22390
rect 508 22338 524 22390
rect 576 22338 592 22390
rect 644 22384 660 22390
rect 712 22384 728 22390
rect 780 22384 796 22390
rect 649 22350 660 22384
rect 727 22350 728 22384
rect 644 22338 660 22350
rect 712 22338 728 22350
rect 780 22338 796 22350
rect 848 22338 850 22390
rect 453 22326 850 22338
rect 453 22274 456 22326
rect 508 22274 524 22326
rect 576 22274 592 22326
rect 644 22311 660 22326
rect 712 22311 728 22326
rect 780 22311 796 22326
rect 649 22277 660 22311
rect 727 22277 728 22311
rect 644 22274 660 22277
rect 712 22274 728 22277
rect 780 22274 796 22277
rect 848 22274 850 22326
rect 453 22262 850 22274
rect 453 22210 456 22262
rect 508 22210 524 22262
rect 576 22210 592 22262
rect 644 22238 660 22262
rect 712 22238 728 22262
rect 780 22238 796 22262
rect 649 22210 660 22238
rect 727 22210 728 22238
rect 848 22210 850 22262
rect 453 22204 459 22210
rect 493 22204 537 22210
rect 571 22204 615 22210
rect 649 22204 693 22210
rect 727 22204 771 22210
rect 805 22204 850 22210
rect 453 22198 850 22204
rect 453 22146 456 22198
rect 508 22146 524 22198
rect 576 22146 592 22198
rect 644 22165 660 22198
rect 712 22165 728 22198
rect 780 22165 796 22198
rect 649 22146 660 22165
rect 727 22146 728 22165
rect 848 22146 850 22198
rect 453 22134 459 22146
rect 493 22134 537 22146
rect 571 22134 615 22146
rect 649 22134 693 22146
rect 727 22134 771 22146
rect 805 22134 850 22146
rect 453 22082 456 22134
rect 508 22082 524 22134
rect 576 22082 592 22134
rect 649 22131 660 22134
rect 727 22131 728 22134
rect 644 22092 660 22131
rect 712 22092 728 22131
rect 780 22092 796 22131
rect 649 22082 660 22092
rect 727 22082 728 22092
rect 848 22082 850 22134
rect 453 22070 459 22082
rect 493 22070 537 22082
rect 571 22070 615 22082
rect 649 22070 693 22082
rect 727 22070 771 22082
rect 805 22070 850 22082
rect 453 22018 456 22070
rect 508 22018 524 22070
rect 576 22018 592 22070
rect 649 22058 660 22070
rect 727 22058 728 22070
rect 644 22019 660 22058
rect 712 22019 728 22058
rect 780 22019 796 22058
rect 649 22018 660 22019
rect 727 22018 728 22019
rect 848 22018 850 22070
rect 453 22006 459 22018
rect 493 22006 537 22018
rect 571 22006 615 22018
rect 649 22006 693 22018
rect 727 22006 771 22018
rect 805 22006 850 22018
rect 453 21954 456 22006
rect 508 21954 524 22006
rect 576 21954 592 22006
rect 649 21985 660 22006
rect 727 21985 728 22006
rect 644 21954 660 21985
rect 712 21954 728 21985
rect 780 21954 796 21985
rect 848 21954 850 22006
rect 453 21946 850 21954
rect 453 21942 459 21946
rect 493 21942 537 21946
rect 571 21942 615 21946
rect 649 21942 693 21946
rect 727 21942 771 21946
rect 805 21942 850 21946
rect 453 21890 456 21942
rect 508 21890 524 21942
rect 576 21890 592 21942
rect 649 21912 660 21942
rect 727 21912 728 21942
rect 644 21890 660 21912
rect 712 21890 728 21912
rect 780 21890 796 21912
rect 848 21890 850 21942
rect 453 21878 850 21890
rect 453 21826 456 21878
rect 508 21826 524 21878
rect 576 21826 592 21878
rect 644 21873 660 21878
rect 712 21873 728 21878
rect 780 21873 796 21878
rect 649 21839 660 21873
rect 727 21839 728 21873
rect 644 21826 660 21839
rect 712 21826 728 21839
rect 780 21826 796 21839
rect 848 21826 850 21878
rect 453 21814 850 21826
rect 453 21762 456 21814
rect 508 21762 524 21814
rect 576 21762 592 21814
rect 644 21800 660 21814
rect 712 21800 728 21814
rect 780 21800 796 21814
rect 649 21766 660 21800
rect 727 21766 728 21800
rect 644 21762 660 21766
rect 712 21762 728 21766
rect 780 21762 796 21766
rect 848 21762 850 21814
rect 453 21750 850 21762
rect 453 21698 456 21750
rect 508 21698 524 21750
rect 576 21698 592 21750
rect 644 21727 660 21750
rect 712 21727 728 21750
rect 780 21727 796 21750
rect 649 21698 660 21727
rect 727 21698 728 21727
rect 848 21698 850 21750
rect 453 21693 459 21698
rect 493 21693 537 21698
rect 571 21693 615 21698
rect 649 21693 693 21698
rect 727 21693 771 21698
rect 805 21693 850 21698
rect 453 21686 850 21693
rect 453 21634 456 21686
rect 508 21634 524 21686
rect 576 21634 592 21686
rect 644 21654 660 21686
rect 712 21654 728 21686
rect 780 21654 796 21686
rect 649 21634 660 21654
rect 727 21634 728 21654
rect 848 21634 850 21686
rect 453 21622 459 21634
rect 493 21622 537 21634
rect 571 21622 615 21634
rect 649 21622 693 21634
rect 727 21622 771 21634
rect 805 21622 850 21634
rect 453 21570 456 21622
rect 508 21570 524 21622
rect 576 21570 592 21622
rect 649 21620 660 21622
rect 727 21620 728 21622
rect 644 21581 660 21620
rect 712 21581 728 21620
rect 780 21581 796 21620
rect 649 21570 660 21581
rect 727 21570 728 21581
rect 848 21570 850 21622
rect 453 21558 459 21570
rect 493 21558 537 21570
rect 571 21558 615 21570
rect 649 21558 693 21570
rect 727 21558 771 21570
rect 805 21558 850 21570
rect 453 21506 456 21558
rect 508 21506 524 21558
rect 576 21506 592 21558
rect 649 21547 660 21558
rect 727 21547 728 21558
rect 644 21508 660 21547
rect 712 21508 728 21547
rect 780 21508 796 21547
rect 649 21506 660 21508
rect 727 21506 728 21508
rect 848 21506 850 21558
rect 453 21494 459 21506
rect 493 21494 537 21506
rect 571 21494 615 21506
rect 649 21494 693 21506
rect 727 21494 771 21506
rect 805 21494 850 21506
rect 453 21442 456 21494
rect 508 21442 524 21494
rect 576 21442 592 21494
rect 649 21474 660 21494
rect 727 21474 728 21494
rect 644 21442 660 21474
rect 712 21442 728 21474
rect 780 21442 796 21474
rect 848 21442 850 21494
rect 453 21435 850 21442
rect 453 21430 459 21435
rect 493 21430 537 21435
rect 571 21430 615 21435
rect 649 21430 693 21435
rect 727 21430 771 21435
rect 805 21430 850 21435
rect 453 21378 456 21430
rect 508 21378 524 21430
rect 576 21378 592 21430
rect 649 21401 660 21430
rect 727 21401 728 21430
rect 644 21378 660 21401
rect 712 21378 728 21401
rect 780 21378 796 21401
rect 848 21378 850 21430
rect 453 21366 850 21378
rect 453 21314 456 21366
rect 508 21314 524 21366
rect 576 21314 592 21366
rect 644 21362 660 21366
rect 712 21362 728 21366
rect 780 21362 796 21366
rect 649 21328 660 21362
rect 727 21328 728 21362
rect 644 21314 660 21328
rect 712 21314 728 21328
rect 780 21314 796 21328
rect 848 21314 850 21366
rect 453 21302 850 21314
rect 453 21250 456 21302
rect 508 21250 524 21302
rect 576 21250 592 21302
rect 644 21289 660 21302
rect 712 21289 728 21302
rect 780 21289 796 21302
rect 649 21255 660 21289
rect 727 21255 728 21289
rect 644 21250 660 21255
rect 712 21250 728 21255
rect 780 21250 796 21255
rect 848 21250 850 21302
rect 453 21238 850 21250
rect 453 21186 456 21238
rect 508 21186 524 21238
rect 576 21186 592 21238
rect 644 21216 660 21238
rect 712 21216 728 21238
rect 780 21216 796 21238
rect 649 21186 660 21216
rect 727 21186 728 21216
rect 848 21186 850 21238
rect 453 21182 459 21186
rect 493 21182 537 21186
rect 571 21182 615 21186
rect 649 21182 693 21186
rect 727 21182 771 21186
rect 805 21182 850 21186
rect 453 21174 850 21182
rect 453 21122 456 21174
rect 508 21122 524 21174
rect 576 21122 592 21174
rect 644 21143 660 21174
rect 712 21143 728 21174
rect 780 21143 796 21174
rect 649 21122 660 21143
rect 727 21122 728 21143
rect 848 21122 850 21174
rect 453 21110 459 21122
rect 493 21110 537 21122
rect 571 21110 615 21122
rect 649 21110 693 21122
rect 727 21110 771 21122
rect 805 21110 850 21122
rect 453 21058 456 21110
rect 508 21058 524 21110
rect 576 21058 592 21110
rect 649 21109 660 21110
rect 727 21109 728 21110
rect 644 21070 660 21109
rect 712 21070 728 21109
rect 780 21070 796 21109
rect 649 21058 660 21070
rect 727 21058 728 21070
rect 848 21058 850 21110
rect 453 21046 459 21058
rect 493 21046 537 21058
rect 571 21046 615 21058
rect 649 21046 693 21058
rect 727 21046 771 21058
rect 805 21046 850 21058
rect 453 20994 456 21046
rect 508 20994 524 21046
rect 576 20994 592 21046
rect 649 21036 660 21046
rect 727 21036 728 21046
rect 644 20997 660 21036
rect 712 20997 728 21036
rect 780 20997 796 21036
rect 649 20994 660 20997
rect 727 20994 728 20997
rect 848 20994 850 21046
rect 453 20982 459 20994
rect 493 20982 537 20994
rect 571 20982 615 20994
rect 649 20982 693 20994
rect 727 20982 771 20994
rect 805 20982 850 20994
rect 453 20930 456 20982
rect 508 20930 524 20982
rect 576 20930 592 20982
rect 649 20963 660 20982
rect 727 20963 728 20982
rect 644 20930 660 20963
rect 712 20930 728 20963
rect 780 20930 796 20963
rect 848 20930 850 20982
rect 453 20924 850 20930
rect 453 20918 459 20924
rect 493 20918 537 20924
rect 571 20918 615 20924
rect 649 20918 693 20924
rect 727 20918 771 20924
rect 805 20918 850 20924
rect 453 20866 456 20918
rect 508 20866 524 20918
rect 576 20866 592 20918
rect 649 20890 660 20918
rect 727 20890 728 20918
rect 644 20866 660 20890
rect 712 20866 728 20890
rect 780 20866 796 20890
rect 848 20866 850 20918
rect 453 20854 850 20866
rect 453 20802 456 20854
rect 508 20802 524 20854
rect 576 20802 592 20854
rect 644 20851 660 20854
rect 712 20851 728 20854
rect 780 20851 796 20854
rect 649 20817 660 20851
rect 727 20817 728 20851
rect 644 20802 660 20817
rect 712 20802 728 20817
rect 780 20802 796 20817
rect 848 20802 850 20854
rect 453 20790 850 20802
rect 453 20738 456 20790
rect 508 20738 524 20790
rect 576 20738 592 20790
rect 644 20778 660 20790
rect 712 20778 728 20790
rect 780 20778 796 20790
rect 649 20744 660 20778
rect 727 20744 728 20778
rect 644 20738 660 20744
rect 712 20738 728 20744
rect 780 20738 796 20744
rect 848 20738 850 20790
rect 453 20726 850 20738
rect 453 20674 456 20726
rect 508 20674 524 20726
rect 576 20674 592 20726
rect 644 20705 660 20726
rect 712 20705 728 20726
rect 780 20705 796 20726
rect 649 20674 660 20705
rect 727 20674 728 20705
rect 848 20674 850 20726
rect 453 20671 459 20674
rect 493 20671 537 20674
rect 571 20671 615 20674
rect 649 20671 693 20674
rect 727 20671 771 20674
rect 805 20671 850 20674
rect 453 20662 850 20671
rect 453 20610 456 20662
rect 508 20610 524 20662
rect 576 20610 592 20662
rect 644 20632 660 20662
rect 712 20632 728 20662
rect 780 20632 796 20662
rect 649 20610 660 20632
rect 727 20610 728 20632
rect 848 20610 850 20662
rect 453 20598 459 20610
rect 493 20598 537 20610
rect 571 20598 615 20610
rect 649 20598 693 20610
rect 727 20598 771 20610
rect 805 20598 850 20610
rect 453 20546 456 20598
rect 508 20546 524 20598
rect 576 20546 592 20598
rect 644 20559 660 20598
rect 712 20559 728 20598
rect 780 20559 796 20598
rect 649 20546 660 20559
rect 727 20546 728 20559
rect 848 20546 850 20598
rect 453 20534 459 20546
rect 493 20534 537 20546
rect 571 20534 615 20546
rect 649 20534 693 20546
rect 727 20534 771 20546
rect 805 20534 850 20546
rect 453 20482 456 20534
rect 508 20482 524 20534
rect 576 20482 592 20534
rect 649 20525 660 20534
rect 727 20525 728 20534
rect 644 20486 660 20525
rect 712 20486 728 20525
rect 780 20486 796 20525
rect 848 20513 850 20534
rect 940 20513 971 25263
rect 649 20482 660 20486
rect 727 20482 728 20486
rect 848 20482 971 20513
rect 453 20470 459 20482
rect 493 20470 537 20482
rect 571 20470 615 20482
rect 649 20470 693 20482
rect 727 20470 771 20482
rect 805 20470 971 20482
rect 453 20418 456 20470
rect 508 20418 524 20470
rect 576 20418 592 20470
rect 649 20452 660 20470
rect 727 20452 728 20470
rect 644 20418 660 20452
rect 712 20418 728 20452
rect 780 20418 796 20452
rect 848 20418 971 20470
rect 453 20413 868 20418
rect 453 20406 459 20413
rect 493 20406 537 20413
rect 571 20406 615 20413
rect 649 20406 693 20413
rect 727 20406 771 20413
rect 805 20406 868 20413
rect 453 20354 456 20406
rect 508 20354 524 20406
rect 576 20354 592 20406
rect 649 20379 660 20406
rect 727 20379 728 20406
rect 848 20384 868 20406
rect 902 20384 971 20418
rect 2778 20519 2784 20571
rect 2836 20519 2853 20571
rect 2905 20519 2922 20571
rect 2974 20519 2991 20571
rect 3043 20519 3060 20571
rect 3112 20519 3128 20571
rect 3180 20519 3196 20571
rect 3248 20519 3264 20571
rect 3316 20519 3332 20571
rect 3384 20519 3400 20571
rect 3452 20519 3468 20571
rect 3520 20519 3536 20571
rect 3588 20519 3604 20571
rect 3656 20519 3672 20571
rect 3724 20519 3730 20571
rect 2778 20459 3730 20519
rect 2778 20407 2784 20459
rect 2836 20407 2853 20459
rect 2905 20407 2922 20459
rect 2974 20407 2991 20459
rect 3043 20407 3060 20459
rect 3112 20407 3128 20459
rect 3180 20407 3196 20459
rect 3248 20407 3264 20459
rect 3316 20407 3332 20459
rect 3384 20407 3400 20459
rect 3452 20407 3468 20459
rect 3520 20407 3536 20459
rect 3588 20407 3604 20459
rect 3656 20407 3672 20459
rect 3724 20407 3730 20459
rect 12199 20566 12251 20572
rect 12199 20496 12251 20514
rect 12199 20425 12251 20444
rect 644 20354 660 20379
rect 712 20354 728 20379
rect 780 20354 796 20379
rect 848 20354 971 20384
rect 453 20343 971 20354
rect 453 20342 868 20343
rect 453 20290 456 20342
rect 508 20290 524 20342
rect 576 20290 592 20342
rect 644 20340 660 20342
rect 712 20340 728 20342
rect 780 20340 796 20342
rect 649 20306 660 20340
rect 727 20306 728 20340
rect 848 20309 868 20342
rect 902 20309 971 20343
rect 644 20290 660 20306
rect 712 20290 728 20306
rect 780 20290 796 20306
rect 848 20290 971 20309
rect 453 20277 971 20290
rect 453 20225 456 20277
rect 508 20225 524 20277
rect 576 20225 592 20277
rect 644 20267 660 20277
rect 712 20267 728 20277
rect 780 20267 796 20277
rect 848 20268 971 20277
rect 649 20233 660 20267
rect 727 20233 728 20267
rect 848 20234 868 20268
rect 902 20234 971 20268
rect 644 20225 660 20233
rect 712 20225 728 20233
rect 780 20225 796 20233
rect 848 20225 971 20234
rect 12199 20354 12251 20373
rect 12199 20283 12251 20302
rect 12199 20225 12251 20231
rect 453 20212 971 20225
rect 453 20160 456 20212
rect 508 20160 524 20212
rect 576 20160 592 20212
rect 644 20194 660 20212
rect 712 20194 728 20212
rect 780 20194 796 20212
rect 649 20160 660 20194
rect 727 20160 728 20194
rect 848 20193 971 20212
rect 848 20160 868 20193
rect 453 20159 868 20160
rect 902 20159 971 20193
rect 453 20147 971 20159
rect 453 20095 456 20147
rect 508 20095 524 20147
rect 576 20095 592 20147
rect 644 20121 660 20147
rect 712 20121 728 20147
rect 780 20121 796 20147
rect 649 20095 660 20121
rect 727 20095 728 20121
rect 848 20117 971 20147
rect 848 20095 868 20117
rect 453 20087 459 20095
rect 493 20087 537 20095
rect 571 20087 615 20095
rect 649 20087 693 20095
rect 727 20087 771 20095
rect 805 20087 868 20095
rect 453 20083 868 20087
rect 902 20083 971 20117
rect 453 20082 971 20083
rect 453 20030 456 20082
rect 508 20030 524 20082
rect 576 20030 592 20082
rect 644 20048 660 20082
rect 712 20048 728 20082
rect 780 20048 796 20082
rect 649 20030 660 20048
rect 727 20030 728 20048
rect 848 20041 971 20082
rect 848 20030 868 20041
rect 453 20017 459 20030
rect 493 20017 537 20030
rect 571 20017 615 20030
rect 649 20017 693 20030
rect 727 20017 771 20030
rect 805 20017 868 20030
rect 453 19965 456 20017
rect 508 19965 524 20017
rect 576 19965 592 20017
rect 649 20014 660 20017
rect 727 20014 728 20017
rect 644 19975 660 20014
rect 712 19975 728 20014
rect 780 19975 796 20014
rect 848 20007 868 20017
rect 902 20007 971 20041
rect 649 19965 660 19975
rect 727 19965 728 19975
rect 848 19965 971 20007
rect 453 19952 459 19965
rect 493 19952 537 19965
rect 571 19952 615 19965
rect 649 19952 693 19965
rect 727 19952 771 19965
rect 805 19952 868 19965
rect 453 19900 456 19952
rect 508 19900 524 19952
rect 576 19900 592 19952
rect 649 19941 660 19952
rect 727 19941 728 19952
rect 644 19902 660 19941
rect 712 19902 728 19941
rect 780 19902 796 19941
rect 848 19931 868 19952
rect 902 19931 971 19965
rect 649 19900 660 19902
rect 727 19900 728 19902
rect 848 19900 971 19931
rect 453 19887 459 19900
rect 493 19887 537 19900
rect 571 19887 615 19900
rect 649 19887 693 19900
rect 727 19887 771 19900
rect 805 19889 971 19900
rect 805 19887 868 19889
rect 453 19835 456 19887
rect 508 19835 524 19887
rect 576 19835 592 19887
rect 649 19868 660 19887
rect 727 19868 728 19887
rect 644 19835 660 19868
rect 712 19835 728 19868
rect 780 19835 796 19868
rect 848 19855 868 19887
rect 902 19855 971 19889
rect 848 19835 971 19855
rect 453 19829 971 19835
rect 453 19822 459 19829
rect 493 19822 537 19829
rect 571 19822 615 19829
rect 649 19822 693 19829
rect 727 19822 771 19829
rect 805 19822 971 19829
rect 453 19770 456 19822
rect 508 19770 524 19822
rect 576 19770 592 19822
rect 649 19795 660 19822
rect 727 19795 728 19822
rect 848 19813 971 19822
rect 644 19770 660 19795
rect 712 19770 728 19795
rect 780 19770 796 19795
rect 848 19779 868 19813
rect 902 19779 971 19813
rect 848 19770 971 19779
rect 453 19757 971 19770
rect 453 19705 456 19757
rect 508 19705 524 19757
rect 576 19705 592 19757
rect 644 19756 660 19757
rect 712 19756 728 19757
rect 780 19756 796 19757
rect 649 19722 660 19756
rect 727 19722 728 19756
rect 848 19737 971 19757
rect 644 19705 660 19722
rect 712 19705 728 19722
rect 780 19705 796 19722
rect 848 19705 868 19737
rect 453 19703 868 19705
rect 902 19703 971 19737
rect 453 19692 971 19703
rect 453 19640 456 19692
rect 508 19640 524 19692
rect 576 19640 592 19692
rect 644 19683 660 19692
rect 712 19683 728 19692
rect 780 19683 796 19692
rect 649 19649 660 19683
rect 727 19649 728 19683
rect 848 19661 971 19692
rect 12199 20110 12251 20116
rect 12199 20046 12251 20058
rect 12199 19982 12251 19994
rect 12199 19918 12251 19930
rect 12199 19854 12251 19866
rect 12199 19790 12251 19802
rect 12199 19725 12251 19738
rect 12199 19667 12251 19673
rect 644 19640 660 19649
rect 712 19640 728 19649
rect 780 19640 796 19649
rect 848 19640 868 19661
rect 453 19627 868 19640
rect 902 19627 971 19661
rect 453 19575 456 19627
rect 508 19575 524 19627
rect 576 19575 592 19627
rect 644 19610 660 19627
rect 712 19610 728 19627
rect 780 19610 796 19627
rect 649 19576 660 19610
rect 727 19576 728 19610
rect 848 19585 971 19627
rect 644 19575 660 19576
rect 712 19575 728 19576
rect 780 19575 796 19576
rect 848 19575 868 19585
rect 453 19562 868 19575
rect 453 19510 456 19562
rect 508 19510 524 19562
rect 576 19510 592 19562
rect 644 19537 660 19562
rect 712 19537 728 19562
rect 780 19537 796 19562
rect 848 19551 868 19562
rect 902 19551 971 19585
rect 649 19510 660 19537
rect 727 19510 728 19537
rect 848 19510 971 19551
rect 453 19503 459 19510
rect 493 19503 537 19510
rect 571 19503 615 19510
rect 649 19503 693 19510
rect 727 19503 771 19510
rect 805 19509 971 19510
rect 805 19503 868 19509
rect 453 19497 868 19503
rect 453 19445 456 19497
rect 508 19445 524 19497
rect 576 19445 592 19497
rect 644 19464 660 19497
rect 712 19464 728 19497
rect 780 19464 796 19497
rect 848 19475 868 19497
rect 902 19475 971 19509
rect 649 19445 660 19464
rect 727 19445 728 19464
rect 848 19445 971 19475
rect 453 19432 459 19445
rect 493 19432 537 19445
rect 571 19432 615 19445
rect 649 19432 693 19445
rect 727 19432 771 19445
rect 805 19433 971 19445
rect 805 19432 868 19433
rect 453 19380 456 19432
rect 508 19380 524 19432
rect 576 19380 592 19432
rect 649 19430 660 19432
rect 727 19430 728 19432
rect 644 19391 660 19430
rect 712 19391 728 19430
rect 780 19391 796 19430
rect 848 19399 868 19432
rect 902 19399 971 19433
rect 649 19380 660 19391
rect 727 19380 728 19391
rect 848 19380 971 19399
rect 453 19367 459 19380
rect 493 19367 537 19380
rect 571 19367 615 19380
rect 649 19367 693 19380
rect 727 19367 771 19380
rect 805 19367 971 19380
rect 453 19315 456 19367
rect 508 19315 524 19367
rect 576 19315 592 19367
rect 649 19357 660 19367
rect 727 19357 728 19367
rect 848 19357 971 19367
rect 644 19318 660 19357
rect 712 19318 728 19357
rect 780 19318 796 19357
rect 848 19323 868 19357
rect 902 19323 971 19357
rect 649 19315 660 19318
rect 727 19315 728 19318
rect 848 19315 971 19323
rect 453 19302 459 19315
rect 493 19302 537 19315
rect 571 19302 615 19315
rect 649 19302 693 19315
rect 727 19302 771 19315
rect 805 19302 971 19315
rect 453 19250 456 19302
rect 508 19250 524 19302
rect 576 19250 592 19302
rect 649 19284 660 19302
rect 727 19284 728 19302
rect 644 19250 660 19284
rect 712 19250 728 19284
rect 780 19250 796 19284
rect 848 19281 971 19302
rect 848 19250 868 19281
rect 453 19247 868 19250
rect 902 19247 971 19281
rect 453 19245 971 19247
rect 453 19237 459 19245
rect 493 19237 537 19245
rect 571 19237 615 19245
rect 649 19237 693 19245
rect 727 19237 771 19245
rect 805 19237 971 19245
rect 453 19185 456 19237
rect 508 19185 524 19237
rect 576 19185 592 19237
rect 649 19211 660 19237
rect 727 19211 728 19237
rect 644 19185 660 19211
rect 712 19185 728 19211
rect 780 19185 796 19211
rect 848 19185 971 19237
tri 2775 19191 2781 19197 ne
rect 2781 19191 2787 19243
rect 2839 19191 2854 19243
rect 2906 19191 2921 19243
rect 2973 19191 2988 19243
rect 3040 19191 3055 19243
rect 3107 19191 3122 19243
rect 3174 19191 3189 19243
rect 3241 19191 3256 19243
rect 3308 19191 3323 19243
rect 3375 19191 3390 19243
rect 3442 19191 3456 19243
rect 3508 19191 3522 19243
rect 3574 19191 3588 19243
rect 3640 19191 3654 19243
rect 3706 19191 3720 19243
rect 3772 19191 3778 19243
tri 3778 19191 3784 19197 nw
rect 453 19180 971 19185
rect 453 19153 1794 19180
rect 453 19119 472 19153
rect 506 19119 545 19153
rect 579 19119 618 19153
rect 652 19119 691 19153
rect 725 19119 764 19153
rect 798 19119 837 19153
rect 871 19119 910 19153
rect 944 19119 983 19153
rect 1017 19119 1056 19153
rect 1090 19119 1129 19153
rect 1163 19119 1202 19153
rect 1236 19119 1275 19153
rect 1309 19119 1348 19153
rect 1382 19119 1420 19153
rect 1454 19119 1492 19153
rect 1526 19119 1564 19153
rect 1598 19119 1636 19153
rect 1670 19119 1708 19153
rect 1742 19119 1794 19153
rect 453 19063 1794 19119
tri 3010 19063 3016 19069 se
rect 453 19029 472 19063
rect 506 19029 545 19063
rect 579 19029 618 19063
rect 652 19029 691 19063
rect 725 19029 764 19063
rect 798 19029 837 19063
rect 871 19029 910 19063
rect 944 19029 983 19063
rect 1017 19029 1056 19063
rect 1090 19029 1129 19063
rect 1163 19029 1202 19063
rect 1236 19029 1275 19063
rect 1309 19029 1348 19063
rect 1382 19029 1420 19063
rect 1454 19029 1492 19063
rect 1526 19029 1564 19063
rect 1598 19029 1636 19063
rect 1670 19029 1708 19063
rect 1742 19029 1794 19063
rect 453 19022 1794 19029
tri 1596 18876 1742 19022 ne
rect 1742 18876 1794 19022
rect 3016 19017 3022 19069
rect 3074 19017 3092 19069
rect 3144 19017 3162 19069
rect 3214 19017 3232 19069
rect 3284 19017 3302 19069
rect 3354 19017 3372 19069
rect 3424 19017 3442 19069
rect 3494 19017 3512 19069
rect 3564 19017 3582 19069
rect 3634 19017 3651 19069
rect 3703 19017 3720 19069
rect 3772 19017 3778 19069
tri 3778 19063 3784 19069 sw
rect 270 18824 276 18876
rect 328 18824 341 18876
rect 393 18824 406 18876
rect 458 18824 471 18876
rect 523 18824 536 18876
rect 588 18824 601 18876
rect 653 18824 666 18876
rect 718 18824 1257 18876
rect 1309 18824 1325 18876
rect 1377 18824 1393 18876
rect 1445 18824 1461 18876
rect 1513 18824 1528 18876
rect 1580 18824 1595 18876
rect 1647 18824 1653 18876
tri 1742 18824 1794 18876 ne
rect 270 18794 1653 18824
rect 270 18742 276 18794
rect 328 18742 341 18794
rect 393 18742 406 18794
rect 458 18742 471 18794
rect 523 18742 536 18794
rect 588 18742 601 18794
rect 653 18742 666 18794
rect 718 18742 1257 18794
rect 1309 18742 1325 18794
rect 1377 18742 1393 18794
rect 1445 18742 1461 18794
rect 1513 18742 1528 18794
rect 1580 18742 1595 18794
rect 1647 18742 1653 18794
rect 270 18712 1653 18742
rect 270 18660 276 18712
rect 328 18660 341 18712
rect 393 18660 406 18712
rect 458 18660 471 18712
rect 523 18660 536 18712
rect 588 18660 601 18712
rect 653 18660 666 18712
rect 718 18660 1257 18712
rect 1309 18660 1325 18712
rect 1377 18660 1393 18712
rect 1445 18660 1461 18712
rect 1513 18660 1528 18712
rect 1580 18660 1595 18712
rect 1647 18660 1653 18712
tri 1578 18174 1788 18384 se
rect 1578 18158 1788 18174
rect 1578 17908 1584 18158
rect 1762 17908 1788 18158
rect 1578 17869 1788 17908
rect 1578 17835 1584 17869
rect 1618 17835 1656 17869
rect 1690 17835 1728 17869
rect 1762 17835 1788 17869
rect 1578 17793 1788 17835
tri 1578 17583 1788 17793 ne
tri 3192 17343 3198 17349 se
rect 3198 17297 3204 17349
rect 3256 17297 3296 17349
rect 3348 17297 3354 17349
tri 3354 17343 3360 17349 sw
rect 5731 16777 9142 16802
rect 5731 16725 5737 16777
rect 5789 16725 5802 16777
rect 5854 16725 5867 16777
rect 5919 16725 5932 16777
rect 5984 16725 5997 16777
rect 6049 16725 6062 16777
rect 6114 16725 6127 16777
rect 6179 16725 6192 16777
rect 6244 16725 6257 16777
rect 6309 16725 6322 16777
rect 6374 16725 6387 16777
rect 6439 16725 6452 16777
rect 6504 16725 6517 16777
rect 6569 16725 6582 16777
rect 6634 16725 6647 16777
rect 6699 16725 6712 16777
rect 6764 16725 6777 16777
rect 6829 16725 6842 16777
rect 6894 16725 6907 16777
rect 6959 16725 6972 16777
rect 7024 16725 7036 16777
rect 7088 16725 7100 16777
rect 7152 16725 7164 16777
rect 7216 16725 7228 16777
rect 7280 16725 7292 16777
rect 7344 16725 7356 16777
rect 7408 16725 7420 16777
rect 7472 16725 7484 16777
rect 7536 16725 7548 16777
rect 7600 16725 7612 16777
rect 7664 16725 7676 16777
rect 7728 16725 7740 16777
rect 7792 16725 7804 16777
rect 7856 16725 7868 16777
rect 7920 16725 7932 16777
rect 7984 16725 7996 16777
rect 8048 16725 8060 16777
rect 8112 16725 8124 16777
rect 8176 16725 8188 16777
rect 8240 16725 8252 16777
rect 8304 16725 8316 16777
rect 8368 16725 8380 16777
rect 8432 16725 8444 16777
rect 8496 16725 8508 16777
rect 8560 16725 8572 16777
rect 8624 16725 8636 16777
rect 8688 16725 8700 16777
rect 8752 16725 8764 16777
rect 8816 16725 8828 16777
rect 8880 16725 8892 16777
rect 8944 16725 8956 16777
rect 9008 16725 9020 16777
rect 9072 16725 9084 16777
rect 9136 16725 9142 16777
rect 5731 16700 9142 16725
rect 7396 16154 7660 16155
rect 7396 16102 7402 16154
rect 7454 16102 7469 16154
rect 7521 16102 7536 16154
rect 7588 16102 7602 16154
rect 7654 16102 7660 16154
rect 7396 16082 7660 16102
rect 7396 16030 7402 16082
rect 7454 16030 7469 16082
rect 7521 16030 7536 16082
rect 7588 16030 7602 16082
rect 7654 16030 7660 16082
rect 7396 16010 7660 16030
rect 7396 15958 7402 16010
rect 7454 15958 7469 16010
rect 7521 15958 7536 16010
rect 7588 15958 7602 16010
rect 7654 15958 7660 16010
rect 7396 15957 7660 15958
rect 9190 16154 9292 16155
rect 9190 16102 9196 16154
rect 9248 16102 9292 16154
rect 9190 16082 9292 16102
rect 9190 16030 9196 16082
rect 9248 16030 9292 16082
rect 9190 16010 9292 16030
rect 9190 15958 9196 16010
rect 9248 15958 9292 16010
rect 9190 15957 9292 15958
tri 1839 15509 1873 15543 sw
rect 1403 15457 1590 15509
rect 1642 15457 1654 15509
rect 1706 15457 1894 15509
rect 5523 13889 5946 13895
rect 5523 13855 5535 13889
rect 5569 13855 5608 13889
rect 5642 13855 5681 13889
rect 5715 13855 5754 13889
rect 5788 13865 5827 13889
rect 5861 13865 5900 13889
rect 5788 13855 5816 13865
rect 5868 13855 5900 13865
rect 5934 13855 5946 13889
rect 5523 13813 5816 13855
rect 5868 13813 5946 13855
rect 5523 13801 5946 13813
rect 5523 13781 5816 13801
rect 5868 13781 5946 13801
rect 5523 13747 5535 13781
rect 5569 13747 5608 13781
rect 5642 13747 5681 13781
rect 5715 13747 5754 13781
rect 5788 13749 5816 13781
rect 5868 13749 5900 13781
rect 5788 13747 5827 13749
rect 5861 13747 5900 13749
rect 5934 13747 5946 13781
rect 5523 13741 5946 13747
rect 9477 13574 9529 13580
rect 5293 13563 5946 13569
rect 5293 13529 5305 13563
rect 5339 13529 5380 13563
rect 5414 13529 5455 13563
rect 5489 13529 5530 13563
rect 5564 13529 5604 13563
rect 5638 13529 5678 13563
rect 5712 13529 5752 13563
rect 5786 13562 5826 13563
rect 5860 13562 5900 13563
rect 5786 13529 5816 13562
rect 5868 13529 5900 13562
rect 5934 13529 5946 13563
rect 5293 13510 5816 13529
rect 5868 13510 5946 13529
rect 5293 13498 5946 13510
rect 5293 13455 5816 13498
rect 5868 13455 5946 13498
rect 5293 13421 5305 13455
rect 5339 13421 5380 13455
rect 5414 13421 5455 13455
rect 5489 13421 5530 13455
rect 5564 13421 5604 13455
rect 5638 13421 5678 13455
rect 5712 13421 5752 13455
rect 5786 13446 5816 13455
rect 5868 13446 5900 13455
rect 5786 13421 5826 13446
rect 5860 13421 5900 13446
rect 5934 13421 5946 13455
rect 6025 13554 6199 13560
rect 6077 13514 6199 13554
tri 9529 13558 9551 13580 sw
rect 9529 13522 9671 13558
rect 6025 13490 6077 13502
rect 6025 13432 6077 13438
tri 6077 13432 6159 13514 nw
rect 9477 13512 9671 13522
rect 9477 13510 9529 13512
tri 9529 13478 9563 13512 nw
rect 9477 13452 9529 13458
rect 5293 13415 5946 13421
rect 9359 13059 9411 13065
rect 9359 12995 9411 13007
rect 7533 12945 7585 12951
rect 5486 12910 5875 12916
rect 5486 12876 5498 12910
rect 5532 12876 5581 12910
rect 5615 12876 5664 12910
rect 5698 12876 5747 12910
rect 5781 12876 5816 12910
rect 5486 12858 5816 12876
rect 5868 12858 5875 12910
rect 5486 12846 5875 12858
rect 5486 12828 5816 12846
rect 5486 12794 5498 12828
rect 5532 12794 5581 12828
rect 5615 12794 5664 12828
rect 5698 12794 5747 12828
rect 5781 12794 5816 12828
rect 5868 12794 5875 12846
rect 9359 12935 9411 12943
tri 9411 12935 9413 12937 sw
rect 9359 12923 9413 12935
tri 9359 12919 9363 12923 ne
rect 9363 12919 9413 12923
tri 9413 12919 9429 12935 sw
rect 7533 12885 7585 12893
tri 7585 12885 7619 12919 sw
tri 9363 12885 9397 12919 ne
rect 9397 12885 9429 12919
tri 9429 12885 9463 12919 sw
rect 7533 12881 7739 12885
rect 7585 12839 7739 12881
tri 9397 12869 9413 12885 ne
rect 9413 12869 9463 12885
tri 9463 12869 9479 12885 sw
tri 9413 12839 9443 12869 ne
rect 9443 12839 9667 12869
rect 7533 12823 7585 12829
tri 7585 12823 7601 12839 nw
tri 9443 12823 9459 12839 ne
rect 9459 12823 9667 12839
rect 5486 12788 5875 12794
tri 5278 12278 5381 12381 se
rect 5381 12288 6267 12381
rect 5381 12278 5394 12288
tri 5394 12278 5404 12288 nw
tri 6155 12278 6165 12288 ne
rect 6165 12278 6267 12288
rect 4715 12272 4767 12278
rect 4715 12208 4767 12220
rect 4715 12150 4767 12156
rect 5163 12272 5266 12278
rect 5215 12220 5266 12272
rect 5163 12208 5266 12220
rect 5215 12156 5266 12208
rect 5163 12150 5266 12156
tri 5266 12150 5394 12278 nw
tri 6165 12176 6267 12278 ne
rect 5172 12025 5633 12037
rect 5172 11991 5186 12025
rect 5220 11991 5266 12025
rect 5300 11991 5346 12025
rect 5380 11991 5426 12025
rect 5460 11991 5506 12025
rect 5540 11991 5586 12025
rect 5620 11991 5633 12025
rect 5172 11954 5633 11991
tri 5633 11954 5716 12037 sw
rect 5172 11942 5716 11954
rect 5172 11939 5668 11942
rect 5172 11905 5186 11939
rect 5220 11905 5266 11939
rect 5300 11905 5346 11939
rect 5380 11905 5426 11939
rect 5460 11905 5506 11939
rect 5540 11905 5586 11939
rect 5620 11908 5668 11939
rect 5702 11910 5716 11942
tri 5716 11910 5760 11954 sw
rect 5702 11908 5760 11910
rect 5620 11905 5760 11908
rect 5172 11904 5760 11905
rect 5172 11870 5705 11904
rect 5172 11853 5668 11870
rect 5172 11819 5186 11853
rect 5220 11819 5266 11853
rect 5300 11819 5346 11853
rect 5380 11819 5426 11853
rect 5460 11819 5506 11853
rect 5540 11819 5586 11853
rect 5620 11836 5668 11853
rect 5702 11852 5705 11870
rect 5757 11852 5760 11904
rect 5702 11836 5760 11852
rect 5620 11834 5760 11836
rect 5620 11819 5705 11834
rect 5172 11782 5705 11819
rect 5757 11782 5760 11834
rect 5172 11779 5760 11782
tri 5760 11779 5891 11910 sw
rect 5172 11773 5891 11779
rect 5172 11739 5187 11773
rect 5221 11739 5260 11773
rect 5294 11739 5333 11773
rect 5367 11739 5406 11773
rect 5440 11739 5479 11773
rect 5513 11739 5552 11773
rect 5586 11739 5624 11773
rect 5658 11739 5696 11773
rect 5730 11764 5768 11773
rect 5757 11739 5768 11764
rect 5802 11739 5840 11773
rect 5874 11739 5891 11773
rect 5172 11712 5705 11739
rect 5757 11712 5891 11739
rect 5172 11699 5891 11712
rect 5172 11665 5187 11699
rect 5221 11665 5260 11699
rect 5294 11665 5333 11699
rect 5367 11665 5406 11699
rect 5440 11665 5479 11699
rect 5513 11665 5552 11699
rect 5586 11665 5624 11699
rect 5658 11665 5696 11699
rect 5730 11694 5768 11699
rect 5757 11665 5768 11694
rect 5802 11665 5840 11699
rect 5874 11665 5891 11699
tri 2838 11625 2839 11626 se
rect 2839 11625 2845 11662
tri 2823 11610 2838 11625 se
rect 2838 11610 2845 11625
rect 2897 11610 2909 11662
rect 2961 11634 2967 11662
rect 5172 11642 5705 11665
rect 5757 11642 5891 11665
rect 2961 11627 2984 11634
tri 2984 11627 2991 11634 nw
rect 5172 11627 5891 11642
tri 5891 11627 6043 11779 sw
rect 7657 11695 7663 11747
rect 7715 11695 7727 11747
rect 7779 11695 7952 11747
rect 8004 11695 8016 11747
rect 8068 11695 8074 11747
rect 2961 11625 2982 11627
tri 2982 11625 2984 11627 nw
rect 5172 11625 6043 11627
rect 2961 11610 2967 11625
tri 2967 11610 2982 11625 nw
rect 5172 11591 5187 11625
rect 5221 11591 5260 11625
rect 5294 11591 5333 11625
rect 5367 11591 5406 11625
rect 5440 11591 5479 11625
rect 5513 11591 5552 11625
rect 5586 11591 5624 11625
rect 5658 11591 5696 11625
rect 5730 11624 5768 11625
rect 5757 11591 5768 11624
rect 5802 11591 5840 11625
rect 5874 11610 6043 11625
tri 6043 11610 6060 11627 sw
rect 5874 11591 6060 11610
rect 5172 11572 5705 11591
rect 5757 11572 6060 11591
rect 5172 11556 6060 11572
tri 6060 11556 6114 11610 sw
rect 5172 11553 6267 11556
rect 5172 11551 5705 11553
rect 5757 11551 6267 11553
rect 5172 11517 5187 11551
rect 5221 11517 5260 11551
rect 5294 11517 5333 11551
rect 5367 11517 5406 11551
rect 5440 11517 5479 11551
rect 5513 11517 5552 11551
rect 5586 11517 5624 11551
rect 5658 11517 5696 11551
rect 5757 11517 5768 11551
rect 5802 11517 5840 11551
rect 5874 11517 6267 11551
rect 5172 11511 5705 11517
tri 5614 11457 5668 11511 ne
rect 5668 11501 5705 11511
rect 5757 11501 6267 11517
rect 5668 11482 6267 11501
rect 5668 11457 5705 11482
tri 5668 11424 5701 11457 ne
rect 5701 11430 5705 11457
rect 5757 11457 6267 11482
rect 5757 11430 5807 11457
rect 5701 11424 5807 11430
tri 5701 11351 5774 11424 ne
rect 5774 11351 5807 11424
rect 5913 11351 6267 11457
tri 5774 11341 5784 11351 ne
rect 5784 11341 6267 11351
rect 2994 10333 3000 10385
rect 3052 10333 3065 10385
rect 3117 10333 3130 10385
rect 3182 10333 3194 10385
rect 3246 10333 3258 10385
rect 3310 10333 3322 10385
rect 3374 10333 3386 10385
rect 3438 10333 3450 10385
rect 3502 10333 3514 10385
rect 3566 10333 3578 10385
rect 3630 10333 3642 10385
rect 3694 10333 3706 10385
rect 3758 10333 3764 10385
rect 2994 10309 3764 10333
rect 2994 10257 3000 10309
rect 3052 10257 3065 10309
rect 3117 10257 3130 10309
rect 3182 10257 3194 10309
rect 3246 10257 3258 10309
rect 3310 10257 3322 10309
rect 3374 10257 3386 10309
rect 3438 10257 3450 10309
rect 3502 10257 3514 10309
rect 3566 10257 3578 10309
rect 3630 10257 3642 10309
rect 3694 10257 3706 10309
rect 3758 10257 3764 10309
tri 9362 10257 9406 10301 sw
rect 11001 10281 11007 10333
rect 11059 10281 11081 10333
rect 11133 10281 11155 10333
rect 11207 10281 11229 10333
rect 11281 10281 11287 10333
rect 11001 10269 11287 10281
tri 9297 10244 9310 10257 se
rect 7400 10192 7406 10244
rect 7458 10192 7487 10244
rect 7539 10192 7567 10244
rect 7619 10192 7625 10244
tri 9296 10243 9297 10244 se
rect 9297 10243 9310 10244
rect 9362 10243 9406 10257
tri 9406 10243 9420 10257 sw
rect 9362 10239 9420 10243
tri 9420 10239 9424 10243 sw
rect 11001 10217 11007 10269
rect 11059 10217 11081 10269
rect 11133 10217 11155 10269
rect 11207 10217 11229 10269
rect 11281 10217 11287 10269
rect 11001 10205 11287 10217
rect 11001 10153 11007 10205
rect 11059 10153 11081 10205
rect 11133 10153 11155 10205
rect 11207 10153 11229 10205
rect 11281 10153 11287 10205
rect 3987 10079 3993 10131
rect 4045 10079 4057 10131
rect 4109 10079 4115 10131
rect 4540 10079 4546 10131
rect 4598 10079 4610 10131
rect 4662 10123 4668 10131
tri 4668 10123 4676 10131 sw
tri 6887 10123 6891 10127 se
rect 6891 10123 6897 10131
rect 4662 10113 5721 10123
tri 5721 10113 5731 10123 sw
tri 5904 10113 5914 10123 se
rect 5914 10113 6897 10123
rect 4662 10085 6897 10113
rect 4662 10079 6609 10085
tri 6609 10079 6615 10085 nw
tri 6885 10079 6891 10085 ne
rect 6891 10079 6897 10085
rect 6949 10079 6961 10131
rect 7013 10079 7019 10131
rect 2225 9999 2231 10051
rect 2283 9999 2299 10051
rect 2351 9999 2367 10051
rect 2419 9999 2435 10051
rect 2487 9999 2503 10051
rect 2555 9999 2571 10051
rect 2623 9999 2638 10051
rect 2690 9999 2696 10051
rect 2225 9977 2696 9999
rect 2225 9925 2231 9977
rect 2283 9925 2299 9977
rect 2351 9925 2367 9977
rect 2419 9925 2435 9977
rect 2487 9925 2503 9977
rect 2555 9925 2571 9977
rect 2623 9925 2638 9977
rect 2690 9925 2696 9977
rect 2225 9903 2696 9925
rect 2225 9851 2231 9903
rect 2283 9851 2299 9903
rect 2351 9851 2367 9903
rect 2419 9851 2435 9903
rect 2487 9851 2503 9903
rect 2555 9851 2571 9903
rect 2623 9851 2638 9903
rect 2690 9851 2696 9903
rect 6943 9977 6995 9983
rect 7214 9976 7220 10028
rect 7272 9976 7284 10028
rect 7336 9976 7822 10028
rect 7874 9976 7886 10028
rect 7938 9976 7944 10028
rect 6943 9913 6995 9925
tri 6995 9907 7029 9941 sw
rect 6995 9861 9654 9907
rect 6943 9855 9654 9861
rect 9706 9855 9718 9907
rect 9770 9855 9776 9907
rect 2225 9829 2696 9851
rect 2225 9777 2231 9829
rect 2283 9777 2299 9829
rect 2351 9777 2367 9829
rect 2419 9777 2435 9829
rect 2487 9777 2503 9829
rect 2555 9777 2571 9829
rect 2623 9777 2638 9829
rect 2690 9777 2696 9829
rect 2225 9755 2696 9777
rect 2225 9703 2231 9755
rect 2283 9703 2299 9755
rect 2351 9703 2367 9755
rect 2419 9703 2435 9755
rect 2487 9703 2503 9755
rect 2555 9703 2571 9755
rect 2623 9703 2638 9755
rect 2690 9703 2696 9755
rect 7403 9635 7625 9666
rect 7403 9583 7409 9635
rect 7461 9583 7488 9635
rect 7540 9583 7567 9635
rect 7619 9583 7625 9635
rect 7403 9552 7625 9583
rect 7403 9543 7517 9549
rect 7403 9491 7434 9543
rect 7486 9491 7517 9543
rect 7403 9467 7517 9491
rect 7403 9415 7434 9467
rect 7486 9415 7517 9467
rect 266 9413 558 9414
rect 266 9361 272 9413
rect 324 9361 348 9413
rect 400 9361 424 9413
rect 476 9361 500 9413
rect 552 9361 558 9413
rect 7403 9409 7517 9415
rect 10896 9500 11287 9501
rect 10896 9448 10902 9500
rect 10954 9448 10968 9500
rect 11020 9448 11034 9500
rect 11086 9448 11099 9500
rect 11151 9448 11164 9500
rect 11216 9448 11229 9500
rect 11281 9448 11287 9500
rect 10896 9426 11287 9448
rect 266 9339 558 9361
rect 266 9287 272 9339
rect 324 9287 348 9339
rect 400 9287 424 9339
rect 476 9287 500 9339
rect 552 9287 558 9339
rect 10896 9374 10902 9426
rect 10954 9374 10968 9426
rect 11020 9374 11034 9426
rect 11086 9374 11099 9426
rect 11151 9374 11164 9426
rect 11216 9374 11229 9426
rect 11281 9374 11287 9426
rect 10896 9352 11287 9374
rect 10896 9300 10902 9352
rect 10954 9300 10968 9352
rect 11020 9300 11034 9352
rect 11086 9300 11099 9352
rect 11151 9300 11164 9352
rect 11216 9300 11229 9352
rect 11281 9300 11287 9352
rect 10896 9299 11287 9300
rect 266 9265 558 9287
rect 266 9260 272 9265
rect 249 9233 272 9260
tri 87 9143 177 9233 ne
rect 177 9213 272 9233
rect 324 9213 348 9265
rect 400 9213 424 9265
rect 476 9213 500 9265
rect 552 9260 558 9265
rect 552 9213 1000 9260
rect 177 9191 1000 9213
rect 177 9143 272 9191
tri 177 9109 211 9143 ne
rect 211 9139 272 9143
rect 324 9139 348 9191
rect 400 9139 424 9191
rect 476 9143 500 9191
rect 552 9143 1000 9191
rect 477 9139 500 9143
rect 211 9114 359 9139
rect 211 9109 277 9114
tri 211 9071 249 9109 ne
rect 249 9062 277 9109
rect 329 9109 359 9114
rect 393 9109 443 9139
rect 477 9109 527 9139
rect 561 9109 611 9143
rect 645 9109 694 9143
rect 728 9109 777 9143
rect 811 9109 860 9143
rect 894 9109 1000 9143
rect 329 9062 1000 9109
rect 249 9058 1000 9062
rect 2778 9259 3778 9260
rect 2778 9207 2784 9259
rect 2836 9207 2851 9259
rect 2903 9207 2918 9259
rect 2970 9207 2985 9259
rect 3037 9207 3052 9259
rect 3104 9207 3119 9259
rect 3171 9207 3186 9259
rect 3238 9207 3253 9259
rect 3305 9207 3320 9259
rect 3372 9207 3387 9259
rect 3439 9207 3454 9259
rect 3506 9207 3521 9259
rect 3573 9207 3588 9259
rect 3640 9207 3654 9259
rect 3706 9207 3720 9259
rect 3772 9207 3778 9259
rect 2778 9185 3778 9207
rect 2778 9133 2784 9185
rect 2836 9133 2851 9185
rect 2903 9133 2918 9185
rect 2970 9133 2985 9185
rect 3037 9133 3052 9185
rect 3104 9133 3119 9185
rect 3171 9133 3186 9185
rect 3238 9133 3253 9185
rect 3305 9133 3320 9185
rect 3372 9133 3387 9185
rect 3439 9133 3454 9185
rect 3506 9133 3521 9185
rect 3573 9133 3588 9185
rect 3640 9133 3654 9185
rect 3706 9133 3720 9185
rect 3772 9133 3778 9185
rect 2778 9111 3778 9133
rect 2778 9059 2784 9111
rect 2836 9059 2851 9111
rect 2903 9059 2918 9111
rect 2970 9059 2985 9111
rect 3037 9059 3052 9111
rect 3104 9059 3119 9111
rect 3171 9059 3186 9111
rect 3238 9059 3253 9111
rect 3305 9059 3320 9111
rect 3372 9059 3387 9111
rect 3439 9059 3454 9111
rect 3506 9059 3521 9111
rect 3573 9059 3588 9111
rect 3640 9059 3654 9111
rect 3706 9059 3720 9111
rect 3772 9059 3778 9111
rect 2778 9058 3778 9059
rect 7399 9254 7571 9260
rect 7451 9202 7519 9254
rect 7399 9185 7571 9202
rect 7451 9133 7519 9185
rect 7399 9116 7571 9133
rect 7451 9064 7519 9116
rect 7399 9058 7571 9064
rect 260 9050 346 9058
rect 260 8998 277 9050
rect 329 8998 346 9050
tri 4016 9020 4022 9026 se
rect 260 8985 346 8998
rect 260 8933 277 8985
rect 329 8933 346 8985
rect 1444 8968 1450 9020
rect 1502 8968 1514 9020
rect 1566 9017 2116 9020
tri 2116 9017 2119 9020 sw
tri 2351 9017 2354 9020 se
rect 2354 9017 4022 9020
rect 1566 8974 4022 9017
rect 1566 8968 1572 8974
tri 1572 8968 1578 8974 nw
tri 3994 8968 4000 8974 ne
rect 4000 8968 4022 8974
tri 4000 8946 4022 8968 ne
rect 260 8927 346 8933
rect 1193 8719 1245 8725
tri 1245 8675 1279 8709 sw
rect 1245 8667 1450 8675
rect 1193 8655 1450 8667
rect 1245 8623 1450 8655
rect 1502 8623 1514 8675
rect 1566 8623 1572 8675
rect 1193 8597 1245 8603
tri 1245 8597 1271 8623 nw
rect 15783 8585 15835 8591
tri 15735 8491 15783 8539 ne
rect 15783 8521 15835 8533
rect 15783 8463 15835 8469
rect 9782 8297 9788 8349
rect 9840 8297 9852 8349
rect 9904 8297 11597 8349
rect 11649 8297 11661 8349
rect 11713 8297 11719 8349
rect 13814 8298 13820 8350
rect 13872 8298 13892 8350
rect 13944 8298 13964 8350
rect 14016 8298 14036 8350
rect 14088 8298 14107 8350
rect 14159 8298 14178 8350
rect 14230 8298 14249 8350
rect 14301 8298 14307 8350
rect 13814 8272 14307 8298
rect 2839 8217 2845 8269
rect 2897 8217 2913 8269
rect 2965 8217 2981 8269
rect 3033 8217 3049 8269
rect 3101 8217 3117 8269
rect 3169 8217 3184 8269
rect 3236 8217 3251 8269
rect 3303 8217 3318 8269
rect 3370 8217 3385 8269
rect 3437 8217 3452 8269
rect 3504 8217 3519 8269
rect 3571 8217 3586 8269
rect 3638 8217 3653 8269
rect 3705 8217 3720 8269
rect 3772 8217 3778 8269
rect 2839 8191 3778 8217
rect 2839 8139 2845 8191
rect 2897 8139 2913 8191
rect 2965 8139 2981 8191
rect 3033 8139 3049 8191
rect 3101 8139 3117 8191
rect 3169 8139 3184 8191
rect 3236 8139 3251 8191
rect 3303 8139 3318 8191
rect 3370 8139 3385 8191
rect 3437 8139 3452 8191
rect 3504 8139 3519 8191
rect 3571 8139 3586 8191
rect 3638 8139 3653 8191
rect 3705 8139 3720 8191
rect 3772 8139 3778 8191
rect 10496 8217 10502 8269
rect 10554 8217 10591 8269
rect 10643 8217 10680 8269
rect 10732 8217 10738 8269
rect 13814 8220 13820 8272
rect 13872 8220 13892 8272
rect 13944 8220 13964 8272
rect 14016 8220 14036 8272
rect 14088 8220 14107 8272
rect 14159 8220 14178 8272
rect 14230 8220 14249 8272
rect 14301 8220 14307 8272
rect 10496 8191 10738 8217
rect 10496 8139 10502 8191
rect 10554 8139 10591 8191
rect 10643 8139 10680 8191
rect 10732 8139 10738 8191
rect 4619 7739 4625 7791
rect 4677 7739 4689 7791
rect 4741 7739 6873 7791
rect 6925 7739 6937 7791
rect 6989 7739 6995 7791
rect 7181 7744 7187 7796
rect 7239 7744 7251 7796
rect 7303 7744 10331 7796
rect 10383 7744 10395 7796
rect 10447 7744 10453 7796
rect 15977 7133 16023 7145
rect 15977 7099 15983 7133
rect 16017 7099 16023 7133
rect 15977 7061 16023 7099
rect 15977 7027 15983 7061
rect 16017 7027 16023 7061
rect 15977 6989 16023 7027
rect 15977 6955 15983 6989
rect 16017 6955 16023 6989
rect 15977 6917 16023 6955
rect 15977 6883 15983 6917
rect 16017 6883 16023 6917
tri 15957 6845 15977 6865 se
rect 15977 6845 16023 6883
tri 15923 6811 15957 6845 se
rect 15957 6811 15983 6845
rect 16017 6811 16023 6845
tri 15885 6773 15923 6811 se
rect 15923 6773 16023 6811
tri 15879 6767 15885 6773 se
rect 15885 6767 15983 6773
rect 15825 6739 15983 6767
rect 16017 6739 16023 6773
rect 15825 6701 16023 6739
rect 15825 6667 15983 6701
rect 16017 6667 16023 6701
rect 15825 6629 16023 6667
rect 15825 6595 15983 6629
rect 16017 6595 16023 6629
rect 15825 6557 16023 6595
rect 15825 6523 15983 6557
rect 16017 6523 16023 6557
rect 15825 6485 16023 6523
rect 15825 6451 15983 6485
rect 16017 6451 16023 6485
rect 15825 6413 16023 6451
rect 15825 6401 15983 6413
tri 15879 6379 15901 6401 ne
rect 15901 6379 15983 6401
rect 16017 6379 16023 6413
tri 15901 6356 15924 6379 ne
rect 15924 6356 16023 6379
rect 10773 6304 10779 6356
rect 10831 6304 10843 6356
rect 10895 6304 12036 6356
rect 12088 6304 12100 6356
rect 12152 6304 12158 6356
tri 15924 6341 15939 6356 ne
rect 15939 6341 16023 6356
tri 15939 6307 15973 6341 ne
rect 15973 6307 15983 6341
rect 16017 6307 16023 6341
tri 15973 6304 15976 6307 ne
rect 15976 6304 16023 6307
tri 15976 6303 15977 6304 ne
rect 15977 6269 16023 6304
rect 15977 6235 15983 6269
rect 16017 6235 16023 6269
rect 15977 6197 16023 6235
rect 15977 6163 15983 6197
rect 16017 6163 16023 6197
rect 15977 6125 16023 6163
rect 15977 6091 15983 6125
rect 16017 6091 16023 6125
rect 11808 5975 11814 6027
rect 11866 5975 11878 6027
rect 11930 5975 12467 6027
rect 12519 5975 12531 6027
rect 12583 5975 12589 6027
rect 15977 6024 16023 6091
rect 15977 4991 16023 5003
rect 15977 4957 15983 4991
rect 16017 4957 16023 4991
rect 15977 4919 16023 4957
rect 15977 4885 15983 4919
rect 16017 4885 16023 4919
rect 15977 4847 16023 4885
rect 15977 4813 15983 4847
rect 16017 4813 16023 4847
rect 15977 4775 16023 4813
tri 15971 4741 15977 4747 se
rect 15977 4741 15983 4775
rect 16017 4741 16023 4775
tri 15934 4704 15971 4741 se
rect 15971 4704 16023 4741
rect 1026 4503 2236 4704
tri 15933 4703 15934 4704 se
rect 15934 4703 16023 4704
tri 15899 4669 15933 4703 se
rect 15933 4669 15983 4703
rect 16017 4669 16023 4703
tri 15861 4631 15899 4669 se
rect 15899 4631 16023 4669
tri 15855 4625 15861 4631 se
rect 15861 4625 15983 4631
rect 15766 4597 15983 4625
rect 16017 4597 16023 4631
rect 15766 4559 16023 4597
rect 15766 4525 15983 4559
rect 16017 4525 16023 4559
rect 15766 4487 16023 4525
rect 15766 4453 15983 4487
rect 16017 4453 16023 4487
rect 15766 4415 16023 4453
rect 15766 4381 15983 4415
rect 16017 4381 16023 4415
rect 15766 4343 16023 4381
rect 15766 4309 15983 4343
rect 16017 4309 16023 4343
tri 8623 4283 8631 4291 se
rect 8631 4283 8637 4291
rect 6852 4231 6858 4283
rect 6910 4231 6922 4283
rect 6974 4275 6980 4283
tri 6980 4275 6988 4283 sw
tri 8615 4275 8623 4283 se
rect 8623 4275 8637 4283
rect 6974 4239 8637 4275
rect 8689 4239 8701 4291
rect 8753 4239 8759 4291
rect 15766 4275 16023 4309
tri 15855 4271 15859 4275 ne
rect 15859 4271 16023 4275
tri 15859 4239 15891 4271 ne
rect 15891 4239 15983 4271
rect 6974 4237 6986 4239
tri 6986 4237 6988 4239 nw
tri 15891 4237 15893 4239 ne
rect 15893 4237 15983 4239
rect 16017 4237 16023 4271
rect 6974 4231 6980 4237
tri 6980 4231 6986 4237 nw
tri 15893 4231 15899 4237 ne
rect 15899 4231 16023 4237
tri 15899 4199 15931 4231 ne
rect 15931 4199 16023 4231
tri 15931 4172 15958 4199 ne
rect 15958 4172 15983 4199
rect 1054 4166 1106 4172
tri 1106 4165 1113 4172 sw
tri 15958 4165 15965 4172 ne
rect 15965 4165 15983 4172
rect 16017 4165 16023 4199
rect 1106 4153 1113 4165
tri 1113 4153 1125 4165 sw
tri 15965 4153 15977 4165 ne
rect 1106 4127 1125 4153
tri 1125 4127 1151 4153 sw
rect 15977 4127 16023 4165
rect 1106 4123 1151 4127
tri 1151 4123 1155 4127 sw
rect 1106 4114 1457 4123
rect 1054 4102 1457 4114
rect 1106 4071 1457 4102
rect 1509 4071 1521 4123
rect 1573 4071 1579 4123
rect 15977 4093 15983 4127
rect 16017 4093 16023 4127
rect 1106 4055 1117 4071
tri 1117 4055 1133 4071 nw
rect 15977 4055 16023 4093
rect 1054 4044 1106 4050
tri 1106 4044 1117 4055 nw
rect 15977 4021 15983 4055
rect 16017 4021 16023 4055
rect 15977 3983 16023 4021
rect 15977 3949 15983 3983
rect 16017 3949 16023 3983
rect 15977 3897 16023 3949
rect 1960 3622 1966 3674
rect 2018 3622 2030 3674
rect 2082 3662 2088 3674
tri 2088 3662 2100 3674 sw
tri 5503 3662 5515 3674 se
rect 5515 3662 5521 3674
rect 2082 3622 5521 3662
rect 5573 3622 5585 3674
rect 5637 3622 5643 3674
rect 14304 3347 14310 3399
rect 14362 3347 14374 3399
rect 14426 3347 15361 3399
rect 15413 3347 15425 3399
rect 15477 3347 15483 3399
rect 6848 3344 7071 3345
rect 5489 3144 5517 3344
rect 6848 3292 6854 3344
rect 6906 3292 6934 3344
rect 6986 3292 7013 3344
rect 7065 3292 7071 3344
rect 6848 3272 7071 3292
rect 6848 3220 6854 3272
rect 6906 3220 6934 3272
rect 6986 3220 7013 3272
rect 7065 3220 7071 3272
rect 6848 3200 7071 3220
rect 6848 3148 6854 3200
rect 6906 3148 6934 3200
rect 6986 3148 7013 3200
rect 7065 3148 7071 3200
rect 6848 3147 7071 3148
rect 8615 3293 8621 3345
rect 8673 3293 8717 3345
rect 8769 3293 8775 3345
rect 8615 3271 8775 3293
rect 8615 3219 8621 3271
rect 8673 3219 8717 3271
rect 8769 3219 8775 3271
rect 8615 3197 8775 3219
rect 8615 3145 8621 3197
rect 8673 3145 8717 3197
rect 8769 3145 8775 3197
rect 42 2802 94 2808
rect 42 2738 94 2750
rect 42 2680 94 2686
rect 2440 2646 2761 2647
rect 2440 2594 2446 2646
rect 2498 2594 2511 2646
rect 2563 2594 2575 2646
rect 2627 2594 2639 2646
rect 2691 2594 2703 2646
rect 2755 2594 2761 2646
rect 2440 2574 2761 2594
rect 2440 2522 2446 2574
rect 2498 2522 2511 2574
rect 2563 2522 2575 2574
rect 2627 2522 2639 2574
rect 2691 2522 2703 2574
rect 2755 2522 2761 2574
rect 2440 2502 2761 2522
rect 2440 2450 2446 2502
rect 2498 2450 2511 2502
rect 2563 2450 2575 2502
rect 2627 2450 2639 2502
rect 2691 2450 2703 2502
rect 2755 2450 2761 2502
rect 2440 2449 2761 2450
rect 3627 2646 4312 2647
rect 3627 2594 3633 2646
rect 3685 2594 3702 2646
rect 3754 2594 3771 2646
rect 3823 2594 3840 2646
rect 3892 2594 3909 2646
rect 3961 2594 3978 2646
rect 4030 2594 4047 2646
rect 4099 2594 4116 2646
rect 4168 2594 4185 2646
rect 4237 2594 4254 2646
rect 4306 2594 4312 2646
rect 3627 2574 4312 2594
rect 3627 2522 3633 2574
rect 3685 2522 3702 2574
rect 3754 2522 3771 2574
rect 3823 2522 3840 2574
rect 3892 2522 3909 2574
rect 3961 2522 3978 2574
rect 4030 2522 4047 2574
rect 4099 2522 4116 2574
rect 4168 2522 4185 2574
rect 4237 2522 4254 2574
rect 4306 2522 4312 2574
rect 3627 2502 4312 2522
rect 3627 2450 3633 2502
rect 3685 2450 3702 2502
rect 3754 2450 3771 2502
rect 3823 2450 3840 2502
rect 3892 2450 3909 2502
rect 3961 2450 3978 2502
rect 4030 2450 4047 2502
rect 4099 2450 4116 2502
rect 4168 2450 4185 2502
rect 4237 2450 4254 2502
rect 4306 2450 4312 2502
rect 10506 2595 10512 2647
rect 10564 2595 10579 2647
rect 10631 2595 10637 2647
rect 10506 2575 10637 2595
rect 10506 2523 10512 2575
rect 10564 2523 10579 2575
rect 10631 2523 10637 2575
rect 10506 2503 10637 2523
rect 10506 2451 10512 2503
rect 10564 2451 10579 2503
rect 10631 2451 10637 2503
rect 10701 2595 10707 2647
rect 10759 2595 10780 2647
rect 10832 2595 10853 2647
rect 10905 2595 10926 2647
rect 10978 2595 10999 2647
rect 11051 2595 11057 2647
rect 10701 2575 11057 2595
rect 10701 2523 10707 2575
rect 10759 2523 10780 2575
rect 10832 2523 10853 2575
rect 10905 2523 10926 2575
rect 10978 2523 10999 2575
rect 11051 2523 11057 2575
rect 10701 2503 11057 2523
rect 10701 2451 10707 2503
rect 10759 2451 10780 2503
rect 10832 2451 10853 2503
rect 10905 2451 10926 2503
rect 10978 2451 10999 2503
rect 11051 2451 11057 2503
rect 3627 2449 4312 2450
rect 15421 2423 15473 2429
rect 15421 2359 15473 2371
rect 15421 2286 15473 2307
rect 324 2123 330 2175
rect 382 2123 394 2175
rect 446 2123 811 2175
rect 863 2123 875 2175
rect 927 2123 933 2175
tri 13834 2099 13839 2104 se
tri 13803 2068 13834 2099 se
rect 13834 2068 13839 2099
tri 13769 2034 13803 2068 se
rect 13803 2034 13839 2068
tri 13765 2030 13769 2034 se
rect 13769 2030 13839 2034
rect 13937 2068 14323 2099
rect 13937 2034 13949 2068
rect 13983 2034 14031 2068
rect 14065 2034 14113 2068
rect 14147 2034 14195 2068
rect 14229 2034 14277 2068
rect 14311 2034 14323 2068
tri 13759 2024 13765 2030 se
rect 13765 2024 13900 2030
tri 13738 2003 13759 2024 se
rect 13759 2003 13782 2024
tri 13725 1990 13738 2003 se
rect 13738 1990 13782 2003
rect 13816 1990 13854 2024
rect 13888 1990 13900 2024
rect 13937 2003 14323 2034
rect 14626 2053 14632 2105
rect 14684 2053 14711 2105
rect 14763 2053 14789 2105
rect 14841 2053 14847 2105
rect 14626 2033 14847 2053
tri 13690 1955 13725 1990 se
rect 13725 1984 13900 1990
rect 13725 1955 13839 1984
rect 14626 1981 14632 2033
rect 14684 1981 14711 2033
rect 14763 1981 14789 2033
rect 14841 1981 14847 2033
rect 14626 1961 14847 1981
rect 13373 1949 13885 1955
rect 13373 1915 13451 1949
rect 13485 1915 13529 1949
rect 13563 1915 13607 1949
rect 13641 1915 13685 1949
rect 13719 1915 13762 1949
rect 13796 1915 13839 1949
rect 13873 1915 13885 1949
rect 13373 1909 13885 1915
rect 14626 1909 14632 1961
rect 14684 1909 14711 1961
rect 14763 1909 14789 1961
rect 14841 1909 14847 1961
rect 15077 2099 15251 2105
rect 15129 2047 15199 2099
rect 15077 2033 15251 2047
rect 15129 1981 15199 2033
rect 15077 1967 15251 1981
rect 15129 1915 15199 1967
rect 15077 1909 15251 1915
rect 13373 1873 13419 1909
rect 13373 1839 13379 1873
rect 13413 1839 13419 1873
rect 1497 1804 1625 1810
rect 1549 1752 1573 1804
rect 1497 1738 1625 1752
rect 1549 1686 1573 1738
rect 1497 1680 1625 1686
rect 6848 1758 6854 1810
rect 6906 1758 6934 1810
rect 6986 1758 7013 1810
rect 7065 1758 7071 1810
rect 6848 1732 7071 1758
rect 6848 1680 6854 1732
rect 6906 1680 6934 1732
rect 6986 1680 7013 1732
rect 7065 1680 7071 1732
rect 8615 1758 8621 1810
rect 8673 1758 8717 1810
rect 8769 1758 8775 1810
rect 8615 1732 8775 1758
rect 8615 1680 8621 1732
rect 8673 1680 8717 1732
rect 8769 1680 8775 1732
rect 13373 1797 13419 1839
tri 13419 1821 13507 1909 nw
rect 13373 1763 13379 1797
rect 13413 1763 13419 1797
rect 13373 1721 13419 1763
rect 13373 1687 13379 1721
rect 13413 1687 13419 1721
rect 13373 1675 13419 1687
rect 1499 1646 1655 1652
rect 1551 1594 1603 1646
rect 1499 1577 1655 1594
rect 1551 1525 1603 1577
rect 1499 1508 1655 1525
rect 1551 1456 1603 1508
rect 1499 1450 1655 1456
rect 1780 1651 1858 1652
rect 1780 1599 1786 1651
rect 1838 1599 1858 1651
rect 1780 1577 1858 1599
rect 1780 1525 1786 1577
rect 1838 1525 1858 1577
rect 1780 1503 1858 1525
rect 1780 1451 1786 1503
rect 1838 1451 1858 1503
rect 1780 1450 1858 1451
rect 3847 1651 4275 1652
rect 3847 1599 3853 1651
rect 3905 1599 3926 1651
rect 3978 1599 3999 1651
rect 4051 1599 4072 1651
rect 4124 1599 4145 1651
rect 4197 1599 4217 1651
rect 4269 1599 4275 1651
rect 3847 1577 4275 1599
rect 3847 1525 3853 1577
rect 3905 1525 3926 1577
rect 3978 1525 3999 1577
rect 4051 1525 4072 1577
rect 4124 1525 4145 1577
rect 4197 1525 4217 1577
rect 4269 1525 4275 1577
rect 3847 1503 4275 1525
rect 3847 1451 3853 1503
rect 3905 1451 3926 1503
rect 3978 1451 3999 1503
rect 4051 1451 4072 1503
rect 4124 1451 4145 1503
rect 4197 1451 4217 1503
rect 4269 1451 4275 1503
rect 3847 1450 4275 1451
rect 4848 1651 5253 1652
rect 4848 1599 4854 1651
rect 4906 1599 4923 1651
rect 4975 1599 4991 1651
rect 5043 1599 5059 1651
rect 5111 1599 5127 1651
rect 5179 1599 5195 1651
rect 5247 1599 5253 1651
rect 4848 1577 5253 1599
rect 4848 1525 4854 1577
rect 4906 1525 4923 1577
rect 4975 1525 4991 1577
rect 5043 1525 5059 1577
rect 5111 1525 5127 1577
rect 5179 1525 5195 1577
rect 5247 1525 5253 1577
rect 4848 1503 5253 1525
rect 4848 1451 4854 1503
rect 4906 1451 4923 1503
rect 4975 1451 4991 1503
rect 5043 1451 5059 1503
rect 5111 1451 5127 1503
rect 5179 1451 5195 1503
rect 5247 1451 5253 1503
rect 4848 1450 5253 1451
rect 6838 1651 7057 1652
rect 6838 1599 6844 1651
rect 6896 1599 6922 1651
rect 6974 1599 6999 1651
rect 7051 1599 7057 1651
rect 6838 1577 7057 1599
rect 6838 1525 6844 1577
rect 6896 1525 6922 1577
rect 6974 1525 6999 1577
rect 7051 1525 7057 1577
rect 6838 1503 7057 1525
rect 6838 1451 6844 1503
rect 6896 1451 6922 1503
rect 6974 1451 6999 1503
rect 7051 1451 7057 1503
rect 6838 1450 7057 1451
rect 14181 1339 15084 1391
tri 15062 1337 15064 1339 ne
rect 15064 1337 15084 1339
tri 15084 1337 15138 1391 sw
rect 1163 1285 1188 1337
rect 1240 1285 1252 1337
rect 1304 1285 1310 1337
tri 15064 1331 15070 1337 ne
rect 15070 1331 15138 1337
tri 15138 1331 15144 1337 sw
tri 15070 1329 15072 1331 ne
rect 15072 1329 15144 1331
rect 5592 1300 5636 1329
tri 15072 1317 15084 1329 ne
rect 15084 1317 15144 1329
tri 15084 1309 15092 1317 ne
tri 15068 1176 15092 1200 se
rect 15092 1178 15144 1317
rect 15092 1176 15127 1178
rect 3208 1124 3214 1176
rect 3266 1124 3278 1176
rect 3330 1124 8938 1176
rect 8990 1124 9002 1176
rect 9054 1124 9060 1176
tri 15053 1161 15068 1176 se
rect 15068 1161 15127 1176
tri 15127 1161 15144 1178 nw
rect 12486 1109 12492 1161
rect 12544 1109 12556 1161
rect 12608 1109 15075 1161
tri 15075 1109 15127 1161 nw
rect 2779 1086 3341 1087
rect 2779 1034 2785 1086
rect 2837 1034 2857 1086
rect 2909 1034 2928 1086
rect 2980 1034 2999 1086
rect 3051 1034 3070 1086
rect 3122 1034 3141 1086
rect 3193 1034 3212 1086
rect 3264 1034 3283 1086
rect 3335 1034 3341 1086
rect 2779 1010 3341 1034
rect 2779 958 2785 1010
rect 2837 958 2857 1010
rect 2909 958 2928 1010
rect 2980 958 2999 1010
rect 3051 958 3070 1010
rect 3122 958 3141 1010
rect 3193 958 3212 1010
rect 3264 958 3283 1010
rect 3335 958 3341 1010
rect 2779 934 3341 958
rect 2779 882 2785 934
rect 2837 882 2857 934
rect 2909 882 2928 934
rect 2980 882 2999 934
rect 3051 882 3070 934
rect 3122 882 3141 934
rect 3193 882 3212 934
rect 3264 882 3283 934
rect 3335 882 3341 934
rect 2779 881 3341 882
rect 6911 877 7555 1091
rect 8215 877 9003 1092
tri 12240 1091 12241 1092 sw
rect 10505 1090 10831 1091
rect 10505 1038 10511 1090
rect 10563 1038 10577 1090
rect 10629 1038 10643 1090
rect 10695 1038 10708 1090
rect 10760 1038 10773 1090
rect 10825 1038 10831 1090
rect 12240 1078 12241 1091
tri 12241 1078 12254 1091 sw
rect 10505 1010 10831 1038
rect 10505 958 10511 1010
rect 10563 958 10577 1010
rect 10629 958 10643 1010
rect 10695 958 10708 1010
rect 10760 958 10773 1010
rect 10825 958 10831 1010
rect 10505 930 10831 958
rect 10505 878 10511 930
rect 10563 878 10577 930
rect 10629 878 10643 930
rect 10695 878 10708 930
rect 10760 878 10773 930
rect 10825 878 10831 930
rect 10505 877 10831 878
rect 12223 1069 13635 1078
rect 12223 1035 12312 1069
rect 12346 1035 12387 1069
rect 12421 1035 12462 1069
rect 12496 1035 12536 1069
rect 12570 1035 12610 1069
rect 12644 1035 12684 1069
rect 12718 1035 12758 1069
rect 12792 1035 12832 1069
rect 12866 1035 12906 1069
rect 12940 1035 12980 1069
rect 13014 1035 13054 1069
rect 13088 1035 13128 1069
rect 13162 1035 13202 1069
rect 13236 1035 13276 1069
rect 13310 1035 13350 1069
rect 13384 1035 13424 1069
rect 13458 1035 13635 1069
rect 12223 987 13635 1035
rect 12223 953 12312 987
rect 12346 953 12387 987
rect 12421 953 12462 987
rect 12496 953 12536 987
rect 12570 953 12610 987
rect 12644 953 12684 987
rect 12718 953 12758 987
rect 12792 953 12832 987
rect 12866 953 12906 987
rect 12940 953 12980 987
rect 13014 953 13054 987
rect 13088 953 13128 987
rect 13162 953 13202 987
rect 13236 953 13276 987
rect 13310 953 13350 987
rect 13384 953 13424 987
rect 13458 980 13635 987
rect 15086 1026 15092 1078
rect 15144 1026 15193 1078
rect 15245 1026 15262 1078
rect 15086 1014 15262 1026
rect 13458 953 13518 980
rect 12223 948 13518 953
tri 13518 948 13550 980 nw
tri 15068 962 15086 980 ne
rect 15086 962 15092 1014
rect 15144 962 15193 1014
rect 15245 962 15262 1014
rect 15433 1046 15561 1047
rect 15433 994 15439 1046
rect 15491 994 15503 1046
rect 15555 994 15561 1046
rect 15433 958 15561 994
rect 12223 947 13517 948
tri 13517 947 13518 948 nw
rect 12223 914 13484 947
tri 13484 914 13517 947 nw
rect 12223 877 13447 914
tri 13447 877 13484 914 nw
rect 15433 906 15439 958
rect 15491 906 15503 958
rect 15555 906 15561 958
rect 15433 870 15561 906
rect 8936 839 8988 845
rect 6363 787 6415 793
tri 8988 828 9005 845 sw
rect 8988 818 9005 828
tri 9005 818 9015 828 sw
rect 15433 818 15439 870
rect 15491 818 15503 870
rect 15555 818 15561 870
rect 8988 787 9371 818
rect 7035 777 7079 782
rect 6363 720 6415 735
rect 6363 663 6415 668
rect 7027 771 7079 777
rect 7027 707 7079 719
rect 8936 776 9371 787
rect 8936 775 9006 776
rect 8988 767 9006 775
tri 9006 767 9015 776 nw
tri 9286 767 9295 776 ne
rect 9295 767 9325 776
rect 8988 764 9003 767
tri 9003 764 9006 767 nw
tri 9295 764 9298 767 ne
rect 9298 764 9325 767
tri 8988 749 9003 764 nw
tri 9298 749 9313 764 ne
rect 9313 749 9325 764
tri 9313 737 9325 749 ne
rect 9776 761 9828 799
rect 13655 786 13785 796
rect 13707 784 13733 786
rect 8936 717 8988 723
rect 6363 662 6427 663
rect 7027 649 7079 655
rect 9776 697 9828 709
rect 9776 639 9828 645
rect 10216 762 10268 768
rect 10309 764 10372 768
rect 10216 692 10268 710
rect 10216 634 10268 640
rect 10320 762 10372 764
rect 11410 724 11416 776
rect 11468 724 11487 776
rect 11539 724 11545 776
rect 12048 718 12054 770
rect 12106 718 12118 770
rect 12170 718 12183 770
rect 10320 692 10372 710
rect 10320 634 10372 640
rect 13655 716 13664 734
rect 13770 716 13785 734
rect 15433 782 15561 818
rect 15433 730 15439 782
rect 15491 730 15503 782
rect 15555 730 15561 782
rect 15433 729 15561 730
rect 13655 646 13664 664
rect 13770 646 13785 664
rect 13707 594 13733 606
rect 13655 576 13785 594
rect 2308 523 2314 575
rect 2366 523 2378 575
rect 2430 570 2436 575
tri 2436 570 2441 575 sw
rect 2430 567 2441 570
tri 2441 567 2444 570 sw
rect 2430 560 2444 567
tri 2444 560 2451 567 sw
rect 11890 564 11942 570
rect 2430 558 2797 560
tri 2797 558 2799 560 sw
rect 2430 557 3677 558
tri 3677 557 3678 558 sw
tri 3897 557 3898 558 se
rect 3898 557 5791 558
tri 5791 557 5792 558 sw
tri 6108 557 6109 558 se
rect 6109 557 7013 558
rect 2430 526 7013 557
tri 7013 526 7045 558 sw
rect 2430 524 7045 526
tri 7045 524 7047 526 sw
rect 2430 523 7047 524
tri 7047 523 7048 524 sw
tri 2751 522 2752 523 ne
rect 2752 522 7048 523
tri 6999 519 7002 522 ne
rect 7002 519 7048 522
tri 7048 519 7052 523 sw
rect 1169 467 1175 519
rect 1227 467 1239 519
rect 1291 467 1902 519
rect 1954 467 1966 519
rect 2018 467 2024 519
tri 7002 494 7027 519 ne
rect 7027 494 7052 519
tri 7052 494 7077 519 sw
rect 11890 498 11942 512
tri 7027 486 7035 494 ne
rect 7035 486 7077 494
tri 7077 486 7085 494 sw
tri 7035 476 7045 486 ne
rect 7045 483 7085 486
tri 7085 483 7088 486 sw
rect 7045 476 7088 483
tri 7088 476 7095 483 sw
tri 8615 476 8622 483 se
rect 8622 476 10182 483
tri 7045 467 7054 476 ne
rect 7054 467 7095 476
tri 7095 467 7104 476 sw
tri 8606 467 8615 476 se
rect 8615 467 10182 476
tri 7054 452 7069 467 ne
rect 7069 452 7104 467
tri 7104 452 7119 467 sw
tri 8591 452 8606 467 se
rect 8606 452 10182 467
tri 7069 426 7095 452 ne
rect 7095 433 7119 452
tri 7119 433 7138 452 sw
tri 8572 433 8591 452 se
rect 8591 447 10182 452
rect 8591 433 8622 447
tri 8622 433 8636 447 nw
tri 10160 433 10174 447 ne
rect 10174 433 10182 447
rect 7095 431 7138 433
tri 7138 431 7140 433 sw
tri 8570 431 8572 433 se
rect 8572 431 8620 433
tri 8620 431 8622 433 nw
tri 10174 431 10176 433 ne
rect 10176 431 10182 433
rect 10234 431 10246 483
rect 10298 431 10304 483
rect 13707 524 13733 576
rect 13655 506 13785 524
rect 13707 454 13733 506
rect 13655 448 13785 454
rect 11890 440 11942 446
rect 7095 426 7140 431
tri 7140 426 7145 431 sw
tri 8565 426 8570 431 se
rect 8570 426 8615 431
tri 8615 426 8620 431 nw
tri 7095 415 7106 426 ne
rect 7106 415 8604 426
tri 8604 415 8615 426 nw
tri 7106 390 7131 415 ne
rect 7131 390 8579 415
tri 8579 390 8604 415 nw
tri 8661 390 8686 415 se
rect 8686 390 9536 415
tri 8620 349 8661 390 se
rect 8661 383 9536 390
tri 9536 383 9568 415 sw
rect 8661 369 9568 383
rect 8661 349 8686 369
tri 8686 349 8706 369 nw
tri 9516 349 9536 369 ne
rect 9536 349 9568 369
tri 9568 349 9602 383 sw
tri 10928 349 10962 383 se
rect 10962 356 10975 383
rect 12486 377 12538 383
rect 10962 349 11008 356
tri 8608 337 8620 349 se
rect 8620 337 8674 349
tri 8674 337 8686 349 nw
tri 9536 337 9548 349 ne
rect 9548 337 11008 349
rect 7878 285 7884 337
rect 7936 285 7948 337
rect 8000 285 8622 337
tri 8622 285 8674 337 nw
tri 9548 303 9582 337 ne
rect 9582 303 11008 337
rect 12486 313 12538 325
rect 4654 256 5253 257
rect 6909 256 7555 257
rect 1434 255 2143 256
rect 1434 203 1440 255
rect 1492 203 1548 255
rect 1600 203 1656 255
rect 1708 203 1764 255
rect 1816 203 1871 255
rect 1923 203 1978 255
rect 2030 203 2085 255
rect 2137 203 2143 255
rect 1434 181 2143 203
rect 1434 129 1440 181
rect 1492 129 1548 181
rect 1600 129 1656 181
rect 1708 129 1764 181
rect 1816 129 1871 181
rect 1923 129 1978 181
rect 2030 129 2085 181
rect 2137 129 2143 181
rect 1434 107 2143 129
rect 1434 55 1440 107
rect 1492 55 1548 107
rect 1600 55 1656 107
rect 1708 55 1764 107
rect 1816 55 1871 107
rect 1923 55 1978 107
rect 2030 55 2085 107
rect 2137 55 2143 107
rect 1434 54 2143 55
rect 3847 255 4275 256
rect 3847 203 3853 255
rect 3905 203 3926 255
rect 3978 203 3999 255
rect 4051 203 4072 255
rect 4124 203 4145 255
rect 4197 203 4217 255
rect 4269 203 4275 255
rect 3847 181 4275 203
rect 3847 129 3853 181
rect 3905 129 3926 181
rect 3978 129 3999 181
rect 4051 129 4072 181
rect 4124 129 4145 181
rect 4197 129 4217 181
rect 4269 129 4275 181
rect 3847 107 4275 129
rect 3847 55 3853 107
rect 3905 55 3926 107
rect 3978 55 3999 107
rect 4051 55 4072 107
rect 4124 55 4145 107
rect 4197 55 4217 107
rect 4269 55 4275 107
rect 4654 204 4660 256
rect 4712 204 4767 256
rect 4819 204 4874 256
rect 4926 204 4981 256
rect 5033 204 5088 256
rect 5140 204 5195 256
rect 5247 204 5253 256
rect 4654 182 5253 204
rect 4654 130 4660 182
rect 4712 130 4767 182
rect 4819 130 4874 182
rect 4926 130 4981 182
rect 5033 130 5088 182
rect 5140 130 5195 182
rect 5247 130 5253 182
rect 4654 108 5253 130
rect 4654 56 4660 108
rect 4712 56 4767 108
rect 4819 56 4874 108
rect 4926 56 4981 108
rect 5033 56 5088 108
rect 5140 56 5195 108
rect 5247 56 5253 108
rect 4654 55 5253 56
rect 6680 255 7555 256
rect 6680 203 6686 255
rect 6738 203 6781 255
rect 6833 203 6876 255
rect 6928 203 7555 255
rect 6680 181 7555 203
rect 6680 129 6686 181
rect 6738 129 6781 181
rect 6833 129 6876 181
rect 6928 129 7555 181
rect 6680 107 7555 129
rect 6680 55 6686 107
rect 6738 55 6781 107
rect 6833 55 6876 107
rect 6928 55 7555 107
rect 3847 54 4275 55
rect 6680 54 7555 55
rect 8213 54 8387 257
rect 12486 0 12538 261
rect 12875 180 13459 182
rect 12875 128 12881 180
rect 12933 171 12982 180
rect 13034 171 13459 180
rect 12933 137 12960 171
rect 13067 137 13105 171
rect 13139 137 13177 171
rect 13211 137 13459 171
rect 12933 128 12982 137
rect 13034 128 13459 137
rect 12875 104 13459 128
rect 12875 52 12881 104
rect 12933 93 12982 104
rect 13034 93 13459 104
rect 12933 59 12960 93
rect 13067 59 13105 93
rect 13139 59 13177 93
rect 13211 59 13459 93
rect 12933 52 12982 59
rect 13034 52 13459 59
<< via1 >>
rect 3160 39942 3212 39994
rect 3225 39942 3277 39994
rect 3290 39942 3342 39994
rect 3355 39942 3407 39994
rect 3420 39942 3472 39994
rect 3485 39942 3537 39994
rect 3550 39942 3602 39994
rect 3615 39942 3667 39994
rect 3680 39942 3732 39994
rect 3745 39942 3797 39994
rect 3810 39942 3862 39994
rect 3875 39942 3927 39994
rect 3940 39942 3992 39994
rect 4005 39942 4057 39994
rect 4070 39942 4122 39994
rect 4135 39942 4187 39994
rect 4200 39942 4252 39994
rect 4265 39942 4317 39994
rect 4330 39942 4382 39994
rect 4395 39942 4447 39994
rect 4460 39942 4512 39994
rect 4525 39942 4577 39994
rect 4590 39942 4642 39994
rect 4655 39942 4707 39994
rect 4720 39942 4772 39994
rect 4785 39942 4837 39994
rect 4850 39942 4902 39994
rect 4915 39942 4967 39994
rect 4980 39942 5032 39994
rect 5045 39942 5097 39994
rect 5110 39942 5162 39994
rect 5175 39942 5227 39994
rect 5240 39942 5292 39994
rect 5305 39942 5357 39994
rect 5370 39942 5422 39994
rect 5435 39942 5487 39994
rect 5500 39942 5552 39994
rect 5565 39942 5617 39994
rect 5630 39942 5682 39994
rect 5695 39942 5747 39994
rect 5760 39942 5812 39994
rect 5825 39942 5877 39994
rect 5890 39942 5942 39994
rect 5955 39942 6007 39994
rect 6020 39942 6072 39994
rect 6085 39942 6137 39994
rect 6150 39942 6202 39994
rect 6215 39942 6267 39994
rect 6280 39942 6332 39994
rect 6345 39942 6397 39994
rect 6410 39942 6462 39994
rect 6475 39942 6527 39994
rect 6540 39942 6592 39994
rect 6605 39942 6657 39994
rect 6670 39942 6722 39994
rect 6735 39942 6787 39994
rect 6800 39942 6852 39994
rect 6865 39942 6917 39994
rect 6930 39942 6982 39994
rect 6995 39942 7047 39994
rect 7060 39942 7112 39994
rect 7125 39942 7177 39994
rect 7189 39942 7241 39994
rect 7253 39942 7305 39994
rect 7317 39942 7369 39994
rect 7381 39942 7433 39994
rect 7445 39942 7497 39994
rect 7509 39942 7561 39994
rect 7573 39942 7625 39994
rect 7637 39942 7689 39994
rect 7701 39942 7753 39994
rect 7765 39942 7817 39994
rect 7829 39942 7881 39994
rect 7893 39942 7945 39994
rect 7957 39942 8009 39994
rect 8021 39942 8073 39994
rect 8085 39942 8137 39994
rect 8149 39942 8201 39994
rect 8213 39942 8265 39994
rect 8277 39942 8329 39994
rect 8341 39942 8393 39994
rect 8405 39942 8457 39994
rect 8469 39942 8521 39994
rect 8533 39942 8585 39994
rect 8597 39942 8649 39994
rect 8661 39942 8713 39994
rect 8725 39942 8777 39994
rect 8789 39942 8841 39994
rect 8853 39942 8905 39994
rect 8917 39942 8969 39994
rect 8981 39942 9033 39994
rect 9045 39942 9097 39994
rect 9109 39942 9161 39994
rect 9173 39942 9225 39994
rect 9237 39942 9289 39994
rect 9301 39942 9353 39994
rect 9365 39942 9417 39994
rect 9429 39942 9481 39994
rect 9493 39942 9545 39994
rect 9557 39942 9609 39994
rect 9621 39942 9673 39994
rect 9685 39942 9737 39994
rect 9749 39942 9801 39994
rect 9813 39942 9865 39994
rect 9877 39942 9929 39994
rect 9941 39942 9993 39994
rect 10005 39942 10057 39994
rect 10069 39942 10121 39994
rect 10133 39942 10185 39994
rect 10197 39942 10249 39994
rect 10261 39942 10313 39994
rect 10325 39942 10377 39994
rect 10389 39942 10441 39994
rect 10453 39942 10505 39994
rect 10517 39942 10569 39994
rect 10581 39942 10633 39994
rect 10645 39942 10697 39994
rect 10709 39942 10761 39994
rect 10773 39942 10825 39994
rect 10837 39942 10889 39994
rect 10901 39942 10953 39994
rect 10965 39942 11017 39994
rect 11029 39942 11081 39994
rect 11093 39942 11145 39994
rect 11157 39942 11209 39994
rect 11221 39942 11273 39994
rect 11285 39942 11337 39994
rect 3160 39874 3212 39926
rect 3225 39874 3277 39926
rect 3290 39874 3342 39926
rect 3355 39874 3407 39926
rect 3420 39874 3472 39926
rect 3485 39874 3537 39926
rect 3550 39874 3602 39926
rect 3615 39874 3667 39926
rect 3680 39874 3732 39926
rect 3745 39874 3797 39926
rect 3810 39874 3862 39926
rect 3875 39874 3927 39926
rect 3940 39874 3992 39926
rect 4005 39874 4057 39926
rect 4070 39874 4122 39926
rect 4135 39874 4187 39926
rect 4200 39874 4252 39926
rect 4265 39874 4317 39926
rect 4330 39874 4382 39926
rect 4395 39874 4447 39926
rect 4460 39874 4512 39926
rect 4525 39874 4577 39926
rect 4590 39874 4642 39926
rect 4655 39874 4707 39926
rect 4720 39874 4772 39926
rect 4785 39874 4837 39926
rect 4850 39874 4902 39926
rect 4915 39874 4967 39926
rect 4980 39874 5032 39926
rect 5045 39874 5097 39926
rect 5110 39874 5162 39926
rect 5175 39874 5227 39926
rect 5240 39874 5292 39926
rect 5305 39874 5357 39926
rect 5370 39874 5422 39926
rect 5435 39874 5487 39926
rect 5500 39874 5552 39926
rect 5565 39874 5617 39926
rect 5630 39874 5682 39926
rect 5695 39874 5747 39926
rect 5760 39874 5812 39926
rect 5825 39874 5877 39926
rect 5890 39874 5942 39926
rect 5955 39874 6007 39926
rect 6020 39874 6072 39926
rect 6085 39874 6137 39926
rect 6150 39874 6202 39926
rect 6215 39874 6267 39926
rect 6280 39874 6332 39926
rect 6345 39874 6397 39926
rect 6410 39874 6462 39926
rect 6475 39874 6527 39926
rect 6540 39874 6592 39926
rect 6605 39874 6657 39926
rect 6670 39874 6722 39926
rect 6735 39874 6787 39926
rect 6800 39874 6852 39926
rect 6865 39874 6917 39926
rect 6930 39874 6982 39926
rect 6995 39874 7047 39926
rect 7060 39874 7112 39926
rect 7125 39874 7177 39926
rect 7189 39874 7241 39926
rect 7253 39874 7305 39926
rect 7317 39874 7369 39926
rect 7381 39874 7433 39926
rect 7445 39874 7497 39926
rect 7509 39874 7561 39926
rect 7573 39874 7625 39926
rect 7637 39874 7689 39926
rect 7701 39874 7753 39926
rect 7765 39874 7817 39926
rect 7829 39874 7881 39926
rect 7893 39874 7945 39926
rect 7957 39874 8009 39926
rect 8021 39874 8073 39926
rect 8085 39874 8137 39926
rect 8149 39874 8201 39926
rect 8213 39874 8265 39926
rect 8277 39874 8329 39926
rect 8341 39874 8393 39926
rect 8405 39874 8457 39926
rect 8469 39874 8521 39926
rect 8533 39874 8585 39926
rect 8597 39874 8649 39926
rect 8661 39874 8713 39926
rect 8725 39874 8777 39926
rect 8789 39874 8841 39926
rect 8853 39874 8905 39926
rect 8917 39874 8969 39926
rect 8981 39874 9033 39926
rect 9045 39874 9097 39926
rect 9109 39874 9161 39926
rect 9173 39874 9225 39926
rect 9237 39874 9289 39926
rect 9301 39874 9353 39926
rect 9365 39874 9417 39926
rect 9429 39874 9481 39926
rect 9493 39874 9545 39926
rect 9557 39874 9609 39926
rect 9621 39874 9673 39926
rect 9685 39874 9737 39926
rect 9749 39874 9801 39926
rect 9813 39874 9865 39926
rect 9877 39874 9929 39926
rect 9941 39874 9993 39926
rect 10005 39874 10057 39926
rect 10069 39874 10121 39926
rect 10133 39874 10185 39926
rect 10197 39874 10249 39926
rect 10261 39874 10313 39926
rect 10325 39874 10377 39926
rect 10389 39874 10441 39926
rect 10453 39874 10505 39926
rect 10517 39874 10569 39926
rect 10581 39874 10633 39926
rect 10645 39874 10697 39926
rect 10709 39874 10761 39926
rect 10773 39874 10825 39926
rect 10837 39874 10889 39926
rect 10901 39874 10953 39926
rect 10965 39874 11017 39926
rect 11029 39874 11081 39926
rect 11093 39874 11145 39926
rect 11157 39874 11209 39926
rect 11221 39874 11273 39926
rect 11285 39874 11337 39926
rect 3160 39806 3212 39858
rect 3225 39806 3277 39858
rect 3290 39806 3342 39858
rect 3355 39806 3407 39858
rect 3420 39806 3472 39858
rect 3485 39806 3537 39858
rect 3550 39806 3602 39858
rect 3615 39806 3667 39858
rect 3680 39806 3732 39858
rect 3745 39806 3797 39858
rect 3810 39806 3862 39858
rect 3875 39806 3927 39858
rect 3940 39806 3992 39858
rect 4005 39806 4057 39858
rect 4070 39806 4122 39858
rect 4135 39806 4187 39858
rect 4200 39806 4252 39858
rect 4265 39806 4317 39858
rect 4330 39806 4382 39858
rect 4395 39806 4447 39858
rect 4460 39806 4512 39858
rect 4525 39806 4577 39858
rect 4590 39806 4642 39858
rect 4655 39806 4707 39858
rect 4720 39806 4772 39858
rect 4785 39806 4837 39858
rect 4850 39806 4902 39858
rect 4915 39806 4967 39858
rect 4980 39806 5032 39858
rect 5045 39806 5097 39858
rect 5110 39806 5162 39858
rect 5175 39806 5227 39858
rect 5240 39806 5292 39858
rect 5305 39806 5357 39858
rect 5370 39806 5422 39858
rect 5435 39806 5487 39858
rect 5500 39806 5552 39858
rect 5565 39806 5617 39858
rect 5630 39806 5682 39858
rect 5695 39806 5747 39858
rect 5760 39806 5812 39858
rect 5825 39806 5877 39858
rect 5890 39806 5942 39858
rect 5955 39806 6007 39858
rect 6020 39806 6072 39858
rect 6085 39806 6137 39858
rect 6150 39806 6202 39858
rect 6215 39806 6267 39858
rect 6280 39806 6332 39858
rect 6345 39806 6397 39858
rect 6410 39806 6462 39858
rect 6475 39806 6527 39858
rect 6540 39806 6592 39858
rect 6605 39806 6657 39858
rect 6670 39806 6722 39858
rect 6735 39806 6787 39858
rect 6800 39806 6852 39858
rect 6865 39806 6917 39858
rect 6930 39806 6982 39858
rect 6995 39806 7047 39858
rect 7060 39806 7112 39858
rect 7125 39806 7177 39858
rect 7189 39806 7241 39858
rect 7253 39806 7305 39858
rect 7317 39806 7369 39858
rect 7381 39806 7433 39858
rect 7445 39806 7497 39858
rect 7509 39806 7561 39858
rect 7573 39806 7625 39858
rect 7637 39806 7689 39858
rect 7701 39806 7753 39858
rect 7765 39806 7817 39858
rect 7829 39806 7881 39858
rect 7893 39806 7945 39858
rect 7957 39806 8009 39858
rect 8021 39806 8073 39858
rect 8085 39806 8137 39858
rect 8149 39806 8201 39858
rect 8213 39806 8265 39858
rect 8277 39806 8329 39858
rect 8341 39806 8393 39858
rect 8405 39806 8457 39858
rect 8469 39806 8521 39858
rect 8533 39806 8585 39858
rect 8597 39806 8649 39858
rect 8661 39806 8713 39858
rect 8725 39806 8777 39858
rect 8789 39806 8841 39858
rect 8853 39806 8905 39858
rect 8917 39806 8969 39858
rect 8981 39806 9033 39858
rect 9045 39806 9097 39858
rect 9109 39806 9161 39858
rect 9173 39806 9225 39858
rect 9237 39806 9289 39858
rect 9301 39806 9353 39858
rect 9365 39806 9417 39858
rect 9429 39806 9481 39858
rect 9493 39806 9545 39858
rect 9557 39806 9609 39858
rect 9621 39806 9673 39858
rect 9685 39806 9737 39858
rect 9749 39806 9801 39858
rect 9813 39806 9865 39858
rect 9877 39806 9929 39858
rect 9941 39806 9993 39858
rect 10005 39806 10057 39858
rect 10069 39806 10121 39858
rect 10133 39806 10185 39858
rect 10197 39806 10249 39858
rect 10261 39806 10313 39858
rect 10325 39806 10377 39858
rect 10389 39806 10441 39858
rect 10453 39806 10505 39858
rect 10517 39806 10569 39858
rect 10581 39806 10633 39858
rect 10645 39806 10697 39858
rect 10709 39806 10761 39858
rect 10773 39806 10825 39858
rect 10837 39806 10889 39858
rect 10901 39806 10953 39858
rect 10965 39806 11017 39858
rect 11029 39806 11081 39858
rect 11093 39806 11145 39858
rect 11157 39806 11209 39858
rect 11221 39806 11273 39858
rect 11285 39806 11337 39858
rect 3160 39738 3212 39790
rect 3225 39738 3277 39790
rect 3290 39738 3342 39790
rect 3355 39738 3407 39790
rect 3420 39738 3472 39790
rect 3485 39738 3537 39790
rect 3550 39738 3602 39790
rect 3615 39738 3667 39790
rect 3680 39738 3732 39790
rect 3745 39738 3797 39790
rect 3810 39738 3862 39790
rect 3875 39738 3927 39790
rect 3940 39738 3992 39790
rect 4005 39738 4057 39790
rect 4070 39738 4122 39790
rect 4135 39738 4187 39790
rect 4200 39738 4252 39790
rect 4265 39738 4317 39790
rect 4330 39738 4382 39790
rect 4395 39738 4447 39790
rect 4460 39738 4512 39790
rect 4525 39738 4577 39790
rect 4590 39738 4642 39790
rect 4655 39738 4707 39790
rect 4720 39738 4772 39790
rect 4785 39738 4837 39790
rect 4850 39738 4902 39790
rect 4915 39738 4967 39790
rect 4980 39738 5032 39790
rect 5045 39738 5097 39790
rect 5110 39738 5162 39790
rect 5175 39738 5227 39790
rect 5240 39738 5292 39790
rect 5305 39738 5357 39790
rect 5370 39738 5422 39790
rect 5435 39738 5487 39790
rect 5500 39738 5552 39790
rect 5565 39738 5617 39790
rect 5630 39738 5682 39790
rect 5695 39738 5747 39790
rect 5760 39738 5812 39790
rect 5825 39738 5877 39790
rect 5890 39738 5942 39790
rect 5955 39738 6007 39790
rect 6020 39738 6072 39790
rect 6085 39738 6137 39790
rect 6150 39738 6202 39790
rect 6215 39738 6267 39790
rect 6280 39738 6332 39790
rect 6345 39738 6397 39790
rect 6410 39738 6462 39790
rect 6475 39738 6527 39790
rect 6540 39738 6592 39790
rect 6605 39738 6657 39790
rect 6670 39738 6722 39790
rect 6735 39738 6787 39790
rect 6800 39738 6852 39790
rect 6865 39738 6917 39790
rect 6930 39738 6982 39790
rect 6995 39738 7047 39790
rect 7060 39738 7112 39790
rect 7125 39738 7177 39790
rect 7189 39738 7241 39790
rect 7253 39738 7305 39790
rect 7317 39738 7369 39790
rect 7381 39738 7433 39790
rect 7445 39738 7497 39790
rect 7509 39738 7561 39790
rect 7573 39738 7625 39790
rect 7637 39738 7689 39790
rect 7701 39738 7753 39790
rect 7765 39738 7817 39790
rect 7829 39738 7881 39790
rect 7893 39738 7945 39790
rect 7957 39738 8009 39790
rect 8021 39738 8073 39790
rect 8085 39738 8137 39790
rect 8149 39738 8201 39790
rect 8213 39738 8265 39790
rect 8277 39738 8329 39790
rect 8341 39738 8393 39790
rect 8405 39738 8457 39790
rect 8469 39738 8521 39790
rect 8533 39738 8585 39790
rect 8597 39738 8649 39790
rect 8661 39738 8713 39790
rect 8725 39738 8777 39790
rect 8789 39738 8841 39790
rect 8853 39738 8905 39790
rect 8917 39738 8969 39790
rect 8981 39738 9033 39790
rect 9045 39738 9097 39790
rect 9109 39738 9161 39790
rect 9173 39738 9225 39790
rect 9237 39738 9289 39790
rect 9301 39738 9353 39790
rect 9365 39738 9417 39790
rect 9429 39738 9481 39790
rect 9493 39738 9545 39790
rect 9557 39738 9609 39790
rect 9621 39738 9673 39790
rect 9685 39738 9737 39790
rect 9749 39738 9801 39790
rect 9813 39738 9865 39790
rect 9877 39738 9929 39790
rect 9941 39738 9993 39790
rect 10005 39738 10057 39790
rect 10069 39738 10121 39790
rect 10133 39738 10185 39790
rect 10197 39738 10249 39790
rect 10261 39738 10313 39790
rect 10325 39738 10377 39790
rect 10389 39738 10441 39790
rect 10453 39738 10505 39790
rect 10517 39738 10569 39790
rect 10581 39738 10633 39790
rect 10645 39738 10697 39790
rect 10709 39738 10761 39790
rect 10773 39738 10825 39790
rect 10837 39738 10889 39790
rect 10901 39738 10953 39790
rect 10965 39738 11017 39790
rect 11029 39738 11081 39790
rect 11093 39738 11145 39790
rect 11157 39738 11209 39790
rect 11221 39738 11273 39790
rect 11285 39738 11337 39790
rect 14405 39946 14457 39998
rect 14470 39946 14522 39998
rect 14535 39946 14587 39998
rect 14600 39946 14652 39998
rect 14665 39946 14717 39998
rect 14730 39946 14782 39998
rect 14795 39946 14847 39998
rect 14860 39946 14912 39998
rect 14925 39946 14977 39998
rect 14990 39946 15042 39998
rect 15055 39946 15107 39998
rect 15120 39946 15172 39998
rect 15185 39946 15237 39998
rect 15249 39946 15301 39998
rect 15313 39946 15365 39998
rect 14405 39878 14457 39930
rect 14470 39878 14522 39930
rect 14535 39878 14587 39930
rect 14600 39878 14652 39930
rect 14665 39878 14717 39930
rect 14730 39878 14782 39930
rect 14795 39878 14847 39930
rect 14860 39878 14912 39930
rect 14925 39878 14977 39930
rect 14990 39878 15042 39930
rect 15055 39878 15107 39930
rect 15120 39878 15172 39930
rect 15185 39878 15237 39930
rect 15249 39878 15301 39930
rect 15313 39878 15365 39930
rect 14405 39810 14457 39862
rect 14470 39810 14522 39862
rect 14535 39810 14587 39862
rect 14600 39810 14652 39862
rect 14665 39810 14717 39862
rect 14730 39810 14782 39862
rect 14795 39810 14847 39862
rect 14860 39810 14912 39862
rect 14925 39810 14977 39862
rect 14990 39810 15042 39862
rect 15055 39810 15107 39862
rect 15120 39810 15172 39862
rect 15185 39810 15237 39862
rect 15249 39810 15301 39862
rect 15313 39810 15365 39862
rect 14405 39742 14457 39794
rect 14470 39742 14522 39794
rect 14535 39742 14587 39794
rect 14600 39742 14652 39794
rect 14665 39742 14717 39794
rect 14730 39742 14782 39794
rect 14795 39742 14847 39794
rect 14860 39742 14912 39794
rect 14925 39742 14977 39794
rect 14990 39742 15042 39794
rect 15055 39742 15107 39794
rect 15120 39742 15172 39794
rect 15185 39742 15237 39794
rect 15249 39742 15301 39794
rect 15313 39742 15365 39794
rect 2792 36027 2844 36079
rect 2858 36027 2910 36079
rect 2924 36027 2976 36079
rect 2990 36027 3042 36079
rect 3056 36027 3108 36079
rect 3122 36027 3174 36079
rect 3188 36027 3240 36079
rect 3254 36027 3306 36079
rect 3320 36027 3372 36079
rect 3386 36027 3438 36079
rect 3452 36027 3504 36079
rect 3518 36027 3570 36079
rect 3584 36027 3636 36079
rect 3650 36027 3702 36079
rect 3715 36027 3767 36079
rect 2792 35949 2844 36001
rect 2858 35949 2910 36001
rect 2924 35949 2976 36001
rect 2990 35949 3042 36001
rect 3056 35949 3108 36001
rect 3122 35996 3174 36001
rect 3188 35996 3240 36001
rect 3254 35996 3306 36001
rect 3320 35996 3372 36001
rect 3386 35996 3438 36001
rect 3452 35996 3504 36001
rect 3122 35962 3157 35996
rect 3157 35962 3174 35996
rect 3188 35962 3191 35996
rect 3191 35962 3230 35996
rect 3230 35962 3240 35996
rect 3254 35962 3264 35996
rect 3264 35962 3303 35996
rect 3303 35962 3306 35996
rect 3320 35962 3337 35996
rect 3337 35962 3372 35996
rect 3386 35962 3410 35996
rect 3410 35962 3438 35996
rect 3452 35962 3483 35996
rect 3483 35962 3504 35996
rect 3122 35949 3174 35962
rect 3188 35949 3240 35962
rect 3254 35949 3306 35962
rect 3320 35949 3372 35962
rect 3386 35949 3438 35962
rect 3452 35949 3504 35962
rect 3518 35996 3570 36001
rect 3518 35962 3522 35996
rect 3522 35962 3556 35996
rect 3556 35962 3570 35996
rect 3518 35949 3570 35962
rect 3584 35996 3636 36001
rect 3584 35962 3595 35996
rect 3595 35962 3629 35996
rect 3629 35962 3636 35996
rect 3584 35949 3636 35962
rect 3650 35996 3702 36001
rect 3650 35962 3668 35996
rect 3668 35962 3702 35996
rect 3650 35949 3702 35962
rect 3715 35996 3767 36001
rect 3715 35962 3741 35996
rect 3741 35962 3767 35996
rect 3715 35949 3767 35962
rect 2792 35871 2844 35923
rect 2858 35871 2910 35923
rect 2924 35871 2976 35923
rect 2990 35871 3042 35923
rect 3056 35871 3108 35923
rect 3122 35890 3157 35923
rect 3157 35890 3174 35923
rect 3188 35890 3191 35923
rect 3191 35890 3230 35923
rect 3230 35890 3240 35923
rect 3254 35890 3264 35923
rect 3264 35890 3303 35923
rect 3303 35890 3306 35923
rect 3320 35890 3337 35923
rect 3337 35890 3372 35923
rect 3386 35890 3410 35923
rect 3410 35890 3438 35923
rect 3452 35890 3483 35923
rect 3483 35890 3504 35923
rect 3122 35871 3174 35890
rect 3188 35871 3240 35890
rect 3254 35871 3306 35890
rect 3320 35871 3372 35890
rect 3386 35871 3438 35890
rect 3452 35871 3504 35890
rect 3518 35890 3522 35923
rect 3522 35890 3556 35923
rect 3556 35890 3570 35923
rect 3518 35871 3570 35890
rect 3584 35890 3595 35923
rect 3595 35890 3629 35923
rect 3629 35890 3636 35923
rect 3584 35871 3636 35890
rect 3650 35890 3668 35923
rect 3668 35890 3702 35923
rect 3650 35871 3702 35890
rect 3715 35890 3741 35923
rect 3741 35890 3767 35923
rect 3715 35871 3767 35890
rect 2792 35793 2844 35845
rect 2858 35793 2910 35845
rect 2924 35793 2976 35845
rect 2990 35793 3042 35845
rect 3056 35793 3108 35845
rect 3122 35793 3174 35845
rect 3188 35793 3240 35845
rect 3254 35793 3306 35845
rect 3320 35793 3372 35845
rect 3386 35793 3438 35845
rect 3452 35793 3504 35845
rect 3518 35793 3570 35845
rect 3584 35793 3636 35845
rect 3650 35793 3702 35845
rect 3715 35793 3767 35845
rect 454 35648 506 35674
rect 528 35648 580 35674
rect 602 35648 654 35674
rect 454 35622 463 35648
rect 463 35622 506 35648
rect 528 35622 580 35648
rect 602 35622 654 35648
rect 454 35558 463 35610
rect 463 35558 506 35610
rect 528 35558 580 35610
rect 602 35558 654 35610
rect 454 35494 463 35546
rect 463 35494 506 35546
rect 528 35494 580 35546
rect 602 35494 654 35546
rect 454 35430 463 35482
rect 463 35430 506 35482
rect 528 35430 580 35482
rect 602 35430 654 35482
rect 454 35366 463 35418
rect 463 35366 506 35418
rect 528 35366 580 35418
rect 602 35366 654 35418
rect 454 35302 463 35354
rect 463 35302 506 35354
rect 528 35302 580 35354
rect 602 35302 654 35354
rect 454 35238 463 35290
rect 463 35238 506 35290
rect 528 35238 580 35290
rect 602 35238 654 35290
rect 454 35174 463 35226
rect 463 35174 506 35226
rect 528 35174 580 35226
rect 602 35174 654 35226
rect 454 35110 463 35162
rect 463 35110 506 35162
rect 528 35110 580 35162
rect 602 35110 654 35162
rect 454 35046 463 35098
rect 463 35046 506 35098
rect 528 35046 580 35098
rect 602 35046 654 35098
rect 454 34982 463 35034
rect 463 34982 506 35034
rect 528 34982 580 35034
rect 602 34982 654 35034
rect 454 34918 463 34970
rect 463 34918 506 34970
rect 528 34918 580 34970
rect 602 34918 654 34970
rect 454 34854 463 34906
rect 463 34854 506 34906
rect 528 34854 580 34906
rect 602 34854 654 34906
rect 454 34790 463 34842
rect 463 34790 506 34842
rect 528 34790 580 34842
rect 602 34790 654 34842
rect 454 34726 463 34778
rect 463 34726 506 34778
rect 528 34726 580 34778
rect 602 34726 654 34778
rect 454 34662 463 34714
rect 463 34662 506 34714
rect 528 34662 580 34714
rect 602 34662 654 34714
rect 454 34598 463 34650
rect 463 34598 506 34650
rect 528 34598 580 34650
rect 602 34598 654 34650
rect 454 34534 463 34586
rect 463 34534 506 34586
rect 528 34534 580 34586
rect 602 34534 654 34586
rect 454 34470 463 34522
rect 463 34470 506 34522
rect 528 34470 580 34522
rect 602 34470 654 34522
rect 454 34406 463 34458
rect 463 34406 506 34458
rect 528 34406 580 34458
rect 602 34406 654 34458
rect 454 34342 463 34394
rect 463 34342 506 34394
rect 528 34342 580 34394
rect 602 34342 654 34394
rect 454 34278 463 34330
rect 463 34278 506 34330
rect 528 34278 580 34330
rect 602 34278 654 34330
rect 454 34246 463 34266
rect 463 34246 506 34266
rect 528 34246 580 34266
rect 602 34246 654 34266
rect 454 34214 506 34246
rect 528 34214 580 34246
rect 602 34214 654 34246
rect 454 34173 463 34202
rect 463 34173 497 34202
rect 497 34173 506 34202
rect 454 34150 506 34173
rect 528 34173 535 34202
rect 535 34173 569 34202
rect 569 34173 580 34202
rect 528 34150 580 34173
rect 602 34173 607 34202
rect 607 34173 641 34202
rect 641 34173 654 34202
rect 602 34150 654 34173
rect 454 34134 506 34138
rect 454 34100 463 34134
rect 463 34100 497 34134
rect 497 34100 506 34134
rect 454 34086 506 34100
rect 528 34134 580 34138
rect 528 34100 535 34134
rect 535 34100 569 34134
rect 569 34100 580 34134
rect 528 34086 580 34100
rect 602 34134 654 34138
rect 602 34100 607 34134
rect 607 34100 641 34134
rect 641 34100 654 34134
rect 602 34086 654 34100
rect 454 34061 506 34074
rect 454 34027 463 34061
rect 463 34027 497 34061
rect 497 34027 506 34061
rect 454 34022 506 34027
rect 528 34061 580 34074
rect 528 34027 535 34061
rect 535 34027 569 34061
rect 569 34027 580 34061
rect 528 34022 580 34027
rect 602 34061 654 34074
rect 602 34027 607 34061
rect 607 34027 641 34061
rect 641 34027 654 34061
rect 602 34022 654 34027
rect 149 33986 201 34012
rect 149 33960 167 33986
rect 167 33960 201 33986
rect 247 33986 299 34012
rect 247 33960 259 33986
rect 259 33960 293 33986
rect 293 33960 299 33986
rect 149 33914 201 33948
rect 149 33896 167 33914
rect 167 33896 201 33914
rect 247 33914 299 33948
rect 247 33896 259 33914
rect 259 33896 293 33914
rect 293 33896 299 33914
rect 149 33880 167 33884
rect 167 33880 201 33884
rect 149 33842 201 33880
rect 149 33832 167 33842
rect 167 33832 201 33842
rect 247 33880 259 33884
rect 259 33880 293 33884
rect 293 33880 299 33884
rect 247 33842 299 33880
rect 247 33832 259 33842
rect 259 33832 293 33842
rect 293 33832 299 33842
rect 149 33808 167 33820
rect 167 33808 201 33820
rect 149 33769 201 33808
rect 149 33768 167 33769
rect 167 33768 201 33769
rect 247 33808 259 33820
rect 259 33808 293 33820
rect 293 33808 299 33820
rect 247 33769 299 33808
rect 247 33768 259 33769
rect 259 33768 293 33769
rect 293 33768 299 33769
rect 149 33735 167 33756
rect 167 33735 201 33756
rect 149 33704 201 33735
rect 247 33735 259 33756
rect 259 33735 293 33756
rect 293 33735 299 33756
rect 247 33704 299 33735
rect 149 33662 167 33692
rect 167 33662 201 33692
rect 149 33640 201 33662
rect 247 33662 259 33692
rect 259 33662 293 33692
rect 293 33662 299 33692
rect 247 33640 299 33662
rect 149 33623 201 33628
rect 149 33589 167 33623
rect 167 33589 201 33623
rect 149 33576 201 33589
rect 247 33623 299 33628
rect 247 33589 259 33623
rect 259 33589 293 33623
rect 293 33589 299 33623
rect 247 33576 299 33589
rect 149 33550 201 33564
rect 149 33516 167 33550
rect 167 33516 201 33550
rect 149 33512 201 33516
rect 247 33550 299 33564
rect 247 33516 259 33550
rect 259 33516 293 33550
rect 293 33516 299 33550
rect 247 33512 299 33516
rect 149 33477 201 33500
rect 149 33448 167 33477
rect 167 33448 201 33477
rect 247 33477 299 33500
rect 247 33448 259 33477
rect 259 33448 293 33477
rect 293 33448 299 33477
rect 149 33404 201 33436
rect 149 33384 167 33404
rect 167 33384 201 33404
rect 247 33404 299 33436
rect 247 33384 259 33404
rect 259 33384 293 33404
rect 293 33384 299 33404
rect 149 33370 167 33372
rect 167 33370 201 33372
rect 149 33331 201 33370
rect 149 33320 167 33331
rect 167 33320 201 33331
rect 247 33370 259 33372
rect 259 33370 293 33372
rect 293 33370 299 33372
rect 247 33331 299 33370
rect 247 33320 259 33331
rect 259 33320 293 33331
rect 293 33320 299 33331
rect 149 33297 167 33308
rect 167 33297 201 33308
rect 149 33258 201 33297
rect 149 33256 167 33258
rect 167 33256 201 33258
rect 247 33297 259 33308
rect 259 33297 293 33308
rect 293 33297 299 33308
rect 247 33258 299 33297
rect 247 33256 259 33258
rect 259 33256 293 33258
rect 293 33256 299 33258
rect 149 33224 167 33244
rect 167 33224 201 33244
rect 149 33192 201 33224
rect 247 33224 259 33244
rect 259 33224 293 33244
rect 293 33224 299 33244
rect 247 33192 299 33224
rect 149 33151 167 33180
rect 167 33151 201 33180
rect 149 33128 201 33151
rect 247 33151 259 33180
rect 259 33151 293 33180
rect 293 33151 299 33180
rect 247 33128 299 33151
rect 149 33112 201 33116
rect 149 33078 167 33112
rect 167 33078 201 33112
rect 149 33064 201 33078
rect 247 33112 299 33116
rect 247 33078 259 33112
rect 259 33078 293 33112
rect 293 33078 299 33112
rect 247 33064 299 33078
rect 149 33039 201 33052
rect 149 33005 167 33039
rect 167 33005 201 33039
rect 149 33000 201 33005
rect 247 33039 299 33052
rect 247 33005 259 33039
rect 259 33005 293 33039
rect 293 33005 299 33039
rect 247 33000 299 33005
rect 149 32966 201 32988
rect 149 32936 167 32966
rect 167 32936 201 32966
rect 247 32966 299 32988
rect 247 32936 259 32966
rect 259 32936 293 32966
rect 293 32936 299 32966
rect 149 32893 201 32924
rect 149 32872 167 32893
rect 167 32872 201 32893
rect 247 32893 299 32924
rect 247 32872 259 32893
rect 259 32872 293 32893
rect 293 32872 299 32893
rect 149 32820 201 32859
rect 149 32807 167 32820
rect 167 32807 201 32820
rect 247 32820 299 32859
rect 247 32807 259 32820
rect 259 32807 293 32820
rect 293 32807 299 32820
rect 149 32786 167 32794
rect 167 32786 201 32794
rect 149 32747 201 32786
rect 149 32742 167 32747
rect 167 32742 201 32747
rect 247 32786 259 32794
rect 259 32786 293 32794
rect 293 32786 299 32794
rect 247 32747 299 32786
rect 247 32742 259 32747
rect 259 32742 293 32747
rect 293 32742 299 32747
rect 149 32713 167 32729
rect 167 32713 201 32729
rect 149 32677 201 32713
rect 247 32713 259 32729
rect 259 32713 293 32729
rect 293 32713 299 32729
rect 247 32677 299 32713
rect 149 32640 167 32664
rect 167 32640 201 32664
rect 149 32612 201 32640
rect 247 32640 259 32664
rect 259 32640 293 32664
rect 293 32640 299 32664
rect 247 32612 299 32640
rect 149 32567 167 32599
rect 167 32567 201 32599
rect 149 32547 201 32567
rect 247 32567 259 32599
rect 259 32567 293 32599
rect 293 32567 299 32599
rect 247 32547 299 32567
rect 149 32528 201 32534
rect 149 32494 167 32528
rect 167 32494 201 32528
rect 149 32482 201 32494
rect 247 32528 299 32534
rect 247 32494 259 32528
rect 259 32494 293 32528
rect 293 32494 299 32528
rect 247 32482 299 32494
rect 149 32455 201 32469
rect 149 32421 167 32455
rect 167 32421 201 32455
rect 149 32417 201 32421
rect 247 32455 299 32469
rect 247 32421 259 32455
rect 259 32421 293 32455
rect 293 32421 299 32455
rect 247 32417 299 32421
rect 149 32382 201 32404
rect 149 32352 167 32382
rect 167 32352 201 32382
rect 247 32382 299 32404
rect 247 32352 259 32382
rect 259 32352 293 32382
rect 293 32352 299 32382
rect 149 32309 201 32339
rect 149 32287 167 32309
rect 167 32287 201 32309
rect 247 32309 299 32339
rect 247 32287 259 32309
rect 259 32287 293 32309
rect 293 32287 299 32309
rect 149 32236 201 32274
rect 149 32222 167 32236
rect 167 32222 201 32236
rect 247 32236 299 32274
rect 247 32222 259 32236
rect 259 32222 293 32236
rect 293 32222 299 32236
rect 149 32202 167 32209
rect 167 32202 201 32209
rect 149 32163 201 32202
rect 149 32157 167 32163
rect 167 32157 201 32163
rect 247 32202 259 32209
rect 259 32202 293 32209
rect 293 32202 299 32209
rect 247 32163 299 32202
rect 247 32157 259 32163
rect 259 32157 293 32163
rect 293 32157 299 32163
rect 149 32129 167 32144
rect 167 32129 201 32144
rect 149 32092 201 32129
rect 247 32129 259 32144
rect 259 32129 293 32144
rect 293 32129 299 32144
rect 247 32092 299 32129
rect 149 32056 167 32079
rect 167 32056 201 32079
rect 149 32027 201 32056
rect 247 32056 259 32079
rect 259 32056 293 32079
rect 293 32056 299 32079
rect 247 32027 299 32056
rect 149 31983 167 32014
rect 167 31983 201 32014
rect 149 31962 201 31983
rect 247 31983 259 32014
rect 259 31983 293 32014
rect 293 31983 299 32014
rect 247 31962 299 31983
rect 149 31944 201 31949
rect 149 31910 167 31944
rect 167 31910 201 31944
rect 149 31897 201 31910
rect 247 31944 299 31949
rect 247 31910 259 31944
rect 259 31910 293 31944
rect 293 31910 299 31944
rect 247 31897 299 31910
rect 149 31871 201 31884
rect 149 31837 167 31871
rect 167 31837 201 31871
rect 149 31832 201 31837
rect 247 31871 299 31884
rect 247 31837 259 31871
rect 259 31837 293 31871
rect 293 31837 299 31871
rect 247 31832 299 31837
rect 149 31798 201 31819
rect 149 31767 167 31798
rect 167 31767 201 31798
rect 247 31798 299 31819
rect 247 31767 259 31798
rect 259 31767 293 31798
rect 293 31767 299 31798
rect 149 31725 201 31754
rect 149 31702 167 31725
rect 167 31702 201 31725
rect 247 31725 299 31754
rect 247 31702 259 31725
rect 259 31702 293 31725
rect 293 31702 299 31725
rect 149 31652 201 31689
rect 149 31637 167 31652
rect 167 31637 201 31652
rect 247 31652 299 31689
rect 247 31637 259 31652
rect 259 31637 293 31652
rect 293 31637 299 31652
rect 149 31618 167 31624
rect 167 31618 201 31624
rect 149 31579 201 31618
rect 149 31572 167 31579
rect 167 31572 201 31579
rect 247 31618 259 31624
rect 259 31618 293 31624
rect 293 31618 299 31624
rect 247 31579 299 31618
rect 247 31572 259 31579
rect 259 31572 293 31579
rect 293 31572 299 31579
rect 149 31545 167 31559
rect 167 31545 201 31559
rect 149 31507 201 31545
rect 247 31545 259 31559
rect 259 31545 293 31559
rect 293 31545 299 31559
rect 247 31507 299 31545
rect 149 31472 167 31494
rect 167 31472 201 31494
rect 149 31442 201 31472
rect 247 31472 259 31494
rect 259 31472 293 31494
rect 293 31472 299 31494
rect 247 31442 299 31472
rect 149 31399 167 31429
rect 167 31399 201 31429
rect 149 31377 201 31399
rect 247 31399 259 31429
rect 259 31399 293 31429
rect 293 31399 299 31429
rect 247 31377 299 31399
rect 149 31360 201 31364
rect 149 31326 167 31360
rect 167 31326 201 31360
rect 149 31312 201 31326
rect 247 31360 299 31364
rect 247 31326 259 31360
rect 259 31326 293 31360
rect 293 31326 299 31360
rect 247 31312 299 31326
rect 149 31287 201 31299
rect 149 31253 167 31287
rect 167 31253 201 31287
rect 149 31247 201 31253
rect 247 31287 299 31299
rect 247 31253 259 31287
rect 259 31253 293 31287
rect 293 31253 299 31287
rect 247 31247 299 31253
rect 149 31214 201 31234
rect 149 31182 167 31214
rect 167 31182 201 31214
rect 247 31214 299 31234
rect 247 31182 259 31214
rect 259 31182 293 31214
rect 293 31182 299 31214
rect 149 31141 201 31169
rect 149 31117 167 31141
rect 167 31117 201 31141
rect 247 31141 299 31169
rect 247 31117 259 31141
rect 259 31117 293 31141
rect 293 31117 299 31141
rect 149 31068 201 31104
rect 149 31052 167 31068
rect 167 31052 201 31068
rect 247 31068 299 31104
rect 247 31052 259 31068
rect 259 31052 293 31068
rect 293 31052 299 31068
rect 149 31034 167 31039
rect 167 31034 201 31039
rect 149 30995 201 31034
rect 149 30987 167 30995
rect 167 30987 201 30995
rect 247 31034 259 31039
rect 259 31034 293 31039
rect 293 31034 299 31039
rect 247 30995 299 31034
rect 247 30987 259 30995
rect 259 30987 293 30995
rect 293 30987 299 30995
rect 149 30961 167 30974
rect 167 30961 201 30974
rect 149 30922 201 30961
rect 247 30961 259 30974
rect 259 30961 293 30974
rect 293 30961 299 30974
rect 247 30922 299 30961
rect 149 30888 167 30909
rect 167 30888 201 30909
rect 149 30857 201 30888
rect 247 30888 259 30909
rect 259 30888 293 30909
rect 293 30888 299 30909
rect 247 30857 299 30888
rect 149 30815 167 30844
rect 167 30815 201 30844
rect 149 30792 201 30815
rect 247 30815 259 30844
rect 259 30815 293 30844
rect 293 30815 299 30844
rect 247 30792 299 30815
rect 149 30776 201 30779
rect 149 30742 167 30776
rect 167 30742 201 30776
rect 149 30727 201 30742
rect 247 30776 299 30779
rect 247 30742 259 30776
rect 259 30742 293 30776
rect 293 30742 299 30776
rect 247 30727 299 30742
rect 149 30703 201 30714
rect 149 30669 167 30703
rect 167 30669 201 30703
rect 149 30662 201 30669
rect 247 30703 299 30714
rect 247 30669 259 30703
rect 259 30669 293 30703
rect 293 30669 299 30703
rect 247 30662 299 30669
rect 149 30630 201 30649
rect 149 30597 167 30630
rect 167 30597 201 30630
rect 247 30630 299 30649
rect 247 30597 259 30630
rect 259 30597 293 30630
rect 293 30597 299 30630
rect 149 30557 201 30584
rect 149 30532 167 30557
rect 167 30532 201 30557
rect 247 30557 299 30584
rect 247 30532 259 30557
rect 259 30532 293 30557
rect 293 30532 299 30557
rect 149 30484 201 30519
rect 149 30467 167 30484
rect 167 30467 201 30484
rect 247 30484 299 30519
rect 247 30467 259 30484
rect 259 30467 293 30484
rect 293 30467 299 30484
rect 149 30450 167 30454
rect 167 30450 201 30454
rect 149 30411 201 30450
rect 149 30402 167 30411
rect 167 30402 201 30411
rect 247 30450 259 30454
rect 259 30450 293 30454
rect 293 30450 299 30454
rect 247 30411 299 30450
rect 247 30402 259 30411
rect 259 30402 293 30411
rect 293 30402 299 30411
rect 149 30377 167 30389
rect 167 30377 201 30389
rect 149 30338 201 30377
rect 149 30337 167 30338
rect 167 30337 201 30338
rect 247 30377 259 30389
rect 259 30377 293 30389
rect 293 30377 299 30389
rect 247 30338 299 30377
rect 247 30337 259 30338
rect 259 30337 293 30338
rect 293 30337 299 30338
rect 149 30304 167 30324
rect 167 30304 201 30324
rect 149 30272 201 30304
rect 247 30304 259 30324
rect 259 30304 293 30324
rect 293 30304 299 30324
rect 247 30272 299 30304
rect 149 30231 167 30259
rect 167 30231 201 30259
rect 149 30207 201 30231
rect 247 30231 259 30259
rect 259 30231 293 30259
rect 293 30231 299 30259
rect 247 30207 299 30231
rect 149 30192 201 30194
rect 149 30158 167 30192
rect 167 30158 201 30192
rect 149 30142 201 30158
rect 247 30192 299 30194
rect 247 30158 259 30192
rect 259 30158 293 30192
rect 293 30158 299 30192
rect 247 30142 299 30158
rect 149 30119 201 30129
rect 149 30085 167 30119
rect 167 30085 201 30119
rect 149 30077 201 30085
rect 247 30119 299 30129
rect 247 30085 259 30119
rect 259 30085 293 30119
rect 293 30085 299 30119
rect 247 30077 299 30085
rect 149 30046 201 30064
rect 149 30012 167 30046
rect 167 30012 201 30046
rect 247 30046 299 30064
rect 247 30012 259 30046
rect 259 30012 293 30046
rect 293 30012 299 30046
rect 149 29973 201 29999
rect 149 29947 167 29973
rect 167 29947 201 29973
rect 247 29973 299 29999
rect 247 29947 259 29973
rect 259 29947 293 29973
rect 293 29947 299 29973
rect 149 29900 201 29934
rect 149 29882 167 29900
rect 167 29882 201 29900
rect 247 29900 299 29934
rect 247 29882 259 29900
rect 259 29882 293 29900
rect 293 29882 299 29900
rect 149 29866 167 29869
rect 167 29866 201 29869
rect 149 29827 201 29866
rect 149 29817 167 29827
rect 167 29817 201 29827
rect 247 29866 259 29869
rect 259 29866 293 29869
rect 293 29866 299 29869
rect 247 29827 299 29866
rect 247 29817 259 29827
rect 259 29817 293 29827
rect 293 29817 299 29827
rect 149 29793 167 29804
rect 167 29793 201 29804
rect 149 29754 201 29793
rect 149 29752 167 29754
rect 167 29752 201 29754
rect 247 29793 259 29804
rect 259 29793 293 29804
rect 293 29793 299 29804
rect 247 29754 299 29793
rect 247 29752 259 29754
rect 259 29752 293 29754
rect 293 29752 299 29754
rect 149 29720 167 29739
rect 167 29720 201 29739
rect 149 29687 201 29720
rect 247 29720 259 29739
rect 259 29720 293 29739
rect 293 29720 299 29739
rect 247 29687 299 29720
rect 149 29647 167 29674
rect 167 29647 201 29674
rect 149 29622 201 29647
rect 247 29647 259 29674
rect 259 29647 293 29674
rect 293 29647 299 29674
rect 247 29622 299 29647
rect 149 29608 201 29609
rect 149 29574 167 29608
rect 167 29574 201 29608
rect 149 29557 201 29574
rect 247 29608 299 29609
rect 247 29574 259 29608
rect 259 29574 293 29608
rect 293 29574 299 29608
rect 247 29557 299 29574
rect 149 29535 201 29544
rect 149 29501 167 29535
rect 167 29501 201 29535
rect 149 29492 201 29501
rect 247 29535 299 29544
rect 247 29501 259 29535
rect 259 29501 293 29535
rect 293 29501 299 29535
rect 247 29492 299 29501
rect 149 29462 201 29479
rect 149 29428 167 29462
rect 167 29428 201 29462
rect 149 29427 201 29428
rect 247 29462 299 29479
rect 247 29428 259 29462
rect 259 29428 293 29462
rect 293 29428 299 29462
rect 247 29427 299 29428
rect 149 29389 201 29414
rect 149 29362 167 29389
rect 167 29362 201 29389
rect 247 29389 299 29414
rect 247 29362 259 29389
rect 259 29362 293 29389
rect 293 29362 299 29389
rect 149 29316 201 29349
rect 149 29297 167 29316
rect 167 29297 201 29316
rect 247 29316 299 29349
rect 247 29297 259 29316
rect 259 29297 293 29316
rect 293 29297 299 29316
rect 149 29282 167 29284
rect 167 29282 201 29284
rect 149 29243 201 29282
rect 149 29232 167 29243
rect 167 29232 201 29243
rect 247 29282 259 29284
rect 259 29282 293 29284
rect 293 29282 299 29284
rect 247 29243 299 29282
rect 247 29232 259 29243
rect 259 29232 293 29243
rect 293 29232 299 29243
rect 149 29209 167 29219
rect 167 29209 201 29219
rect 149 29170 201 29209
rect 149 29167 167 29170
rect 167 29167 201 29170
rect 247 29209 259 29219
rect 259 29209 293 29219
rect 293 29209 299 29219
rect 247 29170 299 29209
rect 247 29167 259 29170
rect 259 29167 293 29170
rect 293 29167 299 29170
rect 149 29136 167 29154
rect 167 29136 201 29154
rect 149 29102 201 29136
rect 247 29136 259 29154
rect 259 29136 293 29154
rect 293 29136 299 29154
rect 247 29102 299 29136
rect 149 29063 167 29089
rect 167 29063 201 29089
rect 149 29037 201 29063
rect 247 29063 259 29089
rect 259 29063 293 29089
rect 293 29063 299 29089
rect 247 29037 299 29063
rect 454 33988 506 34010
rect 454 33958 463 33988
rect 463 33958 497 33988
rect 497 33958 506 33988
rect 528 33988 580 34010
rect 528 33958 535 33988
rect 535 33958 569 33988
rect 569 33958 580 33988
rect 602 33988 654 34010
rect 602 33958 607 33988
rect 607 33958 641 33988
rect 641 33958 654 33988
rect 454 33915 506 33946
rect 454 33894 463 33915
rect 463 33894 497 33915
rect 497 33894 506 33915
rect 528 33915 580 33946
rect 528 33894 535 33915
rect 535 33894 569 33915
rect 569 33894 580 33915
rect 602 33915 654 33946
rect 602 33894 607 33915
rect 607 33894 641 33915
rect 641 33894 654 33915
rect 454 33881 463 33882
rect 463 33881 497 33882
rect 497 33881 506 33882
rect 454 33842 506 33881
rect 454 33830 463 33842
rect 463 33830 497 33842
rect 497 33830 506 33842
rect 528 33881 535 33882
rect 535 33881 569 33882
rect 569 33881 580 33882
rect 528 33842 580 33881
rect 528 33830 535 33842
rect 535 33830 569 33842
rect 569 33830 580 33842
rect 602 33881 607 33882
rect 607 33881 641 33882
rect 641 33881 654 33882
rect 602 33842 654 33881
rect 602 33830 607 33842
rect 607 33830 641 33842
rect 641 33830 654 33842
rect 454 33808 463 33818
rect 463 33808 497 33818
rect 497 33808 506 33818
rect 454 33769 506 33808
rect 454 33766 463 33769
rect 463 33766 497 33769
rect 497 33766 506 33769
rect 528 33808 535 33818
rect 535 33808 569 33818
rect 569 33808 580 33818
rect 528 33769 580 33808
rect 528 33766 535 33769
rect 535 33766 569 33769
rect 569 33766 580 33769
rect 602 33808 607 33818
rect 607 33808 641 33818
rect 641 33808 654 33818
rect 602 33769 654 33808
rect 602 33766 607 33769
rect 607 33766 641 33769
rect 641 33766 654 33769
rect 454 33735 463 33754
rect 463 33735 497 33754
rect 497 33735 506 33754
rect 454 33702 506 33735
rect 528 33735 535 33754
rect 535 33735 569 33754
rect 569 33735 580 33754
rect 528 33702 580 33735
rect 602 33735 607 33754
rect 607 33735 641 33754
rect 641 33735 654 33754
rect 602 33702 654 33735
rect 454 33662 463 33690
rect 463 33662 497 33690
rect 497 33662 506 33690
rect 454 33638 506 33662
rect 528 33662 535 33690
rect 535 33662 569 33690
rect 569 33662 580 33690
rect 528 33638 580 33662
rect 602 33662 607 33690
rect 607 33662 641 33690
rect 641 33662 654 33690
rect 602 33638 654 33662
rect 454 33623 506 33626
rect 454 33589 463 33623
rect 463 33589 497 33623
rect 497 33589 506 33623
rect 454 33574 506 33589
rect 528 33623 580 33626
rect 528 33589 535 33623
rect 535 33589 569 33623
rect 569 33589 580 33623
rect 528 33574 580 33589
rect 602 33623 654 33626
rect 602 33589 607 33623
rect 607 33589 641 33623
rect 641 33589 654 33623
rect 602 33574 654 33589
rect 454 33550 506 33562
rect 454 33516 463 33550
rect 463 33516 497 33550
rect 497 33516 506 33550
rect 454 33510 506 33516
rect 528 33550 580 33562
rect 528 33516 535 33550
rect 535 33516 569 33550
rect 569 33516 580 33550
rect 528 33510 580 33516
rect 602 33550 654 33562
rect 602 33516 607 33550
rect 607 33516 641 33550
rect 641 33516 654 33550
rect 602 33510 654 33516
rect 454 33477 506 33498
rect 454 33446 463 33477
rect 463 33446 497 33477
rect 497 33446 506 33477
rect 528 33477 580 33498
rect 528 33446 535 33477
rect 535 33446 569 33477
rect 569 33446 580 33477
rect 602 33477 654 33498
rect 602 33446 607 33477
rect 607 33446 641 33477
rect 641 33446 654 33477
rect 454 33404 506 33434
rect 454 33382 463 33404
rect 463 33382 497 33404
rect 497 33382 506 33404
rect 528 33404 580 33434
rect 528 33382 535 33404
rect 535 33382 569 33404
rect 569 33382 580 33404
rect 602 33404 654 33434
rect 602 33382 607 33404
rect 607 33382 641 33404
rect 641 33382 654 33404
rect 454 33331 506 33370
rect 454 33318 463 33331
rect 463 33318 497 33331
rect 497 33318 506 33331
rect 528 33331 580 33370
rect 528 33318 535 33331
rect 535 33318 569 33331
rect 569 33318 580 33331
rect 602 33331 654 33370
rect 602 33318 607 33331
rect 607 33318 641 33331
rect 641 33318 654 33331
rect 454 33297 463 33306
rect 463 33297 497 33306
rect 497 33297 506 33306
rect 454 33258 506 33297
rect 454 33254 463 33258
rect 463 33254 497 33258
rect 497 33254 506 33258
rect 528 33297 535 33306
rect 535 33297 569 33306
rect 569 33297 580 33306
rect 528 33258 580 33297
rect 528 33254 535 33258
rect 535 33254 569 33258
rect 569 33254 580 33258
rect 602 33297 607 33306
rect 607 33297 641 33306
rect 641 33297 654 33306
rect 602 33258 654 33297
rect 602 33254 607 33258
rect 607 33254 641 33258
rect 641 33254 654 33258
rect 454 33224 463 33242
rect 463 33224 497 33242
rect 497 33224 506 33242
rect 454 33190 506 33224
rect 528 33224 535 33242
rect 535 33224 569 33242
rect 569 33224 580 33242
rect 528 33190 580 33224
rect 602 33224 607 33242
rect 607 33224 641 33242
rect 641 33224 654 33242
rect 602 33190 654 33224
rect 454 33151 463 33178
rect 463 33151 497 33178
rect 497 33151 506 33178
rect 454 33126 506 33151
rect 528 33151 535 33178
rect 535 33151 569 33178
rect 569 33151 580 33178
rect 528 33126 580 33151
rect 602 33151 607 33178
rect 607 33151 641 33178
rect 641 33151 654 33178
rect 602 33126 654 33151
rect 454 33112 506 33114
rect 454 33078 463 33112
rect 463 33078 497 33112
rect 497 33078 506 33112
rect 454 33062 506 33078
rect 528 33112 580 33114
rect 528 33078 535 33112
rect 535 33078 569 33112
rect 569 33078 580 33112
rect 528 33062 580 33078
rect 602 33112 654 33114
rect 602 33078 607 33112
rect 607 33078 641 33112
rect 641 33078 654 33112
rect 602 33062 654 33078
rect 454 33039 506 33050
rect 454 33005 463 33039
rect 463 33005 497 33039
rect 497 33005 506 33039
rect 454 32998 506 33005
rect 528 33039 580 33050
rect 528 33005 535 33039
rect 535 33005 569 33039
rect 569 33005 580 33039
rect 528 32998 580 33005
rect 602 33039 654 33050
rect 602 33005 607 33039
rect 607 33005 641 33039
rect 641 33005 654 33039
rect 602 32998 654 33005
rect 454 32966 506 32986
rect 454 32934 463 32966
rect 463 32934 497 32966
rect 497 32934 506 32966
rect 528 32966 580 32986
rect 528 32934 535 32966
rect 535 32934 569 32966
rect 569 32934 580 32966
rect 602 32966 654 32986
rect 602 32934 607 32966
rect 607 32934 641 32966
rect 641 32934 654 32966
rect 454 32893 506 32922
rect 454 32870 463 32893
rect 463 32870 497 32893
rect 497 32870 506 32893
rect 528 32893 580 32922
rect 528 32870 535 32893
rect 535 32870 569 32893
rect 569 32870 580 32893
rect 602 32893 654 32922
rect 602 32870 607 32893
rect 607 32870 641 32893
rect 641 32870 654 32893
rect 454 32820 506 32858
rect 454 32806 463 32820
rect 463 32806 497 32820
rect 497 32806 506 32820
rect 528 32820 580 32858
rect 528 32806 535 32820
rect 535 32806 569 32820
rect 569 32806 580 32820
rect 602 32820 654 32858
rect 602 32806 607 32820
rect 607 32806 641 32820
rect 641 32806 654 32820
rect 454 32786 463 32794
rect 463 32786 497 32794
rect 497 32786 506 32794
rect 454 32747 506 32786
rect 454 32742 463 32747
rect 463 32742 497 32747
rect 497 32742 506 32747
rect 528 32786 535 32794
rect 535 32786 569 32794
rect 569 32786 580 32794
rect 528 32747 580 32786
rect 528 32742 535 32747
rect 535 32742 569 32747
rect 569 32742 580 32747
rect 602 32786 607 32794
rect 607 32786 641 32794
rect 641 32786 654 32794
rect 602 32747 654 32786
rect 602 32742 607 32747
rect 607 32742 641 32747
rect 641 32742 654 32747
rect 454 32713 463 32729
rect 463 32713 497 32729
rect 497 32713 506 32729
rect 454 32677 506 32713
rect 528 32713 535 32729
rect 535 32713 569 32729
rect 569 32713 580 32729
rect 528 32677 580 32713
rect 602 32713 607 32729
rect 607 32713 641 32729
rect 641 32713 654 32729
rect 602 32677 654 32713
rect 454 32640 463 32664
rect 463 32640 497 32664
rect 497 32640 506 32664
rect 454 32612 506 32640
rect 528 32640 535 32664
rect 535 32640 569 32664
rect 569 32640 580 32664
rect 528 32612 580 32640
rect 602 32640 607 32664
rect 607 32640 641 32664
rect 641 32640 654 32664
rect 602 32612 654 32640
rect 454 32567 463 32599
rect 463 32567 497 32599
rect 497 32567 506 32599
rect 454 32547 506 32567
rect 528 32567 535 32599
rect 535 32567 569 32599
rect 569 32567 580 32599
rect 528 32547 580 32567
rect 602 32567 607 32599
rect 607 32567 641 32599
rect 641 32567 654 32599
rect 602 32547 654 32567
rect 454 32528 506 32534
rect 454 32494 463 32528
rect 463 32494 497 32528
rect 497 32494 506 32528
rect 454 32482 506 32494
rect 528 32528 580 32534
rect 528 32494 535 32528
rect 535 32494 569 32528
rect 569 32494 580 32528
rect 528 32482 580 32494
rect 602 32528 654 32534
rect 602 32494 607 32528
rect 607 32494 641 32528
rect 641 32494 654 32528
rect 602 32482 654 32494
rect 454 32455 506 32469
rect 454 32421 463 32455
rect 463 32421 497 32455
rect 497 32421 506 32455
rect 454 32417 506 32421
rect 528 32455 580 32469
rect 528 32421 535 32455
rect 535 32421 569 32455
rect 569 32421 580 32455
rect 528 32417 580 32421
rect 602 32455 654 32469
rect 602 32421 607 32455
rect 607 32421 641 32455
rect 641 32421 654 32455
rect 602 32417 654 32421
rect 454 32382 506 32404
rect 454 32352 463 32382
rect 463 32352 497 32382
rect 497 32352 506 32382
rect 528 32382 580 32404
rect 528 32352 535 32382
rect 535 32352 569 32382
rect 569 32352 580 32382
rect 602 32382 654 32404
rect 602 32352 607 32382
rect 607 32352 641 32382
rect 641 32352 654 32382
rect 454 32309 506 32339
rect 454 32287 463 32309
rect 463 32287 497 32309
rect 497 32287 506 32309
rect 528 32309 580 32339
rect 528 32287 535 32309
rect 535 32287 569 32309
rect 569 32287 580 32309
rect 602 32309 654 32339
rect 602 32287 607 32309
rect 607 32287 641 32309
rect 641 32287 654 32309
rect 454 32236 506 32274
rect 454 32222 463 32236
rect 463 32222 497 32236
rect 497 32222 506 32236
rect 528 32236 580 32274
rect 528 32222 535 32236
rect 535 32222 569 32236
rect 569 32222 580 32236
rect 602 32236 654 32274
rect 602 32222 607 32236
rect 607 32222 641 32236
rect 641 32222 654 32236
rect 454 32202 463 32209
rect 463 32202 497 32209
rect 497 32202 506 32209
rect 454 32163 506 32202
rect 454 32157 463 32163
rect 463 32157 497 32163
rect 497 32157 506 32163
rect 528 32202 535 32209
rect 535 32202 569 32209
rect 569 32202 580 32209
rect 528 32163 580 32202
rect 528 32157 535 32163
rect 535 32157 569 32163
rect 569 32157 580 32163
rect 602 32202 607 32209
rect 607 32202 641 32209
rect 641 32202 654 32209
rect 602 32163 654 32202
rect 602 32157 607 32163
rect 607 32157 641 32163
rect 641 32157 654 32163
rect 454 32129 463 32144
rect 463 32129 497 32144
rect 497 32129 506 32144
rect 454 32092 506 32129
rect 528 32129 535 32144
rect 535 32129 569 32144
rect 569 32129 580 32144
rect 528 32092 580 32129
rect 602 32129 607 32144
rect 607 32129 641 32144
rect 641 32129 654 32144
rect 602 32092 654 32129
rect 454 32056 463 32079
rect 463 32056 497 32079
rect 497 32056 506 32079
rect 454 32027 506 32056
rect 528 32056 535 32079
rect 535 32056 569 32079
rect 569 32056 580 32079
rect 528 32027 580 32056
rect 602 32056 607 32079
rect 607 32056 641 32079
rect 641 32056 654 32079
rect 602 32027 654 32056
rect 454 31983 463 32014
rect 463 31983 497 32014
rect 497 31983 506 32014
rect 454 31962 506 31983
rect 528 31983 535 32014
rect 535 31983 569 32014
rect 569 31983 580 32014
rect 528 31962 580 31983
rect 602 31983 607 32014
rect 607 31983 641 32014
rect 641 31983 654 32014
rect 602 31962 654 31983
rect 454 31944 506 31949
rect 454 31910 463 31944
rect 463 31910 497 31944
rect 497 31910 506 31944
rect 454 31897 506 31910
rect 528 31944 580 31949
rect 528 31910 535 31944
rect 535 31910 569 31944
rect 569 31910 580 31944
rect 528 31897 580 31910
rect 602 31944 654 31949
rect 602 31910 607 31944
rect 607 31910 641 31944
rect 641 31910 654 31944
rect 602 31897 654 31910
rect 454 31871 506 31884
rect 454 31837 463 31871
rect 463 31837 497 31871
rect 497 31837 506 31871
rect 454 31832 506 31837
rect 528 31871 580 31884
rect 528 31837 535 31871
rect 535 31837 569 31871
rect 569 31837 580 31871
rect 528 31832 580 31837
rect 602 31871 654 31884
rect 602 31837 607 31871
rect 607 31837 641 31871
rect 641 31837 654 31871
rect 602 31832 654 31837
rect 454 31798 506 31819
rect 454 31767 463 31798
rect 463 31767 497 31798
rect 497 31767 506 31798
rect 528 31798 580 31819
rect 528 31767 535 31798
rect 535 31767 569 31798
rect 569 31767 580 31798
rect 602 31798 654 31819
rect 602 31767 607 31798
rect 607 31767 641 31798
rect 641 31767 654 31798
rect 454 31725 506 31754
rect 454 31702 463 31725
rect 463 31702 497 31725
rect 497 31702 506 31725
rect 528 31725 580 31754
rect 528 31702 535 31725
rect 535 31702 569 31725
rect 569 31702 580 31725
rect 602 31725 654 31754
rect 602 31702 607 31725
rect 607 31702 641 31725
rect 641 31702 654 31725
rect 454 31652 506 31689
rect 454 31637 463 31652
rect 463 31637 497 31652
rect 497 31637 506 31652
rect 528 31652 580 31689
rect 528 31637 535 31652
rect 535 31637 569 31652
rect 569 31637 580 31652
rect 602 31652 654 31689
rect 602 31637 607 31652
rect 607 31637 641 31652
rect 641 31637 654 31652
rect 454 31618 463 31624
rect 463 31618 497 31624
rect 497 31618 506 31624
rect 454 31579 506 31618
rect 454 31572 463 31579
rect 463 31572 497 31579
rect 497 31572 506 31579
rect 528 31618 535 31624
rect 535 31618 569 31624
rect 569 31618 580 31624
rect 528 31579 580 31618
rect 528 31572 535 31579
rect 535 31572 569 31579
rect 569 31572 580 31579
rect 602 31618 607 31624
rect 607 31618 641 31624
rect 641 31618 654 31624
rect 602 31579 654 31618
rect 602 31572 607 31579
rect 607 31572 641 31579
rect 641 31572 654 31579
rect 454 31545 463 31559
rect 463 31545 497 31559
rect 497 31545 506 31559
rect 454 31507 506 31545
rect 528 31545 535 31559
rect 535 31545 569 31559
rect 569 31545 580 31559
rect 528 31507 580 31545
rect 602 31545 607 31559
rect 607 31545 641 31559
rect 641 31545 654 31559
rect 602 31507 654 31545
rect 454 31472 463 31494
rect 463 31472 497 31494
rect 497 31472 506 31494
rect 454 31442 506 31472
rect 528 31472 535 31494
rect 535 31472 569 31494
rect 569 31472 580 31494
rect 528 31442 580 31472
rect 602 31472 607 31494
rect 607 31472 641 31494
rect 641 31472 654 31494
rect 602 31442 654 31472
rect 454 31399 463 31429
rect 463 31399 497 31429
rect 497 31399 506 31429
rect 454 31377 506 31399
rect 528 31399 535 31429
rect 535 31399 569 31429
rect 569 31399 580 31429
rect 528 31377 580 31399
rect 602 31399 607 31429
rect 607 31399 641 31429
rect 641 31399 654 31429
rect 602 31377 654 31399
rect 454 31360 506 31364
rect 454 31326 463 31360
rect 463 31326 497 31360
rect 497 31326 506 31360
rect 454 31312 506 31326
rect 528 31360 580 31364
rect 528 31326 535 31360
rect 535 31326 569 31360
rect 569 31326 580 31360
rect 528 31312 580 31326
rect 602 31360 654 31364
rect 602 31326 607 31360
rect 607 31326 641 31360
rect 641 31326 654 31360
rect 602 31312 654 31326
rect 454 31287 506 31299
rect 454 31253 463 31287
rect 463 31253 497 31287
rect 497 31253 506 31287
rect 454 31247 506 31253
rect 528 31287 580 31299
rect 528 31253 535 31287
rect 535 31253 569 31287
rect 569 31253 580 31287
rect 528 31247 580 31253
rect 602 31287 654 31299
rect 602 31253 607 31287
rect 607 31253 641 31287
rect 641 31253 654 31287
rect 602 31247 654 31253
rect 454 31214 506 31234
rect 454 31182 463 31214
rect 463 31182 497 31214
rect 497 31182 506 31214
rect 528 31214 580 31234
rect 528 31182 535 31214
rect 535 31182 569 31214
rect 569 31182 580 31214
rect 602 31214 654 31234
rect 602 31182 607 31214
rect 607 31182 641 31214
rect 641 31182 654 31214
rect 454 31141 506 31169
rect 454 31117 463 31141
rect 463 31117 497 31141
rect 497 31117 506 31141
rect 528 31141 580 31169
rect 528 31117 535 31141
rect 535 31117 569 31141
rect 569 31117 580 31141
rect 602 31141 654 31169
rect 602 31117 607 31141
rect 607 31117 641 31141
rect 641 31117 654 31141
rect 454 31068 506 31104
rect 454 31052 463 31068
rect 463 31052 497 31068
rect 497 31052 506 31068
rect 528 31068 580 31104
rect 528 31052 535 31068
rect 535 31052 569 31068
rect 569 31052 580 31068
rect 602 31068 654 31104
rect 602 31052 607 31068
rect 607 31052 641 31068
rect 641 31052 654 31068
rect 454 31034 463 31039
rect 463 31034 497 31039
rect 497 31034 506 31039
rect 454 30995 506 31034
rect 454 30987 463 30995
rect 463 30987 497 30995
rect 497 30987 506 30995
rect 528 31034 535 31039
rect 535 31034 569 31039
rect 569 31034 580 31039
rect 528 30995 580 31034
rect 528 30987 535 30995
rect 535 30987 569 30995
rect 569 30987 580 30995
rect 602 31034 607 31039
rect 607 31034 641 31039
rect 641 31034 654 31039
rect 602 30995 654 31034
rect 602 30987 607 30995
rect 607 30987 641 30995
rect 641 30987 654 30995
rect 454 30961 463 30974
rect 463 30961 497 30974
rect 497 30961 506 30974
rect 454 30922 506 30961
rect 528 30961 535 30974
rect 535 30961 569 30974
rect 569 30961 580 30974
rect 528 30922 580 30961
rect 602 30961 607 30974
rect 607 30961 641 30974
rect 641 30961 654 30974
rect 602 30922 654 30961
rect 454 30888 463 30909
rect 463 30888 497 30909
rect 497 30888 506 30909
rect 454 30857 506 30888
rect 528 30888 535 30909
rect 535 30888 569 30909
rect 569 30888 580 30909
rect 528 30857 580 30888
rect 602 30888 607 30909
rect 607 30888 641 30909
rect 641 30888 654 30909
rect 602 30857 654 30888
rect 454 30815 463 30844
rect 463 30815 497 30844
rect 497 30815 506 30844
rect 454 30792 506 30815
rect 528 30815 535 30844
rect 535 30815 569 30844
rect 569 30815 580 30844
rect 528 30792 580 30815
rect 602 30815 607 30844
rect 607 30815 641 30844
rect 641 30815 654 30844
rect 602 30792 654 30815
rect 454 30776 506 30779
rect 454 30742 463 30776
rect 463 30742 497 30776
rect 497 30742 506 30776
rect 454 30727 506 30742
rect 528 30776 580 30779
rect 528 30742 535 30776
rect 535 30742 569 30776
rect 569 30742 580 30776
rect 528 30727 580 30742
rect 602 30776 654 30779
rect 602 30742 607 30776
rect 607 30742 641 30776
rect 641 30742 654 30776
rect 602 30727 654 30742
rect 454 30703 506 30714
rect 454 30669 463 30703
rect 463 30669 497 30703
rect 497 30669 506 30703
rect 454 30662 506 30669
rect 528 30703 580 30714
rect 528 30669 535 30703
rect 535 30669 569 30703
rect 569 30669 580 30703
rect 528 30662 580 30669
rect 602 30703 654 30714
rect 602 30669 607 30703
rect 607 30669 641 30703
rect 641 30669 654 30703
rect 602 30662 654 30669
rect 454 30630 506 30649
rect 454 30597 463 30630
rect 463 30597 497 30630
rect 497 30597 506 30630
rect 528 30630 580 30649
rect 528 30597 535 30630
rect 535 30597 569 30630
rect 569 30597 580 30630
rect 602 30630 654 30649
rect 602 30597 607 30630
rect 607 30597 641 30630
rect 641 30597 654 30630
rect 454 30557 506 30584
rect 454 30532 463 30557
rect 463 30532 497 30557
rect 497 30532 506 30557
rect 528 30557 580 30584
rect 528 30532 535 30557
rect 535 30532 569 30557
rect 569 30532 580 30557
rect 602 30557 654 30584
rect 602 30532 607 30557
rect 607 30532 641 30557
rect 641 30532 654 30557
rect 454 30484 506 30519
rect 454 30467 463 30484
rect 463 30467 497 30484
rect 497 30467 506 30484
rect 528 30484 580 30519
rect 528 30467 535 30484
rect 535 30467 569 30484
rect 569 30467 580 30484
rect 602 30484 654 30519
rect 602 30467 607 30484
rect 607 30467 641 30484
rect 641 30467 654 30484
rect 454 30450 463 30454
rect 463 30450 497 30454
rect 497 30450 506 30454
rect 454 30411 506 30450
rect 454 30402 463 30411
rect 463 30402 497 30411
rect 497 30402 506 30411
rect 528 30450 535 30454
rect 535 30450 569 30454
rect 569 30450 580 30454
rect 528 30411 580 30450
rect 528 30402 535 30411
rect 535 30402 569 30411
rect 569 30402 580 30411
rect 602 30450 607 30454
rect 607 30450 641 30454
rect 641 30450 654 30454
rect 602 30411 654 30450
rect 602 30402 607 30411
rect 607 30402 641 30411
rect 641 30402 654 30411
rect 454 30377 463 30389
rect 463 30377 497 30389
rect 497 30377 506 30389
rect 454 30338 506 30377
rect 454 30337 463 30338
rect 463 30337 497 30338
rect 497 30337 506 30338
rect 528 30377 535 30389
rect 535 30377 569 30389
rect 569 30377 580 30389
rect 528 30338 580 30377
rect 528 30337 535 30338
rect 535 30337 569 30338
rect 569 30337 580 30338
rect 602 30377 607 30389
rect 607 30377 641 30389
rect 641 30377 654 30389
rect 602 30338 654 30377
rect 602 30337 607 30338
rect 607 30337 641 30338
rect 641 30337 654 30338
rect 454 30304 463 30324
rect 463 30304 497 30324
rect 497 30304 506 30324
rect 454 30272 506 30304
rect 528 30304 535 30324
rect 535 30304 569 30324
rect 569 30304 580 30324
rect 528 30272 580 30304
rect 602 30304 607 30324
rect 607 30304 641 30324
rect 641 30304 654 30324
rect 602 30272 654 30304
rect 454 30231 463 30259
rect 463 30231 497 30259
rect 497 30231 506 30259
rect 454 30207 506 30231
rect 528 30231 535 30259
rect 535 30231 569 30259
rect 569 30231 580 30259
rect 528 30207 580 30231
rect 602 30231 607 30259
rect 607 30231 641 30259
rect 641 30231 654 30259
rect 602 30207 654 30231
rect 454 30192 506 30194
rect 454 30158 463 30192
rect 463 30158 497 30192
rect 497 30158 506 30192
rect 454 30142 506 30158
rect 528 30192 580 30194
rect 528 30158 535 30192
rect 535 30158 569 30192
rect 569 30158 580 30192
rect 528 30142 580 30158
rect 602 30192 654 30194
rect 602 30158 607 30192
rect 607 30158 641 30192
rect 641 30158 654 30192
rect 602 30142 654 30158
rect 454 30119 506 30129
rect 454 30085 463 30119
rect 463 30085 497 30119
rect 497 30085 506 30119
rect 454 30077 506 30085
rect 528 30119 580 30129
rect 528 30085 535 30119
rect 535 30085 569 30119
rect 569 30085 580 30119
rect 528 30077 580 30085
rect 602 30119 654 30129
rect 602 30085 607 30119
rect 607 30085 641 30119
rect 641 30085 654 30119
rect 602 30077 654 30085
rect 454 30046 506 30064
rect 454 30012 463 30046
rect 463 30012 497 30046
rect 497 30012 506 30046
rect 528 30046 580 30064
rect 528 30012 535 30046
rect 535 30012 569 30046
rect 569 30012 580 30046
rect 602 30046 654 30064
rect 602 30012 607 30046
rect 607 30012 641 30046
rect 641 30012 654 30046
rect 454 29973 506 29999
rect 454 29947 463 29973
rect 463 29947 497 29973
rect 497 29947 506 29973
rect 528 29973 580 29999
rect 528 29947 535 29973
rect 535 29947 569 29973
rect 569 29947 580 29973
rect 602 29973 654 29999
rect 602 29947 607 29973
rect 607 29947 641 29973
rect 641 29947 654 29973
rect 454 29900 506 29934
rect 454 29882 463 29900
rect 463 29882 497 29900
rect 497 29882 506 29900
rect 528 29900 580 29934
rect 528 29882 535 29900
rect 535 29882 569 29900
rect 569 29882 580 29900
rect 602 29900 654 29934
rect 602 29882 607 29900
rect 607 29882 641 29900
rect 641 29882 654 29900
rect 454 29866 463 29869
rect 463 29866 497 29869
rect 497 29866 506 29869
rect 454 29827 506 29866
rect 454 29817 463 29827
rect 463 29817 497 29827
rect 497 29817 506 29827
rect 528 29866 535 29869
rect 535 29866 569 29869
rect 569 29866 580 29869
rect 528 29827 580 29866
rect 528 29817 535 29827
rect 535 29817 569 29827
rect 569 29817 580 29827
rect 602 29866 607 29869
rect 607 29866 641 29869
rect 641 29866 654 29869
rect 602 29827 654 29866
rect 602 29817 607 29827
rect 607 29817 641 29827
rect 641 29817 654 29827
rect 454 29793 463 29804
rect 463 29793 497 29804
rect 497 29793 506 29804
rect 454 29754 506 29793
rect 454 29752 463 29754
rect 463 29752 497 29754
rect 497 29752 506 29754
rect 528 29793 535 29804
rect 535 29793 569 29804
rect 569 29793 580 29804
rect 528 29754 580 29793
rect 528 29752 535 29754
rect 535 29752 569 29754
rect 569 29752 580 29754
rect 602 29793 607 29804
rect 607 29793 641 29804
rect 641 29793 654 29804
rect 602 29754 654 29793
rect 602 29752 607 29754
rect 607 29752 641 29754
rect 641 29752 654 29754
rect 454 29720 463 29739
rect 463 29720 497 29739
rect 497 29720 506 29739
rect 454 29687 506 29720
rect 528 29720 535 29739
rect 535 29720 569 29739
rect 569 29720 580 29739
rect 528 29687 580 29720
rect 602 29720 607 29739
rect 607 29720 641 29739
rect 641 29720 654 29739
rect 602 29687 654 29720
rect 454 29647 463 29674
rect 463 29647 497 29674
rect 497 29647 506 29674
rect 454 29622 506 29647
rect 528 29647 535 29674
rect 535 29647 569 29674
rect 569 29647 580 29674
rect 528 29622 580 29647
rect 602 29647 607 29674
rect 607 29647 641 29674
rect 641 29647 654 29674
rect 602 29622 654 29647
rect 454 29608 506 29609
rect 454 29574 463 29608
rect 463 29574 497 29608
rect 497 29574 506 29608
rect 454 29557 506 29574
rect 528 29608 580 29609
rect 528 29574 535 29608
rect 535 29574 569 29608
rect 569 29574 580 29608
rect 528 29557 580 29574
rect 602 29608 654 29609
rect 602 29574 607 29608
rect 607 29574 641 29608
rect 641 29574 654 29608
rect 602 29557 654 29574
rect 454 29535 506 29544
rect 454 29501 463 29535
rect 463 29501 497 29535
rect 497 29501 506 29535
rect 454 29492 506 29501
rect 528 29535 580 29544
rect 528 29501 535 29535
rect 535 29501 569 29535
rect 569 29501 580 29535
rect 528 29492 580 29501
rect 602 29535 654 29544
rect 602 29501 607 29535
rect 607 29501 641 29535
rect 641 29501 654 29535
rect 602 29492 654 29501
rect 454 29462 506 29479
rect 454 29428 463 29462
rect 463 29428 497 29462
rect 497 29428 506 29462
rect 454 29427 506 29428
rect 528 29462 580 29479
rect 528 29428 535 29462
rect 535 29428 569 29462
rect 569 29428 580 29462
rect 528 29427 580 29428
rect 602 29462 654 29479
rect 602 29428 607 29462
rect 607 29428 641 29462
rect 641 29428 654 29462
rect 602 29427 654 29428
rect 454 29389 506 29414
rect 454 29362 463 29389
rect 463 29362 497 29389
rect 497 29362 506 29389
rect 528 29389 580 29414
rect 528 29362 535 29389
rect 535 29362 569 29389
rect 569 29362 580 29389
rect 602 29389 654 29414
rect 602 29362 607 29389
rect 607 29362 641 29389
rect 641 29362 654 29389
rect 454 29316 506 29349
rect 454 29297 463 29316
rect 463 29297 497 29316
rect 497 29297 506 29316
rect 528 29316 580 29349
rect 528 29297 535 29316
rect 535 29297 569 29316
rect 569 29297 580 29316
rect 602 29316 654 29349
rect 602 29297 607 29316
rect 607 29297 641 29316
rect 641 29297 654 29316
rect 454 29282 463 29284
rect 463 29282 497 29284
rect 497 29282 506 29284
rect 454 29243 506 29282
rect 454 29232 463 29243
rect 463 29232 497 29243
rect 497 29232 506 29243
rect 528 29282 535 29284
rect 535 29282 569 29284
rect 569 29282 580 29284
rect 528 29243 580 29282
rect 528 29232 535 29243
rect 535 29232 569 29243
rect 569 29232 580 29243
rect 602 29282 607 29284
rect 607 29282 641 29284
rect 641 29282 654 29284
rect 602 29243 654 29282
rect 602 29232 607 29243
rect 607 29232 641 29243
rect 641 29232 654 29243
rect 454 29209 463 29219
rect 463 29209 497 29219
rect 497 29209 506 29219
rect 454 29170 506 29209
rect 454 29167 463 29170
rect 463 29167 497 29170
rect 497 29167 506 29170
rect 528 29209 535 29219
rect 535 29209 569 29219
rect 569 29209 580 29219
rect 528 29170 580 29209
rect 528 29167 535 29170
rect 535 29167 569 29170
rect 569 29167 580 29170
rect 602 29209 607 29219
rect 607 29209 641 29219
rect 641 29209 654 29219
rect 602 29170 654 29209
rect 602 29167 607 29170
rect 607 29167 641 29170
rect 641 29167 654 29170
rect 454 29136 463 29154
rect 463 29136 497 29154
rect 497 29136 506 29154
rect 454 29102 506 29136
rect 528 29136 535 29154
rect 535 29136 569 29154
rect 569 29136 580 29154
rect 528 29102 580 29136
rect 602 29136 607 29154
rect 607 29136 641 29154
rect 641 29136 654 29154
rect 602 29102 654 29136
rect 454 29063 463 29089
rect 463 29063 497 29089
rect 497 29063 506 29089
rect 454 29037 506 29063
rect 528 29063 535 29089
rect 535 29063 569 29089
rect 569 29063 580 29089
rect 528 29037 580 29063
rect 602 29063 607 29089
rect 607 29063 641 29089
rect 641 29063 654 29089
rect 602 29037 654 29063
rect 2788 28509 2840 28561
rect 2854 28509 2906 28561
rect 2919 28509 2971 28561
rect 2984 28509 3036 28561
rect 3049 28509 3101 28561
rect 3114 28509 3166 28561
rect 3179 28509 3231 28561
rect 3244 28509 3296 28561
rect 3309 28509 3361 28561
rect 3374 28509 3426 28561
rect 3439 28509 3491 28561
rect 3504 28509 3556 28561
rect 3569 28509 3621 28561
rect 3634 28509 3686 28561
rect 3699 28509 3751 28561
rect 2788 28439 2840 28491
rect 2854 28439 2906 28491
rect 2919 28439 2971 28491
rect 2984 28439 3036 28491
rect 3049 28439 3101 28491
rect 3114 28439 3166 28491
rect 3179 28439 3231 28491
rect 3244 28439 3296 28491
rect 3309 28439 3361 28491
rect 3374 28439 3426 28491
rect 3439 28439 3491 28491
rect 3504 28439 3556 28491
rect 3569 28439 3621 28491
rect 3634 28439 3686 28491
rect 3699 28439 3751 28491
rect 2788 28369 2840 28421
rect 2854 28369 2906 28421
rect 2919 28369 2971 28421
rect 2984 28369 3036 28421
rect 3049 28369 3101 28421
rect 3114 28369 3166 28421
rect 3179 28369 3231 28421
rect 3244 28369 3296 28421
rect 3309 28369 3361 28421
rect 3374 28369 3426 28421
rect 3439 28369 3491 28421
rect 3504 28369 3556 28421
rect 3569 28369 3621 28421
rect 3634 28369 3686 28421
rect 3699 28369 3751 28421
rect 149 27998 201 28024
rect 149 27972 167 27998
rect 167 27972 201 27998
rect 247 27998 299 28024
rect 247 27972 259 27998
rect 259 27972 293 27998
rect 293 27972 299 27998
rect 149 27925 201 27958
rect 149 27906 167 27925
rect 167 27906 201 27925
rect 247 27925 299 27958
rect 247 27906 259 27925
rect 259 27906 293 27925
rect 293 27906 299 27925
rect 149 27891 167 27892
rect 167 27891 201 27892
rect 149 27852 201 27891
rect 149 27840 167 27852
rect 167 27840 201 27852
rect 247 27891 259 27892
rect 259 27891 293 27892
rect 293 27891 299 27892
rect 247 27852 299 27891
rect 247 27840 259 27852
rect 259 27840 293 27852
rect 293 27840 299 27852
rect 149 27818 167 27826
rect 167 27818 201 27826
rect 149 27779 201 27818
rect 149 27774 167 27779
rect 167 27774 201 27779
rect 247 27818 259 27826
rect 259 27818 293 27826
rect 293 27818 299 27826
rect 247 27779 299 27818
rect 247 27774 259 27779
rect 259 27774 293 27779
rect 293 27774 299 27779
rect 149 27745 167 27760
rect 167 27745 201 27760
rect 149 27708 201 27745
rect 247 27745 259 27760
rect 259 27745 293 27760
rect 293 27745 299 27760
rect 247 27708 299 27745
rect 149 27672 167 27694
rect 167 27672 201 27694
rect 149 27642 201 27672
rect 247 27672 259 27694
rect 259 27672 293 27694
rect 293 27672 299 27694
rect 247 27642 299 27672
rect 149 27599 167 27628
rect 167 27599 201 27628
rect 149 27576 201 27599
rect 247 27599 259 27628
rect 259 27599 293 27628
rect 293 27599 299 27628
rect 247 27576 299 27599
rect 149 27560 201 27562
rect 149 27526 167 27560
rect 167 27526 201 27560
rect 149 27510 201 27526
rect 247 27560 299 27562
rect 247 27526 259 27560
rect 259 27526 293 27560
rect 293 27526 299 27560
rect 247 27510 299 27526
rect 149 27487 201 27496
rect 149 27453 167 27487
rect 167 27453 201 27487
rect 149 27444 201 27453
rect 247 27487 299 27496
rect 247 27453 259 27487
rect 259 27453 293 27487
rect 293 27453 299 27487
rect 247 27444 299 27453
rect 149 27414 201 27430
rect 149 27380 167 27414
rect 167 27380 201 27414
rect 149 27378 201 27380
rect 247 27414 299 27430
rect 247 27380 259 27414
rect 259 27380 293 27414
rect 293 27380 299 27414
rect 247 27378 299 27380
rect 149 27341 201 27364
rect 149 27312 167 27341
rect 167 27312 201 27341
rect 247 27341 299 27364
rect 247 27312 259 27341
rect 259 27312 293 27341
rect 293 27312 299 27341
rect 149 27268 201 27298
rect 149 27246 167 27268
rect 167 27246 201 27268
rect 247 27268 299 27298
rect 247 27246 259 27268
rect 259 27246 293 27268
rect 293 27246 299 27268
rect 149 27195 201 27232
rect 149 27180 167 27195
rect 167 27180 201 27195
rect 247 27195 299 27232
rect 247 27180 259 27195
rect 259 27180 293 27195
rect 293 27180 299 27195
rect 149 27161 167 27166
rect 167 27161 201 27166
rect 149 27122 201 27161
rect 149 27114 167 27122
rect 167 27114 201 27122
rect 247 27161 259 27166
rect 259 27161 293 27166
rect 293 27161 299 27166
rect 247 27122 299 27161
rect 247 27114 259 27122
rect 259 27114 293 27122
rect 293 27114 299 27122
rect 149 27088 167 27100
rect 167 27088 201 27100
rect 149 27049 201 27088
rect 149 27048 167 27049
rect 167 27048 201 27049
rect 247 27088 259 27100
rect 259 27088 293 27100
rect 293 27088 299 27100
rect 247 27049 299 27088
rect 247 27048 259 27049
rect 259 27048 293 27049
rect 293 27048 299 27049
rect 149 27015 167 27034
rect 167 27015 201 27034
rect 149 26982 201 27015
rect 247 27015 259 27034
rect 259 27015 293 27034
rect 293 27015 299 27034
rect 247 26982 299 27015
rect 149 26942 167 26968
rect 167 26942 201 26968
rect 149 26916 201 26942
rect 247 26942 259 26968
rect 259 26942 293 26968
rect 293 26942 299 26968
rect 247 26916 299 26942
rect 149 26869 167 26902
rect 167 26869 201 26902
rect 149 26850 201 26869
rect 247 26869 259 26902
rect 259 26869 293 26902
rect 293 26869 299 26902
rect 247 26850 299 26869
rect 149 26830 201 26836
rect 149 26796 167 26830
rect 167 26796 201 26830
rect 149 26784 201 26796
rect 247 26830 299 26836
rect 247 26796 259 26830
rect 259 26796 293 26830
rect 293 26796 299 26830
rect 247 26784 299 26796
rect 149 26757 201 26770
rect 149 26723 167 26757
rect 167 26723 201 26757
rect 149 26718 201 26723
rect 247 26757 299 26770
rect 247 26723 259 26757
rect 259 26723 293 26757
rect 293 26723 299 26757
rect 247 26718 299 26723
rect 149 26684 201 26704
rect 149 26652 167 26684
rect 167 26652 201 26684
rect 247 26684 299 26704
rect 247 26652 259 26684
rect 259 26652 293 26684
rect 293 26652 299 26684
rect 149 26611 201 26638
rect 149 26586 167 26611
rect 167 26586 201 26611
rect 247 26611 299 26638
rect 247 26586 259 26611
rect 259 26586 293 26611
rect 293 26586 299 26611
rect 149 26538 201 26573
rect 149 26521 167 26538
rect 167 26521 201 26538
rect 247 26538 299 26573
rect 247 26521 259 26538
rect 259 26521 293 26538
rect 293 26521 299 26538
rect 149 26504 167 26508
rect 167 26504 201 26508
rect 149 26465 201 26504
rect 149 26456 167 26465
rect 167 26456 201 26465
rect 247 26504 259 26508
rect 259 26504 293 26508
rect 293 26504 299 26508
rect 247 26465 299 26504
rect 247 26456 259 26465
rect 259 26456 293 26465
rect 293 26456 299 26465
rect 149 26431 167 26443
rect 167 26431 201 26443
rect 149 26393 201 26431
rect 149 26391 167 26393
rect 167 26391 201 26393
rect 247 26431 259 26443
rect 259 26431 293 26443
rect 293 26431 299 26443
rect 247 26393 299 26431
rect 247 26391 259 26393
rect 259 26391 293 26393
rect 293 26391 299 26393
rect 149 26359 167 26378
rect 167 26359 201 26378
rect 149 26326 201 26359
rect 247 26359 259 26378
rect 259 26359 293 26378
rect 293 26359 299 26378
rect 247 26326 299 26359
rect 149 26287 167 26313
rect 167 26287 201 26313
rect 149 26261 201 26287
rect 247 26287 259 26313
rect 259 26287 293 26313
rect 293 26287 299 26313
rect 247 26261 299 26287
rect 454 27978 506 28024
rect 454 27972 463 27978
rect 463 27972 497 27978
rect 497 27972 506 27978
rect 528 27978 580 28024
rect 528 27972 535 27978
rect 535 27972 569 27978
rect 569 27972 580 27978
rect 602 27978 654 28024
rect 602 27972 607 27978
rect 607 27972 641 27978
rect 641 27972 654 27978
rect 454 27944 463 27958
rect 463 27944 497 27958
rect 497 27944 506 27958
rect 454 27906 506 27944
rect 528 27944 535 27958
rect 535 27944 569 27958
rect 569 27944 580 27958
rect 528 27906 580 27944
rect 602 27944 607 27958
rect 607 27944 641 27958
rect 641 27944 654 27958
rect 602 27906 654 27944
rect 454 27869 463 27892
rect 463 27869 497 27892
rect 497 27869 506 27892
rect 454 27840 506 27869
rect 528 27869 535 27892
rect 535 27869 569 27892
rect 569 27869 580 27892
rect 528 27840 580 27869
rect 602 27869 607 27892
rect 607 27869 641 27892
rect 641 27869 654 27892
rect 602 27840 654 27869
rect 454 27794 463 27826
rect 463 27794 497 27826
rect 497 27794 506 27826
rect 454 27774 506 27794
rect 528 27794 535 27826
rect 535 27794 569 27826
rect 569 27794 580 27826
rect 528 27774 580 27794
rect 602 27794 607 27826
rect 607 27794 641 27826
rect 641 27794 654 27826
rect 602 27774 654 27794
rect 454 27753 506 27760
rect 454 27719 463 27753
rect 463 27719 497 27753
rect 497 27719 506 27753
rect 454 27708 506 27719
rect 528 27753 580 27760
rect 528 27719 535 27753
rect 535 27719 569 27753
rect 569 27719 580 27753
rect 528 27708 580 27719
rect 602 27753 654 27760
rect 602 27719 607 27753
rect 607 27719 641 27753
rect 641 27719 654 27753
rect 602 27708 654 27719
rect 454 27678 506 27694
rect 454 27644 463 27678
rect 463 27644 497 27678
rect 497 27644 506 27678
rect 454 27642 506 27644
rect 528 27678 580 27694
rect 528 27644 535 27678
rect 535 27644 569 27678
rect 569 27644 580 27678
rect 528 27642 580 27644
rect 602 27678 654 27694
rect 602 27644 607 27678
rect 607 27644 641 27678
rect 641 27644 654 27678
rect 602 27642 654 27644
rect 454 27603 506 27628
rect 454 27576 463 27603
rect 463 27576 497 27603
rect 497 27576 506 27603
rect 528 27603 580 27628
rect 528 27576 535 27603
rect 535 27576 569 27603
rect 569 27576 580 27603
rect 602 27603 654 27628
rect 602 27576 607 27603
rect 607 27576 641 27603
rect 641 27576 654 27603
rect 454 27528 506 27562
rect 454 27510 463 27528
rect 463 27510 497 27528
rect 497 27510 506 27528
rect 528 27528 580 27562
rect 528 27510 535 27528
rect 535 27510 569 27528
rect 569 27510 580 27528
rect 602 27528 654 27562
rect 602 27510 607 27528
rect 607 27510 641 27528
rect 641 27510 654 27528
rect 454 27494 463 27496
rect 463 27494 497 27496
rect 497 27494 506 27496
rect 454 27453 506 27494
rect 454 27444 463 27453
rect 463 27444 497 27453
rect 497 27444 506 27453
rect 528 27494 535 27496
rect 535 27494 569 27496
rect 569 27494 580 27496
rect 528 27453 580 27494
rect 528 27444 535 27453
rect 535 27444 569 27453
rect 569 27444 580 27453
rect 602 27494 607 27496
rect 607 27494 641 27496
rect 641 27494 654 27496
rect 602 27453 654 27494
rect 602 27444 607 27453
rect 607 27444 641 27453
rect 641 27444 654 27453
rect 454 27419 463 27430
rect 463 27419 497 27430
rect 497 27419 506 27430
rect 454 27378 506 27419
rect 528 27419 535 27430
rect 535 27419 569 27430
rect 569 27419 580 27430
rect 528 27378 580 27419
rect 602 27419 607 27430
rect 607 27419 641 27430
rect 641 27419 654 27430
rect 602 27378 654 27419
rect 454 27344 463 27364
rect 463 27344 497 27364
rect 497 27344 506 27364
rect 454 27312 506 27344
rect 528 27344 535 27364
rect 535 27344 569 27364
rect 569 27344 580 27364
rect 528 27312 580 27344
rect 602 27344 607 27364
rect 607 27344 641 27364
rect 641 27344 654 27364
rect 602 27312 654 27344
rect 454 27269 463 27298
rect 463 27269 497 27298
rect 497 27269 506 27298
rect 454 27246 506 27269
rect 528 27269 535 27298
rect 535 27269 569 27298
rect 569 27269 580 27298
rect 528 27246 580 27269
rect 602 27269 607 27298
rect 607 27269 641 27298
rect 641 27269 654 27298
rect 602 27246 654 27269
rect 454 27228 506 27232
rect 454 27194 463 27228
rect 463 27194 497 27228
rect 497 27194 506 27228
rect 454 27180 506 27194
rect 528 27228 580 27232
rect 528 27194 535 27228
rect 535 27194 569 27228
rect 569 27194 580 27228
rect 528 27180 580 27194
rect 602 27228 654 27232
rect 602 27194 607 27228
rect 607 27194 641 27228
rect 641 27194 654 27228
rect 602 27180 654 27194
rect 454 27153 506 27167
rect 454 27119 463 27153
rect 463 27119 497 27153
rect 497 27119 506 27153
rect 454 27115 506 27119
rect 528 27153 580 27167
rect 528 27119 535 27153
rect 535 27119 569 27153
rect 569 27119 580 27153
rect 528 27115 580 27119
rect 602 27153 654 27167
rect 602 27119 607 27153
rect 607 27119 641 27153
rect 641 27119 654 27153
rect 602 27115 654 27119
rect 454 27079 506 27102
rect 454 27050 463 27079
rect 463 27050 497 27079
rect 497 27050 506 27079
rect 528 27079 580 27102
rect 528 27050 535 27079
rect 535 27050 569 27079
rect 569 27050 580 27079
rect 602 27079 654 27102
rect 14213 27431 14265 27483
rect 14285 27431 14337 27483
rect 14357 27431 14409 27483
rect 14213 27364 14265 27416
rect 14285 27364 14337 27416
rect 14357 27364 14409 27416
rect 14213 27297 14265 27349
rect 14285 27297 14337 27349
rect 14357 27297 14409 27349
rect 14213 27229 14265 27281
rect 14285 27229 14337 27281
rect 14357 27229 14409 27281
rect 14213 27161 14265 27213
rect 14285 27161 14337 27213
rect 14357 27161 14409 27213
rect 14213 27093 14265 27145
rect 14285 27093 14337 27145
rect 14357 27093 14409 27145
rect 602 27050 607 27079
rect 607 27050 641 27079
rect 641 27050 654 27079
rect 454 27005 506 27037
rect 454 26985 463 27005
rect 463 26985 497 27005
rect 497 26985 506 27005
rect 528 27005 580 27037
rect 528 26985 535 27005
rect 535 26985 569 27005
rect 569 26985 580 27005
rect 602 27005 654 27037
rect 602 26985 607 27005
rect 607 26985 641 27005
rect 641 26985 654 27005
rect 454 26971 463 26972
rect 463 26971 497 26972
rect 497 26971 506 26972
rect 454 26931 506 26971
rect 454 26920 463 26931
rect 463 26920 497 26931
rect 497 26920 506 26931
rect 528 26971 535 26972
rect 535 26971 569 26972
rect 569 26971 580 26972
rect 528 26931 580 26971
rect 528 26920 535 26931
rect 535 26920 569 26931
rect 569 26920 580 26931
rect 602 26971 607 26972
rect 607 26971 641 26972
rect 641 26971 654 26972
rect 602 26931 654 26971
rect 602 26920 607 26931
rect 607 26920 641 26931
rect 641 26920 654 26931
rect 454 26897 463 26907
rect 463 26897 497 26907
rect 497 26897 506 26907
rect 454 26857 506 26897
rect 454 26855 463 26857
rect 463 26855 497 26857
rect 497 26855 506 26857
rect 528 26897 535 26907
rect 535 26897 569 26907
rect 569 26897 580 26907
rect 528 26857 580 26897
rect 528 26855 535 26857
rect 535 26855 569 26857
rect 569 26855 580 26857
rect 602 26897 607 26907
rect 607 26897 641 26907
rect 641 26897 654 26907
rect 602 26857 654 26897
rect 602 26855 607 26857
rect 607 26855 641 26857
rect 641 26855 654 26857
rect 454 26823 463 26842
rect 463 26823 497 26842
rect 497 26823 506 26842
rect 454 26790 506 26823
rect 528 26823 535 26842
rect 535 26823 569 26842
rect 569 26823 580 26842
rect 528 26790 580 26823
rect 602 26823 607 26842
rect 607 26823 641 26842
rect 641 26823 654 26842
rect 602 26790 654 26823
rect 454 26749 463 26777
rect 463 26749 497 26777
rect 497 26749 506 26777
rect 454 26725 506 26749
rect 528 26749 535 26777
rect 535 26749 569 26777
rect 569 26749 580 26777
rect 528 26725 580 26749
rect 602 26749 607 26777
rect 607 26749 641 26777
rect 641 26749 654 26777
rect 602 26725 654 26749
rect 454 26709 506 26712
rect 454 26675 463 26709
rect 463 26675 497 26709
rect 497 26675 506 26709
rect 454 26660 506 26675
rect 528 26709 580 26712
rect 528 26675 535 26709
rect 535 26675 569 26709
rect 569 26675 580 26709
rect 528 26660 580 26675
rect 602 26709 654 26712
rect 602 26675 607 26709
rect 607 26675 641 26709
rect 641 26675 654 26709
rect 602 26660 654 26675
rect 454 26635 506 26647
rect 454 26601 463 26635
rect 463 26601 497 26635
rect 497 26601 506 26635
rect 454 26595 506 26601
rect 528 26635 580 26647
rect 528 26601 535 26635
rect 535 26601 569 26635
rect 569 26601 580 26635
rect 528 26595 580 26601
rect 602 26635 654 26647
rect 602 26601 607 26635
rect 607 26601 641 26635
rect 641 26601 654 26635
rect 602 26595 654 26601
rect 454 26561 506 26582
rect 454 26530 463 26561
rect 463 26530 497 26561
rect 497 26530 506 26561
rect 528 26561 580 26582
rect 528 26530 535 26561
rect 535 26530 569 26561
rect 569 26530 580 26561
rect 602 26561 654 26582
rect 602 26530 607 26561
rect 607 26530 641 26561
rect 641 26530 654 26561
rect 454 26487 506 26517
rect 454 26465 463 26487
rect 463 26465 497 26487
rect 497 26465 506 26487
rect 528 26487 580 26517
rect 528 26465 535 26487
rect 535 26465 569 26487
rect 569 26465 580 26487
rect 602 26487 654 26517
rect 602 26465 607 26487
rect 607 26465 641 26487
rect 641 26465 654 26487
rect 454 26413 506 26452
rect 454 26400 463 26413
rect 463 26400 497 26413
rect 497 26400 506 26413
rect 528 26413 580 26452
rect 528 26400 535 26413
rect 535 26400 569 26413
rect 569 26400 580 26413
rect 602 26413 654 26452
rect 602 26400 607 26413
rect 607 26400 641 26413
rect 641 26400 654 26413
rect 454 26379 463 26387
rect 463 26379 497 26387
rect 497 26379 506 26387
rect 454 26339 506 26379
rect 454 26335 463 26339
rect 463 26335 497 26339
rect 497 26335 506 26339
rect 528 26379 535 26387
rect 535 26379 569 26387
rect 569 26379 580 26387
rect 528 26339 580 26379
rect 528 26335 535 26339
rect 535 26335 569 26339
rect 569 26335 580 26339
rect 602 26379 607 26387
rect 607 26379 641 26387
rect 641 26379 654 26387
rect 602 26339 654 26379
rect 602 26335 607 26339
rect 607 26335 641 26339
rect 641 26335 654 26339
rect 454 26305 463 26322
rect 463 26305 497 26322
rect 497 26305 506 26322
rect 454 26270 506 26305
rect 528 26305 535 26322
rect 535 26305 569 26322
rect 569 26305 580 26322
rect 528 26270 580 26305
rect 602 26305 607 26322
rect 607 26305 641 26322
rect 641 26305 654 26322
rect 602 26270 654 26305
rect 454 26231 463 26257
rect 463 26231 497 26257
rect 497 26231 506 26257
rect 454 26205 506 26231
rect 528 26231 535 26257
rect 535 26231 569 26257
rect 569 26231 580 26257
rect 528 26205 580 26231
rect 602 26231 607 26257
rect 607 26231 641 26257
rect 641 26231 654 26257
rect 602 26205 654 26231
rect 149 26012 201 26038
rect 149 25986 167 26012
rect 167 25986 201 26012
rect 247 26012 299 26038
rect 247 25986 259 26012
rect 259 25986 293 26012
rect 293 25986 299 26012
rect 149 25940 201 25974
rect 149 25922 167 25940
rect 167 25922 201 25940
rect 247 25940 299 25974
rect 247 25922 259 25940
rect 259 25922 293 25940
rect 293 25922 299 25940
rect 149 25906 167 25910
rect 167 25906 201 25910
rect 149 25868 201 25906
rect 149 25858 167 25868
rect 167 25858 201 25868
rect 247 25906 259 25910
rect 259 25906 293 25910
rect 293 25906 299 25910
rect 247 25868 299 25906
rect 247 25858 259 25868
rect 259 25858 293 25868
rect 293 25858 299 25868
rect 149 25834 167 25846
rect 167 25834 201 25846
rect 149 25796 201 25834
rect 149 25794 167 25796
rect 167 25794 201 25796
rect 247 25834 259 25846
rect 259 25834 293 25846
rect 293 25834 299 25846
rect 247 25796 299 25834
rect 247 25794 259 25796
rect 259 25794 293 25796
rect 293 25794 299 25796
rect 149 25762 167 25782
rect 167 25762 201 25782
rect 149 25730 201 25762
rect 247 25762 259 25782
rect 259 25762 293 25782
rect 293 25762 299 25782
rect 247 25730 299 25762
rect 149 25690 167 25718
rect 167 25690 201 25718
rect 149 25666 201 25690
rect 247 25690 259 25718
rect 259 25690 293 25718
rect 293 25690 299 25718
rect 247 25666 299 25690
rect 149 25652 201 25654
rect 149 25618 167 25652
rect 167 25618 201 25652
rect 149 25602 201 25618
rect 247 25652 299 25654
rect 247 25618 259 25652
rect 259 25618 293 25652
rect 293 25618 299 25652
rect 247 25602 299 25618
rect 149 25580 201 25590
rect 149 25546 167 25580
rect 167 25546 201 25580
rect 149 25538 201 25546
rect 247 25580 299 25590
rect 247 25546 259 25580
rect 259 25546 293 25580
rect 293 25546 299 25580
rect 247 25538 299 25546
rect 149 25508 201 25526
rect 149 25474 167 25508
rect 167 25474 201 25508
rect 247 25508 299 25526
rect 247 25474 259 25508
rect 259 25474 293 25508
rect 293 25474 299 25508
rect 149 25436 201 25462
rect 149 25410 167 25436
rect 167 25410 201 25436
rect 247 25436 299 25462
rect 247 25410 259 25436
rect 259 25410 293 25436
rect 293 25410 299 25436
rect 149 25364 201 25398
rect 149 25346 167 25364
rect 167 25346 201 25364
rect 247 25364 299 25398
rect 247 25346 259 25364
rect 259 25346 293 25364
rect 293 25346 299 25364
rect 149 25330 167 25334
rect 167 25330 201 25334
rect 149 25292 201 25330
rect 149 25282 167 25292
rect 167 25282 201 25292
rect 247 25330 259 25334
rect 259 25330 293 25334
rect 293 25330 299 25334
rect 247 25292 299 25330
rect 247 25282 259 25292
rect 259 25282 293 25292
rect 293 25282 299 25292
rect 149 25258 167 25270
rect 167 25258 201 25270
rect 149 25220 201 25258
rect 149 25218 167 25220
rect 167 25218 201 25220
rect 247 25258 259 25270
rect 259 25258 293 25270
rect 293 25258 299 25270
rect 247 25220 299 25258
rect 247 25218 259 25220
rect 259 25218 293 25220
rect 293 25218 299 25220
rect 149 25186 167 25206
rect 167 25186 201 25206
rect 149 25154 201 25186
rect 247 25186 259 25206
rect 259 25186 293 25206
rect 293 25186 299 25206
rect 247 25154 299 25186
rect 149 25114 167 25142
rect 167 25114 201 25142
rect 149 25090 201 25114
rect 247 25114 259 25142
rect 259 25114 293 25142
rect 293 25114 299 25142
rect 247 25090 299 25114
rect 149 25076 201 25078
rect 149 25042 167 25076
rect 167 25042 201 25076
rect 149 25026 201 25042
rect 247 25076 299 25078
rect 247 25042 259 25076
rect 259 25042 293 25076
rect 293 25042 299 25076
rect 247 25026 299 25042
rect 149 25004 201 25014
rect 149 24970 167 25004
rect 167 24970 201 25004
rect 149 24962 201 24970
rect 247 25004 299 25014
rect 247 24970 259 25004
rect 259 24970 293 25004
rect 293 24970 299 25004
rect 247 24962 299 24970
rect 149 24932 201 24950
rect 149 24898 167 24932
rect 167 24898 201 24932
rect 247 24932 299 24950
rect 247 24898 259 24932
rect 259 24898 293 24932
rect 293 24898 299 24932
rect 149 24860 201 24886
rect 149 24834 167 24860
rect 167 24834 201 24860
rect 247 24860 299 24886
rect 247 24834 259 24860
rect 259 24834 293 24860
rect 293 24834 299 24860
rect 149 24788 201 24822
rect 149 24770 167 24788
rect 167 24770 201 24788
rect 247 24788 299 24822
rect 247 24770 259 24788
rect 259 24770 293 24788
rect 293 24770 299 24788
rect 149 24754 167 24758
rect 167 24754 201 24758
rect 149 24716 201 24754
rect 149 24706 167 24716
rect 167 24706 201 24716
rect 247 24754 259 24758
rect 259 24754 293 24758
rect 293 24754 299 24758
rect 247 24716 299 24754
rect 247 24706 259 24716
rect 259 24706 293 24716
rect 293 24706 299 24716
rect 149 24682 167 24694
rect 167 24682 201 24694
rect 149 24644 201 24682
rect 149 24642 167 24644
rect 167 24642 201 24644
rect 247 24682 259 24694
rect 259 24682 293 24694
rect 293 24682 299 24694
rect 247 24644 299 24682
rect 247 24642 259 24644
rect 259 24642 293 24644
rect 293 24642 299 24644
rect 149 24610 167 24630
rect 167 24610 201 24630
rect 149 24578 201 24610
rect 247 24610 259 24630
rect 259 24610 293 24630
rect 293 24610 299 24630
rect 247 24578 299 24610
rect 149 24538 167 24566
rect 167 24538 201 24566
rect 149 24514 201 24538
rect 247 24538 259 24566
rect 259 24538 293 24566
rect 293 24538 299 24566
rect 247 24514 299 24538
rect 149 24500 201 24502
rect 149 24466 167 24500
rect 167 24466 201 24500
rect 149 24450 201 24466
rect 247 24500 299 24502
rect 247 24466 259 24500
rect 259 24466 293 24500
rect 293 24466 299 24500
rect 247 24450 299 24466
rect 149 24428 201 24438
rect 149 24394 167 24428
rect 167 24394 201 24428
rect 149 24386 201 24394
rect 247 24428 299 24438
rect 247 24394 259 24428
rect 259 24394 293 24428
rect 293 24394 299 24428
rect 247 24386 299 24394
rect 149 24355 201 24374
rect 149 24322 167 24355
rect 167 24322 201 24355
rect 247 24355 299 24374
rect 247 24322 259 24355
rect 259 24322 293 24355
rect 293 24322 299 24355
rect 149 24282 201 24310
rect 149 24258 167 24282
rect 167 24258 201 24282
rect 247 24282 299 24310
rect 247 24258 259 24282
rect 259 24258 293 24282
rect 293 24258 299 24282
rect 149 24209 201 24246
rect 149 24194 167 24209
rect 167 24194 201 24209
rect 247 24209 299 24246
rect 247 24194 259 24209
rect 259 24194 293 24209
rect 293 24194 299 24209
rect 149 24175 167 24182
rect 167 24175 201 24182
rect 149 24136 201 24175
rect 149 24130 167 24136
rect 167 24130 201 24136
rect 247 24175 259 24182
rect 259 24175 293 24182
rect 293 24175 299 24182
rect 247 24136 299 24175
rect 247 24130 259 24136
rect 259 24130 293 24136
rect 293 24130 299 24136
rect 149 24102 167 24118
rect 167 24102 201 24118
rect 149 24066 201 24102
rect 247 24102 259 24118
rect 259 24102 293 24118
rect 293 24102 299 24118
rect 247 24066 299 24102
rect 149 24029 167 24054
rect 167 24029 201 24054
rect 149 24002 201 24029
rect 247 24029 259 24054
rect 259 24029 293 24054
rect 293 24029 299 24054
rect 247 24002 299 24029
rect 149 23956 167 23990
rect 167 23956 201 23990
rect 149 23938 201 23956
rect 247 23956 259 23990
rect 259 23956 293 23990
rect 293 23956 299 23990
rect 247 23938 299 23956
rect 149 23917 201 23926
rect 149 23883 167 23917
rect 167 23883 201 23917
rect 149 23874 201 23883
rect 247 23917 299 23926
rect 247 23883 259 23917
rect 259 23883 293 23917
rect 293 23883 299 23917
rect 247 23874 299 23883
rect 149 23844 201 23862
rect 149 23810 167 23844
rect 167 23810 201 23844
rect 247 23844 299 23862
rect 247 23810 259 23844
rect 259 23810 293 23844
rect 293 23810 299 23844
rect 149 23771 201 23798
rect 149 23746 167 23771
rect 167 23746 201 23771
rect 247 23771 299 23798
rect 247 23746 259 23771
rect 259 23746 293 23771
rect 293 23746 299 23771
rect 149 23698 201 23734
rect 149 23682 167 23698
rect 167 23682 201 23698
rect 247 23698 299 23734
rect 247 23682 259 23698
rect 259 23682 293 23698
rect 293 23682 299 23698
rect 149 23664 167 23670
rect 167 23664 201 23670
rect 149 23625 201 23664
rect 149 23618 167 23625
rect 167 23618 201 23625
rect 247 23664 259 23670
rect 259 23664 293 23670
rect 293 23664 299 23670
rect 247 23625 299 23664
rect 247 23618 259 23625
rect 259 23618 293 23625
rect 293 23618 299 23625
rect 149 23591 167 23606
rect 167 23591 201 23606
rect 149 23554 201 23591
rect 247 23591 259 23606
rect 259 23591 293 23606
rect 293 23591 299 23606
rect 247 23554 299 23591
rect 149 23518 167 23542
rect 167 23518 201 23542
rect 149 23490 201 23518
rect 247 23518 259 23542
rect 259 23518 293 23542
rect 293 23518 299 23542
rect 247 23490 299 23518
rect 149 23445 167 23478
rect 167 23445 201 23478
rect 149 23426 201 23445
rect 247 23445 259 23478
rect 259 23445 293 23478
rect 293 23445 299 23478
rect 247 23426 299 23445
rect 149 23406 201 23414
rect 149 23372 167 23406
rect 167 23372 201 23406
rect 149 23362 201 23372
rect 247 23406 299 23414
rect 247 23372 259 23406
rect 259 23372 293 23406
rect 293 23372 299 23406
rect 247 23362 299 23372
rect 149 23333 201 23350
rect 149 23299 167 23333
rect 167 23299 201 23333
rect 149 23298 201 23299
rect 247 23333 299 23350
rect 247 23299 259 23333
rect 259 23299 293 23333
rect 293 23299 299 23333
rect 247 23298 299 23299
rect 149 23260 201 23286
rect 149 23234 167 23260
rect 167 23234 201 23260
rect 247 23260 299 23286
rect 247 23234 259 23260
rect 259 23234 293 23260
rect 293 23234 299 23260
rect 149 23187 201 23222
rect 149 23170 167 23187
rect 167 23170 201 23187
rect 247 23187 299 23222
rect 247 23170 259 23187
rect 259 23170 293 23187
rect 293 23170 299 23187
rect 149 23153 167 23158
rect 167 23153 201 23158
rect 149 23114 201 23153
rect 149 23106 167 23114
rect 167 23106 201 23114
rect 247 23153 259 23158
rect 259 23153 293 23158
rect 293 23153 299 23158
rect 247 23114 299 23153
rect 247 23106 259 23114
rect 259 23106 293 23114
rect 293 23106 299 23114
rect 149 23080 167 23094
rect 167 23080 201 23094
rect 149 23042 201 23080
rect 247 23080 259 23094
rect 259 23080 293 23094
rect 293 23080 299 23094
rect 247 23042 299 23080
rect 149 23007 167 23030
rect 167 23007 201 23030
rect 149 22978 201 23007
rect 247 23007 259 23030
rect 259 23007 293 23030
rect 293 23007 299 23030
rect 247 22978 299 23007
rect 149 22934 167 22966
rect 167 22934 201 22966
rect 149 22914 201 22934
rect 247 22934 259 22966
rect 259 22934 293 22966
rect 293 22934 299 22966
rect 247 22914 299 22934
rect 149 22895 201 22902
rect 149 22861 167 22895
rect 167 22861 201 22895
rect 149 22850 201 22861
rect 247 22895 299 22902
rect 247 22861 259 22895
rect 259 22861 293 22895
rect 293 22861 299 22895
rect 247 22850 299 22861
rect 149 22822 201 22838
rect 149 22788 167 22822
rect 167 22788 201 22822
rect 149 22786 201 22788
rect 247 22822 299 22838
rect 247 22788 259 22822
rect 259 22788 293 22822
rect 293 22788 299 22822
rect 247 22786 299 22788
rect 149 22749 201 22774
rect 149 22722 167 22749
rect 167 22722 201 22749
rect 247 22749 299 22774
rect 247 22722 259 22749
rect 259 22722 293 22749
rect 293 22722 299 22749
rect 149 22676 201 22710
rect 149 22658 167 22676
rect 167 22658 201 22676
rect 247 22676 299 22710
rect 247 22658 259 22676
rect 259 22658 293 22676
rect 293 22658 299 22676
rect 149 22642 167 22646
rect 167 22642 201 22646
rect 149 22603 201 22642
rect 149 22594 167 22603
rect 167 22594 201 22603
rect 247 22642 259 22646
rect 259 22642 293 22646
rect 293 22642 299 22646
rect 247 22603 299 22642
rect 247 22594 259 22603
rect 259 22594 293 22603
rect 293 22594 299 22603
rect 149 22569 167 22582
rect 167 22569 201 22582
rect 149 22530 201 22569
rect 247 22569 259 22582
rect 259 22569 293 22582
rect 293 22569 299 22582
rect 247 22530 299 22569
rect 149 22496 167 22518
rect 167 22496 201 22518
rect 149 22466 201 22496
rect 247 22496 259 22518
rect 259 22496 293 22518
rect 293 22496 299 22518
rect 247 22466 299 22496
rect 149 22423 167 22454
rect 167 22423 201 22454
rect 149 22402 201 22423
rect 247 22423 259 22454
rect 259 22423 293 22454
rect 293 22423 299 22454
rect 247 22402 299 22423
rect 149 22384 201 22390
rect 149 22350 167 22384
rect 167 22350 201 22384
rect 149 22338 201 22350
rect 247 22384 299 22390
rect 247 22350 259 22384
rect 259 22350 293 22384
rect 293 22350 299 22384
rect 247 22338 299 22350
rect 149 22311 201 22326
rect 149 22277 167 22311
rect 167 22277 201 22311
rect 149 22274 201 22277
rect 247 22311 299 22326
rect 247 22277 259 22311
rect 259 22277 293 22311
rect 293 22277 299 22311
rect 247 22274 299 22277
rect 149 22238 201 22262
rect 149 22210 167 22238
rect 167 22210 201 22238
rect 247 22238 299 22262
rect 247 22210 259 22238
rect 259 22210 293 22238
rect 293 22210 299 22238
rect 149 22165 201 22198
rect 149 22146 167 22165
rect 167 22146 201 22165
rect 247 22165 299 22198
rect 247 22146 259 22165
rect 259 22146 293 22165
rect 293 22146 299 22165
rect 149 22131 167 22134
rect 167 22131 201 22134
rect 149 22092 201 22131
rect 149 22082 167 22092
rect 167 22082 201 22092
rect 247 22131 259 22134
rect 259 22131 293 22134
rect 293 22131 299 22134
rect 247 22092 299 22131
rect 247 22082 259 22092
rect 259 22082 293 22092
rect 293 22082 299 22092
rect 149 22058 167 22070
rect 167 22058 201 22070
rect 149 22019 201 22058
rect 149 22018 167 22019
rect 167 22018 201 22019
rect 247 22058 259 22070
rect 259 22058 293 22070
rect 293 22058 299 22070
rect 247 22019 299 22058
rect 247 22018 259 22019
rect 259 22018 293 22019
rect 293 22018 299 22019
rect 149 21985 167 22006
rect 167 21985 201 22006
rect 149 21954 201 21985
rect 247 21985 259 22006
rect 259 21985 293 22006
rect 293 21985 299 22006
rect 247 21954 299 21985
rect 149 21912 167 21942
rect 167 21912 201 21942
rect 149 21890 201 21912
rect 247 21912 259 21942
rect 259 21912 293 21942
rect 293 21912 299 21942
rect 247 21890 299 21912
rect 149 21873 201 21878
rect 149 21839 167 21873
rect 167 21839 201 21873
rect 149 21826 201 21839
rect 247 21873 299 21878
rect 247 21839 259 21873
rect 259 21839 293 21873
rect 293 21839 299 21873
rect 247 21826 299 21839
rect 149 21800 201 21814
rect 149 21766 167 21800
rect 167 21766 201 21800
rect 149 21762 201 21766
rect 247 21800 299 21814
rect 247 21766 259 21800
rect 259 21766 293 21800
rect 293 21766 299 21800
rect 247 21762 299 21766
rect 149 21727 201 21750
rect 149 21698 167 21727
rect 167 21698 201 21727
rect 247 21727 299 21750
rect 247 21698 259 21727
rect 259 21698 293 21727
rect 293 21698 299 21727
rect 149 21654 201 21686
rect 149 21634 167 21654
rect 167 21634 201 21654
rect 247 21654 299 21686
rect 247 21634 259 21654
rect 259 21634 293 21654
rect 293 21634 299 21654
rect 149 21620 167 21622
rect 167 21620 201 21622
rect 149 21581 201 21620
rect 149 21570 167 21581
rect 167 21570 201 21581
rect 247 21620 259 21622
rect 259 21620 293 21622
rect 293 21620 299 21622
rect 247 21581 299 21620
rect 247 21570 259 21581
rect 259 21570 293 21581
rect 293 21570 299 21581
rect 149 21547 167 21558
rect 167 21547 201 21558
rect 149 21508 201 21547
rect 149 21506 167 21508
rect 167 21506 201 21508
rect 247 21547 259 21558
rect 259 21547 293 21558
rect 293 21547 299 21558
rect 247 21508 299 21547
rect 247 21506 259 21508
rect 259 21506 293 21508
rect 293 21506 299 21508
rect 149 21474 167 21494
rect 167 21474 201 21494
rect 149 21442 201 21474
rect 247 21474 259 21494
rect 259 21474 293 21494
rect 293 21474 299 21494
rect 247 21442 299 21474
rect 149 21401 167 21430
rect 167 21401 201 21430
rect 149 21378 201 21401
rect 247 21401 259 21430
rect 259 21401 293 21430
rect 293 21401 299 21430
rect 247 21378 299 21401
rect 149 21362 201 21366
rect 149 21328 167 21362
rect 167 21328 201 21362
rect 149 21314 201 21328
rect 247 21362 299 21366
rect 247 21328 259 21362
rect 259 21328 293 21362
rect 293 21328 299 21362
rect 247 21314 299 21328
rect 149 21289 201 21302
rect 149 21255 167 21289
rect 167 21255 201 21289
rect 149 21250 201 21255
rect 247 21289 299 21302
rect 247 21255 259 21289
rect 259 21255 293 21289
rect 293 21255 299 21289
rect 247 21250 299 21255
rect 149 21216 201 21238
rect 149 21186 167 21216
rect 167 21186 201 21216
rect 247 21216 299 21238
rect 247 21186 259 21216
rect 259 21186 293 21216
rect 293 21186 299 21216
rect 149 21143 201 21174
rect 149 21122 167 21143
rect 167 21122 201 21143
rect 247 21143 299 21174
rect 247 21122 259 21143
rect 259 21122 293 21143
rect 293 21122 299 21143
rect 149 21109 167 21110
rect 167 21109 201 21110
rect 149 21070 201 21109
rect 149 21058 167 21070
rect 167 21058 201 21070
rect 247 21109 259 21110
rect 259 21109 293 21110
rect 293 21109 299 21110
rect 247 21070 299 21109
rect 247 21058 259 21070
rect 259 21058 293 21070
rect 293 21058 299 21070
rect 149 21036 167 21046
rect 167 21036 201 21046
rect 149 20997 201 21036
rect 149 20994 167 20997
rect 167 20994 201 20997
rect 247 21036 259 21046
rect 259 21036 293 21046
rect 293 21036 299 21046
rect 247 20997 299 21036
rect 247 20994 259 20997
rect 259 20994 293 20997
rect 293 20994 299 20997
rect 149 20963 167 20982
rect 167 20963 201 20982
rect 149 20930 201 20963
rect 247 20963 259 20982
rect 259 20963 293 20982
rect 293 20963 299 20982
rect 247 20930 299 20963
rect 149 20890 167 20918
rect 167 20890 201 20918
rect 149 20866 201 20890
rect 247 20890 259 20918
rect 259 20890 293 20918
rect 293 20890 299 20918
rect 247 20866 299 20890
rect 149 20851 201 20854
rect 149 20817 167 20851
rect 167 20817 201 20851
rect 149 20802 201 20817
rect 247 20851 299 20854
rect 247 20817 259 20851
rect 259 20817 293 20851
rect 293 20817 299 20851
rect 247 20802 299 20817
rect 149 20778 201 20790
rect 149 20744 167 20778
rect 167 20744 201 20778
rect 149 20738 201 20744
rect 247 20778 299 20790
rect 247 20744 259 20778
rect 259 20744 293 20778
rect 293 20744 299 20778
rect 247 20738 299 20744
rect 149 20705 201 20726
rect 149 20674 167 20705
rect 167 20674 201 20705
rect 247 20705 299 20726
rect 247 20674 259 20705
rect 259 20674 293 20705
rect 293 20674 299 20705
rect 149 20632 201 20662
rect 149 20610 167 20632
rect 167 20610 201 20632
rect 247 20632 299 20662
rect 247 20610 259 20632
rect 259 20610 293 20632
rect 293 20610 299 20632
rect 149 20559 201 20598
rect 149 20546 167 20559
rect 167 20546 201 20559
rect 247 20559 299 20598
rect 247 20546 259 20559
rect 259 20546 293 20559
rect 293 20546 299 20559
rect 149 20525 167 20534
rect 167 20525 201 20534
rect 149 20486 201 20525
rect 149 20482 167 20486
rect 167 20482 201 20486
rect 247 20525 259 20534
rect 259 20525 293 20534
rect 293 20525 299 20534
rect 247 20486 299 20525
rect 247 20482 259 20486
rect 259 20482 293 20486
rect 293 20482 299 20486
rect 149 20452 167 20470
rect 167 20452 201 20470
rect 149 20418 201 20452
rect 247 20452 259 20470
rect 259 20452 293 20470
rect 293 20452 299 20470
rect 247 20418 299 20452
rect 149 20379 167 20406
rect 167 20379 201 20406
rect 149 20354 201 20379
rect 247 20379 259 20406
rect 259 20379 293 20406
rect 293 20379 299 20406
rect 247 20354 299 20379
rect 149 20340 201 20342
rect 149 20306 167 20340
rect 167 20306 201 20340
rect 149 20290 201 20306
rect 247 20340 299 20342
rect 247 20306 259 20340
rect 259 20306 293 20340
rect 293 20306 299 20340
rect 247 20290 299 20306
rect 149 20267 201 20277
rect 149 20233 167 20267
rect 167 20233 201 20267
rect 149 20225 201 20233
rect 247 20267 299 20277
rect 247 20233 259 20267
rect 259 20233 293 20267
rect 293 20233 299 20267
rect 247 20225 299 20233
rect 149 20194 201 20212
rect 149 20160 167 20194
rect 167 20160 201 20194
rect 247 20194 299 20212
rect 247 20160 259 20194
rect 259 20160 293 20194
rect 293 20160 299 20194
rect 149 20121 201 20147
rect 149 20095 167 20121
rect 167 20095 201 20121
rect 247 20121 299 20147
rect 247 20095 259 20121
rect 259 20095 293 20121
rect 293 20095 299 20121
rect 149 20048 201 20082
rect 149 20030 167 20048
rect 167 20030 201 20048
rect 247 20048 299 20082
rect 247 20030 259 20048
rect 259 20030 293 20048
rect 293 20030 299 20048
rect 149 20014 167 20017
rect 167 20014 201 20017
rect 149 19975 201 20014
rect 149 19965 167 19975
rect 167 19965 201 19975
rect 247 20014 259 20017
rect 259 20014 293 20017
rect 293 20014 299 20017
rect 247 19975 299 20014
rect 247 19965 259 19975
rect 259 19965 293 19975
rect 293 19965 299 19975
rect 149 19941 167 19952
rect 167 19941 201 19952
rect 149 19902 201 19941
rect 149 19900 167 19902
rect 167 19900 201 19902
rect 247 19941 259 19952
rect 259 19941 293 19952
rect 293 19941 299 19952
rect 247 19902 299 19941
rect 247 19900 259 19902
rect 259 19900 293 19902
rect 293 19900 299 19902
rect 149 19868 167 19887
rect 167 19868 201 19887
rect 149 19835 201 19868
rect 247 19868 259 19887
rect 259 19868 293 19887
rect 293 19868 299 19887
rect 247 19835 299 19868
rect 149 19795 167 19822
rect 167 19795 201 19822
rect 149 19770 201 19795
rect 247 19795 259 19822
rect 259 19795 293 19822
rect 293 19795 299 19822
rect 247 19770 299 19795
rect 149 19756 201 19757
rect 149 19722 167 19756
rect 167 19722 201 19756
rect 149 19705 201 19722
rect 247 19756 299 19757
rect 247 19722 259 19756
rect 259 19722 293 19756
rect 293 19722 299 19756
rect 247 19705 299 19722
rect 149 19683 201 19692
rect 149 19649 167 19683
rect 167 19649 201 19683
rect 149 19640 201 19649
rect 247 19683 299 19692
rect 247 19649 259 19683
rect 259 19649 293 19683
rect 293 19649 299 19683
rect 247 19640 299 19649
rect 149 19610 201 19627
rect 149 19576 167 19610
rect 167 19576 201 19610
rect 149 19575 201 19576
rect 247 19610 299 19627
rect 247 19576 259 19610
rect 259 19576 293 19610
rect 293 19576 299 19610
rect 247 19575 299 19576
rect 149 19537 201 19562
rect 149 19510 167 19537
rect 167 19510 201 19537
rect 247 19537 299 19562
rect 247 19510 259 19537
rect 259 19510 293 19537
rect 293 19510 299 19537
rect 149 19464 201 19497
rect 149 19445 167 19464
rect 167 19445 201 19464
rect 247 19464 299 19497
rect 247 19445 259 19464
rect 259 19445 293 19464
rect 293 19445 299 19464
rect 149 19430 167 19432
rect 167 19430 201 19432
rect 149 19391 201 19430
rect 149 19380 167 19391
rect 167 19380 201 19391
rect 247 19430 259 19432
rect 259 19430 293 19432
rect 293 19430 299 19432
rect 247 19391 299 19430
rect 247 19380 259 19391
rect 259 19380 293 19391
rect 293 19380 299 19391
rect 149 19357 167 19367
rect 167 19357 201 19367
rect 149 19318 201 19357
rect 149 19315 167 19318
rect 167 19315 201 19318
rect 247 19357 259 19367
rect 259 19357 293 19367
rect 293 19357 299 19367
rect 247 19318 299 19357
rect 247 19315 259 19318
rect 259 19315 293 19318
rect 293 19315 299 19318
rect 149 19284 167 19302
rect 167 19284 201 19302
rect 149 19250 201 19284
rect 247 19284 259 19302
rect 259 19284 293 19302
rect 293 19284 299 19302
rect 247 19250 299 19284
rect 149 19211 167 19237
rect 167 19211 201 19237
rect 149 19185 201 19211
rect 247 19211 259 19237
rect 259 19211 293 19237
rect 293 19211 299 19237
rect 247 19185 299 19211
rect 456 26012 508 26038
rect 456 25986 459 26012
rect 459 25986 493 26012
rect 493 25986 508 26012
rect 524 26012 576 26038
rect 524 25986 537 26012
rect 537 25986 571 26012
rect 571 25986 576 26012
rect 592 26012 644 26038
rect 660 26012 712 26038
rect 728 26012 780 26038
rect 796 26012 848 26038
rect 592 25986 615 26012
rect 615 25986 644 26012
rect 660 25986 693 26012
rect 693 25986 712 26012
rect 728 25986 771 26012
rect 771 25986 780 26012
rect 796 25986 805 26012
rect 805 25986 848 26012
rect 456 25940 508 25974
rect 456 25922 459 25940
rect 459 25922 493 25940
rect 493 25922 508 25940
rect 524 25940 576 25974
rect 524 25922 537 25940
rect 537 25922 571 25940
rect 571 25922 576 25940
rect 592 25940 644 25974
rect 660 25940 712 25974
rect 728 25940 780 25974
rect 796 25940 848 25974
rect 592 25922 615 25940
rect 615 25922 644 25940
rect 660 25922 693 25940
rect 693 25922 712 25940
rect 728 25922 771 25940
rect 771 25922 780 25940
rect 796 25922 805 25940
rect 805 25922 848 25940
rect 456 25906 459 25910
rect 459 25906 493 25910
rect 493 25906 508 25910
rect 456 25868 508 25906
rect 456 25858 459 25868
rect 459 25858 493 25868
rect 493 25858 508 25868
rect 524 25906 537 25910
rect 537 25906 571 25910
rect 571 25906 576 25910
rect 524 25868 576 25906
rect 524 25858 537 25868
rect 537 25858 571 25868
rect 571 25858 576 25868
rect 592 25906 615 25910
rect 615 25906 644 25910
rect 660 25906 693 25910
rect 693 25906 712 25910
rect 728 25906 771 25910
rect 771 25906 780 25910
rect 796 25906 805 25910
rect 805 25906 848 25910
rect 592 25868 644 25906
rect 660 25868 712 25906
rect 728 25868 780 25906
rect 796 25868 848 25906
rect 592 25858 615 25868
rect 615 25858 644 25868
rect 660 25858 693 25868
rect 693 25858 712 25868
rect 728 25858 771 25868
rect 771 25858 780 25868
rect 796 25858 805 25868
rect 805 25858 848 25868
rect 456 25834 459 25846
rect 459 25834 493 25846
rect 493 25834 508 25846
rect 456 25796 508 25834
rect 456 25794 459 25796
rect 459 25794 493 25796
rect 493 25794 508 25796
rect 524 25834 537 25846
rect 537 25834 571 25846
rect 571 25834 576 25846
rect 524 25796 576 25834
rect 524 25794 537 25796
rect 537 25794 571 25796
rect 571 25794 576 25796
rect 592 25834 615 25846
rect 615 25834 644 25846
rect 660 25834 693 25846
rect 693 25834 712 25846
rect 728 25834 771 25846
rect 771 25834 780 25846
rect 796 25834 805 25846
rect 805 25834 848 25846
rect 592 25796 644 25834
rect 660 25796 712 25834
rect 728 25796 780 25834
rect 796 25796 848 25834
rect 592 25794 615 25796
rect 615 25794 644 25796
rect 660 25794 693 25796
rect 693 25794 712 25796
rect 728 25794 771 25796
rect 771 25794 780 25796
rect 796 25794 805 25796
rect 805 25794 848 25796
rect 456 25762 459 25782
rect 459 25762 493 25782
rect 493 25762 508 25782
rect 456 25730 508 25762
rect 524 25762 537 25782
rect 537 25762 571 25782
rect 571 25762 576 25782
rect 524 25730 576 25762
rect 592 25762 615 25782
rect 615 25762 644 25782
rect 660 25762 693 25782
rect 693 25762 712 25782
rect 728 25762 771 25782
rect 771 25762 780 25782
rect 796 25762 805 25782
rect 805 25762 848 25782
rect 592 25730 644 25762
rect 660 25730 712 25762
rect 728 25730 780 25762
rect 796 25730 848 25762
rect 456 25690 459 25718
rect 459 25690 493 25718
rect 493 25690 508 25718
rect 456 25666 508 25690
rect 524 25690 537 25718
rect 537 25690 571 25718
rect 571 25690 576 25718
rect 524 25666 576 25690
rect 592 25690 615 25718
rect 615 25690 644 25718
rect 660 25690 693 25718
rect 693 25690 712 25718
rect 728 25690 771 25718
rect 771 25690 780 25718
rect 796 25690 805 25718
rect 805 25690 848 25718
rect 592 25666 644 25690
rect 660 25666 712 25690
rect 728 25666 780 25690
rect 796 25666 848 25690
rect 456 25652 508 25654
rect 456 25618 459 25652
rect 459 25618 493 25652
rect 493 25618 508 25652
rect 456 25602 508 25618
rect 524 25652 576 25654
rect 524 25618 537 25652
rect 537 25618 571 25652
rect 571 25618 576 25652
rect 524 25602 576 25618
rect 592 25652 644 25654
rect 660 25652 712 25654
rect 728 25652 780 25654
rect 796 25652 848 25654
rect 592 25618 615 25652
rect 615 25618 644 25652
rect 660 25618 693 25652
rect 693 25618 712 25652
rect 728 25618 771 25652
rect 771 25618 780 25652
rect 796 25618 805 25652
rect 805 25618 848 25652
rect 592 25602 644 25618
rect 660 25602 712 25618
rect 728 25602 780 25618
rect 796 25602 848 25618
rect 456 25580 508 25590
rect 456 25546 459 25580
rect 459 25546 493 25580
rect 493 25546 508 25580
rect 456 25538 508 25546
rect 524 25580 576 25590
rect 524 25546 537 25580
rect 537 25546 571 25580
rect 571 25546 576 25580
rect 524 25538 576 25546
rect 592 25580 644 25590
rect 660 25580 712 25590
rect 728 25580 780 25590
rect 796 25580 848 25590
rect 592 25546 615 25580
rect 615 25546 644 25580
rect 660 25546 693 25580
rect 693 25546 712 25580
rect 728 25546 771 25580
rect 771 25546 780 25580
rect 796 25546 805 25580
rect 805 25546 848 25580
rect 592 25538 644 25546
rect 660 25538 712 25546
rect 728 25538 780 25546
rect 796 25538 848 25546
rect 456 25508 508 25526
rect 456 25474 459 25508
rect 459 25474 493 25508
rect 493 25474 508 25508
rect 524 25508 576 25526
rect 524 25474 537 25508
rect 537 25474 571 25508
rect 571 25474 576 25508
rect 592 25508 644 25526
rect 660 25508 712 25526
rect 728 25508 780 25526
rect 796 25508 848 25526
rect 592 25474 615 25508
rect 615 25474 644 25508
rect 660 25474 693 25508
rect 693 25474 712 25508
rect 728 25474 771 25508
rect 771 25474 780 25508
rect 796 25474 805 25508
rect 805 25474 848 25508
rect 456 25436 508 25462
rect 456 25410 459 25436
rect 459 25410 493 25436
rect 493 25410 508 25436
rect 524 25436 576 25462
rect 524 25410 537 25436
rect 537 25410 571 25436
rect 571 25410 576 25436
rect 592 25436 644 25462
rect 660 25436 712 25462
rect 728 25436 780 25462
rect 796 25436 848 25462
rect 592 25410 615 25436
rect 615 25410 644 25436
rect 660 25410 693 25436
rect 693 25410 712 25436
rect 728 25410 771 25436
rect 771 25410 780 25436
rect 796 25410 805 25436
rect 805 25410 848 25436
rect 456 25364 508 25398
rect 456 25346 459 25364
rect 459 25346 493 25364
rect 493 25346 508 25364
rect 524 25364 576 25398
rect 524 25346 537 25364
rect 537 25346 571 25364
rect 571 25346 576 25364
rect 592 25364 644 25398
rect 660 25364 712 25398
rect 728 25364 780 25398
rect 796 25364 848 25398
rect 592 25346 615 25364
rect 615 25346 644 25364
rect 660 25346 693 25364
rect 693 25346 712 25364
rect 728 25346 771 25364
rect 771 25346 780 25364
rect 796 25346 805 25364
rect 805 25346 848 25364
rect 456 25330 459 25334
rect 459 25330 493 25334
rect 493 25330 508 25334
rect 456 25292 508 25330
rect 456 25282 459 25292
rect 459 25282 493 25292
rect 493 25282 508 25292
rect 524 25330 537 25334
rect 537 25330 571 25334
rect 571 25330 576 25334
rect 524 25292 576 25330
rect 524 25282 537 25292
rect 537 25282 571 25292
rect 571 25282 576 25292
rect 592 25330 615 25334
rect 615 25330 644 25334
rect 660 25330 693 25334
rect 693 25330 712 25334
rect 728 25330 771 25334
rect 771 25330 780 25334
rect 796 25330 805 25334
rect 805 25330 848 25334
rect 592 25292 644 25330
rect 660 25292 712 25330
rect 728 25292 780 25330
rect 796 25292 848 25330
rect 592 25282 615 25292
rect 615 25282 644 25292
rect 660 25282 693 25292
rect 693 25282 712 25292
rect 728 25282 771 25292
rect 771 25282 780 25292
rect 796 25282 805 25292
rect 805 25282 848 25292
rect 456 25258 459 25270
rect 459 25258 493 25270
rect 493 25258 508 25270
rect 456 25220 508 25258
rect 456 25218 459 25220
rect 459 25218 493 25220
rect 493 25218 508 25220
rect 524 25258 537 25270
rect 537 25258 571 25270
rect 571 25258 576 25270
rect 524 25220 576 25258
rect 524 25218 537 25220
rect 537 25218 571 25220
rect 571 25218 576 25220
rect 592 25258 615 25270
rect 615 25258 644 25270
rect 660 25258 693 25270
rect 693 25258 712 25270
rect 728 25258 771 25270
rect 771 25258 780 25270
rect 796 25258 805 25270
rect 805 25258 848 25270
rect 592 25220 644 25258
rect 660 25220 712 25258
rect 728 25220 780 25258
rect 796 25220 848 25258
rect 592 25218 615 25220
rect 615 25218 644 25220
rect 660 25218 693 25220
rect 693 25218 712 25220
rect 728 25218 771 25220
rect 771 25218 780 25220
rect 796 25218 805 25220
rect 805 25218 848 25220
rect 456 25186 459 25206
rect 459 25186 493 25206
rect 493 25186 508 25206
rect 456 25154 508 25186
rect 524 25186 537 25206
rect 537 25186 571 25206
rect 571 25186 576 25206
rect 524 25154 576 25186
rect 592 25186 615 25206
rect 615 25186 644 25206
rect 660 25186 693 25206
rect 693 25186 712 25206
rect 728 25186 771 25206
rect 771 25186 780 25206
rect 796 25186 805 25206
rect 805 25186 848 25206
rect 592 25154 644 25186
rect 660 25154 712 25186
rect 728 25154 780 25186
rect 796 25154 848 25186
rect 456 25114 459 25142
rect 459 25114 493 25142
rect 493 25114 508 25142
rect 456 25090 508 25114
rect 524 25114 537 25142
rect 537 25114 571 25142
rect 571 25114 576 25142
rect 524 25090 576 25114
rect 592 25114 615 25142
rect 615 25114 644 25142
rect 660 25114 693 25142
rect 693 25114 712 25142
rect 728 25114 771 25142
rect 771 25114 780 25142
rect 796 25114 805 25142
rect 805 25114 848 25142
rect 592 25090 644 25114
rect 660 25090 712 25114
rect 728 25090 780 25114
rect 796 25090 848 25114
rect 456 25076 508 25078
rect 456 25042 459 25076
rect 459 25042 493 25076
rect 493 25042 508 25076
rect 456 25026 508 25042
rect 524 25076 576 25078
rect 524 25042 537 25076
rect 537 25042 571 25076
rect 571 25042 576 25076
rect 524 25026 576 25042
rect 592 25076 644 25078
rect 660 25076 712 25078
rect 728 25076 780 25078
rect 796 25076 848 25078
rect 592 25042 615 25076
rect 615 25042 644 25076
rect 660 25042 693 25076
rect 693 25042 712 25076
rect 728 25042 771 25076
rect 771 25042 780 25076
rect 796 25042 805 25076
rect 805 25042 848 25076
rect 592 25026 644 25042
rect 660 25026 712 25042
rect 728 25026 780 25042
rect 796 25026 848 25042
rect 456 25004 508 25014
rect 456 24970 459 25004
rect 459 24970 493 25004
rect 493 24970 508 25004
rect 456 24962 508 24970
rect 524 25004 576 25014
rect 524 24970 537 25004
rect 537 24970 571 25004
rect 571 24970 576 25004
rect 524 24962 576 24970
rect 592 25004 644 25014
rect 660 25004 712 25014
rect 728 25004 780 25014
rect 796 25004 848 25014
rect 592 24970 615 25004
rect 615 24970 644 25004
rect 660 24970 693 25004
rect 693 24970 712 25004
rect 728 24970 771 25004
rect 771 24970 780 25004
rect 796 24970 805 25004
rect 805 24970 848 25004
rect 592 24962 644 24970
rect 660 24962 712 24970
rect 728 24962 780 24970
rect 796 24962 848 24970
rect 456 24932 508 24950
rect 456 24898 459 24932
rect 459 24898 493 24932
rect 493 24898 508 24932
rect 524 24932 576 24950
rect 524 24898 537 24932
rect 537 24898 571 24932
rect 571 24898 576 24932
rect 592 24932 644 24950
rect 660 24932 712 24950
rect 728 24932 780 24950
rect 796 24932 848 24950
rect 592 24898 615 24932
rect 615 24898 644 24932
rect 660 24898 693 24932
rect 693 24898 712 24932
rect 728 24898 771 24932
rect 771 24898 780 24932
rect 796 24898 805 24932
rect 805 24898 848 24932
rect 456 24860 508 24886
rect 456 24834 459 24860
rect 459 24834 493 24860
rect 493 24834 508 24860
rect 524 24860 576 24886
rect 524 24834 537 24860
rect 537 24834 571 24860
rect 571 24834 576 24860
rect 592 24860 644 24886
rect 660 24860 712 24886
rect 728 24860 780 24886
rect 796 24860 848 24886
rect 592 24834 615 24860
rect 615 24834 644 24860
rect 660 24834 693 24860
rect 693 24834 712 24860
rect 728 24834 771 24860
rect 771 24834 780 24860
rect 796 24834 805 24860
rect 805 24834 848 24860
rect 456 24788 508 24822
rect 456 24770 459 24788
rect 459 24770 493 24788
rect 493 24770 508 24788
rect 524 24788 576 24822
rect 524 24770 537 24788
rect 537 24770 571 24788
rect 571 24770 576 24788
rect 592 24788 644 24822
rect 660 24788 712 24822
rect 728 24788 780 24822
rect 796 24788 848 24822
rect 592 24770 615 24788
rect 615 24770 644 24788
rect 660 24770 693 24788
rect 693 24770 712 24788
rect 728 24770 771 24788
rect 771 24770 780 24788
rect 796 24770 805 24788
rect 805 24770 848 24788
rect 456 24754 459 24758
rect 459 24754 493 24758
rect 493 24754 508 24758
rect 456 24716 508 24754
rect 456 24706 459 24716
rect 459 24706 493 24716
rect 493 24706 508 24716
rect 524 24754 537 24758
rect 537 24754 571 24758
rect 571 24754 576 24758
rect 524 24716 576 24754
rect 524 24706 537 24716
rect 537 24706 571 24716
rect 571 24706 576 24716
rect 592 24754 615 24758
rect 615 24754 644 24758
rect 660 24754 693 24758
rect 693 24754 712 24758
rect 728 24754 771 24758
rect 771 24754 780 24758
rect 796 24754 805 24758
rect 805 24754 848 24758
rect 592 24716 644 24754
rect 660 24716 712 24754
rect 728 24716 780 24754
rect 796 24716 848 24754
rect 592 24706 615 24716
rect 615 24706 644 24716
rect 660 24706 693 24716
rect 693 24706 712 24716
rect 728 24706 771 24716
rect 771 24706 780 24716
rect 796 24706 805 24716
rect 805 24706 848 24716
rect 456 24682 459 24694
rect 459 24682 493 24694
rect 493 24682 508 24694
rect 456 24644 508 24682
rect 456 24642 459 24644
rect 459 24642 493 24644
rect 493 24642 508 24644
rect 524 24682 537 24694
rect 537 24682 571 24694
rect 571 24682 576 24694
rect 524 24644 576 24682
rect 524 24642 537 24644
rect 537 24642 571 24644
rect 571 24642 576 24644
rect 592 24682 615 24694
rect 615 24682 644 24694
rect 660 24682 693 24694
rect 693 24682 712 24694
rect 728 24682 771 24694
rect 771 24682 780 24694
rect 796 24682 805 24694
rect 805 24682 848 24694
rect 592 24644 644 24682
rect 660 24644 712 24682
rect 728 24644 780 24682
rect 796 24644 848 24682
rect 592 24642 615 24644
rect 615 24642 644 24644
rect 660 24642 693 24644
rect 693 24642 712 24644
rect 728 24642 771 24644
rect 771 24642 780 24644
rect 796 24642 805 24644
rect 805 24642 848 24644
rect 456 24610 459 24630
rect 459 24610 493 24630
rect 493 24610 508 24630
rect 456 24578 508 24610
rect 524 24610 537 24630
rect 537 24610 571 24630
rect 571 24610 576 24630
rect 524 24578 576 24610
rect 592 24610 615 24630
rect 615 24610 644 24630
rect 660 24610 693 24630
rect 693 24610 712 24630
rect 728 24610 771 24630
rect 771 24610 780 24630
rect 796 24610 805 24630
rect 805 24610 848 24630
rect 592 24578 644 24610
rect 660 24578 712 24610
rect 728 24578 780 24610
rect 796 24578 848 24610
rect 456 24538 459 24566
rect 459 24538 493 24566
rect 493 24538 508 24566
rect 456 24514 508 24538
rect 524 24538 537 24566
rect 537 24538 571 24566
rect 571 24538 576 24566
rect 524 24514 576 24538
rect 592 24538 615 24566
rect 615 24538 644 24566
rect 660 24538 693 24566
rect 693 24538 712 24566
rect 728 24538 771 24566
rect 771 24538 780 24566
rect 796 24538 805 24566
rect 805 24538 848 24566
rect 592 24514 644 24538
rect 660 24514 712 24538
rect 728 24514 780 24538
rect 796 24514 848 24538
rect 456 24500 508 24502
rect 456 24466 459 24500
rect 459 24466 493 24500
rect 493 24466 508 24500
rect 456 24450 508 24466
rect 524 24500 576 24502
rect 524 24466 537 24500
rect 537 24466 571 24500
rect 571 24466 576 24500
rect 524 24450 576 24466
rect 592 24500 644 24502
rect 660 24500 712 24502
rect 728 24500 780 24502
rect 796 24500 848 24502
rect 592 24466 615 24500
rect 615 24466 644 24500
rect 660 24466 693 24500
rect 693 24466 712 24500
rect 728 24466 771 24500
rect 771 24466 780 24500
rect 796 24466 805 24500
rect 805 24466 848 24500
rect 592 24450 644 24466
rect 660 24450 712 24466
rect 728 24450 780 24466
rect 796 24450 848 24466
rect 456 24428 508 24438
rect 456 24394 459 24428
rect 459 24394 493 24428
rect 493 24394 508 24428
rect 456 24386 508 24394
rect 524 24428 576 24438
rect 524 24394 537 24428
rect 537 24394 571 24428
rect 571 24394 576 24428
rect 524 24386 576 24394
rect 592 24428 644 24438
rect 660 24428 712 24438
rect 728 24428 780 24438
rect 796 24428 848 24438
rect 592 24394 615 24428
rect 615 24394 644 24428
rect 660 24394 693 24428
rect 693 24394 712 24428
rect 728 24394 771 24428
rect 771 24394 780 24428
rect 796 24394 805 24428
rect 805 24394 848 24428
rect 592 24386 644 24394
rect 660 24386 712 24394
rect 728 24386 780 24394
rect 796 24386 848 24394
rect 456 24355 508 24374
rect 456 24322 459 24355
rect 459 24322 493 24355
rect 493 24322 508 24355
rect 524 24355 576 24374
rect 524 24322 537 24355
rect 537 24322 571 24355
rect 571 24322 576 24355
rect 592 24355 644 24374
rect 660 24355 712 24374
rect 728 24355 780 24374
rect 796 24355 848 24374
rect 592 24322 615 24355
rect 615 24322 644 24355
rect 660 24322 693 24355
rect 693 24322 712 24355
rect 728 24322 771 24355
rect 771 24322 780 24355
rect 796 24322 805 24355
rect 805 24322 848 24355
rect 456 24282 508 24310
rect 456 24258 459 24282
rect 459 24258 493 24282
rect 493 24258 508 24282
rect 524 24282 576 24310
rect 524 24258 537 24282
rect 537 24258 571 24282
rect 571 24258 576 24282
rect 592 24282 644 24310
rect 660 24282 712 24310
rect 728 24282 780 24310
rect 796 24282 848 24310
rect 592 24258 615 24282
rect 615 24258 644 24282
rect 660 24258 693 24282
rect 693 24258 712 24282
rect 728 24258 771 24282
rect 771 24258 780 24282
rect 796 24258 805 24282
rect 805 24258 848 24282
rect 456 24209 508 24246
rect 456 24194 459 24209
rect 459 24194 493 24209
rect 493 24194 508 24209
rect 524 24209 576 24246
rect 524 24194 537 24209
rect 537 24194 571 24209
rect 571 24194 576 24209
rect 592 24209 644 24246
rect 660 24209 712 24246
rect 728 24209 780 24246
rect 796 24209 848 24246
rect 592 24194 615 24209
rect 615 24194 644 24209
rect 660 24194 693 24209
rect 693 24194 712 24209
rect 728 24194 771 24209
rect 771 24194 780 24209
rect 796 24194 805 24209
rect 805 24194 848 24209
rect 456 24175 459 24182
rect 459 24175 493 24182
rect 493 24175 508 24182
rect 456 24136 508 24175
rect 456 24130 459 24136
rect 459 24130 493 24136
rect 493 24130 508 24136
rect 524 24175 537 24182
rect 537 24175 571 24182
rect 571 24175 576 24182
rect 524 24136 576 24175
rect 524 24130 537 24136
rect 537 24130 571 24136
rect 571 24130 576 24136
rect 592 24175 615 24182
rect 615 24175 644 24182
rect 660 24175 693 24182
rect 693 24175 712 24182
rect 728 24175 771 24182
rect 771 24175 780 24182
rect 796 24175 805 24182
rect 805 24175 848 24182
rect 592 24136 644 24175
rect 660 24136 712 24175
rect 728 24136 780 24175
rect 796 24136 848 24175
rect 592 24130 615 24136
rect 615 24130 644 24136
rect 660 24130 693 24136
rect 693 24130 712 24136
rect 728 24130 771 24136
rect 771 24130 780 24136
rect 796 24130 805 24136
rect 805 24130 848 24136
rect 456 24102 459 24118
rect 459 24102 493 24118
rect 493 24102 508 24118
rect 456 24066 508 24102
rect 524 24102 537 24118
rect 537 24102 571 24118
rect 571 24102 576 24118
rect 524 24066 576 24102
rect 592 24102 615 24118
rect 615 24102 644 24118
rect 660 24102 693 24118
rect 693 24102 712 24118
rect 728 24102 771 24118
rect 771 24102 780 24118
rect 796 24102 805 24118
rect 805 24102 848 24118
rect 592 24066 644 24102
rect 660 24066 712 24102
rect 728 24066 780 24102
rect 796 24066 848 24102
rect 456 24029 459 24054
rect 459 24029 493 24054
rect 493 24029 508 24054
rect 456 24002 508 24029
rect 524 24029 537 24054
rect 537 24029 571 24054
rect 571 24029 576 24054
rect 524 24002 576 24029
rect 592 24029 615 24054
rect 615 24029 644 24054
rect 660 24029 693 24054
rect 693 24029 712 24054
rect 728 24029 771 24054
rect 771 24029 780 24054
rect 796 24029 805 24054
rect 805 24029 848 24054
rect 592 24002 644 24029
rect 660 24002 712 24029
rect 728 24002 780 24029
rect 796 24002 848 24029
rect 456 23956 459 23990
rect 459 23956 493 23990
rect 493 23956 508 23990
rect 456 23938 508 23956
rect 524 23956 537 23990
rect 537 23956 571 23990
rect 571 23956 576 23990
rect 524 23938 576 23956
rect 592 23956 615 23990
rect 615 23956 644 23990
rect 660 23956 693 23990
rect 693 23956 712 23990
rect 728 23956 771 23990
rect 771 23956 780 23990
rect 796 23956 805 23990
rect 805 23956 848 23990
rect 592 23938 644 23956
rect 660 23938 712 23956
rect 728 23938 780 23956
rect 796 23938 848 23956
rect 456 23917 508 23926
rect 456 23883 459 23917
rect 459 23883 493 23917
rect 493 23883 508 23917
rect 456 23874 508 23883
rect 524 23917 576 23926
rect 524 23883 537 23917
rect 537 23883 571 23917
rect 571 23883 576 23917
rect 524 23874 576 23883
rect 592 23917 644 23926
rect 660 23917 712 23926
rect 728 23917 780 23926
rect 796 23917 848 23926
rect 592 23883 615 23917
rect 615 23883 644 23917
rect 660 23883 693 23917
rect 693 23883 712 23917
rect 728 23883 771 23917
rect 771 23883 780 23917
rect 796 23883 805 23917
rect 805 23883 848 23917
rect 592 23874 644 23883
rect 660 23874 712 23883
rect 728 23874 780 23883
rect 796 23874 848 23883
rect 456 23844 508 23862
rect 456 23810 459 23844
rect 459 23810 493 23844
rect 493 23810 508 23844
rect 524 23844 576 23862
rect 524 23810 537 23844
rect 537 23810 571 23844
rect 571 23810 576 23844
rect 592 23844 644 23862
rect 660 23844 712 23862
rect 728 23844 780 23862
rect 796 23844 848 23862
rect 592 23810 615 23844
rect 615 23810 644 23844
rect 660 23810 693 23844
rect 693 23810 712 23844
rect 728 23810 771 23844
rect 771 23810 780 23844
rect 796 23810 805 23844
rect 805 23810 848 23844
rect 456 23771 508 23798
rect 456 23746 459 23771
rect 459 23746 493 23771
rect 493 23746 508 23771
rect 524 23771 576 23798
rect 524 23746 537 23771
rect 537 23746 571 23771
rect 571 23746 576 23771
rect 592 23771 644 23798
rect 660 23771 712 23798
rect 728 23771 780 23798
rect 796 23771 848 23798
rect 592 23746 615 23771
rect 615 23746 644 23771
rect 660 23746 693 23771
rect 693 23746 712 23771
rect 728 23746 771 23771
rect 771 23746 780 23771
rect 796 23746 805 23771
rect 805 23746 848 23771
rect 456 23698 508 23734
rect 456 23682 459 23698
rect 459 23682 493 23698
rect 493 23682 508 23698
rect 524 23698 576 23734
rect 524 23682 537 23698
rect 537 23682 571 23698
rect 571 23682 576 23698
rect 592 23698 644 23734
rect 660 23698 712 23734
rect 728 23698 780 23734
rect 796 23698 848 23734
rect 592 23682 615 23698
rect 615 23682 644 23698
rect 660 23682 693 23698
rect 693 23682 712 23698
rect 728 23682 771 23698
rect 771 23682 780 23698
rect 796 23682 805 23698
rect 805 23682 848 23698
rect 456 23664 459 23670
rect 459 23664 493 23670
rect 493 23664 508 23670
rect 456 23625 508 23664
rect 456 23618 459 23625
rect 459 23618 493 23625
rect 493 23618 508 23625
rect 524 23664 537 23670
rect 537 23664 571 23670
rect 571 23664 576 23670
rect 524 23625 576 23664
rect 524 23618 537 23625
rect 537 23618 571 23625
rect 571 23618 576 23625
rect 592 23664 615 23670
rect 615 23664 644 23670
rect 660 23664 693 23670
rect 693 23664 712 23670
rect 728 23664 771 23670
rect 771 23664 780 23670
rect 796 23664 805 23670
rect 805 23664 848 23670
rect 592 23625 644 23664
rect 660 23625 712 23664
rect 728 23625 780 23664
rect 796 23625 848 23664
rect 592 23618 615 23625
rect 615 23618 644 23625
rect 660 23618 693 23625
rect 693 23618 712 23625
rect 728 23618 771 23625
rect 771 23618 780 23625
rect 796 23618 805 23625
rect 805 23618 848 23625
rect 456 23591 459 23606
rect 459 23591 493 23606
rect 493 23591 508 23606
rect 456 23554 508 23591
rect 524 23591 537 23606
rect 537 23591 571 23606
rect 571 23591 576 23606
rect 524 23554 576 23591
rect 592 23591 615 23606
rect 615 23591 644 23606
rect 660 23591 693 23606
rect 693 23591 712 23606
rect 728 23591 771 23606
rect 771 23591 780 23606
rect 796 23591 805 23606
rect 805 23591 848 23606
rect 592 23554 644 23591
rect 660 23554 712 23591
rect 728 23554 780 23591
rect 796 23554 848 23591
rect 456 23518 459 23542
rect 459 23518 493 23542
rect 493 23518 508 23542
rect 456 23490 508 23518
rect 524 23518 537 23542
rect 537 23518 571 23542
rect 571 23518 576 23542
rect 524 23490 576 23518
rect 592 23518 615 23542
rect 615 23518 644 23542
rect 660 23518 693 23542
rect 693 23518 712 23542
rect 728 23518 771 23542
rect 771 23518 780 23542
rect 796 23518 805 23542
rect 805 23518 848 23542
rect 592 23490 644 23518
rect 660 23490 712 23518
rect 728 23490 780 23518
rect 796 23490 848 23518
rect 456 23445 459 23478
rect 459 23445 493 23478
rect 493 23445 508 23478
rect 456 23426 508 23445
rect 524 23445 537 23478
rect 537 23445 571 23478
rect 571 23445 576 23478
rect 524 23426 576 23445
rect 592 23445 615 23478
rect 615 23445 644 23478
rect 660 23445 693 23478
rect 693 23445 712 23478
rect 728 23445 771 23478
rect 771 23445 780 23478
rect 796 23445 805 23478
rect 805 23445 848 23478
rect 592 23426 644 23445
rect 660 23426 712 23445
rect 728 23426 780 23445
rect 796 23426 848 23445
rect 456 23406 508 23414
rect 456 23372 459 23406
rect 459 23372 493 23406
rect 493 23372 508 23406
rect 456 23362 508 23372
rect 524 23406 576 23414
rect 524 23372 537 23406
rect 537 23372 571 23406
rect 571 23372 576 23406
rect 524 23362 576 23372
rect 592 23406 644 23414
rect 660 23406 712 23414
rect 728 23406 780 23414
rect 796 23406 848 23414
rect 592 23372 615 23406
rect 615 23372 644 23406
rect 660 23372 693 23406
rect 693 23372 712 23406
rect 728 23372 771 23406
rect 771 23372 780 23406
rect 796 23372 805 23406
rect 805 23372 848 23406
rect 592 23362 644 23372
rect 660 23362 712 23372
rect 728 23362 780 23372
rect 796 23362 848 23372
rect 456 23333 508 23350
rect 456 23299 459 23333
rect 459 23299 493 23333
rect 493 23299 508 23333
rect 456 23298 508 23299
rect 524 23333 576 23350
rect 524 23299 537 23333
rect 537 23299 571 23333
rect 571 23299 576 23333
rect 524 23298 576 23299
rect 592 23333 644 23350
rect 660 23333 712 23350
rect 728 23333 780 23350
rect 796 23333 848 23350
rect 592 23299 615 23333
rect 615 23299 644 23333
rect 660 23299 693 23333
rect 693 23299 712 23333
rect 728 23299 771 23333
rect 771 23299 780 23333
rect 796 23299 805 23333
rect 805 23299 848 23333
rect 592 23298 644 23299
rect 660 23298 712 23299
rect 728 23298 780 23299
rect 796 23298 848 23299
rect 456 23260 508 23286
rect 456 23234 459 23260
rect 459 23234 493 23260
rect 493 23234 508 23260
rect 524 23260 576 23286
rect 524 23234 537 23260
rect 537 23234 571 23260
rect 571 23234 576 23260
rect 592 23260 644 23286
rect 660 23260 712 23286
rect 728 23260 780 23286
rect 796 23260 848 23286
rect 592 23234 615 23260
rect 615 23234 644 23260
rect 660 23234 693 23260
rect 693 23234 712 23260
rect 728 23234 771 23260
rect 771 23234 780 23260
rect 796 23234 805 23260
rect 805 23234 848 23260
rect 456 23187 508 23222
rect 456 23170 459 23187
rect 459 23170 493 23187
rect 493 23170 508 23187
rect 524 23187 576 23222
rect 524 23170 537 23187
rect 537 23170 571 23187
rect 571 23170 576 23187
rect 592 23187 644 23222
rect 660 23187 712 23222
rect 728 23187 780 23222
rect 796 23187 848 23222
rect 592 23170 615 23187
rect 615 23170 644 23187
rect 660 23170 693 23187
rect 693 23170 712 23187
rect 728 23170 771 23187
rect 771 23170 780 23187
rect 796 23170 805 23187
rect 805 23170 848 23187
rect 456 23153 459 23158
rect 459 23153 493 23158
rect 493 23153 508 23158
rect 456 23114 508 23153
rect 456 23106 459 23114
rect 459 23106 493 23114
rect 493 23106 508 23114
rect 524 23153 537 23158
rect 537 23153 571 23158
rect 571 23153 576 23158
rect 524 23114 576 23153
rect 524 23106 537 23114
rect 537 23106 571 23114
rect 571 23106 576 23114
rect 592 23153 615 23158
rect 615 23153 644 23158
rect 660 23153 693 23158
rect 693 23153 712 23158
rect 728 23153 771 23158
rect 771 23153 780 23158
rect 796 23153 805 23158
rect 805 23153 848 23158
rect 592 23114 644 23153
rect 660 23114 712 23153
rect 728 23114 780 23153
rect 796 23114 848 23153
rect 592 23106 615 23114
rect 615 23106 644 23114
rect 660 23106 693 23114
rect 693 23106 712 23114
rect 728 23106 771 23114
rect 771 23106 780 23114
rect 796 23106 805 23114
rect 805 23106 848 23114
rect 456 23080 459 23094
rect 459 23080 493 23094
rect 493 23080 508 23094
rect 456 23042 508 23080
rect 524 23080 537 23094
rect 537 23080 571 23094
rect 571 23080 576 23094
rect 524 23042 576 23080
rect 592 23080 615 23094
rect 615 23080 644 23094
rect 660 23080 693 23094
rect 693 23080 712 23094
rect 728 23080 771 23094
rect 771 23080 780 23094
rect 796 23080 805 23094
rect 805 23080 848 23094
rect 592 23042 644 23080
rect 660 23042 712 23080
rect 728 23042 780 23080
rect 796 23042 848 23080
rect 456 23007 459 23030
rect 459 23007 493 23030
rect 493 23007 508 23030
rect 456 22978 508 23007
rect 524 23007 537 23030
rect 537 23007 571 23030
rect 571 23007 576 23030
rect 524 22978 576 23007
rect 592 23007 615 23030
rect 615 23007 644 23030
rect 660 23007 693 23030
rect 693 23007 712 23030
rect 728 23007 771 23030
rect 771 23007 780 23030
rect 796 23007 805 23030
rect 805 23007 848 23030
rect 592 22978 644 23007
rect 660 22978 712 23007
rect 728 22978 780 23007
rect 796 22978 848 23007
rect 456 22934 459 22966
rect 459 22934 493 22966
rect 493 22934 508 22966
rect 456 22914 508 22934
rect 524 22934 537 22966
rect 537 22934 571 22966
rect 571 22934 576 22966
rect 524 22914 576 22934
rect 592 22934 615 22966
rect 615 22934 644 22966
rect 660 22934 693 22966
rect 693 22934 712 22966
rect 728 22934 771 22966
rect 771 22934 780 22966
rect 796 22934 805 22966
rect 805 22934 848 22966
rect 592 22914 644 22934
rect 660 22914 712 22934
rect 728 22914 780 22934
rect 796 22914 848 22934
rect 456 22895 508 22902
rect 456 22861 459 22895
rect 459 22861 493 22895
rect 493 22861 508 22895
rect 456 22850 508 22861
rect 524 22895 576 22902
rect 524 22861 537 22895
rect 537 22861 571 22895
rect 571 22861 576 22895
rect 524 22850 576 22861
rect 592 22895 644 22902
rect 660 22895 712 22902
rect 728 22895 780 22902
rect 796 22895 848 22902
rect 592 22861 615 22895
rect 615 22861 644 22895
rect 660 22861 693 22895
rect 693 22861 712 22895
rect 728 22861 771 22895
rect 771 22861 780 22895
rect 796 22861 805 22895
rect 805 22861 848 22895
rect 592 22850 644 22861
rect 660 22850 712 22861
rect 728 22850 780 22861
rect 796 22850 848 22861
rect 456 22822 508 22838
rect 456 22788 459 22822
rect 459 22788 493 22822
rect 493 22788 508 22822
rect 456 22786 508 22788
rect 524 22822 576 22838
rect 524 22788 537 22822
rect 537 22788 571 22822
rect 571 22788 576 22822
rect 524 22786 576 22788
rect 592 22822 644 22838
rect 660 22822 712 22838
rect 728 22822 780 22838
rect 796 22822 848 22838
rect 592 22788 615 22822
rect 615 22788 644 22822
rect 660 22788 693 22822
rect 693 22788 712 22822
rect 728 22788 771 22822
rect 771 22788 780 22822
rect 796 22788 805 22822
rect 805 22788 848 22822
rect 592 22786 644 22788
rect 660 22786 712 22788
rect 728 22786 780 22788
rect 796 22786 848 22788
rect 456 22749 508 22774
rect 456 22722 459 22749
rect 459 22722 493 22749
rect 493 22722 508 22749
rect 524 22749 576 22774
rect 524 22722 537 22749
rect 537 22722 571 22749
rect 571 22722 576 22749
rect 592 22749 644 22774
rect 660 22749 712 22774
rect 728 22749 780 22774
rect 796 22749 848 22774
rect 592 22722 615 22749
rect 615 22722 644 22749
rect 660 22722 693 22749
rect 693 22722 712 22749
rect 728 22722 771 22749
rect 771 22722 780 22749
rect 796 22722 805 22749
rect 805 22722 848 22749
rect 456 22676 508 22710
rect 456 22658 459 22676
rect 459 22658 493 22676
rect 493 22658 508 22676
rect 524 22676 576 22710
rect 524 22658 537 22676
rect 537 22658 571 22676
rect 571 22658 576 22676
rect 592 22676 644 22710
rect 660 22676 712 22710
rect 728 22676 780 22710
rect 796 22676 848 22710
rect 592 22658 615 22676
rect 615 22658 644 22676
rect 660 22658 693 22676
rect 693 22658 712 22676
rect 728 22658 771 22676
rect 771 22658 780 22676
rect 796 22658 805 22676
rect 805 22658 848 22676
rect 456 22642 459 22646
rect 459 22642 493 22646
rect 493 22642 508 22646
rect 456 22603 508 22642
rect 456 22594 459 22603
rect 459 22594 493 22603
rect 493 22594 508 22603
rect 524 22642 537 22646
rect 537 22642 571 22646
rect 571 22642 576 22646
rect 524 22603 576 22642
rect 524 22594 537 22603
rect 537 22594 571 22603
rect 571 22594 576 22603
rect 592 22642 615 22646
rect 615 22642 644 22646
rect 660 22642 693 22646
rect 693 22642 712 22646
rect 728 22642 771 22646
rect 771 22642 780 22646
rect 796 22642 805 22646
rect 805 22642 848 22646
rect 592 22603 644 22642
rect 660 22603 712 22642
rect 728 22603 780 22642
rect 796 22603 848 22642
rect 592 22594 615 22603
rect 615 22594 644 22603
rect 660 22594 693 22603
rect 693 22594 712 22603
rect 728 22594 771 22603
rect 771 22594 780 22603
rect 796 22594 805 22603
rect 805 22594 848 22603
rect 456 22569 459 22582
rect 459 22569 493 22582
rect 493 22569 508 22582
rect 456 22530 508 22569
rect 524 22569 537 22582
rect 537 22569 571 22582
rect 571 22569 576 22582
rect 524 22530 576 22569
rect 592 22569 615 22582
rect 615 22569 644 22582
rect 660 22569 693 22582
rect 693 22569 712 22582
rect 728 22569 771 22582
rect 771 22569 780 22582
rect 796 22569 805 22582
rect 805 22569 848 22582
rect 592 22530 644 22569
rect 660 22530 712 22569
rect 728 22530 780 22569
rect 796 22530 848 22569
rect 456 22496 459 22518
rect 459 22496 493 22518
rect 493 22496 508 22518
rect 456 22466 508 22496
rect 524 22496 537 22518
rect 537 22496 571 22518
rect 571 22496 576 22518
rect 524 22466 576 22496
rect 592 22496 615 22518
rect 615 22496 644 22518
rect 660 22496 693 22518
rect 693 22496 712 22518
rect 728 22496 771 22518
rect 771 22496 780 22518
rect 796 22496 805 22518
rect 805 22496 848 22518
rect 592 22466 644 22496
rect 660 22466 712 22496
rect 728 22466 780 22496
rect 796 22466 848 22496
rect 456 22423 459 22454
rect 459 22423 493 22454
rect 493 22423 508 22454
rect 456 22402 508 22423
rect 524 22423 537 22454
rect 537 22423 571 22454
rect 571 22423 576 22454
rect 524 22402 576 22423
rect 592 22423 615 22454
rect 615 22423 644 22454
rect 660 22423 693 22454
rect 693 22423 712 22454
rect 728 22423 771 22454
rect 771 22423 780 22454
rect 796 22423 805 22454
rect 805 22423 848 22454
rect 592 22402 644 22423
rect 660 22402 712 22423
rect 728 22402 780 22423
rect 796 22402 848 22423
rect 456 22384 508 22390
rect 456 22350 459 22384
rect 459 22350 493 22384
rect 493 22350 508 22384
rect 456 22338 508 22350
rect 524 22384 576 22390
rect 524 22350 537 22384
rect 537 22350 571 22384
rect 571 22350 576 22384
rect 524 22338 576 22350
rect 592 22384 644 22390
rect 660 22384 712 22390
rect 728 22384 780 22390
rect 796 22384 848 22390
rect 592 22350 615 22384
rect 615 22350 644 22384
rect 660 22350 693 22384
rect 693 22350 712 22384
rect 728 22350 771 22384
rect 771 22350 780 22384
rect 796 22350 805 22384
rect 805 22350 848 22384
rect 592 22338 644 22350
rect 660 22338 712 22350
rect 728 22338 780 22350
rect 796 22338 848 22350
rect 456 22311 508 22326
rect 456 22277 459 22311
rect 459 22277 493 22311
rect 493 22277 508 22311
rect 456 22274 508 22277
rect 524 22311 576 22326
rect 524 22277 537 22311
rect 537 22277 571 22311
rect 571 22277 576 22311
rect 524 22274 576 22277
rect 592 22311 644 22326
rect 660 22311 712 22326
rect 728 22311 780 22326
rect 796 22311 848 22326
rect 592 22277 615 22311
rect 615 22277 644 22311
rect 660 22277 693 22311
rect 693 22277 712 22311
rect 728 22277 771 22311
rect 771 22277 780 22311
rect 796 22277 805 22311
rect 805 22277 848 22311
rect 592 22274 644 22277
rect 660 22274 712 22277
rect 728 22274 780 22277
rect 796 22274 848 22277
rect 456 22238 508 22262
rect 456 22210 459 22238
rect 459 22210 493 22238
rect 493 22210 508 22238
rect 524 22238 576 22262
rect 524 22210 537 22238
rect 537 22210 571 22238
rect 571 22210 576 22238
rect 592 22238 644 22262
rect 660 22238 712 22262
rect 728 22238 780 22262
rect 796 22238 848 22262
rect 592 22210 615 22238
rect 615 22210 644 22238
rect 660 22210 693 22238
rect 693 22210 712 22238
rect 728 22210 771 22238
rect 771 22210 780 22238
rect 796 22210 805 22238
rect 805 22210 848 22238
rect 456 22165 508 22198
rect 456 22146 459 22165
rect 459 22146 493 22165
rect 493 22146 508 22165
rect 524 22165 576 22198
rect 524 22146 537 22165
rect 537 22146 571 22165
rect 571 22146 576 22165
rect 592 22165 644 22198
rect 660 22165 712 22198
rect 728 22165 780 22198
rect 796 22165 848 22198
rect 592 22146 615 22165
rect 615 22146 644 22165
rect 660 22146 693 22165
rect 693 22146 712 22165
rect 728 22146 771 22165
rect 771 22146 780 22165
rect 796 22146 805 22165
rect 805 22146 848 22165
rect 456 22131 459 22134
rect 459 22131 493 22134
rect 493 22131 508 22134
rect 456 22092 508 22131
rect 456 22082 459 22092
rect 459 22082 493 22092
rect 493 22082 508 22092
rect 524 22131 537 22134
rect 537 22131 571 22134
rect 571 22131 576 22134
rect 524 22092 576 22131
rect 524 22082 537 22092
rect 537 22082 571 22092
rect 571 22082 576 22092
rect 592 22131 615 22134
rect 615 22131 644 22134
rect 660 22131 693 22134
rect 693 22131 712 22134
rect 728 22131 771 22134
rect 771 22131 780 22134
rect 796 22131 805 22134
rect 805 22131 848 22134
rect 592 22092 644 22131
rect 660 22092 712 22131
rect 728 22092 780 22131
rect 796 22092 848 22131
rect 592 22082 615 22092
rect 615 22082 644 22092
rect 660 22082 693 22092
rect 693 22082 712 22092
rect 728 22082 771 22092
rect 771 22082 780 22092
rect 796 22082 805 22092
rect 805 22082 848 22092
rect 456 22058 459 22070
rect 459 22058 493 22070
rect 493 22058 508 22070
rect 456 22019 508 22058
rect 456 22018 459 22019
rect 459 22018 493 22019
rect 493 22018 508 22019
rect 524 22058 537 22070
rect 537 22058 571 22070
rect 571 22058 576 22070
rect 524 22019 576 22058
rect 524 22018 537 22019
rect 537 22018 571 22019
rect 571 22018 576 22019
rect 592 22058 615 22070
rect 615 22058 644 22070
rect 660 22058 693 22070
rect 693 22058 712 22070
rect 728 22058 771 22070
rect 771 22058 780 22070
rect 796 22058 805 22070
rect 805 22058 848 22070
rect 592 22019 644 22058
rect 660 22019 712 22058
rect 728 22019 780 22058
rect 796 22019 848 22058
rect 592 22018 615 22019
rect 615 22018 644 22019
rect 660 22018 693 22019
rect 693 22018 712 22019
rect 728 22018 771 22019
rect 771 22018 780 22019
rect 796 22018 805 22019
rect 805 22018 848 22019
rect 456 21985 459 22006
rect 459 21985 493 22006
rect 493 21985 508 22006
rect 456 21954 508 21985
rect 524 21985 537 22006
rect 537 21985 571 22006
rect 571 21985 576 22006
rect 524 21954 576 21985
rect 592 21985 615 22006
rect 615 21985 644 22006
rect 660 21985 693 22006
rect 693 21985 712 22006
rect 728 21985 771 22006
rect 771 21985 780 22006
rect 796 21985 805 22006
rect 805 21985 848 22006
rect 592 21954 644 21985
rect 660 21954 712 21985
rect 728 21954 780 21985
rect 796 21954 848 21985
rect 456 21912 459 21942
rect 459 21912 493 21942
rect 493 21912 508 21942
rect 456 21890 508 21912
rect 524 21912 537 21942
rect 537 21912 571 21942
rect 571 21912 576 21942
rect 524 21890 576 21912
rect 592 21912 615 21942
rect 615 21912 644 21942
rect 660 21912 693 21942
rect 693 21912 712 21942
rect 728 21912 771 21942
rect 771 21912 780 21942
rect 796 21912 805 21942
rect 805 21912 848 21942
rect 592 21890 644 21912
rect 660 21890 712 21912
rect 728 21890 780 21912
rect 796 21890 848 21912
rect 456 21873 508 21878
rect 456 21839 459 21873
rect 459 21839 493 21873
rect 493 21839 508 21873
rect 456 21826 508 21839
rect 524 21873 576 21878
rect 524 21839 537 21873
rect 537 21839 571 21873
rect 571 21839 576 21873
rect 524 21826 576 21839
rect 592 21873 644 21878
rect 660 21873 712 21878
rect 728 21873 780 21878
rect 796 21873 848 21878
rect 592 21839 615 21873
rect 615 21839 644 21873
rect 660 21839 693 21873
rect 693 21839 712 21873
rect 728 21839 771 21873
rect 771 21839 780 21873
rect 796 21839 805 21873
rect 805 21839 848 21873
rect 592 21826 644 21839
rect 660 21826 712 21839
rect 728 21826 780 21839
rect 796 21826 848 21839
rect 456 21800 508 21814
rect 456 21766 459 21800
rect 459 21766 493 21800
rect 493 21766 508 21800
rect 456 21762 508 21766
rect 524 21800 576 21814
rect 524 21766 537 21800
rect 537 21766 571 21800
rect 571 21766 576 21800
rect 524 21762 576 21766
rect 592 21800 644 21814
rect 660 21800 712 21814
rect 728 21800 780 21814
rect 796 21800 848 21814
rect 592 21766 615 21800
rect 615 21766 644 21800
rect 660 21766 693 21800
rect 693 21766 712 21800
rect 728 21766 771 21800
rect 771 21766 780 21800
rect 796 21766 805 21800
rect 805 21766 848 21800
rect 592 21762 644 21766
rect 660 21762 712 21766
rect 728 21762 780 21766
rect 796 21762 848 21766
rect 456 21727 508 21750
rect 456 21698 459 21727
rect 459 21698 493 21727
rect 493 21698 508 21727
rect 524 21727 576 21750
rect 524 21698 537 21727
rect 537 21698 571 21727
rect 571 21698 576 21727
rect 592 21727 644 21750
rect 660 21727 712 21750
rect 728 21727 780 21750
rect 796 21727 848 21750
rect 592 21698 615 21727
rect 615 21698 644 21727
rect 660 21698 693 21727
rect 693 21698 712 21727
rect 728 21698 771 21727
rect 771 21698 780 21727
rect 796 21698 805 21727
rect 805 21698 848 21727
rect 456 21654 508 21686
rect 456 21634 459 21654
rect 459 21634 493 21654
rect 493 21634 508 21654
rect 524 21654 576 21686
rect 524 21634 537 21654
rect 537 21634 571 21654
rect 571 21634 576 21654
rect 592 21654 644 21686
rect 660 21654 712 21686
rect 728 21654 780 21686
rect 796 21654 848 21686
rect 592 21634 615 21654
rect 615 21634 644 21654
rect 660 21634 693 21654
rect 693 21634 712 21654
rect 728 21634 771 21654
rect 771 21634 780 21654
rect 796 21634 805 21654
rect 805 21634 848 21654
rect 456 21620 459 21622
rect 459 21620 493 21622
rect 493 21620 508 21622
rect 456 21581 508 21620
rect 456 21570 459 21581
rect 459 21570 493 21581
rect 493 21570 508 21581
rect 524 21620 537 21622
rect 537 21620 571 21622
rect 571 21620 576 21622
rect 524 21581 576 21620
rect 524 21570 537 21581
rect 537 21570 571 21581
rect 571 21570 576 21581
rect 592 21620 615 21622
rect 615 21620 644 21622
rect 660 21620 693 21622
rect 693 21620 712 21622
rect 728 21620 771 21622
rect 771 21620 780 21622
rect 796 21620 805 21622
rect 805 21620 848 21622
rect 592 21581 644 21620
rect 660 21581 712 21620
rect 728 21581 780 21620
rect 796 21581 848 21620
rect 592 21570 615 21581
rect 615 21570 644 21581
rect 660 21570 693 21581
rect 693 21570 712 21581
rect 728 21570 771 21581
rect 771 21570 780 21581
rect 796 21570 805 21581
rect 805 21570 848 21581
rect 456 21547 459 21558
rect 459 21547 493 21558
rect 493 21547 508 21558
rect 456 21508 508 21547
rect 456 21506 459 21508
rect 459 21506 493 21508
rect 493 21506 508 21508
rect 524 21547 537 21558
rect 537 21547 571 21558
rect 571 21547 576 21558
rect 524 21508 576 21547
rect 524 21506 537 21508
rect 537 21506 571 21508
rect 571 21506 576 21508
rect 592 21547 615 21558
rect 615 21547 644 21558
rect 660 21547 693 21558
rect 693 21547 712 21558
rect 728 21547 771 21558
rect 771 21547 780 21558
rect 796 21547 805 21558
rect 805 21547 848 21558
rect 592 21508 644 21547
rect 660 21508 712 21547
rect 728 21508 780 21547
rect 796 21508 848 21547
rect 592 21506 615 21508
rect 615 21506 644 21508
rect 660 21506 693 21508
rect 693 21506 712 21508
rect 728 21506 771 21508
rect 771 21506 780 21508
rect 796 21506 805 21508
rect 805 21506 848 21508
rect 456 21474 459 21494
rect 459 21474 493 21494
rect 493 21474 508 21494
rect 456 21442 508 21474
rect 524 21474 537 21494
rect 537 21474 571 21494
rect 571 21474 576 21494
rect 524 21442 576 21474
rect 592 21474 615 21494
rect 615 21474 644 21494
rect 660 21474 693 21494
rect 693 21474 712 21494
rect 728 21474 771 21494
rect 771 21474 780 21494
rect 796 21474 805 21494
rect 805 21474 848 21494
rect 592 21442 644 21474
rect 660 21442 712 21474
rect 728 21442 780 21474
rect 796 21442 848 21474
rect 456 21401 459 21430
rect 459 21401 493 21430
rect 493 21401 508 21430
rect 456 21378 508 21401
rect 524 21401 537 21430
rect 537 21401 571 21430
rect 571 21401 576 21430
rect 524 21378 576 21401
rect 592 21401 615 21430
rect 615 21401 644 21430
rect 660 21401 693 21430
rect 693 21401 712 21430
rect 728 21401 771 21430
rect 771 21401 780 21430
rect 796 21401 805 21430
rect 805 21401 848 21430
rect 592 21378 644 21401
rect 660 21378 712 21401
rect 728 21378 780 21401
rect 796 21378 848 21401
rect 456 21362 508 21366
rect 456 21328 459 21362
rect 459 21328 493 21362
rect 493 21328 508 21362
rect 456 21314 508 21328
rect 524 21362 576 21366
rect 524 21328 537 21362
rect 537 21328 571 21362
rect 571 21328 576 21362
rect 524 21314 576 21328
rect 592 21362 644 21366
rect 660 21362 712 21366
rect 728 21362 780 21366
rect 796 21362 848 21366
rect 592 21328 615 21362
rect 615 21328 644 21362
rect 660 21328 693 21362
rect 693 21328 712 21362
rect 728 21328 771 21362
rect 771 21328 780 21362
rect 796 21328 805 21362
rect 805 21328 848 21362
rect 592 21314 644 21328
rect 660 21314 712 21328
rect 728 21314 780 21328
rect 796 21314 848 21328
rect 456 21289 508 21302
rect 456 21255 459 21289
rect 459 21255 493 21289
rect 493 21255 508 21289
rect 456 21250 508 21255
rect 524 21289 576 21302
rect 524 21255 537 21289
rect 537 21255 571 21289
rect 571 21255 576 21289
rect 524 21250 576 21255
rect 592 21289 644 21302
rect 660 21289 712 21302
rect 728 21289 780 21302
rect 796 21289 848 21302
rect 592 21255 615 21289
rect 615 21255 644 21289
rect 660 21255 693 21289
rect 693 21255 712 21289
rect 728 21255 771 21289
rect 771 21255 780 21289
rect 796 21255 805 21289
rect 805 21255 848 21289
rect 592 21250 644 21255
rect 660 21250 712 21255
rect 728 21250 780 21255
rect 796 21250 848 21255
rect 456 21216 508 21238
rect 456 21186 459 21216
rect 459 21186 493 21216
rect 493 21186 508 21216
rect 524 21216 576 21238
rect 524 21186 537 21216
rect 537 21186 571 21216
rect 571 21186 576 21216
rect 592 21216 644 21238
rect 660 21216 712 21238
rect 728 21216 780 21238
rect 796 21216 848 21238
rect 592 21186 615 21216
rect 615 21186 644 21216
rect 660 21186 693 21216
rect 693 21186 712 21216
rect 728 21186 771 21216
rect 771 21186 780 21216
rect 796 21186 805 21216
rect 805 21186 848 21216
rect 456 21143 508 21174
rect 456 21122 459 21143
rect 459 21122 493 21143
rect 493 21122 508 21143
rect 524 21143 576 21174
rect 524 21122 537 21143
rect 537 21122 571 21143
rect 571 21122 576 21143
rect 592 21143 644 21174
rect 660 21143 712 21174
rect 728 21143 780 21174
rect 796 21143 848 21174
rect 592 21122 615 21143
rect 615 21122 644 21143
rect 660 21122 693 21143
rect 693 21122 712 21143
rect 728 21122 771 21143
rect 771 21122 780 21143
rect 796 21122 805 21143
rect 805 21122 848 21143
rect 456 21109 459 21110
rect 459 21109 493 21110
rect 493 21109 508 21110
rect 456 21070 508 21109
rect 456 21058 459 21070
rect 459 21058 493 21070
rect 493 21058 508 21070
rect 524 21109 537 21110
rect 537 21109 571 21110
rect 571 21109 576 21110
rect 524 21070 576 21109
rect 524 21058 537 21070
rect 537 21058 571 21070
rect 571 21058 576 21070
rect 592 21109 615 21110
rect 615 21109 644 21110
rect 660 21109 693 21110
rect 693 21109 712 21110
rect 728 21109 771 21110
rect 771 21109 780 21110
rect 796 21109 805 21110
rect 805 21109 848 21110
rect 592 21070 644 21109
rect 660 21070 712 21109
rect 728 21070 780 21109
rect 796 21070 848 21109
rect 592 21058 615 21070
rect 615 21058 644 21070
rect 660 21058 693 21070
rect 693 21058 712 21070
rect 728 21058 771 21070
rect 771 21058 780 21070
rect 796 21058 805 21070
rect 805 21058 848 21070
rect 456 21036 459 21046
rect 459 21036 493 21046
rect 493 21036 508 21046
rect 456 20997 508 21036
rect 456 20994 459 20997
rect 459 20994 493 20997
rect 493 20994 508 20997
rect 524 21036 537 21046
rect 537 21036 571 21046
rect 571 21036 576 21046
rect 524 20997 576 21036
rect 524 20994 537 20997
rect 537 20994 571 20997
rect 571 20994 576 20997
rect 592 21036 615 21046
rect 615 21036 644 21046
rect 660 21036 693 21046
rect 693 21036 712 21046
rect 728 21036 771 21046
rect 771 21036 780 21046
rect 796 21036 805 21046
rect 805 21036 848 21046
rect 592 20997 644 21036
rect 660 20997 712 21036
rect 728 20997 780 21036
rect 796 20997 848 21036
rect 592 20994 615 20997
rect 615 20994 644 20997
rect 660 20994 693 20997
rect 693 20994 712 20997
rect 728 20994 771 20997
rect 771 20994 780 20997
rect 796 20994 805 20997
rect 805 20994 848 20997
rect 456 20963 459 20982
rect 459 20963 493 20982
rect 493 20963 508 20982
rect 456 20930 508 20963
rect 524 20963 537 20982
rect 537 20963 571 20982
rect 571 20963 576 20982
rect 524 20930 576 20963
rect 592 20963 615 20982
rect 615 20963 644 20982
rect 660 20963 693 20982
rect 693 20963 712 20982
rect 728 20963 771 20982
rect 771 20963 780 20982
rect 796 20963 805 20982
rect 805 20963 848 20982
rect 592 20930 644 20963
rect 660 20930 712 20963
rect 728 20930 780 20963
rect 796 20930 848 20963
rect 456 20890 459 20918
rect 459 20890 493 20918
rect 493 20890 508 20918
rect 456 20866 508 20890
rect 524 20890 537 20918
rect 537 20890 571 20918
rect 571 20890 576 20918
rect 524 20866 576 20890
rect 592 20890 615 20918
rect 615 20890 644 20918
rect 660 20890 693 20918
rect 693 20890 712 20918
rect 728 20890 771 20918
rect 771 20890 780 20918
rect 796 20890 805 20918
rect 805 20890 848 20918
rect 592 20866 644 20890
rect 660 20866 712 20890
rect 728 20866 780 20890
rect 796 20866 848 20890
rect 456 20851 508 20854
rect 456 20817 459 20851
rect 459 20817 493 20851
rect 493 20817 508 20851
rect 456 20802 508 20817
rect 524 20851 576 20854
rect 524 20817 537 20851
rect 537 20817 571 20851
rect 571 20817 576 20851
rect 524 20802 576 20817
rect 592 20851 644 20854
rect 660 20851 712 20854
rect 728 20851 780 20854
rect 796 20851 848 20854
rect 592 20817 615 20851
rect 615 20817 644 20851
rect 660 20817 693 20851
rect 693 20817 712 20851
rect 728 20817 771 20851
rect 771 20817 780 20851
rect 796 20817 805 20851
rect 805 20817 848 20851
rect 592 20802 644 20817
rect 660 20802 712 20817
rect 728 20802 780 20817
rect 796 20802 848 20817
rect 456 20778 508 20790
rect 456 20744 459 20778
rect 459 20744 493 20778
rect 493 20744 508 20778
rect 456 20738 508 20744
rect 524 20778 576 20790
rect 524 20744 537 20778
rect 537 20744 571 20778
rect 571 20744 576 20778
rect 524 20738 576 20744
rect 592 20778 644 20790
rect 660 20778 712 20790
rect 728 20778 780 20790
rect 796 20778 848 20790
rect 592 20744 615 20778
rect 615 20744 644 20778
rect 660 20744 693 20778
rect 693 20744 712 20778
rect 728 20744 771 20778
rect 771 20744 780 20778
rect 796 20744 805 20778
rect 805 20744 848 20778
rect 592 20738 644 20744
rect 660 20738 712 20744
rect 728 20738 780 20744
rect 796 20738 848 20744
rect 456 20705 508 20726
rect 456 20674 459 20705
rect 459 20674 493 20705
rect 493 20674 508 20705
rect 524 20705 576 20726
rect 524 20674 537 20705
rect 537 20674 571 20705
rect 571 20674 576 20705
rect 592 20705 644 20726
rect 660 20705 712 20726
rect 728 20705 780 20726
rect 796 20705 848 20726
rect 592 20674 615 20705
rect 615 20674 644 20705
rect 660 20674 693 20705
rect 693 20674 712 20705
rect 728 20674 771 20705
rect 771 20674 780 20705
rect 796 20674 805 20705
rect 805 20674 848 20705
rect 456 20632 508 20662
rect 456 20610 459 20632
rect 459 20610 493 20632
rect 493 20610 508 20632
rect 524 20632 576 20662
rect 524 20610 537 20632
rect 537 20610 571 20632
rect 571 20610 576 20632
rect 592 20632 644 20662
rect 660 20632 712 20662
rect 728 20632 780 20662
rect 796 20632 848 20662
rect 592 20610 615 20632
rect 615 20610 644 20632
rect 660 20610 693 20632
rect 693 20610 712 20632
rect 728 20610 771 20632
rect 771 20610 780 20632
rect 796 20610 805 20632
rect 805 20610 848 20632
rect 456 20559 508 20598
rect 456 20546 459 20559
rect 459 20546 493 20559
rect 493 20546 508 20559
rect 524 20559 576 20598
rect 524 20546 537 20559
rect 537 20546 571 20559
rect 571 20546 576 20559
rect 592 20559 644 20598
rect 660 20559 712 20598
rect 728 20559 780 20598
rect 796 20559 848 20598
rect 592 20546 615 20559
rect 615 20546 644 20559
rect 660 20546 693 20559
rect 693 20546 712 20559
rect 728 20546 771 20559
rect 771 20546 780 20559
rect 796 20546 805 20559
rect 805 20546 848 20559
rect 456 20525 459 20534
rect 459 20525 493 20534
rect 493 20525 508 20534
rect 456 20486 508 20525
rect 456 20482 459 20486
rect 459 20482 493 20486
rect 493 20482 508 20486
rect 524 20525 537 20534
rect 537 20525 571 20534
rect 571 20525 576 20534
rect 524 20486 576 20525
rect 524 20482 537 20486
rect 537 20482 571 20486
rect 571 20482 576 20486
rect 592 20525 615 20534
rect 615 20525 644 20534
rect 660 20525 693 20534
rect 693 20525 712 20534
rect 728 20525 771 20534
rect 771 20525 780 20534
rect 796 20525 805 20534
rect 805 20525 848 20534
rect 592 20486 644 20525
rect 660 20486 712 20525
rect 728 20486 780 20525
rect 796 20486 848 20525
rect 592 20482 615 20486
rect 615 20482 644 20486
rect 660 20482 693 20486
rect 693 20482 712 20486
rect 728 20482 771 20486
rect 771 20482 780 20486
rect 796 20482 805 20486
rect 805 20482 848 20486
rect 456 20452 459 20470
rect 459 20452 493 20470
rect 493 20452 508 20470
rect 456 20418 508 20452
rect 524 20452 537 20470
rect 537 20452 571 20470
rect 571 20452 576 20470
rect 524 20418 576 20452
rect 592 20452 615 20470
rect 615 20452 644 20470
rect 660 20452 693 20470
rect 693 20452 712 20470
rect 728 20452 771 20470
rect 771 20452 780 20470
rect 796 20452 805 20470
rect 805 20452 848 20470
rect 592 20418 644 20452
rect 660 20418 712 20452
rect 728 20418 780 20452
rect 796 20418 848 20452
rect 456 20379 459 20406
rect 459 20379 493 20406
rect 493 20379 508 20406
rect 456 20354 508 20379
rect 524 20379 537 20406
rect 537 20379 571 20406
rect 571 20379 576 20406
rect 524 20354 576 20379
rect 592 20379 615 20406
rect 615 20379 644 20406
rect 660 20379 693 20406
rect 693 20379 712 20406
rect 728 20379 771 20406
rect 771 20379 780 20406
rect 796 20379 805 20406
rect 805 20379 848 20406
rect 2784 20519 2836 20571
rect 2853 20519 2905 20571
rect 2922 20519 2974 20571
rect 2991 20519 3043 20571
rect 3060 20519 3112 20571
rect 3128 20519 3180 20571
rect 3196 20519 3248 20571
rect 3264 20519 3316 20571
rect 3332 20519 3384 20571
rect 3400 20519 3452 20571
rect 3468 20519 3520 20571
rect 3536 20519 3588 20571
rect 3604 20519 3656 20571
rect 3672 20519 3724 20571
rect 2784 20407 2836 20459
rect 2853 20407 2905 20459
rect 2922 20407 2974 20459
rect 2991 20407 3043 20459
rect 3060 20407 3112 20459
rect 3128 20407 3180 20459
rect 3196 20407 3248 20459
rect 3264 20407 3316 20459
rect 3332 20407 3384 20459
rect 3400 20407 3452 20459
rect 3468 20407 3520 20459
rect 3536 20407 3588 20459
rect 3604 20407 3656 20459
rect 3672 20407 3724 20459
rect 12199 20514 12251 20566
rect 12199 20444 12251 20496
rect 592 20354 644 20379
rect 660 20354 712 20379
rect 728 20354 780 20379
rect 796 20354 848 20379
rect 456 20340 508 20342
rect 456 20306 459 20340
rect 459 20306 493 20340
rect 493 20306 508 20340
rect 456 20290 508 20306
rect 524 20340 576 20342
rect 524 20306 537 20340
rect 537 20306 571 20340
rect 571 20306 576 20340
rect 524 20290 576 20306
rect 592 20340 644 20342
rect 660 20340 712 20342
rect 728 20340 780 20342
rect 796 20340 848 20342
rect 592 20306 615 20340
rect 615 20306 644 20340
rect 660 20306 693 20340
rect 693 20306 712 20340
rect 728 20306 771 20340
rect 771 20306 780 20340
rect 796 20306 805 20340
rect 805 20306 848 20340
rect 592 20290 644 20306
rect 660 20290 712 20306
rect 728 20290 780 20306
rect 796 20290 848 20306
rect 456 20267 508 20277
rect 456 20233 459 20267
rect 459 20233 493 20267
rect 493 20233 508 20267
rect 456 20225 508 20233
rect 524 20267 576 20277
rect 524 20233 537 20267
rect 537 20233 571 20267
rect 571 20233 576 20267
rect 524 20225 576 20233
rect 592 20267 644 20277
rect 660 20267 712 20277
rect 728 20267 780 20277
rect 796 20267 848 20277
rect 592 20233 615 20267
rect 615 20233 644 20267
rect 660 20233 693 20267
rect 693 20233 712 20267
rect 728 20233 771 20267
rect 771 20233 780 20267
rect 796 20233 805 20267
rect 805 20233 848 20267
rect 592 20225 644 20233
rect 660 20225 712 20233
rect 728 20225 780 20233
rect 796 20225 848 20233
rect 12199 20373 12251 20425
rect 12199 20302 12251 20354
rect 12199 20231 12251 20283
rect 456 20194 508 20212
rect 456 20160 459 20194
rect 459 20160 493 20194
rect 493 20160 508 20194
rect 524 20194 576 20212
rect 524 20160 537 20194
rect 537 20160 571 20194
rect 571 20160 576 20194
rect 592 20194 644 20212
rect 660 20194 712 20212
rect 728 20194 780 20212
rect 796 20194 848 20212
rect 592 20160 615 20194
rect 615 20160 644 20194
rect 660 20160 693 20194
rect 693 20160 712 20194
rect 728 20160 771 20194
rect 771 20160 780 20194
rect 796 20160 805 20194
rect 805 20160 848 20194
rect 456 20121 508 20147
rect 456 20095 459 20121
rect 459 20095 493 20121
rect 493 20095 508 20121
rect 524 20121 576 20147
rect 524 20095 537 20121
rect 537 20095 571 20121
rect 571 20095 576 20121
rect 592 20121 644 20147
rect 660 20121 712 20147
rect 728 20121 780 20147
rect 796 20121 848 20147
rect 592 20095 615 20121
rect 615 20095 644 20121
rect 660 20095 693 20121
rect 693 20095 712 20121
rect 728 20095 771 20121
rect 771 20095 780 20121
rect 796 20095 805 20121
rect 805 20095 848 20121
rect 456 20048 508 20082
rect 456 20030 459 20048
rect 459 20030 493 20048
rect 493 20030 508 20048
rect 524 20048 576 20082
rect 524 20030 537 20048
rect 537 20030 571 20048
rect 571 20030 576 20048
rect 592 20048 644 20082
rect 660 20048 712 20082
rect 728 20048 780 20082
rect 796 20048 848 20082
rect 592 20030 615 20048
rect 615 20030 644 20048
rect 660 20030 693 20048
rect 693 20030 712 20048
rect 728 20030 771 20048
rect 771 20030 780 20048
rect 796 20030 805 20048
rect 805 20030 848 20048
rect 456 20014 459 20017
rect 459 20014 493 20017
rect 493 20014 508 20017
rect 456 19975 508 20014
rect 456 19965 459 19975
rect 459 19965 493 19975
rect 493 19965 508 19975
rect 524 20014 537 20017
rect 537 20014 571 20017
rect 571 20014 576 20017
rect 524 19975 576 20014
rect 524 19965 537 19975
rect 537 19965 571 19975
rect 571 19965 576 19975
rect 592 20014 615 20017
rect 615 20014 644 20017
rect 660 20014 693 20017
rect 693 20014 712 20017
rect 728 20014 771 20017
rect 771 20014 780 20017
rect 796 20014 805 20017
rect 805 20014 848 20017
rect 592 19975 644 20014
rect 660 19975 712 20014
rect 728 19975 780 20014
rect 796 19975 848 20014
rect 592 19965 615 19975
rect 615 19965 644 19975
rect 660 19965 693 19975
rect 693 19965 712 19975
rect 728 19965 771 19975
rect 771 19965 780 19975
rect 796 19965 805 19975
rect 805 19965 848 19975
rect 456 19941 459 19952
rect 459 19941 493 19952
rect 493 19941 508 19952
rect 456 19902 508 19941
rect 456 19900 459 19902
rect 459 19900 493 19902
rect 493 19900 508 19902
rect 524 19941 537 19952
rect 537 19941 571 19952
rect 571 19941 576 19952
rect 524 19902 576 19941
rect 524 19900 537 19902
rect 537 19900 571 19902
rect 571 19900 576 19902
rect 592 19941 615 19952
rect 615 19941 644 19952
rect 660 19941 693 19952
rect 693 19941 712 19952
rect 728 19941 771 19952
rect 771 19941 780 19952
rect 796 19941 805 19952
rect 805 19941 848 19952
rect 592 19902 644 19941
rect 660 19902 712 19941
rect 728 19902 780 19941
rect 796 19902 848 19941
rect 592 19900 615 19902
rect 615 19900 644 19902
rect 660 19900 693 19902
rect 693 19900 712 19902
rect 728 19900 771 19902
rect 771 19900 780 19902
rect 796 19900 805 19902
rect 805 19900 848 19902
rect 456 19868 459 19887
rect 459 19868 493 19887
rect 493 19868 508 19887
rect 456 19835 508 19868
rect 524 19868 537 19887
rect 537 19868 571 19887
rect 571 19868 576 19887
rect 524 19835 576 19868
rect 592 19868 615 19887
rect 615 19868 644 19887
rect 660 19868 693 19887
rect 693 19868 712 19887
rect 728 19868 771 19887
rect 771 19868 780 19887
rect 796 19868 805 19887
rect 805 19868 848 19887
rect 592 19835 644 19868
rect 660 19835 712 19868
rect 728 19835 780 19868
rect 796 19835 848 19868
rect 456 19795 459 19822
rect 459 19795 493 19822
rect 493 19795 508 19822
rect 456 19770 508 19795
rect 524 19795 537 19822
rect 537 19795 571 19822
rect 571 19795 576 19822
rect 524 19770 576 19795
rect 592 19795 615 19822
rect 615 19795 644 19822
rect 660 19795 693 19822
rect 693 19795 712 19822
rect 728 19795 771 19822
rect 771 19795 780 19822
rect 796 19795 805 19822
rect 805 19795 848 19822
rect 592 19770 644 19795
rect 660 19770 712 19795
rect 728 19770 780 19795
rect 796 19770 848 19795
rect 456 19756 508 19757
rect 456 19722 459 19756
rect 459 19722 493 19756
rect 493 19722 508 19756
rect 456 19705 508 19722
rect 524 19756 576 19757
rect 524 19722 537 19756
rect 537 19722 571 19756
rect 571 19722 576 19756
rect 524 19705 576 19722
rect 592 19756 644 19757
rect 660 19756 712 19757
rect 728 19756 780 19757
rect 796 19756 848 19757
rect 592 19722 615 19756
rect 615 19722 644 19756
rect 660 19722 693 19756
rect 693 19722 712 19756
rect 728 19722 771 19756
rect 771 19722 780 19756
rect 796 19722 805 19756
rect 805 19722 848 19756
rect 592 19705 644 19722
rect 660 19705 712 19722
rect 728 19705 780 19722
rect 796 19705 848 19722
rect 456 19683 508 19692
rect 456 19649 459 19683
rect 459 19649 493 19683
rect 493 19649 508 19683
rect 456 19640 508 19649
rect 524 19683 576 19692
rect 524 19649 537 19683
rect 537 19649 571 19683
rect 571 19649 576 19683
rect 524 19640 576 19649
rect 592 19683 644 19692
rect 660 19683 712 19692
rect 728 19683 780 19692
rect 796 19683 848 19692
rect 592 19649 615 19683
rect 615 19649 644 19683
rect 660 19649 693 19683
rect 693 19649 712 19683
rect 728 19649 771 19683
rect 771 19649 780 19683
rect 796 19649 805 19683
rect 805 19649 848 19683
rect 12199 20058 12251 20110
rect 12199 19994 12251 20046
rect 12199 19930 12251 19982
rect 12199 19866 12251 19918
rect 12199 19802 12251 19854
rect 12199 19738 12251 19790
rect 12199 19673 12251 19725
rect 592 19640 644 19649
rect 660 19640 712 19649
rect 728 19640 780 19649
rect 796 19640 848 19649
rect 456 19610 508 19627
rect 456 19576 459 19610
rect 459 19576 493 19610
rect 493 19576 508 19610
rect 456 19575 508 19576
rect 524 19610 576 19627
rect 524 19576 537 19610
rect 537 19576 571 19610
rect 571 19576 576 19610
rect 524 19575 576 19576
rect 592 19610 644 19627
rect 660 19610 712 19627
rect 728 19610 780 19627
rect 796 19610 848 19627
rect 592 19576 615 19610
rect 615 19576 644 19610
rect 660 19576 693 19610
rect 693 19576 712 19610
rect 728 19576 771 19610
rect 771 19576 780 19610
rect 796 19576 805 19610
rect 805 19576 848 19610
rect 592 19575 644 19576
rect 660 19575 712 19576
rect 728 19575 780 19576
rect 796 19575 848 19576
rect 456 19537 508 19562
rect 456 19510 459 19537
rect 459 19510 493 19537
rect 493 19510 508 19537
rect 524 19537 576 19562
rect 524 19510 537 19537
rect 537 19510 571 19537
rect 571 19510 576 19537
rect 592 19537 644 19562
rect 660 19537 712 19562
rect 728 19537 780 19562
rect 796 19537 848 19562
rect 592 19510 615 19537
rect 615 19510 644 19537
rect 660 19510 693 19537
rect 693 19510 712 19537
rect 728 19510 771 19537
rect 771 19510 780 19537
rect 796 19510 805 19537
rect 805 19510 848 19537
rect 456 19464 508 19497
rect 456 19445 459 19464
rect 459 19445 493 19464
rect 493 19445 508 19464
rect 524 19464 576 19497
rect 524 19445 537 19464
rect 537 19445 571 19464
rect 571 19445 576 19464
rect 592 19464 644 19497
rect 660 19464 712 19497
rect 728 19464 780 19497
rect 796 19464 848 19497
rect 592 19445 615 19464
rect 615 19445 644 19464
rect 660 19445 693 19464
rect 693 19445 712 19464
rect 728 19445 771 19464
rect 771 19445 780 19464
rect 796 19445 805 19464
rect 805 19445 848 19464
rect 456 19430 459 19432
rect 459 19430 493 19432
rect 493 19430 508 19432
rect 456 19391 508 19430
rect 456 19380 459 19391
rect 459 19380 493 19391
rect 493 19380 508 19391
rect 524 19430 537 19432
rect 537 19430 571 19432
rect 571 19430 576 19432
rect 524 19391 576 19430
rect 524 19380 537 19391
rect 537 19380 571 19391
rect 571 19380 576 19391
rect 592 19430 615 19432
rect 615 19430 644 19432
rect 660 19430 693 19432
rect 693 19430 712 19432
rect 728 19430 771 19432
rect 771 19430 780 19432
rect 796 19430 805 19432
rect 805 19430 848 19432
rect 592 19391 644 19430
rect 660 19391 712 19430
rect 728 19391 780 19430
rect 796 19391 848 19430
rect 592 19380 615 19391
rect 615 19380 644 19391
rect 660 19380 693 19391
rect 693 19380 712 19391
rect 728 19380 771 19391
rect 771 19380 780 19391
rect 796 19380 805 19391
rect 805 19380 848 19391
rect 456 19357 459 19367
rect 459 19357 493 19367
rect 493 19357 508 19367
rect 456 19318 508 19357
rect 456 19315 459 19318
rect 459 19315 493 19318
rect 493 19315 508 19318
rect 524 19357 537 19367
rect 537 19357 571 19367
rect 571 19357 576 19367
rect 524 19318 576 19357
rect 524 19315 537 19318
rect 537 19315 571 19318
rect 571 19315 576 19318
rect 592 19357 615 19367
rect 615 19357 644 19367
rect 660 19357 693 19367
rect 693 19357 712 19367
rect 728 19357 771 19367
rect 771 19357 780 19367
rect 796 19357 805 19367
rect 805 19357 848 19367
rect 592 19318 644 19357
rect 660 19318 712 19357
rect 728 19318 780 19357
rect 796 19318 848 19357
rect 592 19315 615 19318
rect 615 19315 644 19318
rect 660 19315 693 19318
rect 693 19315 712 19318
rect 728 19315 771 19318
rect 771 19315 780 19318
rect 796 19315 805 19318
rect 805 19315 848 19318
rect 456 19284 459 19302
rect 459 19284 493 19302
rect 493 19284 508 19302
rect 456 19250 508 19284
rect 524 19284 537 19302
rect 537 19284 571 19302
rect 571 19284 576 19302
rect 524 19250 576 19284
rect 592 19284 615 19302
rect 615 19284 644 19302
rect 660 19284 693 19302
rect 693 19284 712 19302
rect 728 19284 771 19302
rect 771 19284 780 19302
rect 796 19284 805 19302
rect 805 19284 848 19302
rect 592 19250 644 19284
rect 660 19250 712 19284
rect 728 19250 780 19284
rect 796 19250 848 19284
rect 456 19211 459 19237
rect 459 19211 493 19237
rect 493 19211 508 19237
rect 456 19185 508 19211
rect 524 19211 537 19237
rect 537 19211 571 19237
rect 571 19211 576 19237
rect 524 19185 576 19211
rect 592 19211 615 19237
rect 615 19211 644 19237
rect 660 19211 693 19237
rect 693 19211 712 19237
rect 728 19211 771 19237
rect 771 19211 780 19237
rect 796 19211 805 19237
rect 805 19211 848 19237
rect 592 19185 644 19211
rect 660 19185 712 19211
rect 728 19185 780 19211
rect 796 19185 848 19211
rect 2787 19191 2839 19243
rect 2854 19191 2906 19243
rect 2921 19191 2973 19243
rect 2988 19191 3040 19243
rect 3055 19191 3107 19243
rect 3122 19191 3174 19243
rect 3189 19191 3241 19243
rect 3256 19191 3308 19243
rect 3323 19191 3375 19243
rect 3390 19191 3442 19243
rect 3456 19191 3508 19243
rect 3522 19191 3574 19243
rect 3588 19191 3640 19243
rect 3654 19191 3706 19243
rect 3720 19191 3772 19243
rect 3022 19017 3074 19069
rect 3092 19017 3144 19069
rect 3162 19017 3214 19069
rect 3232 19017 3284 19069
rect 3302 19017 3354 19069
rect 3372 19017 3424 19069
rect 3442 19017 3494 19069
rect 3512 19017 3564 19069
rect 3582 19017 3634 19069
rect 3651 19017 3703 19069
rect 3720 19017 3772 19069
rect 276 18824 328 18876
rect 341 18824 393 18876
rect 406 18824 458 18876
rect 471 18824 523 18876
rect 536 18824 588 18876
rect 601 18824 653 18876
rect 666 18824 718 18876
rect 1257 18824 1309 18876
rect 1325 18824 1377 18876
rect 1393 18824 1445 18876
rect 1461 18824 1513 18876
rect 1528 18824 1580 18876
rect 1595 18824 1647 18876
rect 276 18742 328 18794
rect 341 18742 393 18794
rect 406 18742 458 18794
rect 471 18742 523 18794
rect 536 18742 588 18794
rect 601 18742 653 18794
rect 666 18742 718 18794
rect 1257 18742 1309 18794
rect 1325 18742 1377 18794
rect 1393 18742 1445 18794
rect 1461 18742 1513 18794
rect 1528 18742 1580 18794
rect 1595 18742 1647 18794
rect 276 18660 328 18712
rect 341 18660 393 18712
rect 406 18660 458 18712
rect 471 18660 523 18712
rect 536 18660 588 18712
rect 601 18660 653 18712
rect 666 18660 718 18712
rect 1257 18660 1309 18712
rect 1325 18660 1377 18712
rect 1393 18660 1445 18712
rect 1461 18660 1513 18712
rect 1528 18660 1580 18712
rect 1595 18660 1647 18712
rect 3204 17297 3256 17349
rect 3296 17297 3348 17349
rect 5737 16725 5789 16777
rect 5802 16725 5854 16777
rect 5867 16725 5919 16777
rect 5932 16725 5984 16777
rect 5997 16725 6049 16777
rect 6062 16725 6114 16777
rect 6127 16725 6179 16777
rect 6192 16725 6244 16777
rect 6257 16725 6309 16777
rect 6322 16725 6374 16777
rect 6387 16725 6439 16777
rect 6452 16725 6504 16777
rect 6517 16725 6569 16777
rect 6582 16725 6634 16777
rect 6647 16725 6699 16777
rect 6712 16725 6764 16777
rect 6777 16725 6829 16777
rect 6842 16725 6894 16777
rect 6907 16725 6959 16777
rect 6972 16725 7024 16777
rect 7036 16725 7088 16777
rect 7100 16725 7152 16777
rect 7164 16725 7216 16777
rect 7228 16725 7280 16777
rect 7292 16725 7344 16777
rect 7356 16725 7408 16777
rect 7420 16725 7472 16777
rect 7484 16725 7536 16777
rect 7548 16725 7600 16777
rect 7612 16725 7664 16777
rect 7676 16725 7728 16777
rect 7740 16725 7792 16777
rect 7804 16725 7856 16777
rect 7868 16725 7920 16777
rect 7932 16725 7984 16777
rect 7996 16725 8048 16777
rect 8060 16725 8112 16777
rect 8124 16725 8176 16777
rect 8188 16725 8240 16777
rect 8252 16725 8304 16777
rect 8316 16725 8368 16777
rect 8380 16725 8432 16777
rect 8444 16725 8496 16777
rect 8508 16725 8560 16777
rect 8572 16725 8624 16777
rect 8636 16725 8688 16777
rect 8700 16725 8752 16777
rect 8764 16725 8816 16777
rect 8828 16725 8880 16777
rect 8892 16725 8944 16777
rect 8956 16725 9008 16777
rect 9020 16725 9072 16777
rect 9084 16725 9136 16777
rect 7402 16102 7454 16154
rect 7469 16102 7521 16154
rect 7536 16102 7588 16154
rect 7602 16102 7654 16154
rect 7402 16030 7454 16082
rect 7469 16030 7521 16082
rect 7536 16030 7588 16082
rect 7602 16030 7654 16082
rect 7402 15958 7454 16010
rect 7469 15958 7521 16010
rect 7536 15958 7588 16010
rect 7602 15958 7654 16010
rect 9196 16102 9248 16154
rect 9196 16030 9248 16082
rect 9196 15958 9248 16010
rect 1590 15457 1642 15509
rect 1654 15457 1706 15509
rect 5816 13855 5827 13865
rect 5827 13855 5861 13865
rect 5861 13855 5868 13865
rect 5816 13813 5868 13855
rect 5816 13781 5868 13801
rect 5816 13749 5827 13781
rect 5827 13749 5861 13781
rect 5861 13749 5868 13781
rect 5816 13529 5826 13562
rect 5826 13529 5860 13562
rect 5860 13529 5868 13562
rect 5816 13510 5868 13529
rect 5816 13455 5868 13498
rect 5816 13446 5826 13455
rect 5826 13446 5860 13455
rect 5860 13446 5868 13455
rect 6025 13502 6077 13554
rect 9477 13522 9529 13574
rect 6025 13438 6077 13490
rect 9477 13458 9529 13510
rect 9359 13007 9411 13059
rect 5816 12876 5829 12910
rect 5829 12876 5863 12910
rect 5863 12876 5868 12910
rect 5816 12858 5868 12876
rect 5816 12828 5868 12846
rect 5816 12794 5829 12828
rect 5829 12794 5863 12828
rect 5863 12794 5868 12828
rect 7533 12893 7585 12945
rect 9359 12943 9411 12995
rect 7533 12829 7585 12881
rect 4715 12220 4767 12272
rect 4715 12156 4767 12208
rect 5163 12220 5215 12272
rect 5163 12156 5215 12208
rect 5705 11852 5757 11904
rect 5705 11782 5757 11834
rect 5705 11739 5730 11764
rect 5730 11739 5757 11764
rect 5705 11712 5757 11739
rect 5705 11665 5730 11694
rect 5730 11665 5757 11694
rect 2845 11610 2897 11662
rect 2909 11610 2961 11662
rect 5705 11642 5757 11665
rect 7663 11695 7715 11747
rect 7727 11695 7779 11747
rect 7952 11695 8004 11747
rect 8016 11695 8068 11747
rect 5705 11591 5730 11624
rect 5730 11591 5757 11624
rect 5705 11572 5757 11591
rect 5705 11551 5757 11553
rect 5705 11517 5730 11551
rect 5730 11517 5757 11551
rect 5705 11501 5757 11517
rect 5705 11430 5757 11482
rect 3000 10333 3052 10385
rect 3065 10333 3117 10385
rect 3130 10333 3182 10385
rect 3194 10333 3246 10385
rect 3258 10333 3310 10385
rect 3322 10333 3374 10385
rect 3386 10333 3438 10385
rect 3450 10333 3502 10385
rect 3514 10333 3566 10385
rect 3578 10333 3630 10385
rect 3642 10333 3694 10385
rect 3706 10333 3758 10385
rect 3000 10257 3052 10309
rect 3065 10257 3117 10309
rect 3130 10257 3182 10309
rect 3194 10257 3246 10309
rect 3258 10257 3310 10309
rect 3322 10257 3374 10309
rect 3386 10257 3438 10309
rect 3450 10257 3502 10309
rect 3514 10257 3566 10309
rect 3578 10257 3630 10309
rect 3642 10257 3694 10309
rect 3706 10257 3758 10309
rect 11007 10281 11059 10333
rect 11081 10281 11133 10333
rect 11155 10281 11207 10333
rect 11229 10281 11281 10333
rect 7406 10192 7458 10244
rect 7487 10192 7539 10244
rect 7567 10192 7619 10244
rect 11007 10217 11059 10269
rect 11081 10217 11133 10269
rect 11155 10217 11207 10269
rect 11229 10217 11281 10269
rect 11007 10153 11059 10205
rect 11081 10153 11133 10205
rect 11155 10153 11207 10205
rect 11229 10153 11281 10205
rect 3993 10079 4045 10131
rect 4057 10079 4109 10131
rect 4546 10079 4598 10131
rect 4610 10079 4662 10131
rect 6897 10079 6949 10131
rect 6961 10079 7013 10131
rect 2231 9999 2283 10051
rect 2299 9999 2351 10051
rect 2367 9999 2419 10051
rect 2435 9999 2487 10051
rect 2503 9999 2555 10051
rect 2571 9999 2623 10051
rect 2638 9999 2690 10051
rect 2231 9925 2283 9977
rect 2299 9925 2351 9977
rect 2367 9925 2419 9977
rect 2435 9925 2487 9977
rect 2503 9925 2555 9977
rect 2571 9925 2623 9977
rect 2638 9925 2690 9977
rect 2231 9851 2283 9903
rect 2299 9851 2351 9903
rect 2367 9851 2419 9903
rect 2435 9851 2487 9903
rect 2503 9851 2555 9903
rect 2571 9851 2623 9903
rect 2638 9851 2690 9903
rect 6943 9925 6995 9977
rect 7220 9976 7272 10028
rect 7284 9976 7336 10028
rect 7822 9976 7874 10028
rect 7886 9976 7938 10028
rect 6943 9861 6995 9913
rect 9654 9855 9706 9907
rect 9718 9855 9770 9907
rect 2231 9777 2283 9829
rect 2299 9777 2351 9829
rect 2367 9777 2419 9829
rect 2435 9777 2487 9829
rect 2503 9777 2555 9829
rect 2571 9777 2623 9829
rect 2638 9777 2690 9829
rect 2231 9703 2283 9755
rect 2299 9703 2351 9755
rect 2367 9703 2419 9755
rect 2435 9703 2487 9755
rect 2503 9703 2555 9755
rect 2571 9703 2623 9755
rect 2638 9703 2690 9755
rect 7409 9583 7461 9635
rect 7488 9583 7540 9635
rect 7567 9583 7619 9635
rect 7434 9491 7486 9543
rect 7434 9415 7486 9467
rect 272 9361 324 9413
rect 348 9361 400 9413
rect 424 9361 476 9413
rect 500 9361 552 9413
rect 10902 9448 10954 9500
rect 10968 9448 11020 9500
rect 11034 9448 11086 9500
rect 11099 9448 11151 9500
rect 11164 9448 11216 9500
rect 11229 9448 11281 9500
rect 272 9287 324 9339
rect 348 9287 400 9339
rect 424 9287 476 9339
rect 500 9287 552 9339
rect 10902 9374 10954 9426
rect 10968 9374 11020 9426
rect 11034 9374 11086 9426
rect 11099 9374 11151 9426
rect 11164 9374 11216 9426
rect 11229 9374 11281 9426
rect 10902 9300 10954 9352
rect 10968 9300 11020 9352
rect 11034 9300 11086 9352
rect 11099 9300 11151 9352
rect 11164 9300 11216 9352
rect 11229 9300 11281 9352
rect 272 9213 324 9265
rect 348 9213 400 9265
rect 424 9213 476 9265
rect 500 9213 552 9265
rect 272 9139 324 9191
rect 348 9143 400 9191
rect 348 9139 359 9143
rect 359 9139 393 9143
rect 393 9139 400 9143
rect 424 9143 476 9191
rect 500 9143 552 9191
rect 424 9139 443 9143
rect 443 9139 476 9143
rect 500 9139 527 9143
rect 527 9139 552 9143
rect 277 9062 329 9114
rect 2784 9207 2836 9259
rect 2851 9207 2903 9259
rect 2918 9207 2970 9259
rect 2985 9207 3037 9259
rect 3052 9207 3104 9259
rect 3119 9207 3171 9259
rect 3186 9207 3238 9259
rect 3253 9207 3305 9259
rect 3320 9207 3372 9259
rect 3387 9207 3439 9259
rect 3454 9207 3506 9259
rect 3521 9207 3573 9259
rect 3588 9207 3640 9259
rect 3654 9207 3706 9259
rect 3720 9207 3772 9259
rect 2784 9133 2836 9185
rect 2851 9133 2903 9185
rect 2918 9133 2970 9185
rect 2985 9133 3037 9185
rect 3052 9133 3104 9185
rect 3119 9133 3171 9185
rect 3186 9133 3238 9185
rect 3253 9133 3305 9185
rect 3320 9133 3372 9185
rect 3387 9133 3439 9185
rect 3454 9133 3506 9185
rect 3521 9133 3573 9185
rect 3588 9133 3640 9185
rect 3654 9133 3706 9185
rect 3720 9133 3772 9185
rect 2784 9059 2836 9111
rect 2851 9059 2903 9111
rect 2918 9059 2970 9111
rect 2985 9059 3037 9111
rect 3052 9059 3104 9111
rect 3119 9059 3171 9111
rect 3186 9059 3238 9111
rect 3253 9059 3305 9111
rect 3320 9059 3372 9111
rect 3387 9059 3439 9111
rect 3454 9059 3506 9111
rect 3521 9059 3573 9111
rect 3588 9059 3640 9111
rect 3654 9059 3706 9111
rect 3720 9059 3772 9111
rect 7399 9202 7451 9254
rect 7519 9202 7571 9254
rect 7399 9133 7451 9185
rect 7519 9133 7571 9185
rect 7399 9064 7451 9116
rect 7519 9064 7571 9116
rect 277 8998 329 9050
rect 277 8933 329 8985
rect 1450 8968 1502 9020
rect 1514 8968 1566 9020
rect 1193 8667 1245 8719
rect 1193 8603 1245 8655
rect 1450 8623 1502 8675
rect 1514 8623 1566 8675
rect 15783 8533 15835 8585
rect 15783 8469 15835 8521
rect 9788 8297 9840 8349
rect 9852 8297 9904 8349
rect 11597 8297 11649 8349
rect 11661 8297 11713 8349
rect 13820 8298 13872 8350
rect 13892 8298 13944 8350
rect 13964 8298 14016 8350
rect 14036 8298 14088 8350
rect 14107 8298 14159 8350
rect 14178 8298 14230 8350
rect 14249 8298 14301 8350
rect 2845 8217 2897 8269
rect 2913 8217 2965 8269
rect 2981 8217 3033 8269
rect 3049 8217 3101 8269
rect 3117 8217 3169 8269
rect 3184 8217 3236 8269
rect 3251 8217 3303 8269
rect 3318 8217 3370 8269
rect 3385 8217 3437 8269
rect 3452 8217 3504 8269
rect 3519 8217 3571 8269
rect 3586 8217 3638 8269
rect 3653 8217 3705 8269
rect 3720 8217 3772 8269
rect 2845 8139 2897 8191
rect 2913 8139 2965 8191
rect 2981 8139 3033 8191
rect 3049 8139 3101 8191
rect 3117 8139 3169 8191
rect 3184 8139 3236 8191
rect 3251 8139 3303 8191
rect 3318 8139 3370 8191
rect 3385 8139 3437 8191
rect 3452 8139 3504 8191
rect 3519 8139 3571 8191
rect 3586 8139 3638 8191
rect 3653 8139 3705 8191
rect 3720 8139 3772 8191
rect 10502 8217 10554 8269
rect 10591 8217 10643 8269
rect 10680 8217 10732 8269
rect 13820 8220 13872 8272
rect 13892 8220 13944 8272
rect 13964 8220 14016 8272
rect 14036 8220 14088 8272
rect 14107 8220 14159 8272
rect 14178 8220 14230 8272
rect 14249 8220 14301 8272
rect 10502 8139 10554 8191
rect 10591 8139 10643 8191
rect 10680 8139 10732 8191
rect 4625 7739 4677 7791
rect 4689 7739 4741 7791
rect 6873 7739 6925 7791
rect 6937 7739 6989 7791
rect 7187 7744 7239 7796
rect 7251 7744 7303 7796
rect 10331 7744 10383 7796
rect 10395 7744 10447 7796
rect 10779 6304 10831 6356
rect 10843 6304 10895 6356
rect 12036 6304 12088 6356
rect 12100 6304 12152 6356
rect 11814 5975 11866 6027
rect 11878 5975 11930 6027
rect 12467 5975 12519 6027
rect 12531 5975 12583 6027
rect 6858 4231 6910 4283
rect 6922 4231 6974 4283
rect 8637 4239 8689 4291
rect 8701 4239 8753 4291
rect 1054 4114 1106 4166
rect 1054 4050 1106 4102
rect 1457 4071 1509 4123
rect 1521 4071 1573 4123
rect 1966 3622 2018 3674
rect 2030 3622 2082 3674
rect 5521 3622 5573 3674
rect 5585 3622 5637 3674
rect 14310 3347 14362 3399
rect 14374 3347 14426 3399
rect 15361 3347 15413 3399
rect 15425 3347 15477 3399
rect 6854 3292 6906 3344
rect 6934 3292 6986 3344
rect 7013 3292 7065 3344
rect 6854 3220 6906 3272
rect 6934 3220 6986 3272
rect 7013 3220 7065 3272
rect 6854 3148 6906 3200
rect 6934 3148 6986 3200
rect 7013 3148 7065 3200
rect 8621 3293 8673 3345
rect 8717 3293 8769 3345
rect 8621 3219 8673 3271
rect 8717 3219 8769 3271
rect 8621 3145 8673 3197
rect 8717 3145 8769 3197
rect 42 2750 94 2802
rect 42 2686 94 2738
rect 2446 2594 2498 2646
rect 2511 2594 2563 2646
rect 2575 2594 2627 2646
rect 2639 2594 2691 2646
rect 2703 2594 2755 2646
rect 2446 2522 2498 2574
rect 2511 2522 2563 2574
rect 2575 2522 2627 2574
rect 2639 2522 2691 2574
rect 2703 2522 2755 2574
rect 2446 2450 2498 2502
rect 2511 2450 2563 2502
rect 2575 2450 2627 2502
rect 2639 2450 2691 2502
rect 2703 2450 2755 2502
rect 3633 2594 3685 2646
rect 3702 2594 3754 2646
rect 3771 2594 3823 2646
rect 3840 2594 3892 2646
rect 3909 2594 3961 2646
rect 3978 2594 4030 2646
rect 4047 2594 4099 2646
rect 4116 2594 4168 2646
rect 4185 2594 4237 2646
rect 4254 2594 4306 2646
rect 3633 2522 3685 2574
rect 3702 2522 3754 2574
rect 3771 2522 3823 2574
rect 3840 2522 3892 2574
rect 3909 2522 3961 2574
rect 3978 2522 4030 2574
rect 4047 2522 4099 2574
rect 4116 2522 4168 2574
rect 4185 2522 4237 2574
rect 4254 2522 4306 2574
rect 3633 2450 3685 2502
rect 3702 2450 3754 2502
rect 3771 2450 3823 2502
rect 3840 2450 3892 2502
rect 3909 2450 3961 2502
rect 3978 2450 4030 2502
rect 4047 2450 4099 2502
rect 4116 2450 4168 2502
rect 4185 2450 4237 2502
rect 4254 2450 4306 2502
rect 10512 2595 10564 2647
rect 10579 2595 10631 2647
rect 10512 2523 10564 2575
rect 10579 2523 10631 2575
rect 10512 2451 10564 2503
rect 10579 2451 10631 2503
rect 10707 2595 10759 2647
rect 10780 2595 10832 2647
rect 10853 2595 10905 2647
rect 10926 2595 10978 2647
rect 10999 2595 11051 2647
rect 10707 2523 10759 2575
rect 10780 2523 10832 2575
rect 10853 2523 10905 2575
rect 10926 2523 10978 2575
rect 10999 2523 11051 2575
rect 10707 2451 10759 2503
rect 10780 2451 10832 2503
rect 10853 2451 10905 2503
rect 10926 2451 10978 2503
rect 10999 2451 11051 2503
rect 15421 2371 15473 2423
rect 15421 2307 15473 2359
rect 330 2123 382 2175
rect 394 2123 446 2175
rect 811 2123 863 2175
rect 875 2123 927 2175
rect 14632 2053 14684 2105
rect 14711 2053 14763 2105
rect 14789 2053 14841 2105
rect 14632 1981 14684 2033
rect 14711 1981 14763 2033
rect 14789 1981 14841 2033
rect 14632 1909 14684 1961
rect 14711 1909 14763 1961
rect 14789 1909 14841 1961
rect 15077 2047 15129 2099
rect 15199 2047 15251 2099
rect 15077 1981 15129 2033
rect 15199 1981 15251 2033
rect 15077 1915 15129 1967
rect 15199 1915 15251 1967
rect 1497 1752 1549 1804
rect 1573 1752 1625 1804
rect 1497 1686 1549 1738
rect 1573 1686 1625 1738
rect 6854 1758 6906 1810
rect 6934 1758 6986 1810
rect 7013 1758 7065 1810
rect 6854 1680 6906 1732
rect 6934 1680 6986 1732
rect 7013 1680 7065 1732
rect 8621 1758 8673 1810
rect 8717 1758 8769 1810
rect 8621 1680 8673 1732
rect 8717 1680 8769 1732
rect 1499 1594 1551 1646
rect 1603 1594 1655 1646
rect 1499 1525 1551 1577
rect 1603 1525 1655 1577
rect 1499 1456 1551 1508
rect 1603 1456 1655 1508
rect 1786 1599 1838 1651
rect 1786 1525 1838 1577
rect 1786 1451 1838 1503
rect 3853 1599 3905 1651
rect 3926 1599 3978 1651
rect 3999 1599 4051 1651
rect 4072 1599 4124 1651
rect 4145 1599 4197 1651
rect 4217 1599 4269 1651
rect 3853 1525 3905 1577
rect 3926 1525 3978 1577
rect 3999 1525 4051 1577
rect 4072 1525 4124 1577
rect 4145 1525 4197 1577
rect 4217 1525 4269 1577
rect 3853 1451 3905 1503
rect 3926 1451 3978 1503
rect 3999 1451 4051 1503
rect 4072 1451 4124 1503
rect 4145 1451 4197 1503
rect 4217 1451 4269 1503
rect 4854 1599 4906 1651
rect 4923 1599 4975 1651
rect 4991 1599 5043 1651
rect 5059 1599 5111 1651
rect 5127 1599 5179 1651
rect 5195 1599 5247 1651
rect 4854 1525 4906 1577
rect 4923 1525 4975 1577
rect 4991 1525 5043 1577
rect 5059 1525 5111 1577
rect 5127 1525 5179 1577
rect 5195 1525 5247 1577
rect 4854 1451 4906 1503
rect 4923 1451 4975 1503
rect 4991 1451 5043 1503
rect 5059 1451 5111 1503
rect 5127 1451 5179 1503
rect 5195 1451 5247 1503
rect 6844 1599 6896 1651
rect 6922 1599 6974 1651
rect 6999 1599 7051 1651
rect 6844 1525 6896 1577
rect 6922 1525 6974 1577
rect 6999 1525 7051 1577
rect 6844 1451 6896 1503
rect 6922 1451 6974 1503
rect 6999 1451 7051 1503
rect 1188 1285 1240 1337
rect 1252 1285 1304 1337
rect 3214 1124 3266 1176
rect 3278 1124 3330 1176
rect 8938 1124 8990 1176
rect 9002 1124 9054 1176
rect 12492 1109 12544 1161
rect 12556 1109 12608 1161
rect 2785 1034 2837 1086
rect 2857 1034 2909 1086
rect 2928 1034 2980 1086
rect 2999 1034 3051 1086
rect 3070 1034 3122 1086
rect 3141 1034 3193 1086
rect 3212 1034 3264 1086
rect 3283 1034 3335 1086
rect 2785 958 2837 1010
rect 2857 958 2909 1010
rect 2928 958 2980 1010
rect 2999 958 3051 1010
rect 3070 958 3122 1010
rect 3141 958 3193 1010
rect 3212 958 3264 1010
rect 3283 958 3335 1010
rect 2785 882 2837 934
rect 2857 882 2909 934
rect 2928 882 2980 934
rect 2999 882 3051 934
rect 3070 882 3122 934
rect 3141 882 3193 934
rect 3212 882 3264 934
rect 3283 882 3335 934
rect 10511 1038 10563 1090
rect 10577 1038 10629 1090
rect 10643 1038 10695 1090
rect 10708 1038 10760 1090
rect 10773 1038 10825 1090
rect 10511 958 10563 1010
rect 10577 958 10629 1010
rect 10643 958 10695 1010
rect 10708 958 10760 1010
rect 10773 958 10825 1010
rect 10511 878 10563 930
rect 10577 878 10629 930
rect 10643 878 10695 930
rect 10708 878 10760 930
rect 10773 878 10825 930
rect 15092 1026 15144 1078
rect 15193 1026 15245 1078
rect 15092 962 15144 1014
rect 15193 962 15245 1014
rect 15439 1034 15491 1046
rect 15439 1000 15473 1034
rect 15473 1000 15491 1034
rect 15439 994 15491 1000
rect 15503 1034 15555 1046
rect 15503 1000 15521 1034
rect 15521 1000 15555 1034
rect 15503 994 15555 1000
rect 15439 948 15491 958
rect 15439 914 15473 948
rect 15473 914 15491 948
rect 15439 906 15491 914
rect 15503 948 15555 958
rect 15503 914 15521 948
rect 15521 914 15555 948
rect 15503 906 15555 914
rect 6363 735 6415 787
rect 8936 787 8988 839
rect 15439 862 15491 870
rect 15439 828 15473 862
rect 15473 828 15491 862
rect 15439 818 15491 828
rect 15503 862 15555 870
rect 15503 828 15521 862
rect 15521 828 15555 862
rect 15503 818 15555 828
rect 6363 668 6415 720
rect 7027 719 7079 771
rect 8936 723 8988 775
rect 13655 784 13707 786
rect 13733 784 13785 786
rect 7027 655 7079 707
rect 9776 709 9828 761
rect 9776 645 9828 697
rect 10216 710 10268 762
rect 10216 640 10268 692
rect 10320 710 10372 762
rect 11416 724 11468 776
rect 11487 724 11539 776
rect 12054 718 12106 770
rect 12118 718 12170 770
rect 13655 734 13664 784
rect 13664 734 13707 784
rect 13733 734 13770 784
rect 13770 734 13785 784
rect 10320 640 10372 692
rect 15439 775 15491 782
rect 15439 741 15473 775
rect 15473 741 15491 775
rect 15439 730 15491 741
rect 15503 775 15555 782
rect 15503 741 15521 775
rect 15521 741 15555 775
rect 15503 730 15555 741
rect 13655 664 13664 716
rect 13664 664 13707 716
rect 13733 664 13770 716
rect 13770 664 13785 716
rect 13655 606 13664 646
rect 13664 606 13707 646
rect 13733 606 13770 646
rect 13770 606 13785 646
rect 13655 594 13707 606
rect 13733 594 13785 606
rect 2314 523 2366 575
rect 2378 523 2430 575
rect 11890 558 11942 564
rect 11890 524 11899 558
rect 11899 524 11933 558
rect 11933 524 11942 558
rect 1175 467 1227 519
rect 1239 467 1291 519
rect 1902 467 1954 519
rect 1966 467 2018 519
rect 11890 512 11942 524
rect 11890 486 11942 498
rect 10182 431 10234 483
rect 10246 431 10298 483
rect 11890 452 11899 486
rect 11899 452 11933 486
rect 11933 452 11942 486
rect 11890 446 11942 452
rect 13655 567 13707 576
rect 13655 533 13664 567
rect 13664 533 13698 567
rect 13698 533 13707 567
rect 13655 524 13707 533
rect 13733 567 13785 576
rect 13733 533 13736 567
rect 13736 533 13770 567
rect 13770 533 13785 567
rect 13733 524 13785 533
rect 13655 494 13707 506
rect 13655 460 13664 494
rect 13664 460 13698 494
rect 13698 460 13707 494
rect 13655 454 13707 460
rect 13733 494 13785 506
rect 13733 460 13736 494
rect 13736 460 13770 494
rect 13770 460 13785 494
rect 13733 454 13785 460
rect 7884 285 7936 337
rect 7948 285 8000 337
rect 12486 325 12538 377
rect 12486 261 12538 313
rect 1440 203 1492 255
rect 1548 203 1600 255
rect 1656 203 1708 255
rect 1764 203 1816 255
rect 1871 203 1923 255
rect 1978 203 2030 255
rect 2085 203 2137 255
rect 1440 129 1492 181
rect 1548 129 1600 181
rect 1656 129 1708 181
rect 1764 129 1816 181
rect 1871 129 1923 181
rect 1978 129 2030 181
rect 2085 129 2137 181
rect 1440 55 1492 107
rect 1548 55 1600 107
rect 1656 55 1708 107
rect 1764 55 1816 107
rect 1871 55 1923 107
rect 1978 55 2030 107
rect 2085 55 2137 107
rect 3853 203 3905 255
rect 3926 203 3978 255
rect 3999 203 4051 255
rect 4072 203 4124 255
rect 4145 203 4197 255
rect 4217 203 4269 255
rect 3853 129 3905 181
rect 3926 129 3978 181
rect 3999 129 4051 181
rect 4072 129 4124 181
rect 4145 129 4197 181
rect 4217 129 4269 181
rect 3853 55 3905 107
rect 3926 55 3978 107
rect 3999 55 4051 107
rect 4072 55 4124 107
rect 4145 55 4197 107
rect 4217 55 4269 107
rect 4660 204 4712 256
rect 4767 204 4819 256
rect 4874 204 4926 256
rect 4981 204 5033 256
rect 5088 204 5140 256
rect 5195 204 5247 256
rect 4660 130 4712 182
rect 4767 130 4819 182
rect 4874 130 4926 182
rect 4981 130 5033 182
rect 5088 130 5140 182
rect 5195 130 5247 182
rect 4660 56 4712 108
rect 4767 56 4819 108
rect 4874 56 4926 108
rect 4981 56 5033 108
rect 5088 56 5140 108
rect 5195 56 5247 108
rect 6686 203 6738 255
rect 6781 203 6833 255
rect 6876 203 6928 255
rect 6686 129 6738 181
rect 6781 129 6833 181
rect 6876 129 6928 181
rect 6686 55 6738 107
rect 6781 55 6833 107
rect 6876 55 6928 107
rect 12881 171 12933 180
rect 12982 171 13034 180
rect 12881 137 12887 171
rect 12887 137 12921 171
rect 12921 137 12933 171
rect 12982 137 12994 171
rect 12994 137 13033 171
rect 13033 137 13034 171
rect 12881 128 12933 137
rect 12982 128 13034 137
rect 12881 93 12933 104
rect 12982 93 13034 104
rect 12881 59 12887 93
rect 12887 59 12921 93
rect 12921 59 12933 93
rect 12982 59 12994 93
rect 12994 59 13033 93
rect 13033 59 13034 93
rect 12881 52 12933 59
rect 12982 52 13034 59
<< metal2 >>
rect 14399 39998 15371 40000
rect 1351 39950 1903 39995
rect 1351 39894 1361 39950
rect 1417 39894 1443 39950
rect 1499 39894 1525 39950
rect 1581 39894 1607 39950
rect 1663 39894 1689 39950
rect 1745 39939 1903 39950
rect 1959 39939 1984 39995
rect 2040 39939 2065 39995
rect 2121 39939 2146 39995
rect 2202 39939 2227 39995
rect 2283 39939 2308 39995
rect 2364 39939 2389 39995
rect 2445 39939 2470 39995
rect 2526 39939 2551 39995
rect 2607 39939 2632 39995
rect 2688 39939 2713 39995
rect 2769 39939 2794 39995
rect 2850 39939 2875 39995
rect 2931 39939 2956 39995
rect 3012 39939 3037 39995
rect 3093 39939 3118 39995
rect 11334 39994 11343 39995
rect 11337 39942 11343 39994
rect 1745 39915 3118 39939
rect 11334 39926 11343 39942
rect 1745 39894 1903 39915
rect 1351 39868 1903 39894
rect 1351 39812 1361 39868
rect 1417 39812 1443 39868
rect 1499 39812 1525 39868
rect 1581 39812 1607 39868
rect 1663 39812 1689 39868
rect 1745 39859 1903 39868
rect 1959 39859 1984 39915
rect 2040 39859 2065 39915
rect 2121 39859 2146 39915
rect 2202 39859 2227 39915
rect 2283 39859 2308 39915
rect 2364 39859 2389 39915
rect 2445 39859 2470 39915
rect 2526 39859 2551 39915
rect 2607 39859 2632 39915
rect 2688 39859 2713 39915
rect 2769 39859 2794 39915
rect 2850 39859 2875 39915
rect 2931 39859 2956 39915
rect 3012 39859 3037 39915
rect 3093 39859 3118 39915
rect 11337 39874 11343 39926
rect 1745 39835 3118 39859
rect 11334 39858 11343 39874
rect 1745 39812 1903 39835
rect 1351 39786 1903 39812
rect 1351 39730 1361 39786
rect 1417 39730 1443 39786
rect 1499 39730 1525 39786
rect 1581 39730 1607 39786
rect 1663 39730 1689 39786
rect 1745 39779 1903 39786
rect 1959 39779 1984 39835
rect 2040 39779 2065 39835
rect 2121 39779 2146 39835
rect 2202 39779 2227 39835
rect 2283 39779 2308 39835
rect 2364 39779 2389 39835
rect 2445 39779 2470 39835
rect 2526 39779 2551 39835
rect 2607 39779 2632 39835
rect 2688 39779 2713 39835
rect 2769 39779 2794 39835
rect 2850 39779 2875 39835
rect 2931 39779 2956 39835
rect 3012 39779 3037 39835
rect 3093 39779 3118 39835
rect 11337 39806 11343 39858
rect 11334 39790 11343 39806
rect 1745 39755 3118 39779
rect 1745 39730 1903 39755
rect 1351 39704 1903 39730
rect 1351 39648 1361 39704
rect 1417 39648 1443 39704
rect 1499 39648 1525 39704
rect 1581 39648 1607 39704
rect 1663 39648 1689 39704
rect 1745 39699 1903 39704
rect 1959 39699 1984 39755
rect 2040 39699 2065 39755
rect 2121 39699 2146 39755
rect 2202 39699 2227 39755
rect 2283 39699 2308 39755
rect 2364 39699 2389 39755
rect 2445 39699 2470 39755
rect 2526 39699 2551 39755
rect 2607 39699 2632 39755
rect 2688 39699 2713 39755
rect 2769 39699 2794 39755
rect 2850 39699 2875 39755
rect 2931 39699 2956 39755
rect 3012 39699 3037 39755
rect 3093 39699 3118 39755
rect 11337 39738 11343 39790
rect 14399 39946 14405 39998
rect 14457 39995 14470 39998
rect 14522 39995 14535 39998
rect 14587 39995 14600 39998
rect 14652 39995 14665 39998
rect 14467 39946 14470 39995
rect 14652 39946 14654 39995
rect 14717 39946 14730 39998
rect 14782 39995 14795 39998
rect 14847 39995 14860 39998
rect 14912 39995 14925 39998
rect 14977 39995 14990 39998
rect 14791 39946 14795 39995
rect 15042 39946 15055 39998
rect 15107 39995 15120 39998
rect 15172 39995 15185 39998
rect 15237 39995 15249 39998
rect 15301 39995 15313 39998
rect 15113 39946 15120 39995
rect 15365 39946 15371 39998
rect 14399 39939 14411 39946
rect 14467 39939 14492 39946
rect 14548 39939 14573 39946
rect 14629 39939 14654 39946
rect 14710 39939 14735 39946
rect 14791 39939 14816 39946
rect 14872 39939 14897 39946
rect 14953 39939 14977 39946
rect 15033 39939 15057 39946
rect 15113 39939 15137 39946
rect 15193 39939 15217 39946
rect 15273 39939 15297 39946
rect 15353 39939 15371 39946
rect 14399 39930 15371 39939
rect 14399 39878 14405 39930
rect 14457 39899 14470 39930
rect 14522 39899 14535 39930
rect 14587 39899 14600 39930
rect 14652 39899 14665 39930
rect 14467 39878 14470 39899
rect 14652 39878 14654 39899
rect 14717 39878 14730 39930
rect 14782 39899 14795 39930
rect 14847 39899 14860 39930
rect 14912 39899 14925 39930
rect 14977 39899 14990 39930
rect 14791 39878 14795 39899
rect 15042 39878 15055 39930
rect 15107 39899 15120 39930
rect 15172 39899 15185 39930
rect 15237 39899 15249 39930
rect 15301 39899 15313 39930
rect 15113 39878 15120 39899
rect 15365 39878 15371 39930
rect 14399 39862 14411 39878
rect 14467 39862 14492 39878
rect 14548 39862 14573 39878
rect 14629 39862 14654 39878
rect 14710 39862 14735 39878
rect 14791 39862 14816 39878
rect 14872 39862 14897 39878
rect 14953 39862 14977 39878
rect 15033 39862 15057 39878
rect 15113 39862 15137 39878
rect 15193 39862 15217 39878
rect 15273 39862 15297 39878
rect 15353 39862 15371 39878
rect 14399 39810 14405 39862
rect 14467 39843 14470 39862
rect 14652 39843 14654 39862
rect 14457 39810 14470 39843
rect 14522 39810 14535 39843
rect 14587 39810 14600 39843
rect 14652 39810 14665 39843
rect 14717 39810 14730 39862
rect 14791 39843 14795 39862
rect 14782 39810 14795 39843
rect 14847 39810 14860 39843
rect 14912 39810 14925 39843
rect 14977 39810 14990 39843
rect 15042 39810 15055 39862
rect 15113 39843 15120 39862
rect 15107 39810 15120 39843
rect 15172 39810 15185 39843
rect 15237 39810 15249 39843
rect 15301 39810 15313 39843
rect 15365 39810 15371 39862
rect 14399 39803 15371 39810
rect 14399 39794 14411 39803
rect 14467 39794 14492 39803
rect 14548 39794 14573 39803
rect 14629 39794 14654 39803
rect 14710 39794 14735 39803
rect 14791 39794 14816 39803
rect 14872 39794 14897 39803
rect 14953 39794 14977 39803
rect 15033 39794 15057 39803
rect 15113 39794 15137 39803
rect 15193 39794 15217 39803
rect 15273 39794 15297 39803
rect 15353 39794 15371 39803
rect 14399 39742 14405 39794
rect 14467 39747 14470 39794
rect 14652 39747 14654 39794
rect 14457 39742 14470 39747
rect 14522 39742 14535 39747
rect 14587 39742 14600 39747
rect 14652 39742 14665 39747
rect 14717 39742 14730 39794
rect 14791 39747 14795 39794
rect 14782 39742 14795 39747
rect 14847 39742 14860 39747
rect 14912 39742 14925 39747
rect 14977 39742 14990 39747
rect 15042 39742 15055 39794
rect 15113 39747 15120 39794
rect 15107 39742 15120 39747
rect 15172 39742 15185 39747
rect 15237 39742 15249 39747
rect 15301 39742 15313 39747
rect 15365 39742 15371 39794
rect 14399 39740 15371 39742
rect 1745 39675 3118 39699
rect 1745 39648 1903 39675
rect 1351 39622 1903 39648
rect 1351 39566 1361 39622
rect 1417 39566 1443 39622
rect 1499 39566 1525 39622
rect 1581 39566 1607 39622
rect 1663 39566 1689 39622
rect 1745 39619 1903 39622
rect 1959 39619 1984 39675
rect 2040 39619 2065 39675
rect 2121 39619 2146 39675
rect 2202 39619 2227 39675
rect 2283 39619 2308 39675
rect 2364 39619 2389 39675
rect 2445 39619 2470 39675
rect 2526 39619 2551 39675
rect 2607 39619 2632 39675
rect 2688 39619 2713 39675
rect 2769 39619 2794 39675
rect 2850 39619 2875 39675
rect 2931 39619 2956 39675
rect 3012 39619 3037 39675
rect 3093 39619 3118 39675
rect 1745 39595 3118 39619
rect 1745 39566 1903 39595
rect 1351 39543 1903 39566
rect 1361 39540 1903 39543
rect 1417 39484 1443 39540
rect 1499 39484 1525 39540
rect 1581 39484 1607 39540
rect 1663 39484 1689 39540
rect 1745 39539 1903 39540
rect 1959 39539 1984 39595
rect 2040 39539 2065 39595
rect 2121 39539 2146 39595
rect 2202 39539 2227 39595
rect 2283 39539 2308 39595
rect 2364 39539 2389 39595
rect 2445 39539 2470 39595
rect 2526 39539 2551 39595
rect 2607 39539 2632 39595
rect 2688 39539 2713 39595
rect 2769 39539 2794 39595
rect 2850 39539 2875 39595
rect 2931 39539 2956 39595
rect 3012 39539 3037 39595
rect 3093 39539 3118 39595
rect 11334 39539 11343 39738
rect 1361 39458 1745 39484
rect 1417 39402 1443 39458
rect 1499 39402 1525 39458
rect 1581 39402 1607 39458
rect 1663 39402 1689 39458
rect 1361 39376 1745 39402
rect 1417 39320 1443 39376
rect 1499 39320 1525 39376
rect 1581 39320 1607 39376
rect 1663 39320 1689 39376
rect 1361 39294 1745 39320
rect 1417 39238 1443 39294
rect 1499 39238 1525 39294
rect 1581 39238 1607 39294
rect 1663 39238 1689 39294
tri 1745 39246 2038 39539 nw
rect 1361 39212 1745 39238
rect 1417 39156 1443 39212
rect 1499 39156 1525 39212
rect 1581 39156 1607 39212
rect 1663 39156 1689 39212
rect 1361 39130 1745 39156
rect 1417 39074 1443 39130
rect 1499 39074 1525 39130
rect 1581 39074 1607 39130
rect 1663 39074 1689 39130
rect 1361 39048 1745 39074
rect 1417 38992 1443 39048
rect 1499 38992 1525 39048
rect 1581 38992 1607 39048
rect 1663 38992 1689 39048
rect 1361 38966 1745 38992
rect 1417 38910 1443 38966
rect 1499 38910 1525 38966
rect 1581 38910 1607 38966
rect 1663 38910 1689 38966
rect 1361 38884 1745 38910
rect 1417 38828 1443 38884
rect 1499 38828 1525 38884
rect 1581 38828 1607 38884
rect 1663 38828 1689 38884
rect 1361 38802 1745 38828
rect 1417 38746 1443 38802
rect 1499 38746 1525 38802
rect 1581 38746 1607 38802
rect 1663 38746 1689 38802
rect 1361 38720 1745 38746
rect 1417 38664 1443 38720
rect 1499 38664 1525 38720
rect 1581 38664 1607 38720
rect 1663 38664 1689 38720
rect 1361 38638 1745 38664
rect 1417 38582 1443 38638
rect 1499 38582 1525 38638
rect 1581 38582 1607 38638
rect 1663 38582 1689 38638
rect 1361 38556 1745 38582
rect 1417 38500 1443 38556
rect 1499 38500 1525 38556
rect 1581 38500 1607 38556
rect 1663 38500 1689 38556
rect 1361 38474 1745 38500
rect 1417 38418 1443 38474
rect 1499 38418 1525 38474
rect 1581 38418 1607 38474
rect 1663 38418 1689 38474
rect 1361 38392 1745 38418
rect 1417 38336 1443 38392
rect 1499 38336 1525 38392
rect 1581 38336 1607 38392
rect 1663 38336 1689 38392
rect 1361 38310 1745 38336
rect 1417 38254 1443 38310
rect 1499 38254 1525 38310
rect 1581 38254 1607 38310
rect 1663 38254 1689 38310
rect 1361 38228 1745 38254
rect 1417 38172 1443 38228
rect 1499 38172 1525 38228
rect 1581 38172 1607 38228
rect 1663 38172 1689 38228
rect 1361 38146 1745 38172
rect 1417 38090 1443 38146
rect 1499 38090 1525 38146
rect 1581 38090 1607 38146
rect 1663 38090 1689 38146
rect 1361 38064 1745 38090
rect 1417 38008 1443 38064
rect 1499 38008 1525 38064
rect 1581 38008 1607 38064
rect 1663 38008 1689 38064
rect 1361 37981 1745 38008
rect 1417 37925 1443 37981
rect 1499 37925 1525 37981
rect 1581 37925 1607 37981
rect 1663 37925 1689 37981
rect 1361 37898 1745 37925
rect 1417 37842 1443 37898
rect 1499 37842 1525 37898
rect 1581 37842 1607 37898
rect 1663 37842 1689 37898
rect 1361 37815 1745 37842
rect 1417 37759 1443 37815
rect 1499 37759 1525 37815
rect 1581 37759 1607 37815
rect 1663 37759 1689 37815
rect 1361 37732 1745 37759
rect 1417 37676 1443 37732
rect 1499 37676 1525 37732
rect 1581 37676 1607 37732
rect 1663 37676 1689 37732
rect 1361 37649 1745 37676
rect 1417 37593 1443 37649
rect 1499 37593 1525 37649
rect 1581 37593 1607 37649
rect 1663 37593 1689 37649
rect 1361 37566 1745 37593
rect 1417 37510 1443 37566
rect 1499 37510 1525 37566
rect 1581 37510 1607 37566
rect 1663 37510 1689 37566
rect 1361 37483 1745 37510
rect 1417 37427 1443 37483
rect 1499 37427 1525 37483
rect 1581 37427 1607 37483
rect 1663 37427 1689 37483
rect 1361 37400 1745 37427
rect 1417 37344 1443 37400
rect 1499 37344 1525 37400
rect 1581 37344 1607 37400
rect 1663 37344 1689 37400
rect 1361 37317 1745 37344
rect 1417 37261 1443 37317
rect 1499 37261 1525 37317
rect 1581 37261 1607 37317
rect 1663 37261 1689 37317
rect 1361 37234 1745 37261
rect 1417 37178 1443 37234
rect 1499 37178 1525 37234
rect 1581 37178 1607 37234
rect 1663 37178 1689 37234
rect 1361 37169 1745 37178
rect 4080 36310 4089 36366
rect 4145 36310 4231 36366
rect 4287 36310 4372 36366
rect 4428 36310 4513 36366
rect 4569 36310 4654 36366
rect 4710 36310 4719 36366
rect 4080 36266 4719 36310
tri 802 36203 837 36238 se
rect 837 36229 893 36238
tri 893 36210 921 36238 sw
rect 4080 36210 4089 36266
rect 4145 36210 4231 36266
rect 4287 36210 4372 36266
rect 4428 36210 4513 36266
rect 4569 36210 4654 36266
rect 4710 36210 4719 36266
rect 893 36209 921 36210
tri 921 36209 922 36210 sw
rect 893 36203 922 36209
rect 837 36149 893 36173
rect 837 36084 893 36093
rect 2783 36081 3776 36082
rect 2783 36025 2792 36081
rect 2848 36079 2924 36081
rect 2980 36079 3056 36081
rect 3112 36079 3187 36081
rect 3243 36079 3318 36081
rect 3374 36079 3449 36081
rect 3505 36079 3580 36081
rect 3636 36079 3711 36081
rect 2848 36027 2858 36079
rect 2910 36027 2924 36079
rect 2980 36027 2990 36079
rect 3042 36027 3056 36079
rect 3112 36027 3122 36079
rect 3174 36027 3187 36079
rect 3243 36027 3254 36079
rect 3306 36027 3318 36079
rect 3374 36027 3386 36079
rect 3438 36027 3449 36079
rect 3505 36027 3518 36079
rect 3570 36027 3580 36079
rect 3636 36027 3650 36079
rect 3702 36027 3711 36079
rect 2848 36025 2924 36027
rect 2980 36025 3056 36027
rect 3112 36025 3187 36027
rect 3243 36025 3318 36027
rect 3374 36025 3449 36027
rect 3505 36025 3580 36027
rect 3636 36025 3711 36027
rect 3767 36025 3776 36081
rect 2783 36001 3776 36025
rect 2783 35871 2792 36001
rect 2844 35963 2858 36001
rect 2848 35949 2858 35963
rect 2910 35949 2924 36001
rect 2976 35963 2990 36001
rect 2980 35949 2990 35963
rect 3042 35949 3056 36001
rect 3108 35963 3122 36001
rect 3112 35949 3122 35963
rect 3174 35963 3188 36001
rect 3240 35963 3254 36001
rect 3174 35949 3187 35963
rect 3243 35949 3254 35963
rect 3306 35963 3320 36001
rect 3372 35963 3386 36001
rect 3306 35949 3318 35963
rect 3374 35949 3386 35963
rect 3438 35963 3452 36001
rect 3504 35963 3518 36001
rect 3438 35949 3449 35963
rect 3505 35949 3518 35963
rect 3570 35963 3584 36001
rect 3570 35949 3580 35963
rect 3636 35949 3650 36001
rect 3702 35963 3715 36001
rect 3702 35949 3711 35963
rect 2848 35923 2924 35949
rect 2980 35923 3056 35949
rect 3112 35923 3187 35949
rect 3243 35923 3318 35949
rect 3374 35923 3449 35949
rect 3505 35923 3580 35949
rect 3636 35923 3711 35949
rect 2848 35907 2858 35923
rect 2844 35871 2858 35907
rect 2910 35871 2924 35923
rect 2980 35907 2990 35923
rect 2976 35871 2990 35907
rect 3042 35871 3056 35923
rect 3112 35907 3122 35923
rect 3108 35871 3122 35907
rect 3174 35907 3187 35923
rect 3243 35907 3254 35923
rect 3174 35871 3188 35907
rect 3240 35871 3254 35907
rect 3306 35907 3318 35923
rect 3374 35907 3386 35923
rect 3306 35871 3320 35907
rect 3372 35871 3386 35907
rect 3438 35907 3449 35923
rect 3505 35907 3518 35923
rect 3438 35871 3452 35907
rect 3504 35871 3518 35907
rect 3570 35907 3580 35923
rect 3570 35871 3584 35907
rect 3636 35871 3650 35923
rect 3702 35907 3711 35923
rect 3702 35871 3715 35907
rect 3767 35871 3776 36001
rect 2783 35845 3776 35871
rect 2783 35789 2792 35845
rect 2848 35793 2858 35845
rect 2910 35793 2924 35845
rect 2980 35793 2990 35845
rect 3042 35793 3056 35845
rect 3112 35793 3122 35845
rect 3174 35793 3187 35845
rect 3243 35793 3254 35845
rect 3306 35793 3318 35845
rect 3374 35793 3386 35845
rect 3438 35793 3449 35845
rect 3505 35793 3518 35845
rect 3570 35793 3580 35845
rect 3636 35793 3650 35845
rect 3702 35793 3711 35845
rect 2848 35789 2924 35793
rect 2980 35789 3056 35793
rect 3112 35789 3187 35793
rect 3243 35789 3318 35793
rect 3374 35789 3449 35793
rect 3505 35789 3580 35793
rect 3636 35789 3711 35793
rect 3767 35789 3776 35845
rect 2783 35788 3776 35789
rect 148 35674 654 35680
rect 148 35622 454 35674
rect 506 35622 528 35674
rect 580 35622 602 35674
rect 148 35618 654 35622
rect 148 35562 298 35618
rect 354 35562 396 35618
rect 452 35610 494 35618
rect 550 35610 592 35618
rect 648 35610 654 35618
rect 452 35562 454 35610
rect 580 35562 592 35610
rect 148 35558 454 35562
rect 506 35558 528 35562
rect 580 35558 602 35562
rect 148 35546 654 35558
rect 148 35538 454 35546
rect 506 35538 528 35546
rect 580 35538 602 35546
rect 148 35482 298 35538
rect 354 35482 396 35538
rect 452 35494 454 35538
rect 580 35494 592 35538
rect 452 35482 494 35494
rect 550 35482 592 35494
rect 648 35482 654 35494
rect 148 35458 454 35482
rect 506 35458 528 35482
rect 580 35458 602 35482
rect 148 35402 298 35458
rect 354 35402 396 35458
rect 452 35430 454 35458
rect 580 35430 592 35458
rect 452 35418 494 35430
rect 550 35418 592 35430
rect 648 35418 654 35430
rect 452 35402 454 35418
rect 580 35402 592 35418
rect 148 35378 454 35402
rect 506 35378 528 35402
rect 580 35378 602 35402
rect 148 35322 298 35378
rect 354 35322 396 35378
rect 452 35366 454 35378
rect 580 35366 592 35378
rect 452 35354 494 35366
rect 550 35354 592 35366
rect 648 35354 654 35366
rect 452 35322 454 35354
rect 580 35322 592 35354
rect 148 35302 454 35322
rect 506 35302 528 35322
rect 580 35302 602 35322
rect 148 35298 654 35302
rect 148 35242 298 35298
rect 354 35242 396 35298
rect 452 35290 494 35298
rect 550 35290 592 35298
rect 648 35290 654 35298
rect 452 35242 454 35290
rect 580 35242 592 35290
rect 148 35238 454 35242
rect 506 35238 528 35242
rect 580 35238 602 35242
rect 148 35226 654 35238
rect 148 35218 454 35226
rect 506 35218 528 35226
rect 580 35218 602 35226
rect 148 35162 298 35218
rect 354 35162 396 35218
rect 452 35174 454 35218
rect 580 35174 592 35218
rect 452 35162 494 35174
rect 550 35162 592 35174
rect 648 35162 654 35174
rect 148 35138 454 35162
rect 506 35138 528 35162
rect 580 35138 602 35162
rect 148 35082 298 35138
rect 354 35082 396 35138
rect 452 35110 454 35138
rect 580 35110 592 35138
rect 452 35098 494 35110
rect 550 35098 592 35110
rect 648 35098 654 35110
rect 452 35082 454 35098
rect 580 35082 592 35098
rect 148 35058 454 35082
rect 506 35058 528 35082
rect 580 35058 602 35082
rect 148 35002 298 35058
rect 354 35002 396 35058
rect 452 35046 454 35058
rect 580 35046 592 35058
rect 452 35034 494 35046
rect 550 35034 592 35046
rect 648 35034 654 35046
rect 452 35002 454 35034
rect 580 35002 592 35034
rect 148 34982 454 35002
rect 506 34982 528 35002
rect 580 34982 602 35002
rect 148 34978 654 34982
rect 148 34922 298 34978
rect 354 34922 396 34978
rect 452 34970 494 34978
rect 550 34970 592 34978
rect 648 34970 654 34978
rect 452 34922 454 34970
rect 580 34922 592 34970
rect 148 34918 454 34922
rect 506 34918 528 34922
rect 580 34918 602 34922
rect 148 34906 654 34918
rect 148 34898 454 34906
rect 506 34898 528 34906
rect 580 34898 602 34906
rect 148 34842 298 34898
rect 354 34842 396 34898
rect 452 34854 454 34898
rect 580 34854 592 34898
rect 452 34842 494 34854
rect 550 34842 592 34854
rect 648 34842 654 34854
rect 148 34818 454 34842
rect 506 34818 528 34842
rect 580 34818 602 34842
rect 148 34762 298 34818
rect 354 34762 396 34818
rect 452 34790 454 34818
rect 580 34790 592 34818
rect 452 34778 494 34790
rect 550 34778 592 34790
rect 648 34778 654 34790
rect 452 34762 454 34778
rect 580 34762 592 34778
rect 148 34738 454 34762
rect 506 34738 528 34762
rect 580 34738 602 34762
rect 148 34682 298 34738
rect 354 34682 396 34738
rect 452 34726 454 34738
rect 580 34726 592 34738
rect 452 34714 494 34726
rect 550 34714 592 34726
rect 648 34714 654 34726
rect 452 34682 454 34714
rect 580 34682 592 34714
rect 148 34662 454 34682
rect 506 34662 528 34682
rect 580 34662 602 34682
rect 148 34658 654 34662
rect 148 34602 298 34658
rect 354 34602 396 34658
rect 452 34650 494 34658
rect 550 34650 592 34658
rect 648 34650 654 34658
rect 452 34602 454 34650
rect 580 34602 592 34650
rect 148 34598 454 34602
rect 506 34598 528 34602
rect 580 34598 602 34602
rect 148 34586 654 34598
rect 148 34578 454 34586
rect 506 34578 528 34586
rect 580 34578 602 34586
rect 148 34522 298 34578
rect 354 34522 396 34578
rect 452 34534 454 34578
rect 580 34534 592 34578
rect 452 34522 494 34534
rect 550 34522 592 34534
rect 648 34522 654 34534
rect 148 34498 454 34522
rect 506 34498 528 34522
rect 580 34498 602 34522
rect 148 34442 298 34498
rect 354 34442 396 34498
rect 452 34470 454 34498
rect 580 34470 592 34498
rect 452 34458 494 34470
rect 550 34458 592 34470
rect 648 34458 654 34470
rect 452 34442 454 34458
rect 580 34442 592 34458
rect 148 34418 454 34442
rect 506 34418 528 34442
rect 580 34418 602 34442
rect 148 34362 298 34418
rect 354 34362 396 34418
rect 452 34406 454 34418
rect 580 34406 592 34418
rect 452 34394 494 34406
rect 550 34394 592 34406
rect 648 34394 654 34406
rect 452 34362 454 34394
rect 580 34362 592 34394
rect 148 34342 454 34362
rect 506 34342 528 34362
rect 580 34342 602 34362
rect 148 34338 654 34342
rect 148 34282 298 34338
rect 354 34282 396 34338
rect 452 34330 494 34338
rect 550 34330 592 34338
rect 648 34330 654 34338
rect 452 34282 454 34330
rect 580 34282 592 34330
rect 148 34278 454 34282
rect 506 34278 528 34282
rect 580 34278 602 34282
rect 148 34266 654 34278
rect 148 34258 454 34266
rect 506 34258 528 34266
rect 580 34258 602 34266
rect 148 34202 298 34258
rect 354 34202 396 34258
rect 452 34214 454 34258
rect 580 34214 592 34258
rect 452 34202 494 34214
rect 550 34202 592 34214
rect 648 34202 654 34214
rect 148 34178 454 34202
rect 506 34178 528 34202
rect 580 34178 602 34202
rect 148 34122 298 34178
rect 354 34122 396 34178
rect 452 34150 454 34178
rect 580 34150 592 34178
rect 452 34138 494 34150
rect 550 34138 592 34150
rect 648 34138 654 34150
rect 452 34122 454 34138
rect 580 34122 592 34138
rect 148 34098 454 34122
rect 506 34098 528 34122
rect 580 34098 602 34122
rect 148 34042 298 34098
rect 354 34042 396 34098
rect 452 34086 454 34098
rect 580 34086 592 34098
rect 452 34074 494 34086
rect 550 34074 592 34086
rect 648 34074 654 34086
rect 452 34042 454 34074
rect 580 34042 592 34074
rect 148 34022 454 34042
rect 506 34022 528 34042
rect 580 34022 602 34042
rect 148 34018 654 34022
rect 148 34012 298 34018
rect 148 33960 149 34012
rect 201 33960 247 34012
rect 354 33962 396 34018
rect 452 34010 494 34018
rect 550 34010 592 34018
rect 648 34010 654 34018
rect 452 33962 454 34010
rect 580 33962 592 34010
rect 299 33960 454 33962
rect 148 33958 454 33960
rect 506 33958 528 33962
rect 580 33958 602 33962
rect 148 33948 654 33958
rect 148 33896 149 33948
rect 201 33896 247 33948
rect 299 33946 654 33948
rect 299 33938 454 33946
rect 506 33938 528 33946
rect 580 33938 602 33946
rect 148 33884 298 33896
rect 148 33832 149 33884
rect 201 33832 247 33884
rect 354 33882 396 33938
rect 452 33894 454 33938
rect 580 33894 592 33938
rect 452 33882 494 33894
rect 550 33882 592 33894
rect 648 33882 654 33894
rect 299 33858 454 33882
rect 506 33858 528 33882
rect 580 33858 602 33882
rect 148 33820 298 33832
rect 148 33768 149 33820
rect 201 33768 247 33820
rect 354 33802 396 33858
rect 452 33830 454 33858
rect 580 33830 592 33858
rect 452 33818 494 33830
rect 550 33818 592 33830
rect 648 33818 654 33830
rect 452 33802 454 33818
rect 580 33802 592 33818
rect 299 33778 454 33802
rect 506 33778 528 33802
rect 580 33778 602 33802
rect 148 33756 298 33768
rect 148 33704 149 33756
rect 201 33704 247 33756
rect 354 33722 396 33778
rect 452 33766 454 33778
rect 580 33766 592 33778
rect 452 33754 494 33766
rect 550 33754 592 33766
rect 648 33754 654 33766
rect 452 33722 454 33754
rect 580 33722 592 33754
rect 299 33704 454 33722
rect 148 33702 454 33704
rect 506 33702 528 33722
rect 580 33702 602 33722
rect 148 33698 654 33702
rect 148 33692 298 33698
rect 148 33640 149 33692
rect 201 33640 247 33692
rect 354 33642 396 33698
rect 452 33690 494 33698
rect 550 33690 592 33698
rect 648 33690 654 33698
rect 452 33642 454 33690
rect 580 33642 592 33690
rect 299 33640 454 33642
rect 148 33638 454 33640
rect 506 33638 528 33642
rect 580 33638 602 33642
rect 148 33628 654 33638
rect 148 33576 149 33628
rect 201 33576 247 33628
rect 299 33626 654 33628
rect 299 33618 454 33626
rect 506 33618 528 33626
rect 580 33618 602 33626
rect 148 33564 298 33576
rect 148 33512 149 33564
rect 201 33512 247 33564
rect 354 33562 396 33618
rect 452 33574 454 33618
rect 580 33574 592 33618
rect 452 33562 494 33574
rect 550 33562 592 33574
rect 648 33562 654 33574
rect 299 33538 454 33562
rect 506 33538 528 33562
rect 580 33538 602 33562
rect 148 33500 298 33512
rect 148 33448 149 33500
rect 201 33448 247 33500
rect 354 33482 396 33538
rect 452 33510 454 33538
rect 580 33510 592 33538
rect 452 33498 494 33510
rect 550 33498 592 33510
rect 648 33498 654 33510
rect 452 33482 454 33498
rect 580 33482 592 33498
rect 299 33458 454 33482
rect 506 33458 528 33482
rect 580 33458 602 33482
rect 148 33436 298 33448
rect 148 33384 149 33436
rect 201 33384 247 33436
rect 354 33402 396 33458
rect 452 33446 454 33458
rect 580 33446 592 33458
rect 452 33434 494 33446
rect 550 33434 592 33446
rect 648 33434 654 33446
rect 452 33402 454 33434
rect 580 33402 592 33434
rect 299 33384 454 33402
rect 148 33382 454 33384
rect 506 33382 528 33402
rect 580 33382 602 33402
rect 148 33378 654 33382
rect 148 33372 298 33378
rect 148 33320 149 33372
rect 201 33320 247 33372
rect 354 33322 396 33378
rect 452 33370 494 33378
rect 550 33370 592 33378
rect 648 33370 654 33378
rect 452 33322 454 33370
rect 580 33322 592 33370
rect 299 33320 454 33322
rect 148 33318 454 33320
rect 506 33318 528 33322
rect 580 33318 602 33322
rect 148 33308 654 33318
rect 148 33256 149 33308
rect 201 33256 247 33308
rect 299 33306 654 33308
rect 299 33298 454 33306
rect 506 33298 528 33306
rect 580 33298 602 33306
rect 148 33244 298 33256
rect 148 33192 149 33244
rect 201 33192 247 33244
rect 354 33242 396 33298
rect 452 33254 454 33298
rect 580 33254 592 33298
rect 452 33242 494 33254
rect 550 33242 592 33254
rect 648 33242 654 33254
rect 299 33218 454 33242
rect 506 33218 528 33242
rect 580 33218 602 33242
rect 148 33180 298 33192
rect 148 33128 149 33180
rect 201 33128 247 33180
rect 354 33162 396 33218
rect 452 33190 454 33218
rect 580 33190 592 33218
rect 452 33178 494 33190
rect 550 33178 592 33190
rect 648 33178 654 33190
rect 452 33162 454 33178
rect 580 33162 592 33178
rect 299 33138 454 33162
rect 506 33138 528 33162
rect 580 33138 602 33162
rect 148 33116 298 33128
rect 148 33064 149 33116
rect 201 33064 247 33116
rect 354 33082 396 33138
rect 452 33126 454 33138
rect 580 33126 592 33138
rect 452 33114 494 33126
rect 550 33114 592 33126
rect 648 33114 654 33126
rect 452 33082 454 33114
rect 580 33082 592 33114
rect 299 33064 454 33082
rect 148 33062 454 33064
rect 506 33062 528 33082
rect 580 33062 602 33082
rect 148 33058 654 33062
rect 148 33052 298 33058
rect 148 33000 149 33052
rect 201 33000 247 33052
rect 354 33002 396 33058
rect 452 33050 494 33058
rect 550 33050 592 33058
rect 648 33050 654 33058
rect 452 33002 454 33050
rect 580 33002 592 33050
rect 299 33000 454 33002
rect 148 32998 454 33000
rect 506 32998 528 33002
rect 580 32998 602 33002
rect 148 32988 654 32998
rect 148 32936 149 32988
rect 201 32936 247 32988
rect 299 32986 654 32988
rect 299 32978 454 32986
rect 506 32978 528 32986
rect 580 32978 602 32986
rect 148 32924 298 32936
rect 148 32872 149 32924
rect 201 32872 247 32924
rect 354 32922 396 32978
rect 452 32934 454 32978
rect 580 32934 592 32978
rect 452 32922 494 32934
rect 550 32922 592 32934
rect 648 32922 654 32934
rect 299 32898 454 32922
rect 506 32898 528 32922
rect 580 32898 602 32922
rect 148 32859 298 32872
rect 148 32807 149 32859
rect 201 32807 247 32859
rect 354 32842 396 32898
rect 452 32870 454 32898
rect 580 32870 592 32898
rect 452 32858 494 32870
rect 550 32858 592 32870
rect 648 32858 654 32870
rect 452 32842 454 32858
rect 580 32842 592 32858
rect 299 32818 454 32842
rect 506 32818 528 32842
rect 580 32818 602 32842
rect 148 32794 298 32807
rect 148 32742 149 32794
rect 201 32742 247 32794
rect 354 32762 396 32818
rect 452 32806 454 32818
rect 580 32806 592 32818
rect 452 32794 494 32806
rect 550 32794 592 32806
rect 648 32794 654 32806
rect 452 32762 454 32794
rect 580 32762 592 32794
rect 299 32742 454 32762
rect 506 32742 528 32762
rect 580 32742 602 32762
rect 148 32738 654 32742
rect 148 32729 298 32738
rect 148 32677 149 32729
rect 201 32677 247 32729
rect 354 32682 396 32738
rect 452 32729 494 32738
rect 550 32729 592 32738
rect 648 32729 654 32738
rect 452 32682 454 32729
rect 580 32682 592 32729
rect 299 32677 454 32682
rect 506 32677 528 32682
rect 580 32677 602 32682
rect 148 32664 654 32677
rect 148 32612 149 32664
rect 201 32612 247 32664
rect 299 32658 454 32664
rect 506 32658 528 32664
rect 580 32658 602 32664
rect 148 32602 298 32612
rect 354 32602 396 32658
rect 452 32612 454 32658
rect 580 32612 592 32658
rect 452 32602 494 32612
rect 550 32602 592 32612
rect 648 32602 654 32612
rect 148 32599 654 32602
rect 148 32547 149 32599
rect 201 32547 247 32599
rect 299 32578 454 32599
rect 506 32578 528 32599
rect 580 32578 602 32599
rect 148 32534 298 32547
rect 148 32482 149 32534
rect 201 32482 247 32534
rect 354 32522 396 32578
rect 452 32547 454 32578
rect 580 32547 592 32578
rect 452 32534 494 32547
rect 550 32534 592 32547
rect 648 32534 654 32547
rect 452 32522 454 32534
rect 580 32522 592 32534
rect 299 32498 454 32522
rect 506 32498 528 32522
rect 580 32498 602 32522
rect 148 32469 298 32482
rect 148 32417 149 32469
rect 201 32417 247 32469
rect 354 32442 396 32498
rect 452 32482 454 32498
rect 580 32482 592 32498
rect 452 32469 494 32482
rect 550 32469 592 32482
rect 648 32469 654 32482
rect 452 32442 454 32469
rect 580 32442 592 32469
rect 299 32418 454 32442
rect 506 32418 528 32442
rect 580 32418 602 32442
rect 148 32404 298 32417
rect 148 32352 149 32404
rect 201 32352 247 32404
rect 354 32362 396 32418
rect 452 32417 454 32418
rect 580 32417 592 32418
rect 452 32404 494 32417
rect 550 32404 592 32417
rect 648 32404 654 32417
rect 452 32362 454 32404
rect 580 32362 592 32404
rect 299 32352 454 32362
rect 506 32352 528 32362
rect 580 32352 602 32362
rect 148 32339 654 32352
rect 148 32287 149 32339
rect 201 32287 247 32339
rect 299 32338 454 32339
rect 506 32338 528 32339
rect 580 32338 602 32339
rect 148 32282 298 32287
rect 354 32282 396 32338
rect 452 32287 454 32338
rect 580 32287 592 32338
rect 452 32282 494 32287
rect 550 32282 592 32287
rect 648 32282 654 32287
rect 148 32274 654 32282
rect 148 32222 149 32274
rect 201 32222 247 32274
rect 299 32258 454 32274
rect 506 32258 528 32274
rect 580 32258 602 32274
rect 148 32209 298 32222
rect 148 32157 149 32209
rect 201 32157 247 32209
rect 354 32202 396 32258
rect 452 32222 454 32258
rect 580 32222 592 32258
rect 452 32209 494 32222
rect 550 32209 592 32222
rect 648 32209 654 32222
rect 452 32202 454 32209
rect 580 32202 592 32209
rect 299 32177 454 32202
rect 506 32177 528 32202
rect 580 32177 602 32202
rect 148 32144 298 32157
rect 148 32092 149 32144
rect 201 32092 247 32144
rect 354 32121 396 32177
rect 452 32157 454 32177
rect 580 32157 592 32177
rect 452 32144 494 32157
rect 550 32144 592 32157
rect 648 32144 654 32157
rect 452 32121 454 32144
rect 580 32121 592 32144
rect 299 32096 454 32121
rect 506 32096 528 32121
rect 580 32096 602 32121
rect 148 32079 298 32092
rect 148 32027 149 32079
rect 201 32027 247 32079
rect 354 32040 396 32096
rect 452 32092 454 32096
rect 580 32092 592 32096
rect 452 32079 494 32092
rect 550 32079 592 32092
rect 648 32079 654 32092
rect 452 32040 454 32079
rect 580 32040 592 32079
rect 299 32027 454 32040
rect 506 32027 528 32040
rect 580 32027 602 32040
rect 148 32015 654 32027
rect 148 32014 298 32015
rect 148 31962 149 32014
rect 201 31962 247 32014
rect 148 31959 298 31962
rect 354 31959 396 32015
rect 452 32014 494 32015
rect 550 32014 592 32015
rect 648 32014 654 32015
rect 452 31962 454 32014
rect 580 31962 592 32014
rect 452 31959 494 31962
rect 550 31959 592 31962
rect 648 31959 654 31962
rect 148 31949 654 31959
rect 148 31897 149 31949
rect 201 31897 247 31949
rect 299 31934 454 31949
rect 506 31934 528 31949
rect 580 31934 602 31949
rect 148 31884 298 31897
rect 148 31832 149 31884
rect 201 31832 247 31884
rect 354 31878 396 31934
rect 452 31897 454 31934
rect 580 31897 592 31934
rect 452 31884 494 31897
rect 550 31884 592 31897
rect 648 31884 654 31897
rect 452 31878 454 31884
rect 580 31878 592 31884
rect 299 31853 454 31878
rect 506 31853 528 31878
rect 580 31853 602 31878
rect 148 31819 298 31832
rect 148 31767 149 31819
rect 201 31767 247 31819
rect 354 31797 396 31853
rect 452 31832 454 31853
rect 580 31832 592 31853
rect 452 31819 494 31832
rect 550 31819 592 31832
rect 648 31819 654 31832
rect 452 31797 454 31819
rect 580 31797 592 31819
rect 299 31772 454 31797
rect 506 31772 528 31797
rect 580 31772 602 31797
rect 148 31754 298 31767
rect 148 31702 149 31754
rect 201 31702 247 31754
rect 354 31716 396 31772
rect 452 31767 454 31772
rect 580 31767 592 31772
rect 452 31754 494 31767
rect 550 31754 592 31767
rect 648 31754 654 31767
rect 452 31716 454 31754
rect 580 31716 592 31754
rect 299 31702 454 31716
rect 506 31702 528 31716
rect 580 31702 602 31716
rect 148 31691 654 31702
rect 148 31689 298 31691
rect 148 31637 149 31689
rect 201 31637 247 31689
rect 148 31635 298 31637
rect 354 31635 396 31691
rect 452 31689 494 31691
rect 550 31689 592 31691
rect 648 31689 654 31691
rect 452 31637 454 31689
rect 580 31637 592 31689
rect 452 31635 494 31637
rect 550 31635 592 31637
rect 648 31635 654 31637
rect 148 31624 654 31635
rect 148 31572 149 31624
rect 201 31572 247 31624
rect 299 31610 454 31624
rect 506 31610 528 31624
rect 580 31610 602 31624
rect 148 31559 298 31572
rect 148 31507 149 31559
rect 201 31507 247 31559
rect 354 31554 396 31610
rect 452 31572 454 31610
rect 580 31572 592 31610
rect 452 31559 494 31572
rect 550 31559 592 31572
rect 648 31559 654 31572
rect 452 31554 454 31559
rect 580 31554 592 31559
rect 299 31529 454 31554
rect 506 31529 528 31554
rect 580 31529 602 31554
rect 148 31494 298 31507
rect 148 31442 149 31494
rect 201 31442 247 31494
rect 354 31473 396 31529
rect 452 31507 454 31529
rect 580 31507 592 31529
rect 452 31494 494 31507
rect 550 31494 592 31507
rect 648 31494 654 31507
rect 452 31473 454 31494
rect 580 31473 592 31494
rect 5103 32613 6298 32619
rect 5103 32557 5112 32613
rect 5168 32557 5193 32613
rect 5249 32557 5273 32613
rect 5329 32557 5353 32613
rect 5409 32557 5433 32613
rect 5489 32557 5513 32613
rect 5569 32557 5593 32613
rect 5649 32557 5673 32613
rect 5729 32557 5753 32613
rect 5809 32557 5833 32613
rect 5889 32557 5913 32613
rect 5969 32557 5993 32613
rect 6049 32557 6073 32613
rect 6129 32557 6153 32613
rect 6209 32557 6233 32613
rect 6289 32557 6298 32613
rect 5103 32531 6298 32557
rect 5103 32475 5112 32531
rect 5168 32475 5193 32531
rect 5249 32475 5273 32531
rect 5329 32475 5353 32531
rect 5409 32475 5433 32531
rect 5489 32475 5513 32531
rect 5569 32475 5593 32531
rect 5649 32475 5673 32531
rect 5729 32475 5753 32531
rect 5809 32475 5833 32531
rect 5889 32475 5913 32531
rect 5969 32475 5993 32531
rect 6049 32475 6073 32531
rect 6129 32475 6153 32531
rect 6209 32475 6233 32531
rect 6289 32475 6298 32531
rect 5103 32449 6298 32475
rect 5103 32393 5112 32449
rect 5168 32393 5193 32449
rect 5249 32393 5273 32449
rect 5329 32393 5353 32449
rect 5409 32393 5433 32449
rect 5489 32393 5513 32449
rect 5569 32393 5593 32449
rect 5649 32393 5673 32449
rect 5729 32393 5753 32449
rect 5809 32393 5833 32449
rect 5889 32393 5913 32449
rect 5969 32393 5993 32449
rect 6049 32393 6073 32449
rect 6129 32393 6153 32449
rect 6209 32393 6233 32449
rect 6289 32393 6298 32449
rect 5103 32367 6298 32393
rect 5103 32311 5112 32367
rect 5168 32311 5193 32367
rect 5249 32311 5273 32367
rect 5329 32311 5353 32367
rect 5409 32311 5433 32367
rect 5489 32311 5513 32367
rect 5569 32311 5593 32367
rect 5649 32311 5673 32367
rect 5729 32311 5753 32367
rect 5809 32311 5833 32367
rect 5889 32311 5913 32367
rect 5969 32311 5993 32367
rect 6049 32311 6073 32367
rect 6129 32311 6153 32367
rect 6209 32311 6233 32367
rect 6289 32311 6298 32367
rect 5103 32285 6298 32311
rect 5103 32229 5112 32285
rect 5168 32229 5193 32285
rect 5249 32229 5273 32285
rect 5329 32229 5353 32285
rect 5409 32229 5433 32285
rect 5489 32229 5513 32285
rect 5569 32229 5593 32285
rect 5649 32229 5673 32285
rect 5729 32229 5753 32285
rect 5809 32229 5833 32285
rect 5889 32229 5913 32285
rect 5969 32229 5993 32285
rect 6049 32229 6073 32285
rect 6129 32229 6153 32285
rect 6209 32229 6233 32285
rect 6289 32229 6298 32285
rect 5103 32203 6298 32229
rect 5103 32147 5112 32203
rect 5168 32147 5193 32203
rect 5249 32147 5273 32203
rect 5329 32147 5353 32203
rect 5409 32147 5433 32203
rect 5489 32147 5513 32203
rect 5569 32147 5593 32203
rect 5649 32147 5673 32203
rect 5729 32147 5753 32203
rect 5809 32147 5833 32203
rect 5889 32147 5913 32203
rect 5969 32147 5993 32203
rect 6049 32147 6073 32203
rect 6129 32147 6153 32203
rect 6209 32147 6233 32203
rect 6289 32147 6298 32203
rect 5103 32121 6298 32147
rect 5103 32065 5112 32121
rect 5168 32065 5193 32121
rect 5249 32065 5273 32121
rect 5329 32065 5353 32121
rect 5409 32065 5433 32121
rect 5489 32065 5513 32121
rect 5569 32065 5593 32121
rect 5649 32065 5673 32121
rect 5729 32065 5753 32121
rect 5809 32065 5833 32121
rect 5889 32065 5913 32121
rect 5969 32065 5993 32121
rect 6049 32065 6073 32121
rect 6129 32065 6153 32121
rect 6209 32065 6233 32121
rect 6289 32065 6298 32121
rect 5103 32039 6298 32065
rect 5103 31983 5112 32039
rect 5168 31983 5193 32039
rect 5249 31983 5273 32039
rect 5329 31983 5353 32039
rect 5409 31983 5433 32039
rect 5489 31983 5513 32039
rect 5569 31983 5593 32039
rect 5649 31983 5673 32039
rect 5729 31983 5753 32039
rect 5809 31983 5833 32039
rect 5889 31983 5913 32039
rect 5969 31983 5993 32039
rect 6049 31983 6073 32039
rect 6129 31983 6153 32039
rect 6209 31983 6233 32039
rect 6289 31983 6298 32039
rect 5103 31957 6298 31983
rect 5103 31901 5112 31957
rect 5168 31901 5193 31957
rect 5249 31901 5273 31957
rect 5329 31901 5353 31957
rect 5409 31901 5433 31957
rect 5489 31901 5513 31957
rect 5569 31901 5593 31957
rect 5649 31901 5673 31957
rect 5729 31901 5753 31957
rect 5809 31901 5833 31957
rect 5889 31901 5913 31957
rect 5969 31901 5993 31957
rect 6049 31901 6073 31957
rect 6129 31901 6153 31957
rect 6209 31901 6233 31957
rect 6289 31901 6298 31957
rect 5103 31875 6298 31901
rect 5103 31819 5112 31875
rect 5168 31819 5193 31875
rect 5249 31819 5273 31875
rect 5329 31819 5353 31875
rect 5409 31819 5433 31875
rect 5489 31819 5513 31875
rect 5569 31819 5593 31875
rect 5649 31819 5673 31875
rect 5729 31819 5753 31875
rect 5809 31819 5833 31875
rect 5889 31819 5913 31875
rect 5969 31819 5993 31875
rect 6049 31819 6073 31875
rect 6129 31819 6153 31875
rect 6209 31819 6233 31875
rect 6289 31819 6298 31875
rect 5103 31793 6298 31819
rect 5103 31737 5112 31793
rect 5168 31737 5193 31793
rect 5249 31737 5273 31793
rect 5329 31737 5353 31793
rect 5409 31737 5433 31793
rect 5489 31737 5513 31793
rect 5569 31737 5593 31793
rect 5649 31737 5673 31793
rect 5729 31737 5753 31793
rect 5809 31737 5833 31793
rect 5889 31737 5913 31793
rect 5969 31737 5993 31793
rect 6049 31737 6073 31793
rect 6129 31737 6153 31793
rect 6209 31737 6233 31793
rect 6289 31737 6298 31793
rect 5103 31711 6298 31737
rect 5103 31655 5112 31711
rect 5168 31655 5193 31711
rect 5249 31655 5273 31711
rect 5329 31655 5353 31711
rect 5409 31655 5433 31711
rect 5489 31655 5513 31711
rect 5569 31655 5593 31711
rect 5649 31655 5673 31711
rect 5729 31655 5753 31711
rect 5809 31655 5833 31711
rect 5889 31655 5913 31711
rect 5969 31655 5993 31711
rect 6049 31655 6073 31711
rect 6129 31655 6153 31711
rect 6209 31655 6233 31711
rect 6289 31655 6298 31711
rect 5103 31629 6298 31655
rect 5103 31573 5112 31629
rect 5168 31573 5193 31629
rect 5249 31573 5273 31629
rect 5329 31573 5353 31629
rect 5409 31573 5433 31629
rect 5489 31573 5513 31629
rect 5569 31573 5593 31629
rect 5649 31573 5673 31629
rect 5729 31573 5753 31629
rect 5809 31573 5833 31629
rect 5889 31573 5913 31629
rect 5969 31573 5993 31629
rect 6049 31573 6073 31629
rect 6129 31573 6153 31629
rect 6209 31573 6233 31629
rect 6289 31573 6298 31629
rect 5103 31547 6298 31573
rect 5103 31491 5112 31547
rect 5168 31491 5193 31547
rect 5249 31491 5273 31547
rect 5329 31491 5353 31547
rect 5409 31491 5433 31547
rect 5489 31491 5513 31547
rect 5569 31491 5593 31547
rect 5649 31491 5673 31547
rect 5729 31491 5753 31547
rect 5809 31491 5833 31547
rect 5889 31491 5913 31547
rect 5969 31491 5993 31547
rect 6049 31491 6073 31547
rect 6129 31491 6153 31547
rect 6209 31491 6233 31547
rect 6289 31491 6298 31547
rect 5103 31485 6298 31491
rect 6601 32613 7799 32619
rect 6601 32557 6610 32613
rect 6666 32557 6691 32613
rect 6747 32557 6772 32613
rect 6828 32557 6853 32613
rect 6909 32557 6934 32613
rect 6990 32557 7014 32613
rect 7070 32557 7094 32613
rect 7150 32557 7174 32613
rect 7230 32557 7254 32613
rect 7310 32557 7334 32613
rect 7390 32557 7414 32613
rect 7470 32557 7494 32613
rect 7550 32557 7574 32613
rect 7630 32557 7654 32613
rect 7710 32557 7734 32613
rect 7790 32557 7799 32613
rect 6601 32531 7799 32557
rect 6601 32475 6610 32531
rect 6666 32475 6691 32531
rect 6747 32475 6772 32531
rect 6828 32475 6853 32531
rect 6909 32475 6934 32531
rect 6990 32475 7014 32531
rect 7070 32475 7094 32531
rect 7150 32475 7174 32531
rect 7230 32475 7254 32531
rect 7310 32475 7334 32531
rect 7390 32475 7414 32531
rect 7470 32475 7494 32531
rect 7550 32475 7574 32531
rect 7630 32475 7654 32531
rect 7710 32475 7734 32531
rect 7790 32475 7799 32531
rect 6601 32449 7799 32475
rect 6601 32393 6610 32449
rect 6666 32393 6691 32449
rect 6747 32393 6772 32449
rect 6828 32393 6853 32449
rect 6909 32393 6934 32449
rect 6990 32393 7014 32449
rect 7070 32393 7094 32449
rect 7150 32393 7174 32449
rect 7230 32393 7254 32449
rect 7310 32393 7334 32449
rect 7390 32393 7414 32449
rect 7470 32393 7494 32449
rect 7550 32393 7574 32449
rect 7630 32393 7654 32449
rect 7710 32393 7734 32449
rect 7790 32393 7799 32449
rect 6601 32367 7799 32393
rect 6601 32311 6610 32367
rect 6666 32311 6691 32367
rect 6747 32311 6772 32367
rect 6828 32311 6853 32367
rect 6909 32311 6934 32367
rect 6990 32311 7014 32367
rect 7070 32311 7094 32367
rect 7150 32311 7174 32367
rect 7230 32311 7254 32367
rect 7310 32311 7334 32367
rect 7390 32311 7414 32367
rect 7470 32311 7494 32367
rect 7550 32311 7574 32367
rect 7630 32311 7654 32367
rect 7710 32311 7734 32367
rect 7790 32311 7799 32367
rect 6601 32285 7799 32311
rect 6601 32229 6610 32285
rect 6666 32229 6691 32285
rect 6747 32229 6772 32285
rect 6828 32229 6853 32285
rect 6909 32229 6934 32285
rect 6990 32229 7014 32285
rect 7070 32229 7094 32285
rect 7150 32229 7174 32285
rect 7230 32229 7254 32285
rect 7310 32229 7334 32285
rect 7390 32229 7414 32285
rect 7470 32229 7494 32285
rect 7550 32229 7574 32285
rect 7630 32229 7654 32285
rect 7710 32229 7734 32285
rect 7790 32229 7799 32285
rect 6601 32203 7799 32229
rect 6601 32147 6610 32203
rect 6666 32147 6691 32203
rect 6747 32147 6772 32203
rect 6828 32147 6853 32203
rect 6909 32147 6934 32203
rect 6990 32147 7014 32203
rect 7070 32147 7094 32203
rect 7150 32147 7174 32203
rect 7230 32147 7254 32203
rect 7310 32147 7334 32203
rect 7390 32147 7414 32203
rect 7470 32147 7494 32203
rect 7550 32147 7574 32203
rect 7630 32147 7654 32203
rect 7710 32147 7734 32203
rect 7790 32147 7799 32203
rect 6601 32121 7799 32147
rect 6601 32065 6610 32121
rect 6666 32065 6691 32121
rect 6747 32065 6772 32121
rect 6828 32065 6853 32121
rect 6909 32065 6934 32121
rect 6990 32065 7014 32121
rect 7070 32065 7094 32121
rect 7150 32065 7174 32121
rect 7230 32065 7254 32121
rect 7310 32065 7334 32121
rect 7390 32065 7414 32121
rect 7470 32065 7494 32121
rect 7550 32065 7574 32121
rect 7630 32065 7654 32121
rect 7710 32065 7734 32121
rect 7790 32065 7799 32121
rect 6601 32039 7799 32065
rect 6601 31983 6610 32039
rect 6666 31983 6691 32039
rect 6747 31983 6772 32039
rect 6828 31983 6853 32039
rect 6909 31983 6934 32039
rect 6990 31983 7014 32039
rect 7070 31983 7094 32039
rect 7150 31983 7174 32039
rect 7230 31983 7254 32039
rect 7310 31983 7334 32039
rect 7390 31983 7414 32039
rect 7470 31983 7494 32039
rect 7550 31983 7574 32039
rect 7630 31983 7654 32039
rect 7710 31983 7734 32039
rect 7790 31983 7799 32039
rect 6601 31957 7799 31983
rect 6601 31901 6610 31957
rect 6666 31901 6691 31957
rect 6747 31901 6772 31957
rect 6828 31901 6853 31957
rect 6909 31901 6934 31957
rect 6990 31901 7014 31957
rect 7070 31901 7094 31957
rect 7150 31901 7174 31957
rect 7230 31901 7254 31957
rect 7310 31901 7334 31957
rect 7390 31901 7414 31957
rect 7470 31901 7494 31957
rect 7550 31901 7574 31957
rect 7630 31901 7654 31957
rect 7710 31901 7734 31957
rect 7790 31901 7799 31957
rect 6601 31875 7799 31901
rect 6601 31819 6610 31875
rect 6666 31819 6691 31875
rect 6747 31819 6772 31875
rect 6828 31819 6853 31875
rect 6909 31819 6934 31875
rect 6990 31819 7014 31875
rect 7070 31819 7094 31875
rect 7150 31819 7174 31875
rect 7230 31819 7254 31875
rect 7310 31819 7334 31875
rect 7390 31819 7414 31875
rect 7470 31819 7494 31875
rect 7550 31819 7574 31875
rect 7630 31819 7654 31875
rect 7710 31819 7734 31875
rect 7790 31819 7799 31875
rect 6601 31793 7799 31819
rect 6601 31737 6610 31793
rect 6666 31737 6691 31793
rect 6747 31737 6772 31793
rect 6828 31737 6853 31793
rect 6909 31737 6934 31793
rect 6990 31737 7014 31793
rect 7070 31737 7094 31793
rect 7150 31737 7174 31793
rect 7230 31737 7254 31793
rect 7310 31737 7334 31793
rect 7390 31737 7414 31793
rect 7470 31737 7494 31793
rect 7550 31737 7574 31793
rect 7630 31737 7654 31793
rect 7710 31737 7734 31793
rect 7790 31737 7799 31793
rect 6601 31711 7799 31737
rect 6601 31655 6610 31711
rect 6666 31655 6691 31711
rect 6747 31655 6772 31711
rect 6828 31655 6853 31711
rect 6909 31655 6934 31711
rect 6990 31655 7014 31711
rect 7070 31655 7094 31711
rect 7150 31655 7174 31711
rect 7230 31655 7254 31711
rect 7310 31655 7334 31711
rect 7390 31655 7414 31711
rect 7470 31655 7494 31711
rect 7550 31655 7574 31711
rect 7630 31655 7654 31711
rect 7710 31655 7734 31711
rect 7790 31655 7799 31711
rect 6601 31629 7799 31655
rect 6601 31573 6610 31629
rect 6666 31573 6691 31629
rect 6747 31573 6772 31629
rect 6828 31573 6853 31629
rect 6909 31573 6934 31629
rect 6990 31573 7014 31629
rect 7070 31573 7094 31629
rect 7150 31573 7174 31629
rect 7230 31573 7254 31629
rect 7310 31573 7334 31629
rect 7390 31573 7414 31629
rect 7470 31573 7494 31629
rect 7550 31573 7574 31629
rect 7630 31573 7654 31629
rect 7710 31573 7734 31629
rect 7790 31573 7799 31629
rect 6601 31547 7799 31573
rect 6601 31491 6610 31547
rect 6666 31491 6691 31547
rect 6747 31491 6772 31547
rect 6828 31491 6853 31547
rect 6909 31491 6934 31547
rect 6990 31491 7014 31547
rect 7070 31491 7094 31547
rect 7150 31491 7174 31547
rect 7230 31491 7254 31547
rect 7310 31491 7334 31547
rect 7390 31491 7414 31547
rect 7470 31491 7494 31547
rect 7550 31491 7574 31547
rect 7630 31491 7654 31547
rect 7710 31491 7734 31547
rect 7790 31491 7799 31547
rect 6601 31485 7799 31491
rect 8098 32613 9296 32619
rect 8098 32557 8107 32613
rect 8163 32557 8188 32613
rect 8244 32557 8269 32613
rect 8325 32557 8350 32613
rect 8406 32557 8431 32613
rect 8487 32557 8511 32613
rect 8567 32557 8591 32613
rect 8647 32557 8671 32613
rect 8727 32557 8751 32613
rect 8807 32557 8831 32613
rect 8887 32557 8911 32613
rect 8967 32557 8991 32613
rect 9047 32557 9071 32613
rect 9127 32557 9151 32613
rect 9207 32557 9231 32613
rect 9287 32557 9296 32613
rect 8098 32531 9296 32557
rect 8098 32475 8107 32531
rect 8163 32475 8188 32531
rect 8244 32475 8269 32531
rect 8325 32475 8350 32531
rect 8406 32475 8431 32531
rect 8487 32475 8511 32531
rect 8567 32475 8591 32531
rect 8647 32475 8671 32531
rect 8727 32475 8751 32531
rect 8807 32475 8831 32531
rect 8887 32475 8911 32531
rect 8967 32475 8991 32531
rect 9047 32475 9071 32531
rect 9127 32475 9151 32531
rect 9207 32475 9231 32531
rect 9287 32475 9296 32531
rect 8098 32449 9296 32475
rect 8098 32393 8107 32449
rect 8163 32393 8188 32449
rect 8244 32393 8269 32449
rect 8325 32393 8350 32449
rect 8406 32393 8431 32449
rect 8487 32393 8511 32449
rect 8567 32393 8591 32449
rect 8647 32393 8671 32449
rect 8727 32393 8751 32449
rect 8807 32393 8831 32449
rect 8887 32393 8911 32449
rect 8967 32393 8991 32449
rect 9047 32393 9071 32449
rect 9127 32393 9151 32449
rect 9207 32393 9231 32449
rect 9287 32393 9296 32449
rect 8098 32367 9296 32393
rect 8098 32311 8107 32367
rect 8163 32311 8188 32367
rect 8244 32311 8269 32367
rect 8325 32311 8350 32367
rect 8406 32311 8431 32367
rect 8487 32311 8511 32367
rect 8567 32311 8591 32367
rect 8647 32311 8671 32367
rect 8727 32311 8751 32367
rect 8807 32311 8831 32367
rect 8887 32311 8911 32367
rect 8967 32311 8991 32367
rect 9047 32311 9071 32367
rect 9127 32311 9151 32367
rect 9207 32311 9231 32367
rect 9287 32311 9296 32367
rect 8098 32285 9296 32311
rect 8098 32229 8107 32285
rect 8163 32229 8188 32285
rect 8244 32229 8269 32285
rect 8325 32229 8350 32285
rect 8406 32229 8431 32285
rect 8487 32229 8511 32285
rect 8567 32229 8591 32285
rect 8647 32229 8671 32285
rect 8727 32229 8751 32285
rect 8807 32229 8831 32285
rect 8887 32229 8911 32285
rect 8967 32229 8991 32285
rect 9047 32229 9071 32285
rect 9127 32229 9151 32285
rect 9207 32229 9231 32285
rect 9287 32229 9296 32285
rect 8098 32203 9296 32229
rect 8098 32147 8107 32203
rect 8163 32147 8188 32203
rect 8244 32147 8269 32203
rect 8325 32147 8350 32203
rect 8406 32147 8431 32203
rect 8487 32147 8511 32203
rect 8567 32147 8591 32203
rect 8647 32147 8671 32203
rect 8727 32147 8751 32203
rect 8807 32147 8831 32203
rect 8887 32147 8911 32203
rect 8967 32147 8991 32203
rect 9047 32147 9071 32203
rect 9127 32147 9151 32203
rect 9207 32147 9231 32203
rect 9287 32147 9296 32203
rect 8098 32121 9296 32147
rect 8098 32065 8107 32121
rect 8163 32065 8188 32121
rect 8244 32065 8269 32121
rect 8325 32065 8350 32121
rect 8406 32065 8431 32121
rect 8487 32065 8511 32121
rect 8567 32065 8591 32121
rect 8647 32065 8671 32121
rect 8727 32065 8751 32121
rect 8807 32065 8831 32121
rect 8887 32065 8911 32121
rect 8967 32065 8991 32121
rect 9047 32065 9071 32121
rect 9127 32065 9151 32121
rect 9207 32065 9231 32121
rect 9287 32065 9296 32121
rect 8098 32039 9296 32065
rect 8098 31983 8107 32039
rect 8163 31983 8188 32039
rect 8244 31983 8269 32039
rect 8325 31983 8350 32039
rect 8406 31983 8431 32039
rect 8487 31983 8511 32039
rect 8567 31983 8591 32039
rect 8647 31983 8671 32039
rect 8727 31983 8751 32039
rect 8807 31983 8831 32039
rect 8887 31983 8911 32039
rect 8967 31983 8991 32039
rect 9047 31983 9071 32039
rect 9127 31983 9151 32039
rect 9207 31983 9231 32039
rect 9287 31983 9296 32039
rect 8098 31957 9296 31983
rect 8098 31901 8107 31957
rect 8163 31901 8188 31957
rect 8244 31901 8269 31957
rect 8325 31901 8350 31957
rect 8406 31901 8431 31957
rect 8487 31901 8511 31957
rect 8567 31901 8591 31957
rect 8647 31901 8671 31957
rect 8727 31901 8751 31957
rect 8807 31901 8831 31957
rect 8887 31901 8911 31957
rect 8967 31901 8991 31957
rect 9047 31901 9071 31957
rect 9127 31901 9151 31957
rect 9207 31901 9231 31957
rect 9287 31901 9296 31957
rect 8098 31875 9296 31901
rect 8098 31819 8107 31875
rect 8163 31819 8188 31875
rect 8244 31819 8269 31875
rect 8325 31819 8350 31875
rect 8406 31819 8431 31875
rect 8487 31819 8511 31875
rect 8567 31819 8591 31875
rect 8647 31819 8671 31875
rect 8727 31819 8751 31875
rect 8807 31819 8831 31875
rect 8887 31819 8911 31875
rect 8967 31819 8991 31875
rect 9047 31819 9071 31875
rect 9127 31819 9151 31875
rect 9207 31819 9231 31875
rect 9287 31819 9296 31875
rect 8098 31793 9296 31819
rect 8098 31737 8107 31793
rect 8163 31737 8188 31793
rect 8244 31737 8269 31793
rect 8325 31737 8350 31793
rect 8406 31737 8431 31793
rect 8487 31737 8511 31793
rect 8567 31737 8591 31793
rect 8647 31737 8671 31793
rect 8727 31737 8751 31793
rect 8807 31737 8831 31793
rect 8887 31737 8911 31793
rect 8967 31737 8991 31793
rect 9047 31737 9071 31793
rect 9127 31737 9151 31793
rect 9207 31737 9231 31793
rect 9287 31737 9296 31793
rect 8098 31711 9296 31737
rect 8098 31655 8107 31711
rect 8163 31655 8188 31711
rect 8244 31655 8269 31711
rect 8325 31655 8350 31711
rect 8406 31655 8431 31711
rect 8487 31655 8511 31711
rect 8567 31655 8591 31711
rect 8647 31655 8671 31711
rect 8727 31655 8751 31711
rect 8807 31655 8831 31711
rect 8887 31655 8911 31711
rect 8967 31655 8991 31711
rect 9047 31655 9071 31711
rect 9127 31655 9151 31711
rect 9207 31655 9231 31711
rect 9287 31655 9296 31711
rect 8098 31629 9296 31655
rect 8098 31573 8107 31629
rect 8163 31573 8188 31629
rect 8244 31573 8269 31629
rect 8325 31573 8350 31629
rect 8406 31573 8431 31629
rect 8487 31573 8511 31629
rect 8567 31573 8591 31629
rect 8647 31573 8671 31629
rect 8727 31573 8751 31629
rect 8807 31573 8831 31629
rect 8887 31573 8911 31629
rect 8967 31573 8991 31629
rect 9047 31573 9071 31629
rect 9127 31573 9151 31629
rect 9207 31573 9231 31629
rect 9287 31573 9296 31629
rect 8098 31547 9296 31573
rect 8098 31491 8107 31547
rect 8163 31491 8188 31547
rect 8244 31491 8269 31547
rect 8325 31491 8350 31547
rect 8406 31491 8431 31547
rect 8487 31491 8511 31547
rect 8567 31491 8591 31547
rect 8647 31491 8671 31547
rect 8727 31491 8751 31547
rect 8807 31491 8831 31547
rect 8887 31491 8911 31547
rect 8967 31491 8991 31547
rect 9047 31491 9071 31547
rect 9127 31491 9151 31547
rect 9207 31491 9231 31547
rect 9287 31491 9296 31547
rect 8098 31485 9296 31491
rect 9595 32613 10793 32619
rect 9595 32557 9604 32613
rect 9660 32557 9685 32613
rect 9741 32557 9766 32613
rect 9822 32557 9847 32613
rect 9903 32557 9928 32613
rect 9984 32557 10008 32613
rect 10064 32557 10088 32613
rect 10144 32557 10168 32613
rect 10224 32557 10248 32613
rect 10304 32557 10328 32613
rect 10384 32557 10408 32613
rect 10464 32557 10488 32613
rect 10544 32557 10568 32613
rect 10624 32557 10648 32613
rect 10704 32557 10728 32613
rect 10784 32557 10793 32613
rect 9595 32531 10793 32557
rect 9595 32475 9604 32531
rect 9660 32475 9685 32531
rect 9741 32475 9766 32531
rect 9822 32475 9847 32531
rect 9903 32475 9928 32531
rect 9984 32475 10008 32531
rect 10064 32475 10088 32531
rect 10144 32475 10168 32531
rect 10224 32475 10248 32531
rect 10304 32475 10328 32531
rect 10384 32475 10408 32531
rect 10464 32475 10488 32531
rect 10544 32475 10568 32531
rect 10624 32475 10648 32531
rect 10704 32475 10728 32531
rect 10784 32475 10793 32531
rect 9595 32449 10793 32475
rect 9595 32393 9604 32449
rect 9660 32393 9685 32449
rect 9741 32393 9766 32449
rect 9822 32393 9847 32449
rect 9903 32393 9928 32449
rect 9984 32393 10008 32449
rect 10064 32393 10088 32449
rect 10144 32393 10168 32449
rect 10224 32393 10248 32449
rect 10304 32393 10328 32449
rect 10384 32393 10408 32449
rect 10464 32393 10488 32449
rect 10544 32393 10568 32449
rect 10624 32393 10648 32449
rect 10704 32393 10728 32449
rect 10784 32393 10793 32449
rect 9595 32367 10793 32393
rect 9595 32311 9604 32367
rect 9660 32311 9685 32367
rect 9741 32311 9766 32367
rect 9822 32311 9847 32367
rect 9903 32311 9928 32367
rect 9984 32311 10008 32367
rect 10064 32311 10088 32367
rect 10144 32311 10168 32367
rect 10224 32311 10248 32367
rect 10304 32311 10328 32367
rect 10384 32311 10408 32367
rect 10464 32311 10488 32367
rect 10544 32311 10568 32367
rect 10624 32311 10648 32367
rect 10704 32311 10728 32367
rect 10784 32311 10793 32367
rect 9595 32285 10793 32311
rect 9595 32229 9604 32285
rect 9660 32229 9685 32285
rect 9741 32229 9766 32285
rect 9822 32229 9847 32285
rect 9903 32229 9928 32285
rect 9984 32229 10008 32285
rect 10064 32229 10088 32285
rect 10144 32229 10168 32285
rect 10224 32229 10248 32285
rect 10304 32229 10328 32285
rect 10384 32229 10408 32285
rect 10464 32229 10488 32285
rect 10544 32229 10568 32285
rect 10624 32229 10648 32285
rect 10704 32229 10728 32285
rect 10784 32229 10793 32285
rect 9595 32203 10793 32229
rect 9595 32147 9604 32203
rect 9660 32147 9685 32203
rect 9741 32147 9766 32203
rect 9822 32147 9847 32203
rect 9903 32147 9928 32203
rect 9984 32147 10008 32203
rect 10064 32147 10088 32203
rect 10144 32147 10168 32203
rect 10224 32147 10248 32203
rect 10304 32147 10328 32203
rect 10384 32147 10408 32203
rect 10464 32147 10488 32203
rect 10544 32147 10568 32203
rect 10624 32147 10648 32203
rect 10704 32147 10728 32203
rect 10784 32147 10793 32203
rect 9595 32121 10793 32147
rect 9595 32065 9604 32121
rect 9660 32065 9685 32121
rect 9741 32065 9766 32121
rect 9822 32065 9847 32121
rect 9903 32065 9928 32121
rect 9984 32065 10008 32121
rect 10064 32065 10088 32121
rect 10144 32065 10168 32121
rect 10224 32065 10248 32121
rect 10304 32065 10328 32121
rect 10384 32065 10408 32121
rect 10464 32065 10488 32121
rect 10544 32065 10568 32121
rect 10624 32065 10648 32121
rect 10704 32065 10728 32121
rect 10784 32065 10793 32121
rect 9595 32039 10793 32065
rect 9595 31983 9604 32039
rect 9660 31983 9685 32039
rect 9741 31983 9766 32039
rect 9822 31983 9847 32039
rect 9903 31983 9928 32039
rect 9984 31983 10008 32039
rect 10064 31983 10088 32039
rect 10144 31983 10168 32039
rect 10224 31983 10248 32039
rect 10304 31983 10328 32039
rect 10384 31983 10408 32039
rect 10464 31983 10488 32039
rect 10544 31983 10568 32039
rect 10624 31983 10648 32039
rect 10704 31983 10728 32039
rect 10784 31983 10793 32039
rect 9595 31957 10793 31983
rect 9595 31901 9604 31957
rect 9660 31901 9685 31957
rect 9741 31901 9766 31957
rect 9822 31901 9847 31957
rect 9903 31901 9928 31957
rect 9984 31901 10008 31957
rect 10064 31901 10088 31957
rect 10144 31901 10168 31957
rect 10224 31901 10248 31957
rect 10304 31901 10328 31957
rect 10384 31901 10408 31957
rect 10464 31901 10488 31957
rect 10544 31901 10568 31957
rect 10624 31901 10648 31957
rect 10704 31901 10728 31957
rect 10784 31901 10793 31957
rect 9595 31875 10793 31901
rect 9595 31819 9604 31875
rect 9660 31819 9685 31875
rect 9741 31819 9766 31875
rect 9822 31819 9847 31875
rect 9903 31819 9928 31875
rect 9984 31819 10008 31875
rect 10064 31819 10088 31875
rect 10144 31819 10168 31875
rect 10224 31819 10248 31875
rect 10304 31819 10328 31875
rect 10384 31819 10408 31875
rect 10464 31819 10488 31875
rect 10544 31819 10568 31875
rect 10624 31819 10648 31875
rect 10704 31819 10728 31875
rect 10784 31819 10793 31875
rect 9595 31793 10793 31819
rect 9595 31737 9604 31793
rect 9660 31737 9685 31793
rect 9741 31737 9766 31793
rect 9822 31737 9847 31793
rect 9903 31737 9928 31793
rect 9984 31737 10008 31793
rect 10064 31737 10088 31793
rect 10144 31737 10168 31793
rect 10224 31737 10248 31793
rect 10304 31737 10328 31793
rect 10384 31737 10408 31793
rect 10464 31737 10488 31793
rect 10544 31737 10568 31793
rect 10624 31737 10648 31793
rect 10704 31737 10728 31793
rect 10784 31737 10793 31793
rect 9595 31711 10793 31737
rect 9595 31655 9604 31711
rect 9660 31655 9685 31711
rect 9741 31655 9766 31711
rect 9822 31655 9847 31711
rect 9903 31655 9928 31711
rect 9984 31655 10008 31711
rect 10064 31655 10088 31711
rect 10144 31655 10168 31711
rect 10224 31655 10248 31711
rect 10304 31655 10328 31711
rect 10384 31655 10408 31711
rect 10464 31655 10488 31711
rect 10544 31655 10568 31711
rect 10624 31655 10648 31711
rect 10704 31655 10728 31711
rect 10784 31655 10793 31711
rect 9595 31629 10793 31655
rect 9595 31573 9604 31629
rect 9660 31573 9685 31629
rect 9741 31573 9766 31629
rect 9822 31573 9847 31629
rect 9903 31573 9928 31629
rect 9984 31573 10008 31629
rect 10064 31573 10088 31629
rect 10144 31573 10168 31629
rect 10224 31573 10248 31629
rect 10304 31573 10328 31629
rect 10384 31573 10408 31629
rect 10464 31573 10488 31629
rect 10544 31573 10568 31629
rect 10624 31573 10648 31629
rect 10704 31573 10728 31629
rect 10784 31573 10793 31629
rect 9595 31547 10793 31573
rect 9595 31491 9604 31547
rect 9660 31491 9685 31547
rect 9741 31491 9766 31547
rect 9822 31491 9847 31547
rect 9903 31491 9928 31547
rect 9984 31491 10008 31547
rect 10064 31491 10088 31547
rect 10144 31491 10168 31547
rect 10224 31491 10248 31547
rect 10304 31491 10328 31547
rect 10384 31491 10408 31547
rect 10464 31491 10488 31547
rect 10544 31491 10568 31547
rect 10624 31491 10648 31547
rect 10704 31491 10728 31547
rect 10784 31491 10793 31547
rect 9595 31485 10793 31491
rect 11092 32613 12290 32619
rect 11092 32557 11101 32613
rect 11157 32557 11182 32613
rect 11238 32557 11263 32613
rect 11319 32557 11344 32613
rect 11400 32557 11425 32613
rect 11481 32557 11505 32613
rect 11561 32557 11585 32613
rect 11641 32557 11665 32613
rect 11721 32557 11745 32613
rect 11801 32557 11825 32613
rect 11881 32557 11905 32613
rect 11961 32557 11985 32613
rect 12041 32557 12065 32613
rect 12121 32557 12145 32613
rect 12201 32557 12225 32613
rect 12281 32557 12290 32613
rect 11092 32531 12290 32557
rect 11092 32475 11101 32531
rect 11157 32475 11182 32531
rect 11238 32475 11263 32531
rect 11319 32475 11344 32531
rect 11400 32475 11425 32531
rect 11481 32475 11505 32531
rect 11561 32475 11585 32531
rect 11641 32475 11665 32531
rect 11721 32475 11745 32531
rect 11801 32475 11825 32531
rect 11881 32475 11905 32531
rect 11961 32475 11985 32531
rect 12041 32475 12065 32531
rect 12121 32475 12145 32531
rect 12201 32475 12225 32531
rect 12281 32475 12290 32531
rect 11092 32449 12290 32475
rect 11092 32393 11101 32449
rect 11157 32393 11182 32449
rect 11238 32393 11263 32449
rect 11319 32393 11344 32449
rect 11400 32393 11425 32449
rect 11481 32393 11505 32449
rect 11561 32393 11585 32449
rect 11641 32393 11665 32449
rect 11721 32393 11745 32449
rect 11801 32393 11825 32449
rect 11881 32393 11905 32449
rect 11961 32393 11985 32449
rect 12041 32393 12065 32449
rect 12121 32393 12145 32449
rect 12201 32393 12225 32449
rect 12281 32393 12290 32449
rect 11092 32367 12290 32393
rect 11092 32311 11101 32367
rect 11157 32311 11182 32367
rect 11238 32311 11263 32367
rect 11319 32311 11344 32367
rect 11400 32311 11425 32367
rect 11481 32311 11505 32367
rect 11561 32311 11585 32367
rect 11641 32311 11665 32367
rect 11721 32311 11745 32367
rect 11801 32311 11825 32367
rect 11881 32311 11905 32367
rect 11961 32311 11985 32367
rect 12041 32311 12065 32367
rect 12121 32311 12145 32367
rect 12201 32311 12225 32367
rect 12281 32311 12290 32367
rect 11092 32285 12290 32311
rect 11092 32229 11101 32285
rect 11157 32229 11182 32285
rect 11238 32229 11263 32285
rect 11319 32229 11344 32285
rect 11400 32229 11425 32285
rect 11481 32229 11505 32285
rect 11561 32229 11585 32285
rect 11641 32229 11665 32285
rect 11721 32229 11745 32285
rect 11801 32229 11825 32285
rect 11881 32229 11905 32285
rect 11961 32229 11985 32285
rect 12041 32229 12065 32285
rect 12121 32229 12145 32285
rect 12201 32229 12225 32285
rect 12281 32229 12290 32285
rect 11092 32203 12290 32229
rect 11092 32147 11101 32203
rect 11157 32147 11182 32203
rect 11238 32147 11263 32203
rect 11319 32147 11344 32203
rect 11400 32147 11425 32203
rect 11481 32147 11505 32203
rect 11561 32147 11585 32203
rect 11641 32147 11665 32203
rect 11721 32147 11745 32203
rect 11801 32147 11825 32203
rect 11881 32147 11905 32203
rect 11961 32147 11985 32203
rect 12041 32147 12065 32203
rect 12121 32147 12145 32203
rect 12201 32147 12225 32203
rect 12281 32147 12290 32203
rect 11092 32121 12290 32147
rect 11092 32065 11101 32121
rect 11157 32065 11182 32121
rect 11238 32065 11263 32121
rect 11319 32065 11344 32121
rect 11400 32065 11425 32121
rect 11481 32065 11505 32121
rect 11561 32065 11585 32121
rect 11641 32065 11665 32121
rect 11721 32065 11745 32121
rect 11801 32065 11825 32121
rect 11881 32065 11905 32121
rect 11961 32065 11985 32121
rect 12041 32065 12065 32121
rect 12121 32065 12145 32121
rect 12201 32065 12225 32121
rect 12281 32065 12290 32121
rect 11092 32039 12290 32065
rect 11092 31983 11101 32039
rect 11157 31983 11182 32039
rect 11238 31983 11263 32039
rect 11319 31983 11344 32039
rect 11400 31983 11425 32039
rect 11481 31983 11505 32039
rect 11561 31983 11585 32039
rect 11641 31983 11665 32039
rect 11721 31983 11745 32039
rect 11801 31983 11825 32039
rect 11881 31983 11905 32039
rect 11961 31983 11985 32039
rect 12041 31983 12065 32039
rect 12121 31983 12145 32039
rect 12201 31983 12225 32039
rect 12281 31983 12290 32039
rect 11092 31957 12290 31983
rect 11092 31901 11101 31957
rect 11157 31901 11182 31957
rect 11238 31901 11263 31957
rect 11319 31901 11344 31957
rect 11400 31901 11425 31957
rect 11481 31901 11505 31957
rect 11561 31901 11585 31957
rect 11641 31901 11665 31957
rect 11721 31901 11745 31957
rect 11801 31901 11825 31957
rect 11881 31901 11905 31957
rect 11961 31901 11985 31957
rect 12041 31901 12065 31957
rect 12121 31901 12145 31957
rect 12201 31901 12225 31957
rect 12281 31901 12290 31957
rect 11092 31875 12290 31901
rect 11092 31819 11101 31875
rect 11157 31819 11182 31875
rect 11238 31819 11263 31875
rect 11319 31819 11344 31875
rect 11400 31819 11425 31875
rect 11481 31819 11505 31875
rect 11561 31819 11585 31875
rect 11641 31819 11665 31875
rect 11721 31819 11745 31875
rect 11801 31819 11825 31875
rect 11881 31819 11905 31875
rect 11961 31819 11985 31875
rect 12041 31819 12065 31875
rect 12121 31819 12145 31875
rect 12201 31819 12225 31875
rect 12281 31819 12290 31875
rect 11092 31793 12290 31819
rect 11092 31737 11101 31793
rect 11157 31737 11182 31793
rect 11238 31737 11263 31793
rect 11319 31737 11344 31793
rect 11400 31737 11425 31793
rect 11481 31737 11505 31793
rect 11561 31737 11585 31793
rect 11641 31737 11665 31793
rect 11721 31737 11745 31793
rect 11801 31737 11825 31793
rect 11881 31737 11905 31793
rect 11961 31737 11985 31793
rect 12041 31737 12065 31793
rect 12121 31737 12145 31793
rect 12201 31737 12225 31793
rect 12281 31737 12290 31793
rect 11092 31711 12290 31737
rect 11092 31655 11101 31711
rect 11157 31655 11182 31711
rect 11238 31655 11263 31711
rect 11319 31655 11344 31711
rect 11400 31655 11425 31711
rect 11481 31655 11505 31711
rect 11561 31655 11585 31711
rect 11641 31655 11665 31711
rect 11721 31655 11745 31711
rect 11801 31655 11825 31711
rect 11881 31655 11905 31711
rect 11961 31655 11985 31711
rect 12041 31655 12065 31711
rect 12121 31655 12145 31711
rect 12201 31655 12225 31711
rect 12281 31655 12290 31711
rect 11092 31629 12290 31655
rect 11092 31573 11101 31629
rect 11157 31573 11182 31629
rect 11238 31573 11263 31629
rect 11319 31573 11344 31629
rect 11400 31573 11425 31629
rect 11481 31573 11505 31629
rect 11561 31573 11585 31629
rect 11641 31573 11665 31629
rect 11721 31573 11745 31629
rect 11801 31573 11825 31629
rect 11881 31573 11905 31629
rect 11961 31573 11985 31629
rect 12041 31573 12065 31629
rect 12121 31573 12145 31629
rect 12201 31573 12225 31629
rect 12281 31573 12290 31629
rect 11092 31547 12290 31573
rect 11092 31491 11101 31547
rect 11157 31491 11182 31547
rect 11238 31491 11263 31547
rect 11319 31491 11344 31547
rect 11400 31491 11425 31547
rect 11481 31491 11505 31547
rect 11561 31491 11585 31547
rect 11641 31491 11665 31547
rect 11721 31491 11745 31547
rect 11801 31491 11825 31547
rect 11881 31491 11905 31547
rect 11961 31491 11985 31547
rect 12041 31491 12065 31547
rect 12121 31491 12145 31547
rect 12201 31491 12225 31547
rect 12281 31491 12290 31547
rect 11092 31485 12290 31491
rect 12589 32613 13268 32619
rect 12589 32557 12598 32613
rect 12654 32557 12685 32613
rect 12741 32557 12772 32613
rect 12828 32557 12859 32613
rect 12915 32557 12945 32613
rect 13001 32557 13031 32613
rect 13087 32557 13117 32613
rect 13173 32557 13203 32613
rect 13259 32557 13268 32613
rect 12589 32531 13268 32557
rect 12589 32475 12598 32531
rect 12654 32475 12685 32531
rect 12741 32475 12772 32531
rect 12828 32475 12859 32531
rect 12915 32475 12945 32531
rect 13001 32475 13031 32531
rect 13087 32475 13117 32531
rect 13173 32475 13203 32531
rect 13259 32475 13268 32531
rect 12589 32449 13268 32475
rect 12589 32393 12598 32449
rect 12654 32393 12685 32449
rect 12741 32393 12772 32449
rect 12828 32393 12859 32449
rect 12915 32393 12945 32449
rect 13001 32393 13031 32449
rect 13087 32393 13117 32449
rect 13173 32393 13203 32449
rect 13259 32393 13268 32449
rect 12589 32367 13268 32393
rect 12589 32311 12598 32367
rect 12654 32311 12685 32367
rect 12741 32311 12772 32367
rect 12828 32311 12859 32367
rect 12915 32311 12945 32367
rect 13001 32311 13031 32367
rect 13087 32311 13117 32367
rect 13173 32311 13203 32367
rect 13259 32311 13268 32367
rect 12589 32285 13268 32311
rect 12589 32229 12598 32285
rect 12654 32229 12685 32285
rect 12741 32229 12772 32285
rect 12828 32229 12859 32285
rect 12915 32229 12945 32285
rect 13001 32229 13031 32285
rect 13087 32229 13117 32285
rect 13173 32229 13203 32285
rect 13259 32229 13268 32285
rect 12589 32203 13268 32229
rect 12589 32147 12598 32203
rect 12654 32147 12685 32203
rect 12741 32147 12772 32203
rect 12828 32147 12859 32203
rect 12915 32147 12945 32203
rect 13001 32147 13031 32203
rect 13087 32147 13117 32203
rect 13173 32147 13203 32203
rect 13259 32147 13268 32203
rect 12589 32121 13268 32147
rect 12589 32065 12598 32121
rect 12654 32065 12685 32121
rect 12741 32065 12772 32121
rect 12828 32065 12859 32121
rect 12915 32065 12945 32121
rect 13001 32065 13031 32121
rect 13087 32065 13117 32121
rect 13173 32065 13203 32121
rect 13259 32065 13268 32121
rect 12589 32039 13268 32065
rect 12589 31983 12598 32039
rect 12654 31983 12685 32039
rect 12741 31983 12772 32039
rect 12828 31983 12859 32039
rect 12915 31983 12945 32039
rect 13001 31983 13031 32039
rect 13087 31983 13117 32039
rect 13173 31983 13203 32039
rect 13259 31983 13268 32039
rect 12589 31957 13268 31983
rect 12589 31901 12598 31957
rect 12654 31901 12685 31957
rect 12741 31901 12772 31957
rect 12828 31901 12859 31957
rect 12915 31901 12945 31957
rect 13001 31901 13031 31957
rect 13087 31901 13117 31957
rect 13173 31901 13203 31957
rect 13259 31901 13268 31957
rect 12589 31875 13268 31901
rect 12589 31819 12598 31875
rect 12654 31819 12685 31875
rect 12741 31819 12772 31875
rect 12828 31819 12859 31875
rect 12915 31819 12945 31875
rect 13001 31819 13031 31875
rect 13087 31819 13117 31875
rect 13173 31819 13203 31875
rect 13259 31819 13268 31875
rect 12589 31793 13268 31819
rect 12589 31737 12598 31793
rect 12654 31737 12685 31793
rect 12741 31737 12772 31793
rect 12828 31737 12859 31793
rect 12915 31737 12945 31793
rect 13001 31737 13031 31793
rect 13087 31737 13117 31793
rect 13173 31737 13203 31793
rect 13259 31737 13268 31793
rect 12589 31711 13268 31737
rect 12589 31655 12598 31711
rect 12654 31655 12685 31711
rect 12741 31655 12772 31711
rect 12828 31655 12859 31711
rect 12915 31655 12945 31711
rect 13001 31655 13031 31711
rect 13087 31655 13117 31711
rect 13173 31655 13203 31711
rect 13259 31655 13268 31711
rect 12589 31629 13268 31655
rect 12589 31573 12598 31629
rect 12654 31573 12685 31629
rect 12741 31573 12772 31629
rect 12828 31573 12859 31629
rect 12915 31573 12945 31629
rect 13001 31573 13031 31629
rect 13087 31573 13117 31629
rect 13173 31573 13203 31629
rect 13259 31573 13268 31629
rect 12589 31547 13268 31573
rect 12589 31491 12598 31547
rect 12654 31491 12685 31547
rect 12741 31491 12772 31547
rect 12828 31491 12859 31547
rect 12915 31491 12945 31547
rect 13001 31491 13031 31547
rect 13087 31491 13117 31547
rect 13173 31491 13203 31547
rect 13259 31491 13268 31547
rect 12589 31485 13268 31491
rect 299 31448 454 31473
rect 506 31448 528 31473
rect 580 31448 602 31473
rect 148 31429 298 31442
rect 148 31377 149 31429
rect 201 31377 247 31429
rect 354 31392 396 31448
rect 452 31442 454 31448
rect 580 31442 592 31448
rect 452 31429 494 31442
rect 550 31429 592 31442
rect 648 31429 654 31442
rect 452 31392 454 31429
rect 580 31392 592 31429
rect 299 31377 454 31392
rect 506 31377 528 31392
rect 580 31377 602 31392
rect 148 31367 654 31377
rect 148 31364 298 31367
rect 148 31312 149 31364
rect 201 31312 247 31364
rect 148 31311 298 31312
rect 354 31311 396 31367
rect 452 31364 494 31367
rect 550 31364 592 31367
rect 648 31364 654 31367
rect 452 31312 454 31364
rect 580 31312 592 31364
rect 452 31311 494 31312
rect 550 31311 592 31312
rect 648 31311 654 31312
rect 148 31299 654 31311
rect 148 31247 149 31299
rect 201 31247 247 31299
rect 299 31286 454 31299
rect 506 31286 528 31299
rect 580 31286 602 31299
rect 148 31234 298 31247
rect 148 31182 149 31234
rect 201 31182 247 31234
rect 354 31230 396 31286
rect 452 31247 454 31286
rect 580 31247 592 31286
rect 452 31234 494 31247
rect 550 31234 592 31247
rect 648 31234 654 31247
rect 452 31230 454 31234
rect 580 31230 592 31234
rect 299 31205 454 31230
rect 506 31205 528 31230
rect 580 31205 602 31230
rect 148 31169 298 31182
rect 148 31117 149 31169
rect 201 31117 247 31169
rect 354 31149 396 31205
rect 452 31182 454 31205
rect 580 31182 592 31205
rect 452 31169 494 31182
rect 550 31169 592 31182
rect 648 31169 654 31182
rect 452 31149 454 31169
rect 580 31149 592 31169
rect 299 31124 454 31149
rect 506 31124 528 31149
rect 580 31124 602 31149
rect 148 31104 298 31117
rect 148 31052 149 31104
rect 201 31052 247 31104
rect 354 31068 396 31124
rect 452 31117 454 31124
rect 580 31117 592 31124
rect 452 31104 494 31117
rect 550 31104 592 31117
rect 648 31104 654 31117
rect 452 31068 454 31104
rect 580 31068 592 31104
rect 299 31052 454 31068
rect 506 31052 528 31068
rect 580 31052 602 31068
rect 148 31043 654 31052
rect 148 31039 298 31043
rect 148 30987 149 31039
rect 201 30987 247 31039
rect 354 30987 396 31043
rect 452 31039 494 31043
rect 550 31039 592 31043
rect 648 31039 654 31043
rect 452 30987 454 31039
rect 580 30987 592 31039
rect 148 30974 654 30987
rect 148 30922 149 30974
rect 201 30922 247 30974
rect 299 30962 454 30974
rect 506 30962 528 30974
rect 580 30962 602 30974
rect 148 30909 298 30922
rect 148 30857 149 30909
rect 201 30857 247 30909
rect 354 30906 396 30962
rect 452 30922 454 30962
rect 580 30922 592 30962
rect 452 30909 494 30922
rect 550 30909 592 30922
rect 648 30909 654 30922
rect 452 30906 454 30909
rect 580 30906 592 30909
rect 299 30881 454 30906
rect 506 30881 528 30906
rect 580 30881 602 30906
rect 148 30844 298 30857
rect 148 30792 149 30844
rect 201 30792 247 30844
rect 354 30825 396 30881
rect 452 30857 454 30881
rect 580 30857 592 30881
rect 452 30844 494 30857
rect 550 30844 592 30857
rect 648 30844 654 30857
rect 452 30825 454 30844
rect 580 30825 592 30844
rect 299 30800 454 30825
rect 506 30800 528 30825
rect 580 30800 602 30825
rect 148 30779 298 30792
rect 148 30727 149 30779
rect 201 30727 247 30779
rect 354 30744 396 30800
rect 452 30792 454 30800
rect 580 30792 592 30800
rect 452 30779 494 30792
rect 550 30779 592 30792
rect 648 30779 654 30792
rect 452 30744 454 30779
rect 580 30744 592 30779
rect 299 30727 454 30744
rect 506 30727 528 30744
rect 580 30727 602 30744
rect 148 30719 654 30727
rect 148 30714 298 30719
rect 148 30662 149 30714
rect 201 30662 247 30714
rect 354 30663 396 30719
rect 452 30714 494 30719
rect 550 30714 592 30719
rect 648 30714 654 30719
rect 452 30663 454 30714
rect 580 30663 592 30714
rect 299 30662 454 30663
rect 506 30662 528 30663
rect 580 30662 602 30663
rect 148 30649 654 30662
rect 148 30597 149 30649
rect 201 30597 247 30649
rect 299 30638 454 30649
rect 506 30638 528 30649
rect 580 30638 602 30649
rect 148 30584 298 30597
rect 148 30532 149 30584
rect 201 30532 247 30584
rect 354 30582 396 30638
rect 452 30597 454 30638
rect 580 30597 592 30638
rect 452 30584 494 30597
rect 550 30584 592 30597
rect 648 30584 654 30597
rect 452 30582 454 30584
rect 580 30582 592 30584
rect 299 30557 454 30582
rect 506 30557 528 30582
rect 580 30557 602 30582
rect 148 30519 298 30532
rect 148 30467 149 30519
rect 201 30467 247 30519
rect 354 30501 396 30557
rect 452 30532 454 30557
rect 580 30532 592 30557
rect 452 30519 494 30532
rect 550 30519 592 30532
rect 648 30519 654 30532
rect 452 30501 454 30519
rect 580 30501 592 30519
rect 299 30476 454 30501
rect 506 30476 528 30501
rect 580 30476 602 30501
rect 148 30454 298 30467
rect 148 30402 149 30454
rect 201 30402 247 30454
rect 354 30420 396 30476
rect 452 30467 454 30476
rect 580 30467 592 30476
rect 452 30454 494 30467
rect 550 30454 592 30467
rect 648 30454 654 30467
rect 452 30420 454 30454
rect 580 30420 592 30454
rect 299 30402 454 30420
rect 506 30402 528 30420
rect 580 30402 602 30420
rect 148 30395 654 30402
rect 148 30389 298 30395
rect 148 30337 149 30389
rect 201 30337 247 30389
rect 354 30339 396 30395
rect 452 30389 494 30395
rect 550 30389 592 30395
rect 648 30389 654 30395
rect 452 30339 454 30389
rect 580 30339 592 30389
rect 299 30337 454 30339
rect 506 30337 528 30339
rect 580 30337 602 30339
rect 148 30324 654 30337
rect 148 30272 149 30324
rect 201 30272 247 30324
rect 299 30314 454 30324
rect 506 30314 528 30324
rect 580 30314 602 30324
rect 148 30259 298 30272
rect 148 30207 149 30259
rect 201 30207 247 30259
rect 354 30258 396 30314
rect 452 30272 454 30314
rect 580 30272 592 30314
rect 452 30259 494 30272
rect 550 30259 592 30272
rect 648 30259 654 30272
rect 452 30258 454 30259
rect 580 30258 592 30259
rect 299 30233 454 30258
rect 506 30233 528 30258
rect 580 30233 602 30258
rect 148 30194 298 30207
rect 148 30142 149 30194
rect 201 30142 247 30194
rect 354 30177 396 30233
rect 452 30207 454 30233
rect 580 30207 592 30233
rect 452 30194 494 30207
rect 550 30194 592 30207
rect 648 30194 654 30207
rect 452 30177 454 30194
rect 580 30177 592 30194
rect 299 30152 454 30177
rect 506 30152 528 30177
rect 580 30152 602 30177
rect 148 30129 298 30142
rect 148 30077 149 30129
rect 201 30077 247 30129
rect 354 30096 396 30152
rect 452 30142 454 30152
rect 580 30142 592 30152
rect 452 30129 494 30142
rect 550 30129 592 30142
rect 648 30129 654 30142
rect 452 30096 454 30129
rect 580 30096 592 30129
rect 299 30077 454 30096
rect 506 30077 528 30096
rect 580 30077 602 30096
rect 148 30071 654 30077
rect 148 30064 298 30071
rect 148 30012 149 30064
rect 201 30012 247 30064
rect 354 30015 396 30071
rect 452 30064 494 30071
rect 550 30064 592 30071
rect 648 30064 654 30071
rect 452 30015 454 30064
rect 580 30015 592 30064
rect 299 30012 454 30015
rect 506 30012 528 30015
rect 580 30012 602 30015
rect 148 29999 654 30012
rect 148 29947 149 29999
rect 201 29947 247 29999
rect 299 29990 454 29999
rect 506 29990 528 29999
rect 580 29990 602 29999
rect 148 29934 298 29947
rect 354 29934 396 29990
rect 452 29947 454 29990
rect 580 29947 592 29990
rect 452 29934 494 29947
rect 550 29934 592 29947
rect 648 29934 654 29947
rect 148 29882 149 29934
rect 201 29882 247 29934
rect 299 29909 454 29934
rect 506 29909 528 29934
rect 580 29909 602 29934
rect 148 29869 298 29882
rect 148 29817 149 29869
rect 201 29817 247 29869
rect 354 29853 396 29909
rect 452 29882 454 29909
rect 580 29882 592 29909
rect 452 29869 494 29882
rect 550 29869 592 29882
rect 648 29869 654 29882
rect 452 29853 454 29869
rect 580 29853 592 29869
rect 299 29828 454 29853
rect 506 29828 528 29853
rect 580 29828 602 29853
rect 148 29804 298 29817
rect 148 29752 149 29804
rect 201 29752 247 29804
rect 354 29772 396 29828
rect 452 29817 454 29828
rect 580 29817 592 29828
rect 452 29804 494 29817
rect 550 29804 592 29817
rect 648 29804 654 29817
rect 452 29772 454 29804
rect 580 29772 592 29804
rect 299 29752 454 29772
rect 506 29752 528 29772
rect 580 29752 602 29772
rect 148 29747 654 29752
rect 148 29739 298 29747
rect 148 29687 149 29739
rect 201 29687 247 29739
rect 354 29691 396 29747
rect 452 29739 494 29747
rect 550 29739 592 29747
rect 648 29739 654 29747
rect 452 29691 454 29739
rect 580 29691 592 29739
rect 299 29687 454 29691
rect 506 29687 528 29691
rect 580 29687 602 29691
rect 148 29674 654 29687
rect 148 29622 149 29674
rect 201 29622 247 29674
rect 299 29666 454 29674
rect 506 29666 528 29674
rect 580 29666 602 29674
rect 148 29610 298 29622
rect 354 29610 396 29666
rect 452 29622 454 29666
rect 580 29622 592 29666
rect 452 29610 494 29622
rect 550 29610 592 29622
rect 648 29610 654 29622
rect 148 29609 654 29610
rect 148 29557 149 29609
rect 201 29557 247 29609
rect 299 29585 454 29609
rect 506 29585 528 29609
rect 580 29585 602 29609
rect 148 29544 298 29557
rect 148 29492 149 29544
rect 201 29492 247 29544
rect 354 29529 396 29585
rect 452 29557 454 29585
rect 580 29557 592 29585
rect 452 29544 494 29557
rect 550 29544 592 29557
rect 648 29544 654 29557
rect 452 29529 454 29544
rect 580 29529 592 29544
rect 299 29504 454 29529
rect 506 29504 528 29529
rect 580 29504 602 29529
rect 148 29479 298 29492
rect 148 29427 149 29479
rect 201 29427 247 29479
rect 354 29448 396 29504
rect 452 29492 454 29504
rect 580 29492 592 29504
rect 452 29479 494 29492
rect 550 29479 592 29492
rect 648 29479 654 29492
rect 452 29448 454 29479
rect 580 29448 592 29479
rect 299 29427 454 29448
rect 506 29427 528 29448
rect 580 29427 602 29448
rect 1694 31164 15298 31173
rect 1694 31160 14514 31164
rect 1694 31159 6182 31160
rect 1694 31103 2139 31159
rect 2195 31103 2237 31159
rect 2293 31103 2335 31159
rect 2391 31103 2433 31159
rect 2489 31104 6182 31159
rect 6238 31104 6263 31160
rect 6319 31104 6344 31160
rect 6400 31104 6425 31160
rect 6481 31104 6506 31160
rect 6562 31104 6587 31160
rect 6643 31104 6668 31160
rect 6724 31104 6749 31160
rect 6805 31104 6830 31160
rect 6886 31104 6911 31160
rect 6967 31104 6992 31160
rect 7048 31104 7073 31160
rect 7129 31104 7154 31160
rect 7210 31104 7235 31160
rect 7291 31104 7316 31160
rect 7372 31104 7397 31160
rect 7453 31104 7478 31160
rect 7534 31104 7559 31160
rect 7615 31104 7640 31160
rect 7696 31104 7721 31160
rect 7777 31104 7802 31160
rect 7858 31104 7883 31160
rect 7939 31104 7964 31160
rect 8020 31104 8045 31160
rect 8101 31104 8126 31160
rect 8182 31104 8207 31160
rect 8263 31104 8288 31160
rect 8344 31104 8369 31160
rect 8425 31104 8450 31160
rect 8506 31104 8531 31160
rect 8587 31104 8612 31160
rect 8668 31104 8693 31160
rect 8749 31104 8774 31160
rect 8830 31104 8855 31160
rect 8911 31104 8936 31160
rect 8992 31104 9017 31160
rect 9073 31104 9098 31160
rect 9154 31104 9179 31160
rect 9235 31104 9260 31160
rect 9316 31104 9340 31160
rect 9396 31104 9420 31160
rect 9476 31104 9500 31160
rect 9556 31104 9580 31160
rect 9636 31104 9660 31160
rect 9716 31104 9740 31160
rect 9796 31104 9820 31160
rect 9876 31104 9900 31160
rect 9956 31104 9980 31160
rect 10036 31104 10060 31160
rect 10116 31104 10140 31160
rect 10196 31104 10220 31160
rect 10276 31104 10300 31160
rect 10356 31104 10380 31160
rect 10436 31104 10460 31160
rect 10516 31104 10540 31160
rect 10596 31104 10620 31160
rect 10676 31104 10700 31160
rect 10756 31104 10780 31160
rect 10836 31104 10860 31160
rect 10916 31104 10940 31160
rect 10996 31104 11020 31160
rect 11076 31104 11100 31160
rect 11156 31104 11180 31160
rect 11236 31104 11260 31160
rect 11316 31104 11340 31160
rect 11396 31104 11420 31160
rect 11476 31104 11500 31160
rect 11556 31104 11580 31160
rect 11636 31104 11660 31160
rect 11716 31104 11740 31160
rect 11796 31104 11820 31160
rect 11876 31104 11900 31160
rect 11956 31104 11980 31160
rect 12036 31104 12060 31160
rect 12116 31104 12140 31160
rect 12196 31104 12220 31160
rect 12276 31104 12300 31160
rect 12356 31104 12380 31160
rect 12436 31104 12460 31160
rect 12516 31104 12540 31160
rect 12596 31104 12620 31160
rect 12676 31104 12700 31160
rect 12756 31104 12780 31160
rect 12836 31104 12860 31160
rect 12916 31104 12940 31160
rect 12996 31104 13020 31160
rect 13076 31108 14514 31160
rect 14570 31108 14594 31164
rect 14650 31108 14674 31164
rect 14730 31108 14754 31164
rect 14810 31108 14834 31164
rect 14890 31108 14914 31164
rect 14970 31108 14994 31164
rect 15050 31108 15074 31164
rect 15130 31108 15154 31164
rect 15210 31108 15234 31164
rect 15290 31108 15298 31164
rect 13076 31104 15298 31108
rect 2489 31103 15298 31104
rect 1694 31082 15298 31103
rect 1694 31078 14514 31082
rect 1694 31077 6182 31078
rect 1694 31021 2139 31077
rect 2195 31021 2237 31077
rect 2293 31021 2335 31077
rect 2391 31021 2433 31077
rect 2489 31022 6182 31077
rect 6238 31022 6263 31078
rect 6319 31022 6344 31078
rect 6400 31022 6425 31078
rect 6481 31022 6506 31078
rect 6562 31022 6587 31078
rect 6643 31022 6668 31078
rect 6724 31022 6749 31078
rect 6805 31022 6830 31078
rect 6886 31022 6911 31078
rect 6967 31022 6992 31078
rect 7048 31022 7073 31078
rect 7129 31022 7154 31078
rect 7210 31022 7235 31078
rect 7291 31022 7316 31078
rect 7372 31022 7397 31078
rect 7453 31022 7478 31078
rect 7534 31022 7559 31078
rect 7615 31022 7640 31078
rect 7696 31022 7721 31078
rect 7777 31022 7802 31078
rect 7858 31022 7883 31078
rect 7939 31022 7964 31078
rect 8020 31022 8045 31078
rect 8101 31022 8126 31078
rect 8182 31022 8207 31078
rect 8263 31022 8288 31078
rect 8344 31022 8369 31078
rect 8425 31022 8450 31078
rect 8506 31022 8531 31078
rect 8587 31022 8612 31078
rect 8668 31022 8693 31078
rect 8749 31022 8774 31078
rect 8830 31022 8855 31078
rect 8911 31022 8936 31078
rect 8992 31022 9017 31078
rect 9073 31022 9098 31078
rect 9154 31022 9179 31078
rect 9235 31022 9260 31078
rect 9316 31022 9340 31078
rect 9396 31022 9420 31078
rect 9476 31022 9500 31078
rect 9556 31022 9580 31078
rect 9636 31022 9660 31078
rect 9716 31022 9740 31078
rect 9796 31022 9820 31078
rect 9876 31022 9900 31078
rect 9956 31022 9980 31078
rect 10036 31022 10060 31078
rect 10116 31022 10140 31078
rect 10196 31022 10220 31078
rect 10276 31022 10300 31078
rect 10356 31022 10380 31078
rect 10436 31022 10460 31078
rect 10516 31022 10540 31078
rect 10596 31022 10620 31078
rect 10676 31022 10700 31078
rect 10756 31022 10780 31078
rect 10836 31022 10860 31078
rect 10916 31022 10940 31078
rect 10996 31022 11020 31078
rect 11076 31022 11100 31078
rect 11156 31022 11180 31078
rect 11236 31022 11260 31078
rect 11316 31022 11340 31078
rect 11396 31022 11420 31078
rect 11476 31022 11500 31078
rect 11556 31022 11580 31078
rect 11636 31022 11660 31078
rect 11716 31022 11740 31078
rect 11796 31022 11820 31078
rect 11876 31022 11900 31078
rect 11956 31022 11980 31078
rect 12036 31022 12060 31078
rect 12116 31022 12140 31078
rect 12196 31022 12220 31078
rect 12276 31022 12300 31078
rect 12356 31022 12380 31078
rect 12436 31022 12460 31078
rect 12516 31022 12540 31078
rect 12596 31022 12620 31078
rect 12676 31022 12700 31078
rect 12756 31022 12780 31078
rect 12836 31022 12860 31078
rect 12916 31022 12940 31078
rect 12996 31022 13020 31078
rect 13076 31026 14514 31078
rect 14570 31026 14594 31082
rect 14650 31026 14674 31082
rect 14730 31026 14754 31082
rect 14810 31026 14834 31082
rect 14890 31026 14914 31082
rect 14970 31026 14994 31082
rect 15050 31026 15074 31082
rect 15130 31026 15154 31082
rect 15210 31026 15234 31082
rect 15290 31026 15298 31082
rect 13076 31022 15298 31026
rect 2489 31021 15298 31022
rect 1694 31000 15298 31021
rect 1694 30996 14514 31000
rect 1694 30995 6182 30996
rect 1694 30939 2139 30995
rect 2195 30939 2237 30995
rect 2293 30939 2335 30995
rect 2391 30939 2433 30995
rect 2489 30993 6182 30995
rect 2489 30939 5803 30993
rect 1694 30937 5803 30939
rect 5859 30937 5895 30993
rect 5951 30937 5987 30993
rect 6043 30937 6079 30993
rect 6135 30940 6182 30993
rect 6238 30940 6263 30996
rect 6319 30940 6344 30996
rect 6400 30940 6425 30996
rect 6481 30940 6506 30996
rect 6562 30940 6587 30996
rect 6643 30940 6668 30996
rect 6724 30940 6749 30996
rect 6805 30940 6830 30996
rect 6886 30940 6911 30996
rect 6967 30940 6992 30996
rect 7048 30940 7073 30996
rect 7129 30940 7154 30996
rect 7210 30940 7235 30996
rect 7291 30940 7316 30996
rect 7372 30940 7397 30996
rect 7453 30940 7478 30996
rect 7534 30940 7559 30996
rect 7615 30940 7640 30996
rect 7696 30940 7721 30996
rect 7777 30940 7802 30996
rect 7858 30940 7883 30996
rect 7939 30940 7964 30996
rect 8020 30940 8045 30996
rect 8101 30940 8126 30996
rect 8182 30940 8207 30996
rect 8263 30940 8288 30996
rect 8344 30940 8369 30996
rect 8425 30940 8450 30996
rect 8506 30940 8531 30996
rect 8587 30940 8612 30996
rect 8668 30940 8693 30996
rect 8749 30940 8774 30996
rect 8830 30940 8855 30996
rect 8911 30940 8936 30996
rect 8992 30940 9017 30996
rect 9073 30940 9098 30996
rect 9154 30940 9179 30996
rect 9235 30940 9260 30996
rect 9316 30940 9340 30996
rect 9396 30940 9420 30996
rect 9476 30940 9500 30996
rect 9556 30940 9580 30996
rect 9636 30940 9660 30996
rect 9716 30940 9740 30996
rect 9796 30940 9820 30996
rect 9876 30940 9900 30996
rect 9956 30940 9980 30996
rect 10036 30940 10060 30996
rect 10116 30940 10140 30996
rect 10196 30940 10220 30996
rect 10276 30940 10300 30996
rect 10356 30940 10380 30996
rect 10436 30940 10460 30996
rect 10516 30940 10540 30996
rect 10596 30940 10620 30996
rect 10676 30940 10700 30996
rect 10756 30940 10780 30996
rect 10836 30940 10860 30996
rect 10916 30940 10940 30996
rect 10996 30940 11020 30996
rect 11076 30940 11100 30996
rect 11156 30940 11180 30996
rect 11236 30940 11260 30996
rect 11316 30940 11340 30996
rect 11396 30940 11420 30996
rect 11476 30940 11500 30996
rect 11556 30940 11580 30996
rect 11636 30940 11660 30996
rect 11716 30940 11740 30996
rect 11796 30940 11820 30996
rect 11876 30940 11900 30996
rect 11956 30940 11980 30996
rect 12036 30940 12060 30996
rect 12116 30940 12140 30996
rect 12196 30940 12220 30996
rect 12276 30940 12300 30996
rect 12356 30940 12380 30996
rect 12436 30940 12460 30996
rect 12516 30940 12540 30996
rect 12596 30940 12620 30996
rect 12676 30940 12700 30996
rect 12756 30940 12780 30996
rect 12836 30940 12860 30996
rect 12916 30940 12940 30996
rect 12996 30940 13020 30996
rect 13076 30944 14514 30996
rect 14570 30944 14594 31000
rect 14650 30944 14674 31000
rect 14730 30944 14754 31000
rect 14810 30944 14834 31000
rect 14890 30944 14914 31000
rect 14970 30944 14994 31000
rect 15050 30944 15074 31000
rect 15130 30944 15154 31000
rect 15210 30944 15234 31000
rect 15290 30944 15298 31000
rect 13076 30940 15298 30944
rect 6135 30937 15298 30940
rect 1694 30918 15298 30937
rect 1694 30914 14514 30918
rect 1694 30913 6182 30914
rect 1694 30857 2139 30913
rect 2195 30857 2237 30913
rect 2293 30857 2335 30913
rect 2391 30857 2433 30913
rect 2489 30910 6182 30913
rect 2489 30857 5803 30910
rect 1694 30854 5803 30857
rect 5859 30854 5895 30910
rect 5951 30854 5987 30910
rect 6043 30854 6079 30910
rect 6135 30858 6182 30910
rect 6238 30858 6263 30914
rect 6319 30858 6344 30914
rect 6400 30858 6425 30914
rect 6481 30858 6506 30914
rect 6562 30858 6587 30914
rect 6643 30858 6668 30914
rect 6724 30858 6749 30914
rect 6805 30858 6830 30914
rect 6886 30858 6911 30914
rect 6967 30858 6992 30914
rect 7048 30858 7073 30914
rect 7129 30858 7154 30914
rect 7210 30858 7235 30914
rect 7291 30858 7316 30914
rect 7372 30858 7397 30914
rect 7453 30858 7478 30914
rect 7534 30858 7559 30914
rect 7615 30858 7640 30914
rect 7696 30858 7721 30914
rect 7777 30858 7802 30914
rect 7858 30858 7883 30914
rect 7939 30858 7964 30914
rect 8020 30858 8045 30914
rect 8101 30858 8126 30914
rect 8182 30858 8207 30914
rect 8263 30858 8288 30914
rect 8344 30858 8369 30914
rect 8425 30858 8450 30914
rect 8506 30858 8531 30914
rect 8587 30858 8612 30914
rect 8668 30858 8693 30914
rect 8749 30858 8774 30914
rect 8830 30858 8855 30914
rect 8911 30858 8936 30914
rect 8992 30858 9017 30914
rect 9073 30858 9098 30914
rect 9154 30858 9179 30914
rect 9235 30858 9260 30914
rect 9316 30858 9340 30914
rect 9396 30858 9420 30914
rect 9476 30858 9500 30914
rect 9556 30858 9580 30914
rect 9636 30858 9660 30914
rect 9716 30858 9740 30914
rect 9796 30858 9820 30914
rect 9876 30858 9900 30914
rect 9956 30858 9980 30914
rect 10036 30858 10060 30914
rect 10116 30858 10140 30914
rect 10196 30858 10220 30914
rect 10276 30858 10300 30914
rect 10356 30858 10380 30914
rect 10436 30858 10460 30914
rect 10516 30858 10540 30914
rect 10596 30858 10620 30914
rect 10676 30858 10700 30914
rect 10756 30858 10780 30914
rect 10836 30858 10860 30914
rect 10916 30858 10940 30914
rect 10996 30858 11020 30914
rect 11076 30858 11100 30914
rect 11156 30858 11180 30914
rect 11236 30858 11260 30914
rect 11316 30858 11340 30914
rect 11396 30858 11420 30914
rect 11476 30858 11500 30914
rect 11556 30858 11580 30914
rect 11636 30858 11660 30914
rect 11716 30858 11740 30914
rect 11796 30858 11820 30914
rect 11876 30858 11900 30914
rect 11956 30858 11980 30914
rect 12036 30858 12060 30914
rect 12116 30858 12140 30914
rect 12196 30858 12220 30914
rect 12276 30858 12300 30914
rect 12356 30858 12380 30914
rect 12436 30858 12460 30914
rect 12516 30858 12540 30914
rect 12596 30858 12620 30914
rect 12676 30858 12700 30914
rect 12756 30858 12780 30914
rect 12836 30858 12860 30914
rect 12916 30858 12940 30914
rect 12996 30858 13020 30914
rect 13076 30862 14514 30914
rect 14570 30862 14594 30918
rect 14650 30862 14674 30918
rect 14730 30862 14754 30918
rect 14810 30862 14834 30918
rect 14890 30862 14914 30918
rect 14970 30862 14994 30918
rect 15050 30862 15074 30918
rect 15130 30862 15154 30918
rect 15210 30862 15234 30918
rect 15290 30862 15298 30918
rect 13076 30858 15298 30862
rect 6135 30854 15298 30858
rect 1694 30836 15298 30854
rect 1694 30832 14514 30836
rect 1694 30831 6182 30832
rect 1694 30775 2139 30831
rect 2195 30775 2237 30831
rect 2293 30775 2335 30831
rect 2391 30775 2433 30831
rect 2489 30827 6182 30831
rect 2489 30775 5803 30827
rect 1694 30771 5803 30775
rect 5859 30771 5895 30827
rect 5951 30771 5987 30827
rect 6043 30771 6079 30827
rect 6135 30776 6182 30827
rect 6238 30776 6263 30832
rect 6319 30776 6344 30832
rect 6400 30776 6425 30832
rect 6481 30776 6506 30832
rect 6562 30776 6587 30832
rect 6643 30776 6668 30832
rect 6724 30776 6749 30832
rect 6805 30776 6830 30832
rect 6886 30776 6911 30832
rect 6967 30776 6992 30832
rect 7048 30776 7073 30832
rect 7129 30776 7154 30832
rect 7210 30776 7235 30832
rect 7291 30776 7316 30832
rect 7372 30776 7397 30832
rect 7453 30776 7478 30832
rect 7534 30776 7559 30832
rect 7615 30776 7640 30832
rect 7696 30776 7721 30832
rect 7777 30776 7802 30832
rect 7858 30776 7883 30832
rect 7939 30776 7964 30832
rect 8020 30776 8045 30832
rect 8101 30776 8126 30832
rect 8182 30776 8207 30832
rect 8263 30776 8288 30832
rect 8344 30776 8369 30832
rect 8425 30776 8450 30832
rect 8506 30776 8531 30832
rect 8587 30776 8612 30832
rect 8668 30776 8693 30832
rect 8749 30776 8774 30832
rect 8830 30776 8855 30832
rect 8911 30776 8936 30832
rect 8992 30776 9017 30832
rect 9073 30776 9098 30832
rect 9154 30776 9179 30832
rect 9235 30776 9260 30832
rect 9316 30776 9340 30832
rect 9396 30776 9420 30832
rect 9476 30776 9500 30832
rect 9556 30776 9580 30832
rect 9636 30776 9660 30832
rect 9716 30776 9740 30832
rect 9796 30776 9820 30832
rect 9876 30776 9900 30832
rect 9956 30776 9980 30832
rect 10036 30776 10060 30832
rect 10116 30776 10140 30832
rect 10196 30776 10220 30832
rect 10276 30776 10300 30832
rect 10356 30776 10380 30832
rect 10436 30776 10460 30832
rect 10516 30776 10540 30832
rect 10596 30776 10620 30832
rect 10676 30776 10700 30832
rect 10756 30776 10780 30832
rect 10836 30776 10860 30832
rect 10916 30776 10940 30832
rect 10996 30776 11020 30832
rect 11076 30776 11100 30832
rect 11156 30776 11180 30832
rect 11236 30776 11260 30832
rect 11316 30776 11340 30832
rect 11396 30776 11420 30832
rect 11476 30776 11500 30832
rect 11556 30776 11580 30832
rect 11636 30776 11660 30832
rect 11716 30776 11740 30832
rect 11796 30776 11820 30832
rect 11876 30776 11900 30832
rect 11956 30776 11980 30832
rect 12036 30776 12060 30832
rect 12116 30776 12140 30832
rect 12196 30776 12220 30832
rect 12276 30776 12300 30832
rect 12356 30776 12380 30832
rect 12436 30776 12460 30832
rect 12516 30776 12540 30832
rect 12596 30776 12620 30832
rect 12676 30776 12700 30832
rect 12756 30776 12780 30832
rect 12836 30776 12860 30832
rect 12916 30776 12940 30832
rect 12996 30776 13020 30832
rect 13076 30780 14514 30832
rect 14570 30780 14594 30836
rect 14650 30780 14674 30836
rect 14730 30780 14754 30836
rect 14810 30780 14834 30836
rect 14890 30780 14914 30836
rect 14970 30780 14994 30836
rect 15050 30780 15074 30836
rect 15130 30780 15154 30836
rect 15210 30780 15234 30836
rect 15290 30780 15298 30836
rect 13076 30776 15298 30780
rect 6135 30771 15298 30776
rect 1694 30753 15298 30771
rect 1694 30750 14514 30753
rect 1694 30749 6182 30750
rect 1694 30693 2139 30749
rect 2195 30693 2237 30749
rect 2293 30693 2335 30749
rect 2391 30693 2433 30749
rect 2489 30744 6182 30749
rect 2489 30693 5803 30744
rect 1694 30688 5803 30693
rect 5859 30688 5895 30744
rect 5951 30688 5987 30744
rect 6043 30688 6079 30744
rect 6135 30694 6182 30744
rect 6238 30694 6263 30750
rect 6319 30694 6344 30750
rect 6400 30694 6425 30750
rect 6481 30694 6506 30750
rect 6562 30694 6587 30750
rect 6643 30694 6668 30750
rect 6724 30694 6749 30750
rect 6805 30694 6830 30750
rect 6886 30694 6911 30750
rect 6967 30694 6992 30750
rect 7048 30694 7073 30750
rect 7129 30694 7154 30750
rect 7210 30694 7235 30750
rect 7291 30694 7316 30750
rect 7372 30694 7397 30750
rect 7453 30694 7478 30750
rect 7534 30694 7559 30750
rect 7615 30694 7640 30750
rect 7696 30694 7721 30750
rect 7777 30694 7802 30750
rect 7858 30694 7883 30750
rect 7939 30694 7964 30750
rect 8020 30694 8045 30750
rect 8101 30694 8126 30750
rect 8182 30694 8207 30750
rect 8263 30694 8288 30750
rect 8344 30694 8369 30750
rect 8425 30694 8450 30750
rect 8506 30694 8531 30750
rect 8587 30694 8612 30750
rect 8668 30694 8693 30750
rect 8749 30694 8774 30750
rect 8830 30694 8855 30750
rect 8911 30694 8936 30750
rect 8992 30694 9017 30750
rect 9073 30694 9098 30750
rect 9154 30694 9179 30750
rect 9235 30694 9260 30750
rect 9316 30694 9340 30750
rect 9396 30694 9420 30750
rect 9476 30694 9500 30750
rect 9556 30694 9580 30750
rect 9636 30694 9660 30750
rect 9716 30694 9740 30750
rect 9796 30694 9820 30750
rect 9876 30694 9900 30750
rect 9956 30694 9980 30750
rect 10036 30694 10060 30750
rect 10116 30694 10140 30750
rect 10196 30694 10220 30750
rect 10276 30694 10300 30750
rect 10356 30694 10380 30750
rect 10436 30694 10460 30750
rect 10516 30694 10540 30750
rect 10596 30694 10620 30750
rect 10676 30694 10700 30750
rect 10756 30694 10780 30750
rect 10836 30694 10860 30750
rect 10916 30694 10940 30750
rect 10996 30694 11020 30750
rect 11076 30694 11100 30750
rect 11156 30694 11180 30750
rect 11236 30694 11260 30750
rect 11316 30694 11340 30750
rect 11396 30694 11420 30750
rect 11476 30694 11500 30750
rect 11556 30694 11580 30750
rect 11636 30694 11660 30750
rect 11716 30694 11740 30750
rect 11796 30694 11820 30750
rect 11876 30694 11900 30750
rect 11956 30694 11980 30750
rect 12036 30694 12060 30750
rect 12116 30694 12140 30750
rect 12196 30694 12220 30750
rect 12276 30694 12300 30750
rect 12356 30694 12380 30750
rect 12436 30694 12460 30750
rect 12516 30694 12540 30750
rect 12596 30694 12620 30750
rect 12676 30694 12700 30750
rect 12756 30694 12780 30750
rect 12836 30694 12860 30750
rect 12916 30694 12940 30750
rect 12996 30694 13020 30750
rect 13076 30697 14514 30750
rect 14570 30697 14594 30753
rect 14650 30697 14674 30753
rect 14730 30697 14754 30753
rect 14810 30697 14834 30753
rect 14890 30697 14914 30753
rect 14970 30697 14994 30753
rect 15050 30697 15074 30753
rect 15130 30697 15154 30753
rect 15210 30697 15234 30753
rect 15290 30697 15298 30753
rect 13076 30694 15298 30697
rect 6135 30688 15298 30694
rect 1694 30670 15298 30688
rect 1694 30668 14514 30670
rect 1694 30667 6182 30668
rect 1694 30611 2139 30667
rect 2195 30611 2237 30667
rect 2293 30611 2335 30667
rect 2391 30611 2433 30667
rect 2489 30661 6182 30667
rect 2489 30611 5803 30661
rect 1694 30605 5803 30611
rect 5859 30605 5895 30661
rect 5951 30605 5987 30661
rect 6043 30605 6079 30661
rect 6135 30612 6182 30661
rect 6238 30612 6263 30668
rect 6319 30612 6344 30668
rect 6400 30612 6425 30668
rect 6481 30612 6506 30668
rect 6562 30612 6587 30668
rect 6643 30612 6668 30668
rect 6724 30612 6749 30668
rect 6805 30612 6830 30668
rect 6886 30612 6911 30668
rect 6967 30612 6992 30668
rect 7048 30612 7073 30668
rect 7129 30612 7154 30668
rect 7210 30612 7235 30668
rect 7291 30612 7316 30668
rect 7372 30612 7397 30668
rect 7453 30612 7478 30668
rect 7534 30612 7559 30668
rect 7615 30612 7640 30668
rect 7696 30612 7721 30668
rect 7777 30612 7802 30668
rect 7858 30612 7883 30668
rect 7939 30612 7964 30668
rect 8020 30612 8045 30668
rect 8101 30612 8126 30668
rect 8182 30612 8207 30668
rect 8263 30612 8288 30668
rect 8344 30612 8369 30668
rect 8425 30612 8450 30668
rect 8506 30612 8531 30668
rect 8587 30612 8612 30668
rect 8668 30612 8693 30668
rect 8749 30612 8774 30668
rect 8830 30612 8855 30668
rect 8911 30612 8936 30668
rect 8992 30612 9017 30668
rect 9073 30612 9098 30668
rect 9154 30612 9179 30668
rect 9235 30612 9260 30668
rect 9316 30612 9340 30668
rect 9396 30612 9420 30668
rect 9476 30612 9500 30668
rect 9556 30612 9580 30668
rect 9636 30612 9660 30668
rect 9716 30612 9740 30668
rect 9796 30612 9820 30668
rect 9876 30612 9900 30668
rect 9956 30612 9980 30668
rect 10036 30612 10060 30668
rect 10116 30612 10140 30668
rect 10196 30612 10220 30668
rect 10276 30612 10300 30668
rect 10356 30612 10380 30668
rect 10436 30612 10460 30668
rect 10516 30612 10540 30668
rect 10596 30612 10620 30668
rect 10676 30612 10700 30668
rect 10756 30612 10780 30668
rect 10836 30612 10860 30668
rect 10916 30612 10940 30668
rect 10996 30612 11020 30668
rect 11076 30612 11100 30668
rect 11156 30612 11180 30668
rect 11236 30612 11260 30668
rect 11316 30612 11340 30668
rect 11396 30612 11420 30668
rect 11476 30612 11500 30668
rect 11556 30612 11580 30668
rect 11636 30612 11660 30668
rect 11716 30612 11740 30668
rect 11796 30612 11820 30668
rect 11876 30612 11900 30668
rect 11956 30612 11980 30668
rect 12036 30612 12060 30668
rect 12116 30612 12140 30668
rect 12196 30612 12220 30668
rect 12276 30612 12300 30668
rect 12356 30612 12380 30668
rect 12436 30612 12460 30668
rect 12516 30612 12540 30668
rect 12596 30612 12620 30668
rect 12676 30612 12700 30668
rect 12756 30612 12780 30668
rect 12836 30612 12860 30668
rect 12916 30612 12940 30668
rect 12996 30612 13020 30668
rect 13076 30614 14514 30668
rect 14570 30614 14594 30670
rect 14650 30614 14674 30670
rect 14730 30614 14754 30670
rect 14810 30614 14834 30670
rect 14890 30614 14914 30670
rect 14970 30614 14994 30670
rect 15050 30614 15074 30670
rect 15130 30614 15154 30670
rect 15210 30614 15234 30670
rect 15290 30614 15298 30670
rect 13076 30612 15298 30614
rect 6135 30605 15298 30612
rect 1694 30587 15298 30605
rect 1694 30586 14514 30587
rect 1694 30585 6182 30586
rect 1694 30529 2139 30585
rect 2195 30529 2237 30585
rect 2293 30529 2335 30585
rect 2391 30529 2433 30585
rect 2489 30578 6182 30585
rect 2489 30529 5803 30578
rect 1694 30522 5803 30529
rect 5859 30522 5895 30578
rect 5951 30522 5987 30578
rect 6043 30522 6079 30578
rect 6135 30530 6182 30578
rect 6238 30530 6263 30586
rect 6319 30530 6344 30586
rect 6400 30530 6425 30586
rect 6481 30530 6506 30586
rect 6562 30530 6587 30586
rect 6643 30530 6668 30586
rect 6724 30530 6749 30586
rect 6805 30530 6830 30586
rect 6886 30530 6911 30586
rect 6967 30530 6992 30586
rect 7048 30530 7073 30586
rect 7129 30530 7154 30586
rect 7210 30530 7235 30586
rect 7291 30530 7316 30586
rect 7372 30530 7397 30586
rect 7453 30530 7478 30586
rect 7534 30530 7559 30586
rect 7615 30530 7640 30586
rect 7696 30530 7721 30586
rect 7777 30530 7802 30586
rect 7858 30530 7883 30586
rect 7939 30530 7964 30586
rect 8020 30530 8045 30586
rect 8101 30530 8126 30586
rect 8182 30530 8207 30586
rect 8263 30530 8288 30586
rect 8344 30530 8369 30586
rect 8425 30530 8450 30586
rect 8506 30530 8531 30586
rect 8587 30530 8612 30586
rect 8668 30530 8693 30586
rect 8749 30530 8774 30586
rect 8830 30530 8855 30586
rect 8911 30530 8936 30586
rect 8992 30530 9017 30586
rect 9073 30530 9098 30586
rect 9154 30530 9179 30586
rect 9235 30530 9260 30586
rect 9316 30530 9340 30586
rect 9396 30530 9420 30586
rect 9476 30530 9500 30586
rect 9556 30530 9580 30586
rect 9636 30530 9660 30586
rect 9716 30530 9740 30586
rect 9796 30530 9820 30586
rect 9876 30530 9900 30586
rect 9956 30530 9980 30586
rect 10036 30530 10060 30586
rect 10116 30530 10140 30586
rect 10196 30530 10220 30586
rect 10276 30530 10300 30586
rect 10356 30530 10380 30586
rect 10436 30530 10460 30586
rect 10516 30530 10540 30586
rect 10596 30530 10620 30586
rect 10676 30530 10700 30586
rect 10756 30530 10780 30586
rect 10836 30530 10860 30586
rect 10916 30530 10940 30586
rect 10996 30530 11020 30586
rect 11076 30530 11100 30586
rect 11156 30530 11180 30586
rect 11236 30530 11260 30586
rect 11316 30530 11340 30586
rect 11396 30530 11420 30586
rect 11476 30530 11500 30586
rect 11556 30530 11580 30586
rect 11636 30530 11660 30586
rect 11716 30530 11740 30586
rect 11796 30530 11820 30586
rect 11876 30530 11900 30586
rect 11956 30530 11980 30586
rect 12036 30530 12060 30586
rect 12116 30530 12140 30586
rect 12196 30530 12220 30586
rect 12276 30530 12300 30586
rect 12356 30530 12380 30586
rect 12436 30530 12460 30586
rect 12516 30530 12540 30586
rect 12596 30530 12620 30586
rect 12676 30530 12700 30586
rect 12756 30530 12780 30586
rect 12836 30530 12860 30586
rect 12916 30530 12940 30586
rect 12996 30530 13020 30586
rect 13076 30531 14514 30586
rect 14570 30531 14594 30587
rect 14650 30531 14674 30587
rect 14730 30531 14754 30587
rect 14810 30531 14834 30587
rect 14890 30531 14914 30587
rect 14970 30531 14994 30587
rect 15050 30531 15074 30587
rect 15130 30531 15154 30587
rect 15210 30531 15234 30587
rect 15290 30531 15298 30587
rect 13076 30530 15298 30531
rect 6135 30522 15298 30530
rect 1694 30504 15298 30522
rect 1694 30503 6182 30504
rect 1694 30447 2139 30503
rect 2195 30447 2237 30503
rect 2293 30447 2335 30503
rect 2391 30447 2433 30503
rect 2489 30496 6182 30503
rect 2489 30447 5803 30496
rect 1694 30440 5803 30447
rect 5859 30440 5895 30496
rect 5951 30440 5987 30496
rect 6043 30440 6079 30496
rect 6135 30448 6182 30496
rect 6238 30448 6263 30504
rect 6319 30448 6344 30504
rect 6400 30448 6425 30504
rect 6481 30448 6506 30504
rect 6562 30448 6587 30504
rect 6643 30448 6668 30504
rect 6724 30448 6749 30504
rect 6805 30448 6830 30504
rect 6886 30448 6911 30504
rect 6967 30448 6992 30504
rect 7048 30448 7073 30504
rect 7129 30448 7154 30504
rect 7210 30448 7235 30504
rect 7291 30448 7316 30504
rect 7372 30448 7397 30504
rect 7453 30448 7478 30504
rect 7534 30448 7559 30504
rect 7615 30448 7640 30504
rect 7696 30448 7721 30504
rect 7777 30448 7802 30504
rect 7858 30448 7883 30504
rect 7939 30448 7964 30504
rect 8020 30448 8045 30504
rect 8101 30448 8126 30504
rect 8182 30448 8207 30504
rect 8263 30448 8288 30504
rect 8344 30448 8369 30504
rect 8425 30448 8450 30504
rect 8506 30448 8531 30504
rect 8587 30448 8612 30504
rect 8668 30448 8693 30504
rect 8749 30448 8774 30504
rect 8830 30448 8855 30504
rect 8911 30448 8936 30504
rect 8992 30448 9017 30504
rect 9073 30448 9098 30504
rect 9154 30448 9179 30504
rect 9235 30448 9260 30504
rect 9316 30448 9340 30504
rect 9396 30448 9420 30504
rect 9476 30448 9500 30504
rect 9556 30448 9580 30504
rect 9636 30448 9660 30504
rect 9716 30448 9740 30504
rect 9796 30448 9820 30504
rect 9876 30448 9900 30504
rect 9956 30448 9980 30504
rect 10036 30448 10060 30504
rect 10116 30448 10140 30504
rect 10196 30448 10220 30504
rect 10276 30448 10300 30504
rect 10356 30448 10380 30504
rect 10436 30448 10460 30504
rect 10516 30448 10540 30504
rect 10596 30448 10620 30504
rect 10676 30448 10700 30504
rect 10756 30448 10780 30504
rect 10836 30448 10860 30504
rect 10916 30448 10940 30504
rect 10996 30448 11020 30504
rect 11076 30448 11100 30504
rect 11156 30448 11180 30504
rect 11236 30448 11260 30504
rect 11316 30448 11340 30504
rect 11396 30448 11420 30504
rect 11476 30448 11500 30504
rect 11556 30448 11580 30504
rect 11636 30448 11660 30504
rect 11716 30448 11740 30504
rect 11796 30448 11820 30504
rect 11876 30448 11900 30504
rect 11956 30448 11980 30504
rect 12036 30448 12060 30504
rect 12116 30448 12140 30504
rect 12196 30448 12220 30504
rect 12276 30448 12300 30504
rect 12356 30448 12380 30504
rect 12436 30448 12460 30504
rect 12516 30448 12540 30504
rect 12596 30448 12620 30504
rect 12676 30448 12700 30504
rect 12756 30448 12780 30504
rect 12836 30448 12860 30504
rect 12916 30448 12940 30504
rect 12996 30448 13020 30504
rect 13076 30448 14514 30504
rect 14570 30448 14594 30504
rect 14650 30448 14674 30504
rect 14730 30448 14754 30504
rect 14810 30448 14834 30504
rect 14890 30448 14914 30504
rect 14970 30448 14994 30504
rect 15050 30448 15074 30504
rect 15130 30448 15154 30504
rect 15210 30448 15234 30504
rect 15290 30448 15298 30504
rect 6135 30440 15298 30448
rect 1694 30422 15298 30440
rect 1694 30421 6182 30422
rect 1694 30365 2139 30421
rect 2195 30365 2237 30421
rect 2293 30365 2335 30421
rect 2391 30365 2433 30421
rect 2489 30414 6182 30421
rect 2489 30365 5803 30414
rect 1694 30358 5803 30365
rect 5859 30358 5895 30414
rect 5951 30358 5987 30414
rect 6043 30358 6079 30414
rect 6135 30366 6182 30414
rect 6238 30366 6263 30422
rect 6319 30366 6344 30422
rect 6400 30366 6425 30422
rect 6481 30366 6506 30422
rect 6562 30366 6587 30422
rect 6643 30366 6668 30422
rect 6724 30366 6749 30422
rect 6805 30366 6830 30422
rect 6886 30366 6911 30422
rect 6967 30366 6992 30422
rect 7048 30366 7073 30422
rect 7129 30366 7154 30422
rect 7210 30366 7235 30422
rect 7291 30366 7316 30422
rect 7372 30366 7397 30422
rect 7453 30366 7478 30422
rect 7534 30366 7559 30422
rect 7615 30366 7640 30422
rect 7696 30366 7721 30422
rect 7777 30366 7802 30422
rect 7858 30366 7883 30422
rect 7939 30366 7964 30422
rect 8020 30366 8045 30422
rect 8101 30366 8126 30422
rect 8182 30366 8207 30422
rect 8263 30366 8288 30422
rect 8344 30366 8369 30422
rect 8425 30366 8450 30422
rect 8506 30366 8531 30422
rect 8587 30366 8612 30422
rect 8668 30366 8693 30422
rect 8749 30366 8774 30422
rect 8830 30366 8855 30422
rect 8911 30366 8936 30422
rect 8992 30366 9017 30422
rect 9073 30366 9098 30422
rect 9154 30366 9179 30422
rect 9235 30366 9260 30422
rect 9316 30366 9340 30422
rect 9396 30366 9420 30422
rect 9476 30366 9500 30422
rect 9556 30366 9580 30422
rect 9636 30366 9660 30422
rect 9716 30366 9740 30422
rect 9796 30366 9820 30422
rect 9876 30366 9900 30422
rect 9956 30366 9980 30422
rect 10036 30366 10060 30422
rect 10116 30366 10140 30422
rect 10196 30366 10220 30422
rect 10276 30366 10300 30422
rect 10356 30366 10380 30422
rect 10436 30366 10460 30422
rect 10516 30366 10540 30422
rect 10596 30366 10620 30422
rect 10676 30366 10700 30422
rect 10756 30366 10780 30422
rect 10836 30366 10860 30422
rect 10916 30366 10940 30422
rect 10996 30366 11020 30422
rect 11076 30366 11100 30422
rect 11156 30366 11180 30422
rect 11236 30366 11260 30422
rect 11316 30366 11340 30422
rect 11396 30366 11420 30422
rect 11476 30366 11500 30422
rect 11556 30366 11580 30422
rect 11636 30366 11660 30422
rect 11716 30366 11740 30422
rect 11796 30366 11820 30422
rect 11876 30366 11900 30422
rect 11956 30366 11980 30422
rect 12036 30366 12060 30422
rect 12116 30366 12140 30422
rect 12196 30366 12220 30422
rect 12276 30366 12300 30422
rect 12356 30366 12380 30422
rect 12436 30366 12460 30422
rect 12516 30366 12540 30422
rect 12596 30366 12620 30422
rect 12676 30366 12700 30422
rect 12756 30366 12780 30422
rect 12836 30366 12860 30422
rect 12916 30366 12940 30422
rect 12996 30366 13020 30422
rect 13076 30421 15298 30422
rect 13076 30366 14514 30421
rect 6135 30365 14514 30366
rect 14570 30365 14594 30421
rect 14650 30365 14674 30421
rect 14730 30365 14754 30421
rect 14810 30365 14834 30421
rect 14890 30365 14914 30421
rect 14970 30365 14994 30421
rect 15050 30365 15074 30421
rect 15130 30365 15154 30421
rect 15210 30365 15234 30421
rect 15290 30365 15298 30421
rect 6135 30358 15298 30365
rect 1694 30340 15298 30358
rect 1694 30338 6182 30340
rect 1694 30282 2139 30338
rect 2195 30282 2237 30338
rect 2293 30282 2335 30338
rect 2391 30282 2433 30338
rect 2489 30332 6182 30338
rect 2489 30282 5803 30332
rect 1694 30276 5803 30282
rect 5859 30276 5895 30332
rect 5951 30276 5987 30332
rect 6043 30276 6079 30332
rect 6135 30284 6182 30332
rect 6238 30284 6263 30340
rect 6319 30284 6344 30340
rect 6400 30284 6425 30340
rect 6481 30284 6506 30340
rect 6562 30284 6587 30340
rect 6643 30284 6668 30340
rect 6724 30284 6749 30340
rect 6805 30284 6830 30340
rect 6886 30284 6911 30340
rect 6967 30284 6992 30340
rect 7048 30284 7073 30340
rect 7129 30284 7154 30340
rect 7210 30284 7235 30340
rect 7291 30284 7316 30340
rect 7372 30284 7397 30340
rect 7453 30284 7478 30340
rect 7534 30284 7559 30340
rect 7615 30284 7640 30340
rect 7696 30284 7721 30340
rect 7777 30284 7802 30340
rect 7858 30284 7883 30340
rect 7939 30284 7964 30340
rect 8020 30284 8045 30340
rect 8101 30284 8126 30340
rect 8182 30284 8207 30340
rect 8263 30284 8288 30340
rect 8344 30284 8369 30340
rect 8425 30284 8450 30340
rect 8506 30284 8531 30340
rect 8587 30284 8612 30340
rect 8668 30284 8693 30340
rect 8749 30284 8774 30340
rect 8830 30284 8855 30340
rect 8911 30284 8936 30340
rect 8992 30284 9017 30340
rect 9073 30284 9098 30340
rect 9154 30284 9179 30340
rect 9235 30284 9260 30340
rect 9316 30284 9340 30340
rect 9396 30284 9420 30340
rect 9476 30284 9500 30340
rect 9556 30284 9580 30340
rect 9636 30284 9660 30340
rect 9716 30284 9740 30340
rect 9796 30284 9820 30340
rect 9876 30284 9900 30340
rect 9956 30284 9980 30340
rect 10036 30284 10060 30340
rect 10116 30284 10140 30340
rect 10196 30284 10220 30340
rect 10276 30284 10300 30340
rect 10356 30284 10380 30340
rect 10436 30284 10460 30340
rect 10516 30284 10540 30340
rect 10596 30284 10620 30340
rect 10676 30284 10700 30340
rect 10756 30284 10780 30340
rect 10836 30284 10860 30340
rect 10916 30284 10940 30340
rect 10996 30284 11020 30340
rect 11076 30284 11100 30340
rect 11156 30284 11180 30340
rect 11236 30284 11260 30340
rect 11316 30284 11340 30340
rect 11396 30284 11420 30340
rect 11476 30284 11500 30340
rect 11556 30284 11580 30340
rect 11636 30284 11660 30340
rect 11716 30284 11740 30340
rect 11796 30284 11820 30340
rect 11876 30284 11900 30340
rect 11956 30284 11980 30340
rect 12036 30284 12060 30340
rect 12116 30284 12140 30340
rect 12196 30284 12220 30340
rect 12276 30284 12300 30340
rect 12356 30284 12380 30340
rect 12436 30284 12460 30340
rect 12516 30284 12540 30340
rect 12596 30284 12620 30340
rect 12676 30284 12700 30340
rect 12756 30284 12780 30340
rect 12836 30284 12860 30340
rect 12916 30284 12940 30340
rect 12996 30284 13020 30340
rect 13076 30338 15298 30340
rect 13076 30284 14514 30338
rect 6135 30282 14514 30284
rect 14570 30282 14594 30338
rect 14650 30282 14674 30338
rect 14730 30282 14754 30338
rect 14810 30282 14834 30338
rect 14890 30282 14914 30338
rect 14970 30282 14994 30338
rect 15050 30282 15074 30338
rect 15130 30282 15154 30338
rect 15210 30282 15234 30338
rect 15290 30282 15298 30338
rect 6135 30276 15298 30282
rect 1694 30258 15298 30276
rect 1694 30255 6182 30258
rect 1694 30199 2139 30255
rect 2195 30199 2237 30255
rect 2293 30199 2335 30255
rect 2391 30199 2433 30255
rect 2489 30250 6182 30255
rect 2489 30199 5803 30250
rect 1694 30194 5803 30199
rect 5859 30194 5895 30250
rect 5951 30194 5987 30250
rect 6043 30194 6079 30250
rect 6135 30202 6182 30250
rect 6238 30202 6263 30258
rect 6319 30202 6344 30258
rect 6400 30202 6425 30258
rect 6481 30202 6506 30258
rect 6562 30202 6587 30258
rect 6643 30202 6668 30258
rect 6724 30202 6749 30258
rect 6805 30202 6830 30258
rect 6886 30202 6911 30258
rect 6967 30202 6992 30258
rect 7048 30202 7073 30258
rect 7129 30202 7154 30258
rect 7210 30202 7235 30258
rect 7291 30202 7316 30258
rect 7372 30202 7397 30258
rect 7453 30202 7478 30258
rect 7534 30202 7559 30258
rect 7615 30202 7640 30258
rect 7696 30202 7721 30258
rect 7777 30202 7802 30258
rect 7858 30202 7883 30258
rect 7939 30202 7964 30258
rect 8020 30202 8045 30258
rect 8101 30202 8126 30258
rect 8182 30202 8207 30258
rect 8263 30202 8288 30258
rect 8344 30202 8369 30258
rect 8425 30202 8450 30258
rect 8506 30202 8531 30258
rect 8587 30202 8612 30258
rect 8668 30202 8693 30258
rect 8749 30202 8774 30258
rect 8830 30202 8855 30258
rect 8911 30202 8936 30258
rect 8992 30202 9017 30258
rect 9073 30202 9098 30258
rect 9154 30202 9179 30258
rect 9235 30202 9260 30258
rect 9316 30202 9340 30258
rect 9396 30202 9420 30258
rect 9476 30202 9500 30258
rect 9556 30202 9580 30258
rect 9636 30202 9660 30258
rect 9716 30202 9740 30258
rect 9796 30202 9820 30258
rect 9876 30202 9900 30258
rect 9956 30202 9980 30258
rect 10036 30202 10060 30258
rect 10116 30202 10140 30258
rect 10196 30202 10220 30258
rect 10276 30202 10300 30258
rect 10356 30202 10380 30258
rect 10436 30202 10460 30258
rect 10516 30202 10540 30258
rect 10596 30202 10620 30258
rect 10676 30202 10700 30258
rect 10756 30202 10780 30258
rect 10836 30202 10860 30258
rect 10916 30202 10940 30258
rect 10996 30202 11020 30258
rect 11076 30202 11100 30258
rect 11156 30202 11180 30258
rect 11236 30202 11260 30258
rect 11316 30202 11340 30258
rect 11396 30202 11420 30258
rect 11476 30202 11500 30258
rect 11556 30202 11580 30258
rect 11636 30202 11660 30258
rect 11716 30202 11740 30258
rect 11796 30202 11820 30258
rect 11876 30202 11900 30258
rect 11956 30202 11980 30258
rect 12036 30202 12060 30258
rect 12116 30202 12140 30258
rect 12196 30202 12220 30258
rect 12276 30202 12300 30258
rect 12356 30202 12380 30258
rect 12436 30202 12460 30258
rect 12516 30202 12540 30258
rect 12596 30202 12620 30258
rect 12676 30202 12700 30258
rect 12756 30202 12780 30258
rect 12836 30202 12860 30258
rect 12916 30202 12940 30258
rect 12996 30202 13020 30258
rect 13076 30255 15298 30258
rect 13076 30202 14514 30255
rect 6135 30199 14514 30202
rect 14570 30199 14594 30255
rect 14650 30199 14674 30255
rect 14730 30199 14754 30255
rect 14810 30199 14834 30255
rect 14890 30199 14914 30255
rect 14970 30199 14994 30255
rect 15050 30199 15074 30255
rect 15130 30199 15154 30255
rect 15210 30199 15234 30255
rect 15290 30199 15298 30255
rect 6135 30194 15298 30199
rect 1694 30172 15298 30194
rect 1694 30116 2139 30172
rect 2195 30116 2237 30172
rect 2293 30116 2335 30172
rect 2391 30116 2433 30172
rect 2489 30116 14514 30172
rect 14570 30116 14594 30172
rect 14650 30116 14674 30172
rect 14730 30116 14754 30172
rect 14810 30116 14834 30172
rect 14890 30116 14914 30172
rect 14970 30116 14994 30172
rect 15050 30116 15074 30172
rect 15130 30116 15154 30172
rect 15210 30116 15234 30172
rect 15290 30116 15298 30172
rect 1694 30089 15298 30116
rect 1694 30033 2139 30089
rect 2195 30033 2237 30089
rect 2293 30033 2335 30089
rect 2391 30033 2433 30089
rect 2489 30033 14514 30089
rect 14570 30033 14594 30089
rect 14650 30033 14674 30089
rect 14730 30033 14754 30089
rect 14810 30033 14834 30089
rect 14890 30033 14914 30089
rect 14970 30033 14994 30089
rect 15050 30033 15074 30089
rect 15130 30033 15154 30089
rect 15210 30033 15234 30089
rect 15290 30033 15298 30089
rect 1694 30006 15298 30033
rect 1694 29950 2139 30006
rect 2195 29950 2237 30006
rect 2293 29950 2335 30006
rect 2391 29950 2433 30006
rect 2489 29950 14514 30006
rect 14570 29950 14594 30006
rect 14650 29950 14674 30006
rect 14730 29950 14754 30006
rect 14810 29950 14834 30006
rect 14890 29950 14914 30006
rect 14970 29950 14994 30006
rect 15050 29950 15074 30006
rect 15130 29950 15154 30006
rect 15210 29950 15234 30006
rect 15290 29950 15298 30006
rect 1694 29923 15298 29950
rect 1694 29891 2139 29923
tri 1694 29447 2138 29891 ne
rect 2138 29867 2139 29891
rect 2195 29867 2237 29923
rect 2293 29867 2335 29923
rect 2391 29867 2433 29923
rect 2489 29883 14514 29923
rect 2489 29867 5803 29883
rect 2138 29840 5803 29867
rect 2138 29784 2139 29840
rect 2195 29784 2237 29840
rect 2293 29784 2335 29840
rect 2391 29784 2433 29840
rect 2489 29827 5803 29840
rect 5859 29827 5895 29883
rect 5951 29827 5987 29883
rect 6043 29827 6079 29883
rect 6135 29880 14514 29883
rect 6135 29827 6182 29880
rect 2489 29824 6182 29827
rect 6238 29824 6263 29880
rect 6319 29824 6344 29880
rect 6400 29824 6425 29880
rect 6481 29824 6506 29880
rect 6562 29824 6587 29880
rect 6643 29824 6668 29880
rect 6724 29824 6749 29880
rect 6805 29824 6830 29880
rect 6886 29824 6911 29880
rect 6967 29824 6992 29880
rect 7048 29824 7073 29880
rect 7129 29824 7154 29880
rect 7210 29824 7235 29880
rect 7291 29824 7316 29880
rect 7372 29824 7397 29880
rect 7453 29824 7478 29880
rect 7534 29824 7559 29880
rect 7615 29824 7640 29880
rect 7696 29824 7721 29880
rect 7777 29824 7802 29880
rect 7858 29824 7883 29880
rect 7939 29824 7964 29880
rect 8020 29824 8045 29880
rect 8101 29824 8126 29880
rect 8182 29824 8207 29880
rect 8263 29824 8288 29880
rect 8344 29824 8369 29880
rect 8425 29824 8450 29880
rect 8506 29824 8531 29880
rect 8587 29824 8612 29880
rect 8668 29824 8693 29880
rect 8749 29824 8774 29880
rect 8830 29824 8855 29880
rect 8911 29824 8936 29880
rect 8992 29824 9017 29880
rect 9073 29824 9098 29880
rect 9154 29824 9179 29880
rect 9235 29824 9260 29880
rect 2489 29801 9260 29824
rect 2489 29784 5803 29801
rect 2138 29757 5803 29784
rect 2138 29701 2139 29757
rect 2195 29701 2237 29757
rect 2293 29701 2335 29757
rect 2391 29701 2433 29757
rect 2489 29745 5803 29757
rect 5859 29745 5895 29801
rect 5951 29745 5987 29801
rect 6043 29745 6079 29801
rect 6135 29800 9260 29801
rect 6135 29745 6182 29800
rect 2489 29744 6182 29745
rect 6238 29744 6263 29800
rect 6319 29744 6344 29800
rect 6400 29744 6425 29800
rect 6481 29744 6506 29800
rect 6562 29744 6587 29800
rect 6643 29744 6668 29800
rect 6724 29744 6749 29800
rect 6805 29744 6830 29800
rect 6886 29744 6911 29800
rect 6967 29744 6992 29800
rect 7048 29744 7073 29800
rect 7129 29744 7154 29800
rect 7210 29744 7235 29800
rect 7291 29744 7316 29800
rect 7372 29744 7397 29800
rect 7453 29744 7478 29800
rect 7534 29744 7559 29800
rect 7615 29744 7640 29800
rect 7696 29744 7721 29800
rect 7777 29744 7802 29800
rect 7858 29744 7883 29800
rect 7939 29744 7964 29800
rect 8020 29744 8045 29800
rect 8101 29744 8126 29800
rect 8182 29744 8207 29800
rect 8263 29744 8288 29800
rect 8344 29744 8369 29800
rect 8425 29744 8450 29800
rect 8506 29744 8531 29800
rect 8587 29744 8612 29800
rect 8668 29744 8693 29800
rect 8749 29744 8774 29800
rect 8830 29744 8855 29800
rect 8911 29744 8936 29800
rect 8992 29744 9017 29800
rect 9073 29744 9098 29800
rect 9154 29744 9179 29800
rect 9235 29744 9260 29800
rect 2489 29720 9260 29744
rect 2489 29719 6182 29720
rect 2489 29701 5803 29719
rect 2138 29674 5803 29701
rect 2138 29618 2139 29674
rect 2195 29618 2237 29674
rect 2293 29618 2335 29674
rect 2391 29618 2433 29674
rect 2489 29663 5803 29674
rect 5859 29663 5895 29719
rect 5951 29663 5987 29719
rect 6043 29663 6079 29719
rect 6135 29664 6182 29719
rect 6238 29664 6263 29720
rect 6319 29664 6344 29720
rect 6400 29664 6425 29720
rect 6481 29664 6506 29720
rect 6562 29664 6587 29720
rect 6643 29664 6668 29720
rect 6724 29664 6749 29720
rect 6805 29664 6830 29720
rect 6886 29664 6911 29720
rect 6967 29664 6992 29720
rect 7048 29664 7073 29720
rect 7129 29664 7154 29720
rect 7210 29664 7235 29720
rect 7291 29664 7316 29720
rect 7372 29664 7397 29720
rect 7453 29664 7478 29720
rect 7534 29664 7559 29720
rect 7615 29664 7640 29720
rect 7696 29664 7721 29720
rect 7777 29664 7802 29720
rect 7858 29664 7883 29720
rect 7939 29664 7964 29720
rect 8020 29664 8045 29720
rect 8101 29664 8126 29720
rect 8182 29664 8207 29720
rect 8263 29664 8288 29720
rect 8344 29664 8369 29720
rect 8425 29664 8450 29720
rect 8506 29664 8531 29720
rect 8587 29664 8612 29720
rect 8668 29664 8693 29720
rect 8749 29664 8774 29720
rect 8830 29664 8855 29720
rect 8911 29664 8936 29720
rect 8992 29664 9017 29720
rect 9073 29664 9098 29720
rect 9154 29664 9179 29720
rect 9235 29664 9260 29720
rect 6135 29663 9260 29664
rect 2489 29640 9260 29663
rect 2489 29637 6182 29640
rect 2489 29618 5803 29637
rect 2138 29591 5803 29618
rect 2138 29535 2139 29591
rect 2195 29535 2237 29591
rect 2293 29535 2335 29591
rect 2391 29535 2433 29591
rect 2489 29581 5803 29591
rect 5859 29581 5895 29637
rect 5951 29581 5987 29637
rect 6043 29581 6079 29637
rect 6135 29584 6182 29637
rect 6238 29584 6263 29640
rect 6319 29584 6344 29640
rect 6400 29584 6425 29640
rect 6481 29584 6506 29640
rect 6562 29584 6587 29640
rect 6643 29584 6668 29640
rect 6724 29584 6749 29640
rect 6805 29584 6830 29640
rect 6886 29584 6911 29640
rect 6967 29584 6992 29640
rect 7048 29584 7073 29640
rect 7129 29584 7154 29640
rect 7210 29584 7235 29640
rect 7291 29584 7316 29640
rect 7372 29584 7397 29640
rect 7453 29584 7478 29640
rect 7534 29584 7559 29640
rect 7615 29584 7640 29640
rect 7696 29584 7721 29640
rect 7777 29584 7802 29640
rect 7858 29584 7883 29640
rect 7939 29584 7964 29640
rect 8020 29584 8045 29640
rect 8101 29584 8126 29640
rect 8182 29584 8207 29640
rect 8263 29584 8288 29640
rect 8344 29584 8369 29640
rect 8425 29584 8450 29640
rect 8506 29584 8531 29640
rect 8587 29584 8612 29640
rect 8668 29584 8693 29640
rect 8749 29584 8774 29640
rect 8830 29584 8855 29640
rect 8911 29584 8936 29640
rect 8992 29584 9017 29640
rect 9073 29584 9098 29640
rect 9154 29584 9179 29640
rect 9235 29584 9260 29640
rect 6135 29581 9260 29584
rect 2489 29560 9260 29581
rect 2489 29555 6182 29560
rect 2489 29535 5803 29555
rect 2138 29508 5803 29535
rect 2138 29452 2139 29508
rect 2195 29452 2237 29508
rect 2293 29452 2335 29508
rect 2391 29452 2433 29508
rect 2489 29499 5803 29508
rect 5859 29499 5895 29555
rect 5951 29499 5987 29555
rect 6043 29499 6079 29555
rect 6135 29504 6182 29555
rect 6238 29504 6263 29560
rect 6319 29504 6344 29560
rect 6400 29504 6425 29560
rect 6481 29504 6506 29560
rect 6562 29504 6587 29560
rect 6643 29504 6668 29560
rect 6724 29504 6749 29560
rect 6805 29504 6830 29560
rect 6886 29504 6911 29560
rect 6967 29504 6992 29560
rect 7048 29504 7073 29560
rect 7129 29504 7154 29560
rect 7210 29504 7235 29560
rect 7291 29504 7316 29560
rect 7372 29504 7397 29560
rect 7453 29504 7478 29560
rect 7534 29504 7559 29560
rect 7615 29504 7640 29560
rect 7696 29504 7721 29560
rect 7777 29504 7802 29560
rect 7858 29504 7883 29560
rect 7939 29504 7964 29560
rect 8020 29504 8045 29560
rect 8101 29504 8126 29560
rect 8182 29504 8207 29560
rect 8263 29504 8288 29560
rect 8344 29504 8369 29560
rect 8425 29504 8450 29560
rect 8506 29504 8531 29560
rect 8587 29504 8612 29560
rect 8668 29504 8693 29560
rect 8749 29504 8774 29560
rect 8830 29504 8855 29560
rect 8911 29504 8936 29560
rect 8992 29504 9017 29560
rect 9073 29504 9098 29560
rect 9154 29504 9179 29560
rect 9235 29504 9260 29560
rect 6135 29499 9260 29504
rect 2489 29480 9260 29499
rect 2489 29472 6182 29480
rect 2489 29452 5803 29472
rect 148 29423 654 29427
rect 148 29414 298 29423
rect 148 29362 149 29414
rect 201 29362 247 29414
rect 354 29367 396 29423
rect 452 29414 494 29423
rect 550 29414 592 29423
rect 648 29414 654 29423
rect 452 29367 454 29414
rect 580 29367 592 29414
rect 299 29362 454 29367
rect 506 29362 528 29367
rect 580 29362 602 29367
rect 148 29349 654 29362
rect 148 29297 149 29349
rect 201 29297 247 29349
rect 299 29342 454 29349
rect 506 29342 528 29349
rect 580 29342 602 29349
rect 148 29286 298 29297
rect 354 29286 396 29342
rect 452 29297 454 29342
rect 580 29297 592 29342
rect 452 29286 494 29297
rect 550 29286 592 29297
rect 648 29286 654 29297
rect 148 29284 654 29286
rect 148 29232 149 29284
rect 201 29232 247 29284
rect 299 29261 454 29284
rect 506 29261 528 29284
rect 580 29261 602 29284
rect 148 29219 298 29232
rect 148 29167 149 29219
rect 201 29167 247 29219
rect 354 29205 396 29261
rect 452 29232 454 29261
rect 580 29232 592 29261
rect 452 29219 494 29232
rect 550 29219 592 29232
rect 648 29219 654 29232
rect 452 29205 454 29219
rect 580 29205 592 29219
rect 299 29180 454 29205
rect 506 29180 528 29205
rect 580 29180 602 29205
rect 148 29154 298 29167
rect 148 29102 149 29154
rect 201 29102 247 29154
rect 354 29124 396 29180
rect 452 29167 454 29180
rect 580 29167 592 29180
rect 452 29154 494 29167
rect 550 29154 592 29167
rect 648 29154 654 29167
rect 452 29124 454 29154
rect 580 29124 592 29154
rect 299 29102 454 29124
rect 506 29102 528 29124
rect 580 29102 602 29124
rect 148 29099 654 29102
rect 148 29089 298 29099
rect 148 29037 149 29089
rect 201 29037 247 29089
rect 354 29043 396 29099
rect 452 29089 494 29099
rect 550 29089 592 29099
rect 648 29089 654 29099
rect 452 29043 454 29089
rect 580 29043 592 29089
rect 299 29037 454 29043
rect 506 29037 528 29043
rect 580 29037 602 29043
rect 148 28024 654 29037
rect 2138 29425 5803 29452
rect 2138 29369 2139 29425
rect 2195 29369 2237 29425
rect 2293 29369 2335 29425
rect 2391 29369 2433 29425
rect 2489 29416 5803 29425
rect 5859 29416 5895 29472
rect 5951 29416 5987 29472
rect 6043 29416 6079 29472
rect 6135 29424 6182 29472
rect 6238 29424 6263 29480
rect 6319 29424 6344 29480
rect 6400 29424 6425 29480
rect 6481 29424 6506 29480
rect 6562 29424 6587 29480
rect 6643 29424 6668 29480
rect 6724 29424 6749 29480
rect 6805 29424 6830 29480
rect 6886 29424 6911 29480
rect 6967 29424 6992 29480
rect 7048 29424 7073 29480
rect 7129 29424 7154 29480
rect 7210 29424 7235 29480
rect 7291 29424 7316 29480
rect 7372 29424 7397 29480
rect 7453 29424 7478 29480
rect 7534 29424 7559 29480
rect 7615 29424 7640 29480
rect 7696 29424 7721 29480
rect 7777 29424 7802 29480
rect 7858 29424 7883 29480
rect 7939 29424 7964 29480
rect 8020 29424 8045 29480
rect 8101 29424 8126 29480
rect 8182 29424 8207 29480
rect 8263 29424 8288 29480
rect 8344 29424 8369 29480
rect 8425 29424 8450 29480
rect 8506 29424 8531 29480
rect 8587 29424 8612 29480
rect 8668 29424 8693 29480
rect 8749 29424 8774 29480
rect 8830 29424 8855 29480
rect 8911 29424 8936 29480
rect 8992 29424 9017 29480
rect 9073 29424 9098 29480
rect 9154 29424 9179 29480
rect 9235 29424 9260 29480
rect 6135 29416 9260 29424
rect 2489 29400 9260 29416
rect 2489 29389 6182 29400
rect 2489 29369 5803 29389
rect 2138 29342 5803 29369
rect 2138 29286 2139 29342
rect 2195 29286 2237 29342
rect 2293 29286 2335 29342
rect 2391 29286 2433 29342
rect 2489 29333 5803 29342
rect 5859 29333 5895 29389
rect 5951 29333 5987 29389
rect 6043 29333 6079 29389
rect 6135 29344 6182 29389
rect 6238 29344 6263 29400
rect 6319 29344 6344 29400
rect 6400 29344 6425 29400
rect 6481 29344 6506 29400
rect 6562 29344 6587 29400
rect 6643 29344 6668 29400
rect 6724 29344 6749 29400
rect 6805 29344 6830 29400
rect 6886 29344 6911 29400
rect 6967 29344 6992 29400
rect 7048 29344 7073 29400
rect 7129 29344 7154 29400
rect 7210 29344 7235 29400
rect 7291 29344 7316 29400
rect 7372 29344 7397 29400
rect 7453 29344 7478 29400
rect 7534 29344 7559 29400
rect 7615 29344 7640 29400
rect 7696 29344 7721 29400
rect 7777 29344 7802 29400
rect 7858 29344 7883 29400
rect 7939 29344 7964 29400
rect 8020 29344 8045 29400
rect 8101 29344 8126 29400
rect 8182 29344 8207 29400
rect 8263 29344 8288 29400
rect 8344 29344 8369 29400
rect 8425 29344 8450 29400
rect 8506 29344 8531 29400
rect 8587 29344 8612 29400
rect 8668 29344 8693 29400
rect 8749 29344 8774 29400
rect 8830 29344 8855 29400
rect 8911 29344 8936 29400
rect 8992 29344 9017 29400
rect 9073 29344 9098 29400
rect 9154 29344 9179 29400
rect 9235 29344 9260 29400
rect 6135 29333 9260 29344
rect 2489 29320 9260 29333
rect 2489 29306 6182 29320
rect 2489 29286 5803 29306
rect 2138 29259 5803 29286
rect 2138 29203 2139 29259
rect 2195 29203 2237 29259
rect 2293 29203 2335 29259
rect 2391 29203 2433 29259
rect 2489 29250 5803 29259
rect 5859 29250 5895 29306
rect 5951 29250 5987 29306
rect 6043 29250 6079 29306
rect 6135 29264 6182 29306
rect 6238 29264 6263 29320
rect 6319 29264 6344 29320
rect 6400 29264 6425 29320
rect 6481 29264 6506 29320
rect 6562 29264 6587 29320
rect 6643 29264 6668 29320
rect 6724 29264 6749 29320
rect 6805 29264 6830 29320
rect 6886 29264 6911 29320
rect 6967 29264 6992 29320
rect 7048 29264 7073 29320
rect 7129 29264 7154 29320
rect 7210 29264 7235 29320
rect 7291 29264 7316 29320
rect 7372 29264 7397 29320
rect 7453 29264 7478 29320
rect 7534 29264 7559 29320
rect 7615 29264 7640 29320
rect 7696 29264 7721 29320
rect 7777 29264 7802 29320
rect 7858 29264 7883 29320
rect 7939 29264 7964 29320
rect 8020 29264 8045 29320
rect 8101 29264 8126 29320
rect 8182 29264 8207 29320
rect 8263 29264 8288 29320
rect 8344 29264 8369 29320
rect 8425 29264 8450 29320
rect 8506 29264 8531 29320
rect 8587 29264 8612 29320
rect 8668 29264 8693 29320
rect 8749 29264 8774 29320
rect 8830 29264 8855 29320
rect 8911 29264 8936 29320
rect 8992 29264 9017 29320
rect 9073 29264 9098 29320
rect 9154 29264 9179 29320
rect 9235 29264 9260 29320
rect 6135 29250 9260 29264
rect 2489 29240 9260 29250
rect 2489 29223 6182 29240
rect 2489 29203 5803 29223
rect 2138 29176 5803 29203
rect 2138 29120 2139 29176
rect 2195 29120 2237 29176
rect 2293 29120 2335 29176
rect 2391 29120 2433 29176
rect 2489 29167 5803 29176
rect 5859 29167 5895 29223
rect 5951 29167 5987 29223
rect 6043 29167 6079 29223
rect 6135 29184 6182 29223
rect 6238 29184 6263 29240
rect 6319 29184 6344 29240
rect 6400 29184 6425 29240
rect 6481 29184 6506 29240
rect 6562 29184 6587 29240
rect 6643 29184 6668 29240
rect 6724 29184 6749 29240
rect 6805 29184 6830 29240
rect 6886 29184 6911 29240
rect 6967 29184 6992 29240
rect 7048 29184 7073 29240
rect 7129 29184 7154 29240
rect 7210 29184 7235 29240
rect 7291 29184 7316 29240
rect 7372 29184 7397 29240
rect 7453 29184 7478 29240
rect 7534 29184 7559 29240
rect 7615 29184 7640 29240
rect 7696 29184 7721 29240
rect 7777 29184 7802 29240
rect 7858 29184 7883 29240
rect 7939 29184 7964 29240
rect 8020 29184 8045 29240
rect 8101 29184 8126 29240
rect 8182 29184 8207 29240
rect 8263 29184 8288 29240
rect 8344 29184 8369 29240
rect 8425 29184 8450 29240
rect 8506 29184 8531 29240
rect 8587 29184 8612 29240
rect 8668 29184 8693 29240
rect 8749 29184 8774 29240
rect 8830 29184 8855 29240
rect 8911 29184 8936 29240
rect 8992 29184 9017 29240
rect 9073 29184 9098 29240
rect 9154 29184 9179 29240
rect 9235 29184 9260 29240
rect 6135 29167 9260 29184
rect 2489 29160 9260 29167
rect 2489 29140 6182 29160
rect 2489 29120 5803 29140
rect 2138 29093 5803 29120
rect 2138 29037 2139 29093
rect 2195 29037 2237 29093
rect 2293 29037 2335 29093
rect 2391 29037 2433 29093
rect 2489 29084 5803 29093
rect 5859 29084 5895 29140
rect 5951 29084 5987 29140
rect 6043 29084 6079 29140
rect 6135 29104 6182 29140
rect 6238 29104 6263 29160
rect 6319 29104 6344 29160
rect 6400 29104 6425 29160
rect 6481 29104 6506 29160
rect 6562 29104 6587 29160
rect 6643 29104 6668 29160
rect 6724 29104 6749 29160
rect 6805 29104 6830 29160
rect 6886 29104 6911 29160
rect 6967 29104 6992 29160
rect 7048 29104 7073 29160
rect 7129 29104 7154 29160
rect 7210 29104 7235 29160
rect 7291 29104 7316 29160
rect 7372 29104 7397 29160
rect 7453 29104 7478 29160
rect 7534 29104 7559 29160
rect 7615 29104 7640 29160
rect 7696 29104 7721 29160
rect 7777 29104 7802 29160
rect 7858 29104 7883 29160
rect 7939 29104 7964 29160
rect 8020 29104 8045 29160
rect 8101 29104 8126 29160
rect 8182 29104 8207 29160
rect 8263 29104 8288 29160
rect 8344 29104 8369 29160
rect 8425 29104 8450 29160
rect 8506 29104 8531 29160
rect 8587 29104 8612 29160
rect 8668 29104 8693 29160
rect 8749 29104 8774 29160
rect 8830 29104 8855 29160
rect 8911 29104 8936 29160
rect 8992 29104 9017 29160
rect 9073 29104 9098 29160
rect 9154 29104 9179 29160
rect 9235 29104 9260 29160
rect 6135 29084 9260 29104
rect 2489 29080 9260 29084
rect 2489 29037 6182 29080
rect 2138 29024 6182 29037
rect 6238 29024 6263 29080
rect 6319 29024 6344 29080
rect 6400 29024 6425 29080
rect 6481 29024 6506 29080
rect 6562 29024 6587 29080
rect 6643 29024 6668 29080
rect 6724 29024 6749 29080
rect 6805 29024 6830 29080
rect 6886 29024 6911 29080
rect 6967 29024 6992 29080
rect 7048 29024 7073 29080
rect 7129 29024 7154 29080
rect 7210 29024 7235 29080
rect 7291 29024 7316 29080
rect 7372 29024 7397 29080
rect 7453 29024 7478 29080
rect 7534 29024 7559 29080
rect 7615 29024 7640 29080
rect 7696 29024 7721 29080
rect 7777 29024 7802 29080
rect 7858 29024 7883 29080
rect 7939 29024 7964 29080
rect 8020 29024 8045 29080
rect 8101 29024 8126 29080
rect 8182 29024 8207 29080
rect 8263 29024 8288 29080
rect 8344 29024 8369 29080
rect 8425 29024 8450 29080
rect 8506 29024 8531 29080
rect 8587 29024 8612 29080
rect 8668 29024 8693 29080
rect 8749 29024 8774 29080
rect 8830 29024 8855 29080
rect 8911 29024 8936 29080
rect 8992 29024 9017 29080
rect 9073 29024 9098 29080
rect 9154 29024 9179 29080
rect 9235 29024 9260 29080
rect 2138 29010 9260 29024
rect 2138 28954 2139 29010
rect 2195 28954 2237 29010
rect 2293 28954 2335 29010
rect 2391 28954 2433 29010
rect 2489 29000 9260 29010
rect 2489 28954 6182 29000
rect 2138 28944 6182 28954
rect 6238 28944 6263 29000
rect 6319 28944 6344 29000
rect 6400 28944 6425 29000
rect 6481 28944 6506 29000
rect 6562 28944 6587 29000
rect 6643 28944 6668 29000
rect 6724 28944 6749 29000
rect 6805 28944 6830 29000
rect 6886 28944 6911 29000
rect 6967 28944 6992 29000
rect 7048 28944 7073 29000
rect 7129 28944 7154 29000
rect 7210 28944 7235 29000
rect 7291 28944 7316 29000
rect 7372 28944 7397 29000
rect 7453 28944 7478 29000
rect 7534 28944 7559 29000
rect 7615 28944 7640 29000
rect 7696 28944 7721 29000
rect 7777 28944 7802 29000
rect 7858 28944 7883 29000
rect 7939 28944 7964 29000
rect 8020 28944 8045 29000
rect 8101 28944 8126 29000
rect 8182 28944 8207 29000
rect 8263 28944 8288 29000
rect 8344 28944 8369 29000
rect 8425 28944 8450 29000
rect 8506 28944 8531 29000
rect 8587 28944 8612 29000
rect 8668 28944 8693 29000
rect 8749 28944 8774 29000
rect 8830 28944 8855 29000
rect 8911 28944 8936 29000
rect 8992 28944 9017 29000
rect 9073 28944 9098 29000
rect 9154 28944 9179 29000
rect 9235 28944 9260 29000
rect 2138 28927 9260 28944
rect 2138 28871 2139 28927
rect 2195 28871 2237 28927
rect 2293 28871 2335 28927
rect 2391 28871 2433 28927
rect 2489 28920 9260 28927
rect 2489 28871 6182 28920
rect 2138 28864 6182 28871
rect 6238 28864 6263 28920
rect 6319 28864 6344 28920
rect 6400 28864 6425 28920
rect 6481 28864 6506 28920
rect 6562 28864 6587 28920
rect 6643 28864 6668 28920
rect 6724 28864 6749 28920
rect 6805 28864 6830 28920
rect 6886 28864 6911 28920
rect 6967 28864 6992 28920
rect 7048 28864 7073 28920
rect 7129 28864 7154 28920
rect 7210 28864 7235 28920
rect 7291 28864 7316 28920
rect 7372 28864 7397 28920
rect 7453 28864 7478 28920
rect 7534 28864 7559 28920
rect 7615 28864 7640 28920
rect 7696 28864 7721 28920
rect 7777 28864 7802 28920
rect 7858 28864 7883 28920
rect 7939 28864 7964 28920
rect 8020 28864 8045 28920
rect 8101 28864 8126 28920
rect 8182 28864 8207 28920
rect 8263 28864 8288 28920
rect 8344 28864 8369 28920
rect 8425 28864 8450 28920
rect 8506 28864 8531 28920
rect 8587 28864 8612 28920
rect 8668 28864 8693 28920
rect 8749 28864 8774 28920
rect 8830 28864 8855 28920
rect 8911 28864 8936 28920
rect 8992 28864 9017 28920
rect 9073 28864 9098 28920
rect 9154 28864 9179 28920
rect 9235 28864 9260 28920
rect 13076 29867 14514 29880
rect 14570 29867 14594 29923
rect 14650 29867 14674 29923
rect 14730 29867 14754 29923
rect 14810 29867 14834 29923
rect 14890 29867 14914 29923
rect 14970 29867 14994 29923
rect 15050 29867 15074 29923
rect 15130 29867 15154 29923
rect 15210 29867 15234 29923
rect 15290 29867 15298 29923
rect 13076 29840 15298 29867
rect 13076 29784 14514 29840
rect 14570 29784 14594 29840
rect 14650 29784 14674 29840
rect 14730 29784 14754 29840
rect 14810 29784 14834 29840
rect 14890 29784 14914 29840
rect 14970 29784 14994 29840
rect 15050 29784 15074 29840
rect 15130 29784 15154 29840
rect 15210 29784 15234 29840
rect 15290 29784 15298 29840
rect 13076 29757 15298 29784
rect 13076 29701 14514 29757
rect 14570 29701 14594 29757
rect 14650 29701 14674 29757
rect 14730 29701 14754 29757
rect 14810 29701 14834 29757
rect 14890 29701 14914 29757
rect 14970 29701 14994 29757
rect 15050 29701 15074 29757
rect 15130 29701 15154 29757
rect 15210 29701 15234 29757
rect 15290 29701 15298 29757
rect 13076 29674 15298 29701
rect 13076 29618 14514 29674
rect 14570 29618 14594 29674
rect 14650 29618 14674 29674
rect 14730 29618 14754 29674
rect 14810 29618 14834 29674
rect 14890 29618 14914 29674
rect 14970 29618 14994 29674
rect 15050 29618 15074 29674
rect 15130 29618 15154 29674
rect 15210 29618 15234 29674
rect 15290 29618 15298 29674
rect 13076 29591 15298 29618
rect 13076 29535 14514 29591
rect 14570 29535 14594 29591
rect 14650 29535 14674 29591
rect 14730 29535 14754 29591
rect 14810 29535 14834 29591
rect 14890 29535 14914 29591
rect 14970 29535 14994 29591
rect 15050 29535 15074 29591
rect 15130 29535 15154 29591
rect 15210 29535 15234 29591
rect 15290 29535 15298 29591
rect 13076 29508 15298 29535
rect 13076 29452 14514 29508
rect 14570 29452 14594 29508
rect 14650 29452 14674 29508
rect 14730 29452 14754 29508
rect 14810 29452 14834 29508
rect 14890 29452 14914 29508
rect 14970 29452 14994 29508
rect 15050 29452 15074 29508
rect 15130 29452 15154 29508
rect 15210 29452 15234 29508
rect 15290 29452 15298 29508
rect 13076 29425 15298 29452
rect 13076 29369 14514 29425
rect 14570 29369 14594 29425
rect 14650 29369 14674 29425
rect 14730 29369 14754 29425
rect 14810 29369 14834 29425
rect 14890 29369 14914 29425
rect 14970 29369 14994 29425
rect 15050 29369 15074 29425
rect 15130 29369 15154 29425
rect 15210 29369 15234 29425
rect 15290 29369 15298 29425
rect 13076 29342 15298 29369
rect 13076 29286 14514 29342
rect 14570 29286 14594 29342
rect 14650 29286 14674 29342
rect 14730 29286 14754 29342
rect 14810 29286 14834 29342
rect 14890 29286 14914 29342
rect 14970 29286 14994 29342
rect 15050 29286 15074 29342
rect 15130 29286 15154 29342
rect 15210 29286 15234 29342
rect 15290 29286 15298 29342
rect 13076 29259 15298 29286
rect 13076 29203 14514 29259
rect 14570 29203 14594 29259
rect 14650 29203 14674 29259
rect 14730 29203 14754 29259
rect 14810 29203 14834 29259
rect 14890 29203 14914 29259
rect 14970 29203 14994 29259
rect 15050 29203 15074 29259
rect 15130 29203 15154 29259
rect 15210 29203 15234 29259
rect 15290 29203 15298 29259
rect 13076 29176 15298 29203
rect 13076 29120 14514 29176
rect 14570 29120 14594 29176
rect 14650 29120 14674 29176
rect 14730 29120 14754 29176
rect 14810 29120 14834 29176
rect 14890 29120 14914 29176
rect 14970 29120 14994 29176
rect 15050 29120 15074 29176
rect 15130 29120 15154 29176
rect 15210 29120 15234 29176
rect 15290 29120 15298 29176
rect 13076 29093 15298 29120
rect 13076 29037 14514 29093
rect 14570 29037 14594 29093
rect 14650 29037 14674 29093
rect 14730 29037 14754 29093
rect 14810 29037 14834 29093
rect 14890 29037 14914 29093
rect 14970 29037 14994 29093
rect 15050 29037 15074 29093
rect 15130 29037 15154 29093
rect 15210 29037 15234 29093
rect 15290 29037 15298 29093
rect 13076 29010 15298 29037
rect 13076 28954 14514 29010
rect 14570 28954 14594 29010
rect 14650 28954 14674 29010
rect 14730 28954 14754 29010
rect 14810 28954 14834 29010
rect 14890 28954 14914 29010
rect 14970 28954 14994 29010
rect 15050 28954 15074 29010
rect 15130 28954 15154 29010
rect 15210 28954 15234 29010
rect 15290 28954 15298 29010
rect 13076 28927 15298 28954
rect 13076 28871 14514 28927
rect 14570 28871 14594 28927
rect 14650 28871 14674 28927
rect 14730 28871 14754 28927
rect 14810 28871 14834 28927
rect 14890 28871 14914 28927
rect 14970 28871 14994 28927
rect 15050 28871 15074 28927
rect 15130 28871 15154 28927
rect 15210 28871 15234 28927
rect 15290 28871 15298 28927
rect 13076 28864 15298 28871
rect 2138 28862 15298 28864
tri 7253 28562 7553 28862 ne
rect 7553 28562 10580 28862
tri 10580 28562 10880 28862 nw
rect 2781 28561 2790 28562
rect 2846 28561 2874 28562
rect 2930 28561 2958 28562
rect 3014 28561 3042 28562
rect 3098 28561 3126 28562
rect 3182 28561 3210 28562
rect 3266 28561 3294 28562
rect 3350 28561 3378 28562
rect 3434 28561 3462 28562
rect 3518 28561 3545 28562
rect 3601 28561 3628 28562
rect 3684 28561 3711 28562
rect 2781 28509 2788 28561
rect 2846 28509 2854 28561
rect 3036 28509 3042 28561
rect 3101 28509 3114 28561
rect 3361 28509 3374 28561
rect 3434 28509 3439 28561
rect 3621 28509 3628 28561
rect 3686 28509 3699 28561
rect 2781 28506 2790 28509
rect 2846 28506 2874 28509
rect 2930 28506 2958 28509
rect 3014 28506 3042 28509
rect 3098 28506 3126 28509
rect 3182 28506 3210 28509
rect 3266 28506 3294 28509
rect 3350 28506 3378 28509
rect 3434 28506 3462 28509
rect 3518 28506 3545 28509
rect 3601 28506 3628 28509
rect 3684 28506 3711 28509
rect 3767 28506 3776 28562
rect 2781 28491 3776 28506
rect 2781 28439 2788 28491
rect 2840 28439 2854 28491
rect 2906 28439 2919 28491
rect 2971 28439 2984 28491
rect 3036 28439 3049 28491
rect 3101 28439 3114 28491
rect 3166 28439 3179 28491
rect 3231 28439 3244 28491
rect 3296 28439 3309 28491
rect 3361 28439 3374 28491
rect 3426 28439 3439 28491
rect 3491 28439 3504 28491
rect 3556 28439 3569 28491
rect 3621 28439 3634 28491
rect 3686 28439 3699 28491
rect 3751 28439 3776 28491
rect 2781 28424 3776 28439
rect 2781 28421 2790 28424
rect 2846 28421 2874 28424
rect 2930 28421 2958 28424
rect 3014 28421 3042 28424
rect 3098 28421 3126 28424
rect 3182 28421 3210 28424
rect 3266 28421 3294 28424
rect 3350 28421 3378 28424
rect 3434 28421 3462 28424
rect 3518 28421 3545 28424
rect 3601 28421 3628 28424
rect 3684 28421 3711 28424
rect 2781 28369 2788 28421
rect 2846 28369 2854 28421
rect 3036 28369 3042 28421
rect 3101 28369 3114 28421
rect 3361 28369 3374 28421
rect 3434 28369 3439 28421
rect 3621 28369 3628 28421
rect 3686 28369 3699 28421
rect 2781 28368 2790 28369
rect 2846 28368 2874 28369
rect 2930 28368 2958 28369
rect 3014 28368 3042 28369
rect 3098 28368 3126 28369
rect 3182 28368 3210 28369
rect 3266 28368 3294 28369
rect 3350 28368 3378 28369
rect 3434 28368 3462 28369
rect 3518 28368 3545 28369
rect 3601 28368 3628 28369
rect 3684 28368 3711 28369
rect 3767 28368 3776 28424
tri 7553 28368 7747 28562 ne
rect 7747 28368 10386 28562
tri 10386 28368 10580 28562 nw
tri 7747 28066 8049 28368 ne
rect 8049 28066 10050 28368
rect 148 27972 149 28024
rect 201 27972 247 28024
rect 299 28015 454 28024
rect 506 28015 528 28024
rect 580 28015 602 28024
rect 148 27959 299 27972
rect 355 27959 393 28015
rect 449 27972 454 28015
rect 580 27972 581 28015
rect 449 27959 487 27972
rect 543 27959 581 27972
rect 637 27959 654 27972
rect 148 27958 654 27959
rect 148 27906 149 27958
rect 201 27906 247 27958
rect 299 27933 454 27958
rect 506 27933 528 27958
rect 580 27933 602 27958
rect 148 27892 299 27906
rect 148 27840 149 27892
rect 201 27840 247 27892
rect 355 27877 393 27933
rect 449 27906 454 27933
rect 580 27906 581 27933
rect 449 27892 487 27906
rect 543 27892 581 27906
rect 637 27892 654 27906
rect 449 27877 454 27892
rect 580 27877 581 27892
rect 299 27851 454 27877
rect 506 27851 528 27877
rect 580 27851 602 27877
rect 148 27826 299 27840
rect 148 27774 149 27826
rect 201 27774 247 27826
rect 355 27795 393 27851
rect 449 27840 454 27851
rect 580 27840 581 27851
rect 449 27826 487 27840
rect 543 27826 581 27840
rect 637 27826 654 27840
rect 449 27795 454 27826
rect 580 27795 581 27826
rect 299 27774 454 27795
rect 506 27774 528 27795
rect 580 27774 602 27795
rect 148 27769 654 27774
rect 148 27760 299 27769
rect 148 27708 149 27760
rect 201 27708 247 27760
rect 355 27713 393 27769
rect 449 27760 487 27769
rect 543 27760 581 27769
rect 637 27760 654 27769
rect 449 27713 454 27760
rect 580 27713 581 27760
rect 299 27708 454 27713
rect 506 27708 528 27713
rect 580 27708 602 27713
rect 148 27694 654 27708
rect 148 27642 149 27694
rect 201 27642 247 27694
rect 299 27687 454 27694
rect 506 27687 528 27694
rect 580 27687 602 27694
rect 148 27631 299 27642
rect 355 27631 393 27687
rect 449 27642 454 27687
rect 580 27642 581 27687
rect 449 27631 487 27642
rect 543 27631 581 27642
rect 637 27631 654 27642
rect 148 27628 654 27631
rect 148 27576 149 27628
rect 201 27576 247 27628
rect 299 27605 454 27628
rect 506 27605 528 27628
rect 580 27605 602 27628
rect 148 27562 299 27576
rect 148 27510 149 27562
rect 201 27510 247 27562
rect 355 27549 393 27605
rect 449 27576 454 27605
rect 580 27576 581 27605
rect 449 27562 487 27576
rect 543 27562 581 27576
rect 637 27562 654 27576
rect 449 27549 454 27562
rect 580 27549 581 27562
rect 299 27523 454 27549
rect 506 27523 528 27549
rect 580 27523 602 27549
rect 148 27496 299 27510
rect 148 27444 149 27496
rect 201 27444 247 27496
rect 355 27467 393 27523
rect 449 27510 454 27523
rect 580 27510 581 27523
rect 449 27496 487 27510
rect 543 27496 581 27510
rect 637 27496 654 27510
rect 449 27467 454 27496
rect 580 27467 581 27496
rect 299 27444 454 27467
rect 506 27444 528 27467
rect 580 27444 602 27467
rect 148 27441 654 27444
rect 148 27430 299 27441
rect 148 27378 149 27430
rect 201 27378 247 27430
rect 355 27385 393 27441
rect 449 27430 487 27441
rect 543 27430 581 27441
rect 637 27430 654 27441
rect 449 27385 454 27430
rect 580 27385 581 27430
rect 299 27378 454 27385
rect 506 27378 528 27385
rect 580 27378 602 27385
rect 148 27364 654 27378
rect 148 27312 149 27364
rect 201 27312 247 27364
rect 299 27359 454 27364
rect 506 27359 528 27364
rect 580 27359 602 27364
rect 148 27303 299 27312
rect 355 27303 393 27359
rect 449 27312 454 27359
rect 580 27312 581 27359
rect 449 27303 487 27312
rect 543 27303 581 27312
rect 637 27303 654 27312
rect 148 27298 654 27303
rect 148 27246 149 27298
rect 201 27246 247 27298
rect 299 27277 454 27298
rect 506 27277 528 27298
rect 580 27277 602 27298
rect 148 27232 299 27246
rect 148 27180 149 27232
rect 201 27180 247 27232
rect 355 27221 393 27277
rect 449 27246 454 27277
rect 580 27246 581 27277
rect 449 27232 487 27246
rect 543 27232 581 27246
rect 637 27232 654 27246
rect 449 27221 454 27232
rect 580 27221 581 27232
rect 299 27195 454 27221
rect 506 27195 528 27221
rect 580 27195 602 27221
rect 148 27166 299 27180
rect 148 27114 149 27166
rect 201 27114 247 27166
rect 355 27139 393 27195
rect 449 27180 454 27195
rect 580 27180 581 27195
rect 449 27167 487 27180
rect 543 27167 581 27180
rect 637 27167 654 27180
rect 449 27139 454 27167
rect 580 27139 581 27167
rect 299 27115 454 27139
rect 506 27115 528 27139
rect 580 27115 602 27139
rect 299 27114 654 27115
rect 148 27112 654 27114
rect 148 27100 299 27112
rect 148 27048 149 27100
rect 201 27048 247 27100
rect 355 27056 393 27112
rect 449 27102 487 27112
rect 543 27102 581 27112
rect 637 27102 654 27112
rect 449 27056 454 27102
rect 580 27056 581 27102
rect 299 27050 454 27056
rect 506 27050 528 27056
rect 580 27050 602 27056
rect 299 27048 654 27050
rect 148 27037 654 27048
rect 148 27034 454 27037
rect 148 26982 149 27034
rect 201 26982 247 27034
rect 299 27029 454 27034
rect 506 27029 528 27037
rect 580 27029 602 27037
rect 148 26973 299 26982
rect 355 26973 393 27029
rect 449 26985 454 27029
rect 580 26985 581 27029
rect 449 26973 487 26985
rect 543 26973 581 26985
rect 637 26973 654 26985
rect 148 26972 654 26973
rect 148 26968 454 26972
rect 148 26916 149 26968
rect 201 26916 247 26968
rect 299 26946 454 26968
rect 506 26946 528 26972
rect 580 26946 602 26972
rect 148 26902 299 26916
rect 148 26850 149 26902
rect 201 26850 247 26902
rect 355 26890 393 26946
rect 449 26920 454 26946
rect 580 26920 581 26946
rect 449 26907 487 26920
rect 543 26907 581 26920
rect 637 26907 654 26920
rect 449 26890 454 26907
rect 580 26890 581 26907
rect 299 26863 454 26890
rect 506 26863 528 26890
rect 580 26863 602 26890
rect 148 26836 299 26850
rect 148 26784 149 26836
rect 201 26784 247 26836
rect 355 26807 393 26863
rect 449 26855 454 26863
rect 580 26855 581 26863
rect 449 26842 487 26855
rect 543 26842 581 26855
rect 637 26842 654 26855
rect 449 26807 454 26842
rect 580 26807 581 26842
rect 299 26790 454 26807
rect 506 26790 528 26807
rect 580 26790 602 26807
rect 299 26784 654 26790
rect 148 26780 654 26784
rect 148 26770 299 26780
rect 148 26718 149 26770
rect 201 26718 247 26770
rect 355 26724 393 26780
rect 449 26777 487 26780
rect 543 26777 581 26780
rect 637 26777 654 26780
rect 449 26725 454 26777
rect 580 26725 581 26777
rect 449 26724 487 26725
rect 543 26724 581 26725
rect 637 26724 654 26725
rect 299 26718 654 26724
rect 148 26712 654 26718
rect 148 26704 454 26712
rect 148 26652 149 26704
rect 201 26652 247 26704
rect 299 26697 454 26704
rect 506 26697 528 26712
rect 580 26697 602 26712
rect 148 26641 299 26652
rect 355 26641 393 26697
rect 449 26660 454 26697
rect 580 26660 581 26697
rect 449 26647 487 26660
rect 543 26647 581 26660
rect 637 26647 654 26660
rect 449 26641 454 26647
rect 580 26641 581 26647
rect 148 26638 454 26641
rect 148 26586 149 26638
rect 201 26586 247 26638
rect 299 26614 454 26638
rect 506 26614 528 26641
rect 580 26614 602 26641
rect 148 26573 299 26586
rect 148 26521 149 26573
rect 201 26521 247 26573
rect 355 26558 393 26614
rect 449 26595 454 26614
rect 580 26595 581 26614
rect 449 26582 487 26595
rect 543 26582 581 26595
rect 637 26582 654 26595
rect 449 26558 454 26582
rect 580 26558 581 26582
rect 299 26531 454 26558
rect 506 26531 528 26558
rect 580 26531 602 26558
rect 148 26508 299 26521
rect 148 26456 149 26508
rect 201 26456 247 26508
rect 355 26475 393 26531
rect 449 26530 454 26531
rect 580 26530 581 26531
rect 449 26517 487 26530
rect 543 26517 581 26530
rect 637 26517 654 26530
rect 449 26475 454 26517
rect 580 26475 581 26517
rect 299 26465 454 26475
rect 506 26465 528 26475
rect 580 26465 602 26475
rect 299 26456 654 26465
rect 148 26452 654 26456
rect 148 26448 454 26452
rect 506 26448 528 26452
rect 580 26448 602 26452
rect 148 26443 299 26448
rect 148 26391 149 26443
rect 201 26391 247 26443
rect 355 26392 393 26448
rect 449 26400 454 26448
rect 580 26400 581 26448
rect 449 26392 487 26400
rect 543 26392 581 26400
rect 637 26392 654 26400
rect 299 26391 654 26392
rect 148 26387 654 26391
rect 148 26378 454 26387
rect 148 26326 149 26378
rect 201 26326 247 26378
rect 299 26365 454 26378
rect 506 26365 528 26387
rect 580 26365 602 26387
rect 2163 28057 5086 28066
rect 2163 28001 2165 28057
rect 2221 28001 2255 28057
rect 2311 28001 2345 28057
rect 2401 28001 2435 28057
rect 2491 28001 4105 28057
rect 4161 28001 4189 28057
rect 4245 28001 4273 28057
rect 4329 28001 4357 28057
rect 4413 28001 4441 28057
rect 4497 28001 4525 28057
rect 4581 28001 4609 28057
rect 4665 28001 4693 28057
rect 4749 28001 4777 28057
rect 4833 28001 4861 28057
rect 4917 28001 4945 28057
rect 5001 28001 5029 28057
rect 5085 28001 5086 28057
tri 8049 28032 8083 28066 ne
rect 2163 27977 5086 28001
rect 2163 27921 2165 27977
rect 2221 27921 2255 27977
rect 2311 27921 2345 27977
rect 2401 27921 2435 27977
rect 2491 27921 4105 27977
rect 4161 27921 4189 27977
rect 4245 27921 4273 27977
rect 4329 27921 4357 27977
rect 4413 27921 4441 27977
rect 4497 27921 4525 27977
rect 4581 27921 4609 27977
rect 4665 27921 4693 27977
rect 4749 27921 4777 27977
rect 4833 27921 4861 27977
rect 4917 27921 4945 27977
rect 5001 27921 5029 27977
rect 5085 27921 5086 27977
rect 2163 27897 5086 27921
rect 2163 27841 2165 27897
rect 2221 27841 2255 27897
rect 2311 27841 2345 27897
rect 2401 27841 2435 27897
rect 2491 27841 4105 27897
rect 4161 27841 4189 27897
rect 4245 27841 4273 27897
rect 4329 27841 4357 27897
rect 4413 27841 4441 27897
rect 4497 27841 4525 27897
rect 4581 27841 4609 27897
rect 4665 27841 4693 27897
rect 4749 27841 4777 27897
rect 4833 27841 4861 27897
rect 4917 27841 4945 27897
rect 5001 27841 5029 27897
rect 5085 27841 5086 27897
rect 2163 27817 5086 27841
rect 2163 27761 2165 27817
rect 2221 27761 2255 27817
rect 2311 27761 2345 27817
rect 2401 27761 2435 27817
rect 2491 27761 4105 27817
rect 4161 27761 4189 27817
rect 4245 27761 4273 27817
rect 4329 27761 4357 27817
rect 4413 27761 4441 27817
rect 4497 27761 4525 27817
rect 4581 27761 4609 27817
rect 4665 27761 4693 27817
rect 4749 27761 4777 27817
rect 4833 27761 4861 27817
rect 4917 27761 4945 27817
rect 5001 27761 5029 27817
rect 5085 27761 5086 27817
rect 2163 27737 5086 27761
rect 2163 27681 2165 27737
rect 2221 27681 2255 27737
rect 2311 27681 2345 27737
rect 2401 27681 2435 27737
rect 2491 27681 4105 27737
rect 4161 27681 4189 27737
rect 4245 27681 4273 27737
rect 4329 27681 4357 27737
rect 4413 27681 4441 27737
rect 4497 27681 4525 27737
rect 4581 27681 4609 27737
rect 4665 27681 4693 27737
rect 4749 27681 4777 27737
rect 4833 27681 4861 27737
rect 4917 27681 4945 27737
rect 5001 27681 5029 27737
rect 5085 27681 5086 27737
rect 2163 27657 5086 27681
rect 2163 27601 2165 27657
rect 2221 27601 2255 27657
rect 2311 27601 2345 27657
rect 2401 27601 2435 27657
rect 2491 27601 4105 27657
rect 4161 27601 4189 27657
rect 4245 27601 4273 27657
rect 4329 27601 4357 27657
rect 4413 27601 4441 27657
rect 4497 27601 4525 27657
rect 4581 27601 4609 27657
rect 4665 27601 4693 27657
rect 4749 27601 4777 27657
rect 4833 27601 4861 27657
rect 4917 27601 4945 27657
rect 5001 27601 5029 27657
rect 5085 27601 5086 27657
rect 2163 27577 5086 27601
rect 2163 27521 2165 27577
rect 2221 27521 2255 27577
rect 2311 27521 2345 27577
rect 2401 27521 2435 27577
rect 2491 27521 4105 27577
rect 4161 27521 4189 27577
rect 4245 27521 4273 27577
rect 4329 27521 4357 27577
rect 4413 27521 4441 27577
rect 4497 27521 4525 27577
rect 4581 27521 4609 27577
rect 4665 27521 4693 27577
rect 4749 27521 4777 27577
rect 4833 27521 4861 27577
rect 4917 27521 4945 27577
rect 5001 27521 5029 27577
rect 5085 27521 5086 27577
rect 2163 27497 5086 27521
rect 2163 27441 2165 27497
rect 2221 27441 2255 27497
rect 2311 27441 2345 27497
rect 2401 27441 2435 27497
rect 2491 27441 4105 27497
rect 4161 27441 4189 27497
rect 4245 27441 4273 27497
rect 4329 27441 4357 27497
rect 4413 27441 4441 27497
rect 4497 27441 4525 27497
rect 4581 27441 4609 27497
rect 4665 27441 4693 27497
rect 4749 27441 4777 27497
rect 4833 27441 4861 27497
rect 4917 27441 4945 27497
rect 5001 27441 5029 27497
rect 5085 27441 5086 27497
rect 2163 27417 5086 27441
rect 2163 27361 2165 27417
rect 2221 27361 2255 27417
rect 2311 27361 2345 27417
rect 2401 27361 2435 27417
rect 2491 27361 4105 27417
rect 4161 27361 4189 27417
rect 4245 27361 4273 27417
rect 4329 27361 4357 27417
rect 4413 27361 4441 27417
rect 4497 27361 4525 27417
rect 4581 27361 4609 27417
rect 4665 27361 4693 27417
rect 4749 27361 4777 27417
rect 4833 27361 4861 27417
rect 4917 27361 4945 27417
rect 5001 27361 5029 27417
rect 5085 27361 5086 27417
rect 2163 27337 5086 27361
rect 2163 27281 2165 27337
rect 2221 27281 2255 27337
rect 2311 27281 2345 27337
rect 2401 27281 2435 27337
rect 2491 27281 4105 27337
rect 4161 27281 4189 27337
rect 4245 27281 4273 27337
rect 4329 27281 4357 27337
rect 4413 27281 4441 27337
rect 4497 27281 4525 27337
rect 4581 27281 4609 27337
rect 4665 27281 4693 27337
rect 4749 27281 4777 27337
rect 4833 27281 4861 27337
rect 4917 27281 4945 27337
rect 5001 27281 5029 27337
rect 5085 27281 5086 27337
rect 2163 27257 5086 27281
rect 2163 27201 2165 27257
rect 2221 27201 2255 27257
rect 2311 27201 2345 27257
rect 2401 27201 2435 27257
rect 2491 27201 4105 27257
rect 4161 27201 4189 27257
rect 4245 27201 4273 27257
rect 4329 27201 4357 27257
rect 4413 27201 4441 27257
rect 4497 27201 4525 27257
rect 4581 27201 4609 27257
rect 4665 27201 4693 27257
rect 4749 27201 4777 27257
rect 4833 27201 4861 27257
rect 4917 27201 4945 27257
rect 5001 27201 5029 27257
rect 5085 27201 5086 27257
rect 2163 27177 5086 27201
rect 2163 27121 2165 27177
rect 2221 27121 2255 27177
rect 2311 27121 2345 27177
rect 2401 27121 2435 27177
rect 2491 27121 4105 27177
rect 4161 27121 4189 27177
rect 4245 27121 4273 27177
rect 4329 27121 4357 27177
rect 4413 27121 4441 27177
rect 4497 27121 4525 27177
rect 4581 27121 4609 27177
rect 4665 27121 4693 27177
rect 4749 27121 4777 27177
rect 4833 27121 4861 27177
rect 4917 27121 4945 27177
rect 5001 27121 5029 27177
rect 5085 27121 5086 27177
rect 2163 27097 5086 27121
rect 2163 27041 2165 27097
rect 2221 27041 2255 27097
rect 2311 27041 2345 27097
rect 2401 27041 2435 27097
rect 2491 27041 4105 27097
rect 4161 27041 4189 27097
rect 4245 27041 4273 27097
rect 4329 27041 4357 27097
rect 4413 27041 4441 27097
rect 4497 27041 4525 27097
rect 4581 27041 4609 27097
rect 4665 27041 4693 27097
rect 4749 27041 4777 27097
rect 4833 27041 4861 27097
rect 4917 27041 4945 27097
rect 5001 27041 5029 27097
rect 5085 27041 5086 27097
rect 2163 27017 5086 27041
rect 2163 26961 2165 27017
rect 2221 26961 2255 27017
rect 2311 26961 2345 27017
rect 2401 26961 2435 27017
rect 2491 26961 4105 27017
rect 4161 26961 4189 27017
rect 4245 26961 4273 27017
rect 4329 26961 4357 27017
rect 4413 26961 4441 27017
rect 4497 26961 4525 27017
rect 4581 26961 4609 27017
rect 4665 26961 4693 27017
rect 4749 26961 4777 27017
rect 4833 26961 4861 27017
rect 4917 26961 4945 27017
rect 5001 26961 5029 27017
rect 5085 26961 5086 27017
rect 2163 26936 5086 26961
rect 2163 26880 2165 26936
rect 2221 26880 2255 26936
rect 2311 26880 2345 26936
rect 2401 26880 2435 26936
rect 2491 26880 4105 26936
rect 4161 26880 4189 26936
rect 4245 26880 4273 26936
rect 4329 26880 4357 26936
rect 4413 26880 4441 26936
rect 4497 26880 4525 26936
rect 4581 26880 4609 26936
rect 4665 26880 4693 26936
rect 4749 26880 4777 26936
rect 4833 26880 4861 26936
rect 4917 26880 4945 26936
rect 5001 26880 5029 26936
rect 5085 26880 5086 26936
rect 2163 26855 5086 26880
rect 2163 26799 2165 26855
rect 2221 26799 2255 26855
rect 2311 26799 2345 26855
rect 2401 26799 2435 26855
rect 2491 26799 4105 26855
rect 4161 26799 4189 26855
rect 4245 26799 4273 26855
rect 4329 26799 4357 26855
rect 4413 26799 4441 26855
rect 4497 26799 4525 26855
rect 4581 26799 4609 26855
rect 4665 26799 4693 26855
rect 4749 26799 4777 26855
rect 4833 26799 4861 26855
rect 4917 26799 4945 26855
rect 5001 26799 5029 26855
rect 5085 26799 5086 26855
rect 2163 26774 5086 26799
rect 2163 26718 2165 26774
rect 2221 26718 2255 26774
rect 2311 26718 2345 26774
rect 2401 26718 2435 26774
rect 2491 26718 4105 26774
rect 4161 26718 4189 26774
rect 4245 26718 4273 26774
rect 4329 26718 4357 26774
rect 4413 26718 4441 26774
rect 4497 26718 4525 26774
rect 4581 26718 4609 26774
rect 4665 26718 4693 26774
rect 4749 26718 4777 26774
rect 4833 26718 4861 26774
rect 4917 26718 4945 26774
rect 5001 26718 5029 26774
rect 5085 26718 5086 26774
rect 2163 26693 5086 26718
rect 2163 26637 2165 26693
rect 2221 26637 2255 26693
rect 2311 26637 2345 26693
rect 2401 26637 2435 26693
rect 2491 26637 4105 26693
rect 4161 26637 4189 26693
rect 4245 26637 4273 26693
rect 4329 26637 4357 26693
rect 4413 26637 4441 26693
rect 4497 26637 4525 26693
rect 4581 26637 4609 26693
rect 4665 26637 4693 26693
rect 4749 26637 4777 26693
rect 4833 26637 4861 26693
rect 4917 26637 4945 26693
rect 5001 26637 5029 26693
rect 5085 26637 5086 26693
rect 2163 26612 5086 26637
rect 2163 26556 2165 26612
rect 2221 26556 2255 26612
rect 2311 26556 2345 26612
rect 2401 26556 2435 26612
rect 2491 26556 4105 26612
rect 4161 26556 4189 26612
rect 4245 26556 4273 26612
rect 4329 26556 4357 26612
rect 4413 26556 4441 26612
rect 4497 26556 4525 26612
rect 4581 26556 4609 26612
rect 4665 26556 4693 26612
rect 4749 26556 4777 26612
rect 4833 26556 4861 26612
rect 4917 26556 4945 26612
rect 5001 26556 5029 26612
rect 5085 26556 5086 26612
rect 2163 26531 5086 26556
rect 2163 26475 2165 26531
rect 2221 26475 2255 26531
rect 2311 26475 2345 26531
rect 2401 26475 2435 26531
rect 2491 26475 4105 26531
rect 4161 26475 4189 26531
rect 4245 26475 4273 26531
rect 4329 26475 4357 26531
rect 4413 26475 4441 26531
rect 4497 26475 4525 26531
rect 4581 26475 4609 26531
rect 4665 26475 4693 26531
rect 4749 26475 4777 26531
rect 4833 26475 4861 26531
rect 4917 26475 4945 26531
rect 5001 26475 5029 26531
rect 5085 26475 5086 26531
rect 2163 26450 5086 26475
rect 2163 26394 2165 26450
rect 2221 26394 2255 26450
rect 2311 26394 2345 26450
rect 2401 26394 2435 26450
rect 2491 26394 4105 26450
rect 4161 26394 4189 26450
rect 4245 26394 4273 26450
rect 4329 26394 4357 26450
rect 4413 26394 4441 26450
rect 4497 26394 4525 26450
rect 4581 26394 4609 26450
rect 4665 26394 4693 26450
rect 4749 26394 4777 26450
rect 4833 26394 4861 26450
rect 4917 26394 4945 26450
rect 5001 26394 5029 26450
rect 5085 26394 5086 26450
rect 2163 26385 5086 26394
tri 7695 26385 8083 26773 se
rect 8083 26385 10050 28066
tri 10050 28032 10386 28368 nw
rect 14213 27574 15034 27579
rect 14213 27518 14522 27574
rect 14578 27518 14612 27574
rect 14668 27518 14702 27574
rect 14758 27518 14791 27574
rect 14847 27518 14880 27574
rect 14936 27518 14969 27574
rect 15025 27518 15034 27574
rect 14213 27488 15034 27518
rect 14213 27483 14522 27488
rect 14265 27431 14285 27483
rect 14337 27431 14357 27483
rect 14409 27432 14522 27483
rect 14578 27432 14612 27488
rect 14668 27432 14702 27488
rect 14758 27432 14791 27488
rect 14847 27432 14880 27488
rect 14936 27432 14969 27488
rect 15025 27432 15034 27488
rect 14409 27431 15034 27432
rect 14213 27416 15034 27431
rect 14265 27364 14285 27416
rect 14337 27364 14357 27416
rect 14409 27402 15034 27416
rect 14409 27364 14522 27402
rect 14213 27349 14522 27364
rect 14265 27297 14285 27349
rect 14337 27297 14357 27349
rect 14409 27346 14522 27349
rect 14578 27346 14612 27402
rect 14668 27346 14702 27402
rect 14758 27346 14791 27402
rect 14847 27346 14880 27402
rect 14936 27346 14969 27402
rect 15025 27346 15034 27402
rect 14409 27316 15034 27346
rect 14409 27297 14522 27316
rect 14213 27281 14522 27297
rect 14265 27229 14285 27281
rect 14337 27229 14357 27281
rect 14409 27260 14522 27281
rect 14578 27260 14612 27316
rect 14668 27260 14702 27316
rect 14758 27260 14791 27316
rect 14847 27260 14880 27316
rect 14936 27260 14969 27316
rect 15025 27260 15034 27316
rect 14409 27230 15034 27260
rect 14409 27229 14522 27230
rect 14213 27213 14522 27229
rect 14265 27161 14285 27213
rect 14337 27161 14357 27213
rect 14409 27174 14522 27213
rect 14578 27174 14612 27230
rect 14668 27174 14702 27230
rect 14758 27174 14791 27230
rect 14847 27174 14880 27230
rect 14936 27174 14969 27230
rect 15025 27174 15034 27230
rect 14409 27161 15034 27174
rect 14213 27145 15034 27161
rect 14265 27093 14285 27145
rect 14337 27093 14357 27145
rect 14409 27144 15034 27145
rect 14409 27093 14522 27144
rect 14213 27088 14522 27093
rect 14578 27088 14612 27144
rect 14668 27088 14702 27144
rect 14758 27088 14791 27144
rect 14847 27088 14880 27144
rect 14936 27088 14969 27144
rect 15025 27088 15034 27144
rect 14213 27087 15034 27088
rect 148 26313 299 26326
rect 148 26261 149 26313
rect 201 26261 247 26313
rect 355 26309 393 26365
rect 449 26335 454 26365
rect 580 26335 581 26365
rect 449 26322 487 26335
rect 543 26322 581 26335
rect 637 26322 654 26335
rect 449 26309 454 26322
rect 580 26309 581 26322
rect 299 26282 454 26309
rect 506 26282 528 26309
rect 580 26282 602 26309
rect 148 26226 299 26261
rect 355 26226 393 26282
rect 449 26270 454 26282
rect 580 26270 581 26282
rect 449 26257 487 26270
rect 543 26257 581 26270
rect 637 26257 654 26270
rect 449 26226 454 26257
rect 580 26226 581 26257
rect 148 26205 454 26226
rect 506 26205 528 26226
rect 580 26205 602 26226
rect 148 26199 654 26205
tri 7509 26199 7695 26385 se
rect 7695 26199 10050 26385
tri 7354 26044 7509 26199 se
rect 7509 26044 10050 26199
rect 148 26038 850 26044
rect 148 25986 149 26038
rect 201 25986 247 26038
rect 299 25986 456 26038
rect 508 25986 524 26038
rect 576 25986 592 26038
rect 644 25986 660 26038
rect 712 25986 728 26038
rect 780 25986 796 26038
rect 848 25986 850 26038
rect 148 25974 850 25986
rect 148 25922 149 25974
rect 201 25922 247 25974
rect 299 25922 456 25974
rect 508 25922 524 25974
rect 576 25922 592 25974
rect 644 25922 660 25974
rect 712 25922 728 25974
rect 780 25922 796 25974
rect 848 25922 850 25974
rect 148 25910 850 25922
rect 148 25858 149 25910
rect 201 25858 247 25910
rect 299 25858 456 25910
rect 508 25858 524 25910
rect 576 25858 592 25910
rect 644 25858 660 25910
rect 712 25858 728 25910
rect 780 25858 796 25910
rect 848 25858 850 25910
rect 148 25846 850 25858
rect 148 25794 149 25846
rect 201 25794 247 25846
rect 299 25794 456 25846
rect 508 25794 524 25846
rect 576 25794 592 25846
rect 644 25794 660 25846
rect 712 25794 728 25846
rect 780 25794 796 25846
rect 848 25794 850 25846
tri 7149 25839 7354 26044 se
rect 7354 25839 10050 26044
tri 10050 25839 10984 26773 sw
rect 148 25782 850 25794
rect 148 25730 149 25782
rect 201 25730 247 25782
rect 299 25730 456 25782
rect 508 25730 524 25782
rect 576 25730 592 25782
rect 644 25730 660 25782
rect 712 25730 728 25782
rect 780 25730 796 25782
rect 848 25730 850 25782
rect 148 25718 850 25730
rect 148 25666 149 25718
rect 201 25666 247 25718
rect 299 25666 456 25718
rect 508 25666 524 25718
rect 576 25666 592 25718
rect 644 25666 660 25718
rect 712 25666 728 25718
rect 780 25666 796 25718
rect 848 25666 850 25718
rect 148 25654 850 25666
rect 148 25602 149 25654
rect 201 25602 247 25654
rect 299 25602 456 25654
rect 508 25602 524 25654
rect 576 25602 592 25654
rect 644 25602 660 25654
rect 712 25602 728 25654
rect 780 25602 796 25654
rect 848 25602 850 25654
rect 148 25590 850 25602
rect 148 25538 149 25590
rect 201 25538 247 25590
rect 299 25538 456 25590
rect 508 25538 524 25590
rect 576 25538 592 25590
rect 644 25538 660 25590
rect 712 25538 728 25590
rect 780 25538 796 25590
rect 848 25538 850 25590
rect 148 25526 850 25538
rect 148 25474 149 25526
rect 201 25474 247 25526
rect 299 25474 456 25526
rect 508 25474 524 25526
rect 576 25474 592 25526
rect 644 25474 660 25526
rect 712 25474 728 25526
rect 780 25474 796 25526
rect 848 25474 850 25526
rect 148 25462 850 25474
rect 148 25410 149 25462
rect 201 25410 247 25462
rect 299 25410 456 25462
rect 508 25410 524 25462
rect 576 25410 592 25462
rect 644 25410 660 25462
rect 712 25410 728 25462
rect 780 25410 796 25462
rect 848 25410 850 25462
rect 148 25398 850 25410
rect 148 25346 149 25398
rect 201 25346 247 25398
rect 299 25346 456 25398
rect 508 25346 524 25398
rect 576 25346 592 25398
rect 644 25346 660 25398
rect 712 25346 728 25398
rect 780 25346 796 25398
rect 848 25346 850 25398
rect 148 25334 850 25346
rect 148 25282 149 25334
rect 201 25282 247 25334
rect 299 25282 456 25334
rect 508 25282 524 25334
rect 576 25282 592 25334
rect 644 25282 660 25334
rect 712 25282 728 25334
rect 780 25282 796 25334
rect 848 25282 850 25334
rect 148 25270 850 25282
rect 148 25218 149 25270
rect 201 25218 247 25270
rect 299 25218 456 25270
rect 508 25218 524 25270
rect 576 25218 592 25270
rect 644 25218 660 25270
rect 712 25218 728 25270
rect 780 25218 796 25270
rect 848 25218 850 25270
rect 148 25206 850 25218
rect 148 25154 149 25206
rect 201 25154 247 25206
rect 299 25154 456 25206
rect 508 25154 524 25206
rect 576 25154 592 25206
rect 644 25154 660 25206
rect 712 25154 728 25206
rect 780 25154 796 25206
rect 848 25154 850 25206
rect 148 25142 850 25154
rect 148 25090 149 25142
rect 201 25090 247 25142
rect 299 25090 456 25142
rect 508 25090 524 25142
rect 576 25090 592 25142
rect 644 25090 660 25142
rect 712 25090 728 25142
rect 780 25090 796 25142
rect 848 25090 850 25142
rect 148 25078 850 25090
rect 148 25026 149 25078
rect 201 25026 247 25078
rect 299 25026 456 25078
rect 508 25026 524 25078
rect 576 25026 592 25078
rect 644 25026 660 25078
rect 712 25026 728 25078
rect 780 25026 796 25078
rect 848 25026 850 25078
rect 148 25014 850 25026
rect 148 24962 149 25014
rect 201 24962 247 25014
rect 299 24962 456 25014
rect 508 24962 524 25014
rect 576 24962 592 25014
rect 644 24962 660 25014
rect 712 24962 728 25014
rect 780 24962 796 25014
rect 848 24962 850 25014
rect 148 24950 850 24962
rect 148 24898 149 24950
rect 201 24898 247 24950
rect 299 24898 456 24950
rect 508 24898 524 24950
rect 576 24898 592 24950
rect 644 24898 660 24950
rect 712 24898 728 24950
rect 780 24898 796 24950
rect 848 24898 850 24950
rect 148 24886 850 24898
rect 148 24834 149 24886
rect 201 24834 247 24886
rect 299 24834 456 24886
rect 508 24834 524 24886
rect 576 24834 592 24886
rect 644 24834 660 24886
rect 712 24834 728 24886
rect 780 24834 796 24886
rect 848 24834 850 24886
rect 148 24822 850 24834
rect 148 24770 149 24822
rect 201 24770 247 24822
rect 299 24770 456 24822
rect 508 24770 524 24822
rect 576 24770 592 24822
rect 644 24770 660 24822
rect 712 24770 728 24822
rect 780 24770 796 24822
rect 848 24770 850 24822
rect 148 24758 850 24770
rect 148 24706 149 24758
rect 201 24706 247 24758
rect 299 24706 456 24758
rect 508 24706 524 24758
rect 576 24706 592 24758
rect 644 24706 660 24758
rect 712 24706 728 24758
rect 780 24706 796 24758
rect 848 24706 850 24758
rect 148 24694 850 24706
rect 148 24642 149 24694
rect 201 24642 247 24694
rect 299 24642 456 24694
rect 508 24642 524 24694
rect 576 24642 592 24694
rect 644 24642 660 24694
rect 712 24642 728 24694
rect 780 24642 796 24694
rect 848 24642 850 24694
rect 148 24630 850 24642
rect 148 24578 149 24630
rect 201 24578 247 24630
rect 299 24578 456 24630
rect 508 24578 524 24630
rect 576 24578 592 24630
rect 644 24578 660 24630
rect 712 24578 728 24630
rect 780 24578 796 24630
rect 848 24578 850 24630
rect 148 24566 850 24578
rect 148 24514 149 24566
rect 201 24514 247 24566
rect 299 24514 456 24566
rect 508 24514 524 24566
rect 576 24514 592 24566
rect 644 24514 660 24566
rect 712 24514 728 24566
rect 780 24514 796 24566
rect 848 24514 850 24566
rect 148 24502 850 24514
rect 148 24450 149 24502
rect 201 24450 247 24502
rect 299 24450 456 24502
rect 508 24450 524 24502
rect 576 24450 592 24502
rect 644 24450 660 24502
rect 712 24450 728 24502
rect 780 24450 796 24502
rect 848 24450 850 24502
rect 148 24438 850 24450
rect 148 24386 149 24438
rect 201 24386 247 24438
rect 299 24386 456 24438
rect 508 24386 524 24438
rect 576 24386 592 24438
rect 644 24386 660 24438
rect 712 24386 728 24438
rect 780 24386 796 24438
rect 848 24386 850 24438
rect 148 24374 850 24386
rect 148 24322 149 24374
rect 201 24322 247 24374
rect 299 24322 456 24374
rect 508 24322 524 24374
rect 576 24322 592 24374
rect 644 24322 660 24374
rect 712 24322 728 24374
rect 780 24322 796 24374
rect 848 24322 850 24374
rect 148 24310 850 24322
rect 148 24258 149 24310
rect 201 24258 247 24310
rect 299 24258 456 24310
rect 508 24258 524 24310
rect 576 24258 592 24310
rect 644 24258 660 24310
rect 712 24258 728 24310
rect 780 24258 796 24310
rect 848 24258 850 24310
rect 148 24246 850 24258
rect 148 24194 149 24246
rect 201 24194 247 24246
rect 299 24194 456 24246
rect 508 24194 524 24246
rect 576 24194 592 24246
rect 644 24194 660 24246
rect 712 24194 728 24246
rect 780 24194 796 24246
rect 848 24194 850 24246
rect 148 24182 850 24194
rect 148 24130 149 24182
rect 201 24130 247 24182
rect 299 24130 456 24182
rect 508 24130 524 24182
rect 576 24130 592 24182
rect 644 24130 660 24182
rect 712 24130 728 24182
rect 780 24130 796 24182
rect 848 24130 850 24182
rect 148 24118 850 24130
rect 148 24066 149 24118
rect 201 24066 247 24118
rect 299 24066 456 24118
rect 508 24066 524 24118
rect 576 24066 592 24118
rect 644 24066 660 24118
rect 712 24066 728 24118
rect 780 24066 796 24118
rect 848 24066 850 24118
rect 148 24054 850 24066
rect 148 24002 149 24054
rect 201 24002 247 24054
rect 299 24002 456 24054
rect 508 24002 524 24054
rect 576 24002 592 24054
rect 644 24002 660 24054
rect 712 24002 728 24054
rect 780 24002 796 24054
rect 848 24002 850 24054
rect 148 23990 850 24002
rect 148 23938 149 23990
rect 201 23938 247 23990
rect 299 23938 456 23990
rect 508 23938 524 23990
rect 576 23938 592 23990
rect 644 23938 660 23990
rect 712 23938 728 23990
rect 780 23938 796 23990
rect 848 23938 850 23990
rect 148 23926 850 23938
rect 148 23874 149 23926
rect 201 23874 247 23926
rect 299 23874 456 23926
rect 508 23874 524 23926
rect 576 23874 592 23926
rect 644 23874 660 23926
rect 712 23874 728 23926
rect 780 23874 796 23926
rect 848 23874 850 23926
rect 148 23862 850 23874
rect 148 23810 149 23862
rect 201 23810 247 23862
rect 299 23810 456 23862
rect 508 23810 524 23862
rect 576 23810 592 23862
rect 644 23810 660 23862
rect 712 23810 728 23862
rect 780 23810 796 23862
rect 848 23810 850 23862
rect 148 23798 850 23810
rect 148 23746 149 23798
rect 201 23746 247 23798
rect 299 23746 456 23798
rect 508 23746 524 23798
rect 576 23746 592 23798
rect 644 23746 660 23798
rect 712 23746 728 23798
rect 780 23746 796 23798
rect 848 23746 850 23798
rect 148 23734 850 23746
rect 148 23682 149 23734
rect 201 23682 247 23734
rect 299 23682 456 23734
rect 508 23682 524 23734
rect 576 23682 592 23734
rect 644 23682 660 23734
rect 712 23682 728 23734
rect 780 23682 796 23734
rect 848 23682 850 23734
rect 148 23670 850 23682
rect 148 23618 149 23670
rect 201 23618 247 23670
rect 299 23618 456 23670
rect 508 23618 524 23670
rect 576 23618 592 23670
rect 644 23618 660 23670
rect 712 23618 728 23670
rect 780 23618 796 23670
rect 848 23618 850 23670
rect 148 23606 850 23618
rect 148 23554 149 23606
rect 201 23554 247 23606
rect 299 23554 456 23606
rect 508 23554 524 23606
rect 576 23554 592 23606
rect 644 23554 660 23606
rect 712 23554 728 23606
rect 780 23554 796 23606
rect 848 23554 850 23606
rect 148 23542 850 23554
rect 148 23490 149 23542
rect 201 23490 247 23542
rect 299 23490 456 23542
rect 508 23490 524 23542
rect 576 23490 592 23542
rect 644 23490 660 23542
rect 712 23490 728 23542
rect 780 23490 796 23542
rect 848 23490 850 23542
rect 148 23478 850 23490
rect 148 23426 149 23478
rect 201 23426 247 23478
rect 299 23426 456 23478
rect 508 23426 524 23478
rect 576 23426 592 23478
rect 644 23426 660 23478
rect 712 23426 728 23478
rect 780 23426 796 23478
rect 848 23426 850 23478
rect 148 23414 850 23426
rect 148 23362 149 23414
rect 201 23362 247 23414
rect 299 23362 456 23414
rect 508 23362 524 23414
rect 576 23362 592 23414
rect 644 23362 660 23414
rect 712 23362 728 23414
rect 780 23362 796 23414
rect 848 23362 850 23414
rect 148 23350 850 23362
rect 148 23298 149 23350
rect 201 23298 247 23350
rect 299 23298 456 23350
rect 508 23298 524 23350
rect 576 23298 592 23350
rect 644 23298 660 23350
rect 712 23298 728 23350
rect 780 23298 796 23350
rect 848 23298 850 23350
rect 148 23286 850 23298
rect 148 23234 149 23286
rect 201 23234 247 23286
rect 299 23234 456 23286
rect 508 23234 524 23286
rect 576 23234 592 23286
rect 644 23234 660 23286
rect 712 23234 728 23286
rect 780 23234 796 23286
rect 848 23234 850 23286
rect 148 23222 850 23234
rect 148 23170 149 23222
rect 201 23170 247 23222
rect 299 23170 456 23222
rect 508 23170 524 23222
rect 576 23170 592 23222
rect 644 23170 660 23222
rect 712 23170 728 23222
rect 780 23170 796 23222
rect 848 23170 850 23222
rect 148 23158 850 23170
rect 148 23106 149 23158
rect 201 23106 247 23158
rect 299 23106 456 23158
rect 508 23106 524 23158
rect 576 23106 592 23158
rect 644 23106 660 23158
rect 712 23106 728 23158
rect 780 23106 796 23158
rect 848 23106 850 23158
rect 1852 25828 15047 25839
rect 1852 25820 5425 25828
rect 1852 25764 2170 25820
rect 2226 25764 2252 25820
rect 2308 25764 2334 25820
rect 2390 25764 2416 25820
rect 2472 25772 5425 25820
rect 5481 25772 5506 25828
rect 5562 25772 5587 25828
rect 5643 25772 5668 25828
rect 5724 25772 5749 25828
rect 5805 25772 5830 25828
rect 5886 25772 5911 25828
rect 5967 25772 5992 25828
rect 6048 25772 6073 25828
rect 6129 25772 6154 25828
rect 6210 25772 6235 25828
rect 6291 25772 6316 25828
rect 6372 25772 6397 25828
rect 6453 25772 6478 25828
rect 6534 25772 6559 25828
rect 6615 25772 6640 25828
rect 6696 25772 6721 25828
rect 6777 25772 6802 25828
rect 6858 25772 6883 25828
rect 6939 25772 6964 25828
rect 7020 25772 7045 25828
rect 7101 25772 7126 25828
rect 7182 25772 7207 25828
rect 7263 25772 7288 25828
rect 7344 25772 7369 25828
rect 7425 25772 7450 25828
rect 7506 25772 7531 25828
rect 7587 25772 7612 25828
rect 7668 25772 7693 25828
rect 7749 25772 7774 25828
rect 7830 25772 7855 25828
rect 7911 25772 7936 25828
rect 7992 25772 8017 25828
rect 8073 25772 8098 25828
rect 8154 25772 8179 25828
rect 8235 25772 8260 25828
rect 8316 25772 8341 25828
rect 8397 25772 8422 25828
rect 8478 25772 8503 25828
rect 8559 25772 8584 25828
rect 8640 25772 8665 25828
rect 8721 25772 8746 25828
rect 8802 25772 8827 25828
rect 8883 25772 8908 25828
rect 8964 25772 8989 25828
rect 9045 25772 9070 25828
rect 9126 25772 9151 25828
rect 9207 25772 9232 25828
rect 9288 25772 9313 25828
rect 9369 25772 9394 25828
rect 9450 25772 9475 25828
rect 9531 25772 9556 25828
rect 9612 25772 9637 25828
rect 9693 25772 9718 25828
rect 9774 25772 9799 25828
rect 9855 25772 9880 25828
rect 9936 25772 9961 25828
rect 10017 25772 10042 25828
rect 10098 25772 10123 25828
rect 10179 25772 10204 25828
rect 10260 25772 10285 25828
rect 10341 25772 10366 25828
rect 10422 25772 10447 25828
rect 10503 25772 10528 25828
rect 10584 25772 10609 25828
rect 10665 25772 10690 25828
rect 10746 25772 10771 25828
rect 10827 25772 10852 25828
rect 10908 25772 10933 25828
rect 10989 25772 11014 25828
rect 11070 25772 11095 25828
rect 11151 25772 11176 25828
rect 11232 25772 11257 25828
rect 11313 25772 11338 25828
rect 11394 25772 11419 25828
rect 11475 25772 11500 25828
rect 2472 25764 11500 25772
rect 1852 25748 11500 25764
rect 1852 25739 5425 25748
rect 1852 25683 2170 25739
rect 2226 25683 2252 25739
rect 2308 25683 2334 25739
rect 2390 25683 2416 25739
rect 2472 25692 5425 25739
rect 5481 25692 5506 25748
rect 5562 25692 5587 25748
rect 5643 25692 5668 25748
rect 5724 25692 5749 25748
rect 5805 25692 5830 25748
rect 5886 25692 5911 25748
rect 5967 25692 5992 25748
rect 6048 25692 6073 25748
rect 6129 25692 6154 25748
rect 6210 25692 6235 25748
rect 6291 25692 6316 25748
rect 6372 25692 6397 25748
rect 6453 25692 6478 25748
rect 6534 25692 6559 25748
rect 6615 25692 6640 25748
rect 6696 25692 6721 25748
rect 6777 25692 6802 25748
rect 6858 25692 6883 25748
rect 6939 25692 6964 25748
rect 7020 25692 7045 25748
rect 7101 25692 7126 25748
rect 7182 25692 7207 25748
rect 7263 25692 7288 25748
rect 7344 25692 7369 25748
rect 7425 25692 7450 25748
rect 7506 25692 7531 25748
rect 7587 25692 7612 25748
rect 7668 25692 7693 25748
rect 7749 25692 7774 25748
rect 7830 25692 7855 25748
rect 7911 25692 7936 25748
rect 7992 25692 8017 25748
rect 8073 25692 8098 25748
rect 8154 25692 8179 25748
rect 8235 25692 8260 25748
rect 8316 25692 8341 25748
rect 8397 25692 8422 25748
rect 8478 25692 8503 25748
rect 8559 25692 8584 25748
rect 8640 25692 8665 25748
rect 8721 25692 8746 25748
rect 8802 25692 8827 25748
rect 8883 25692 8908 25748
rect 8964 25692 8989 25748
rect 9045 25692 9070 25748
rect 9126 25692 9151 25748
rect 9207 25692 9232 25748
rect 9288 25692 9313 25748
rect 9369 25692 9394 25748
rect 9450 25692 9475 25748
rect 9531 25692 9556 25748
rect 9612 25692 9637 25748
rect 9693 25692 9718 25748
rect 9774 25692 9799 25748
rect 9855 25692 9880 25748
rect 9936 25692 9961 25748
rect 10017 25692 10042 25748
rect 10098 25692 10123 25748
rect 10179 25692 10204 25748
rect 10260 25692 10285 25748
rect 10341 25692 10366 25748
rect 10422 25692 10447 25748
rect 10503 25692 10528 25748
rect 10584 25692 10609 25748
rect 10665 25692 10690 25748
rect 10746 25692 10771 25748
rect 10827 25692 10852 25748
rect 10908 25692 10933 25748
rect 10989 25692 11014 25748
rect 11070 25692 11095 25748
rect 11151 25692 11176 25748
rect 11232 25692 11257 25748
rect 11313 25692 11338 25748
rect 11394 25692 11419 25748
rect 11475 25692 11500 25748
rect 2472 25683 11500 25692
rect 1852 25668 11500 25683
rect 1852 25658 5425 25668
rect 1852 25602 2170 25658
rect 2226 25602 2252 25658
rect 2308 25602 2334 25658
rect 2390 25602 2416 25658
rect 2472 25612 5425 25658
rect 5481 25612 5506 25668
rect 5562 25612 5587 25668
rect 5643 25612 5668 25668
rect 5724 25612 5749 25668
rect 5805 25612 5830 25668
rect 5886 25612 5911 25668
rect 5967 25612 5992 25668
rect 6048 25612 6073 25668
rect 6129 25612 6154 25668
rect 6210 25612 6235 25668
rect 6291 25612 6316 25668
rect 6372 25612 6397 25668
rect 6453 25612 6478 25668
rect 6534 25612 6559 25668
rect 6615 25612 6640 25668
rect 6696 25612 6721 25668
rect 6777 25612 6802 25668
rect 6858 25612 6883 25668
rect 6939 25612 6964 25668
rect 7020 25612 7045 25668
rect 7101 25612 7126 25668
rect 7182 25612 7207 25668
rect 7263 25612 7288 25668
rect 7344 25612 7369 25668
rect 7425 25612 7450 25668
rect 7506 25612 7531 25668
rect 7587 25612 7612 25668
rect 7668 25612 7693 25668
rect 7749 25612 7774 25668
rect 7830 25612 7855 25668
rect 7911 25612 7936 25668
rect 7992 25612 8017 25668
rect 8073 25612 8098 25668
rect 8154 25612 8179 25668
rect 8235 25612 8260 25668
rect 8316 25612 8341 25668
rect 8397 25612 8422 25668
rect 8478 25612 8503 25668
rect 8559 25612 8584 25668
rect 8640 25612 8665 25668
rect 8721 25612 8746 25668
rect 8802 25612 8827 25668
rect 8883 25612 8908 25668
rect 8964 25612 8989 25668
rect 9045 25612 9070 25668
rect 9126 25612 9151 25668
rect 9207 25612 9232 25668
rect 9288 25612 9313 25668
rect 9369 25612 9394 25668
rect 9450 25612 9475 25668
rect 9531 25612 9556 25668
rect 9612 25612 9637 25668
rect 9693 25612 9718 25668
rect 9774 25612 9799 25668
rect 9855 25612 9880 25668
rect 9936 25612 9961 25668
rect 10017 25612 10042 25668
rect 10098 25612 10123 25668
rect 10179 25612 10204 25668
rect 10260 25612 10285 25668
rect 10341 25612 10366 25668
rect 10422 25612 10447 25668
rect 10503 25612 10528 25668
rect 10584 25612 10609 25668
rect 10665 25612 10690 25668
rect 10746 25612 10771 25668
rect 10827 25612 10852 25668
rect 10908 25612 10933 25668
rect 10989 25612 11014 25668
rect 11070 25612 11095 25668
rect 11151 25612 11176 25668
rect 11232 25612 11257 25668
rect 11313 25612 11338 25668
rect 11394 25612 11419 25668
rect 11475 25612 11500 25668
rect 2472 25602 11500 25612
rect 1852 25588 11500 25602
rect 1852 25577 5425 25588
rect 1852 25521 2170 25577
rect 2226 25521 2252 25577
rect 2308 25521 2334 25577
rect 2390 25521 2416 25577
rect 2472 25532 5425 25577
rect 5481 25532 5506 25588
rect 5562 25532 5587 25588
rect 5643 25532 5668 25588
rect 5724 25532 5749 25588
rect 5805 25532 5830 25588
rect 5886 25532 5911 25588
rect 5967 25532 5992 25588
rect 6048 25532 6073 25588
rect 6129 25532 6154 25588
rect 6210 25532 6235 25588
rect 6291 25532 6316 25588
rect 6372 25532 6397 25588
rect 6453 25532 6478 25588
rect 6534 25532 6559 25588
rect 6615 25532 6640 25588
rect 6696 25532 6721 25588
rect 6777 25532 6802 25588
rect 6858 25532 6883 25588
rect 6939 25532 6964 25588
rect 7020 25532 7045 25588
rect 7101 25532 7126 25588
rect 7182 25532 7207 25588
rect 7263 25532 7288 25588
rect 7344 25532 7369 25588
rect 7425 25532 7450 25588
rect 7506 25532 7531 25588
rect 7587 25532 7612 25588
rect 7668 25532 7693 25588
rect 7749 25532 7774 25588
rect 7830 25532 7855 25588
rect 7911 25532 7936 25588
rect 7992 25532 8017 25588
rect 8073 25532 8098 25588
rect 8154 25532 8179 25588
rect 8235 25532 8260 25588
rect 8316 25532 8341 25588
rect 8397 25532 8422 25588
rect 8478 25532 8503 25588
rect 8559 25532 8584 25588
rect 8640 25532 8665 25588
rect 8721 25532 8746 25588
rect 8802 25532 8827 25588
rect 8883 25532 8908 25588
rect 8964 25532 8989 25588
rect 9045 25532 9070 25588
rect 9126 25532 9151 25588
rect 9207 25532 9232 25588
rect 9288 25532 9313 25588
rect 9369 25532 9394 25588
rect 9450 25532 9475 25588
rect 9531 25532 9556 25588
rect 9612 25532 9637 25588
rect 9693 25532 9718 25588
rect 9774 25532 9799 25588
rect 9855 25532 9880 25588
rect 9936 25532 9961 25588
rect 10017 25532 10042 25588
rect 10098 25532 10123 25588
rect 10179 25532 10204 25588
rect 10260 25532 10285 25588
rect 10341 25532 10366 25588
rect 10422 25532 10447 25588
rect 10503 25532 10528 25588
rect 10584 25532 10609 25588
rect 10665 25532 10690 25588
rect 10746 25532 10771 25588
rect 10827 25532 10852 25588
rect 10908 25532 10933 25588
rect 10989 25532 11014 25588
rect 11070 25532 11095 25588
rect 11151 25532 11176 25588
rect 11232 25532 11257 25588
rect 11313 25532 11338 25588
rect 11394 25532 11419 25588
rect 11475 25532 11500 25588
rect 2472 25521 11500 25532
rect 1852 25508 11500 25521
rect 1852 25496 5425 25508
rect 1852 25440 2170 25496
rect 2226 25440 2252 25496
rect 2308 25440 2334 25496
rect 2390 25440 2416 25496
rect 2472 25452 5425 25496
rect 5481 25452 5506 25508
rect 5562 25452 5587 25508
rect 5643 25452 5668 25508
rect 5724 25452 5749 25508
rect 5805 25452 5830 25508
rect 5886 25452 5911 25508
rect 5967 25452 5992 25508
rect 6048 25452 6073 25508
rect 6129 25452 6154 25508
rect 6210 25452 6235 25508
rect 6291 25452 6316 25508
rect 6372 25452 6397 25508
rect 6453 25452 6478 25508
rect 6534 25452 6559 25508
rect 6615 25452 6640 25508
rect 6696 25452 6721 25508
rect 6777 25452 6802 25508
rect 6858 25452 6883 25508
rect 6939 25452 6964 25508
rect 7020 25452 7045 25508
rect 7101 25452 7126 25508
rect 7182 25452 7207 25508
rect 7263 25452 7288 25508
rect 7344 25452 7369 25508
rect 7425 25452 7450 25508
rect 7506 25452 7531 25508
rect 7587 25452 7612 25508
rect 7668 25452 7693 25508
rect 7749 25452 7774 25508
rect 7830 25452 7855 25508
rect 7911 25452 7936 25508
rect 7992 25452 8017 25508
rect 8073 25452 8098 25508
rect 8154 25452 8179 25508
rect 8235 25452 8260 25508
rect 8316 25452 8341 25508
rect 8397 25452 8422 25508
rect 8478 25452 8503 25508
rect 8559 25452 8584 25508
rect 8640 25452 8665 25508
rect 8721 25452 8746 25508
rect 8802 25452 8827 25508
rect 8883 25452 8908 25508
rect 8964 25452 8989 25508
rect 9045 25452 9070 25508
rect 9126 25452 9151 25508
rect 9207 25452 9232 25508
rect 9288 25452 9313 25508
rect 9369 25452 9394 25508
rect 9450 25452 9475 25508
rect 9531 25452 9556 25508
rect 9612 25452 9637 25508
rect 9693 25452 9718 25508
rect 9774 25452 9799 25508
rect 9855 25452 9880 25508
rect 9936 25452 9961 25508
rect 10017 25452 10042 25508
rect 10098 25452 10123 25508
rect 10179 25452 10204 25508
rect 10260 25452 10285 25508
rect 10341 25452 10366 25508
rect 10422 25452 10447 25508
rect 10503 25452 10528 25508
rect 10584 25452 10609 25508
rect 10665 25452 10690 25508
rect 10746 25452 10771 25508
rect 10827 25452 10852 25508
rect 10908 25452 10933 25508
rect 10989 25452 11014 25508
rect 11070 25452 11095 25508
rect 11151 25452 11176 25508
rect 11232 25452 11257 25508
rect 11313 25452 11338 25508
rect 11394 25452 11419 25508
rect 11475 25452 11500 25508
rect 2472 25440 11500 25452
rect 1852 25428 11500 25440
rect 1852 25415 5425 25428
rect 1852 25359 2170 25415
rect 2226 25359 2252 25415
rect 2308 25359 2334 25415
rect 2390 25359 2416 25415
rect 2472 25372 5425 25415
rect 5481 25372 5506 25428
rect 5562 25372 5587 25428
rect 5643 25372 5668 25428
rect 5724 25372 5749 25428
rect 5805 25372 5830 25428
rect 5886 25372 5911 25428
rect 5967 25372 5992 25428
rect 6048 25372 6073 25428
rect 6129 25372 6154 25428
rect 6210 25372 6235 25428
rect 6291 25372 6316 25428
rect 6372 25372 6397 25428
rect 6453 25372 6478 25428
rect 6534 25372 6559 25428
rect 6615 25372 6640 25428
rect 6696 25372 6721 25428
rect 6777 25372 6802 25428
rect 6858 25372 6883 25428
rect 6939 25372 6964 25428
rect 7020 25372 7045 25428
rect 7101 25372 7126 25428
rect 7182 25372 7207 25428
rect 7263 25372 7288 25428
rect 7344 25372 7369 25428
rect 7425 25372 7450 25428
rect 7506 25372 7531 25428
rect 7587 25372 7612 25428
rect 7668 25372 7693 25428
rect 7749 25372 7774 25428
rect 7830 25372 7855 25428
rect 7911 25372 7936 25428
rect 7992 25372 8017 25428
rect 8073 25372 8098 25428
rect 8154 25372 8179 25428
rect 8235 25372 8260 25428
rect 8316 25372 8341 25428
rect 8397 25372 8422 25428
rect 8478 25372 8503 25428
rect 8559 25372 8584 25428
rect 8640 25372 8665 25428
rect 8721 25372 8746 25428
rect 8802 25372 8827 25428
rect 8883 25372 8908 25428
rect 8964 25372 8989 25428
rect 9045 25372 9070 25428
rect 9126 25372 9151 25428
rect 9207 25372 9232 25428
rect 9288 25372 9313 25428
rect 9369 25372 9394 25428
rect 9450 25372 9475 25428
rect 9531 25372 9556 25428
rect 9612 25372 9637 25428
rect 9693 25372 9718 25428
rect 9774 25372 9799 25428
rect 9855 25372 9880 25428
rect 9936 25372 9961 25428
rect 10017 25372 10042 25428
rect 10098 25372 10123 25428
rect 10179 25372 10204 25428
rect 10260 25372 10285 25428
rect 10341 25372 10366 25428
rect 10422 25372 10447 25428
rect 10503 25372 10528 25428
rect 10584 25372 10609 25428
rect 10665 25372 10690 25428
rect 10746 25372 10771 25428
rect 10827 25372 10852 25428
rect 10908 25372 10933 25428
rect 10989 25372 11014 25428
rect 11070 25372 11095 25428
rect 11151 25372 11176 25428
rect 11232 25372 11257 25428
rect 11313 25372 11338 25428
rect 11394 25372 11419 25428
rect 11475 25372 11500 25428
rect 2472 25359 11500 25372
rect 1852 25348 11500 25359
rect 1852 25334 5425 25348
rect 1852 25278 2170 25334
rect 2226 25278 2252 25334
rect 2308 25278 2334 25334
rect 2390 25278 2416 25334
rect 2472 25292 5425 25334
rect 5481 25292 5506 25348
rect 5562 25292 5587 25348
rect 5643 25292 5668 25348
rect 5724 25292 5749 25348
rect 5805 25292 5830 25348
rect 5886 25292 5911 25348
rect 5967 25292 5992 25348
rect 6048 25292 6073 25348
rect 6129 25292 6154 25348
rect 6210 25292 6235 25348
rect 6291 25292 6316 25348
rect 6372 25292 6397 25348
rect 6453 25292 6478 25348
rect 6534 25292 6559 25348
rect 6615 25292 6640 25348
rect 6696 25292 6721 25348
rect 6777 25292 6802 25348
rect 6858 25292 6883 25348
rect 6939 25292 6964 25348
rect 7020 25292 7045 25348
rect 7101 25292 7126 25348
rect 7182 25292 7207 25348
rect 7263 25292 7288 25348
rect 7344 25292 7369 25348
rect 7425 25292 7450 25348
rect 7506 25292 7531 25348
rect 7587 25292 7612 25348
rect 7668 25292 7693 25348
rect 7749 25292 7774 25348
rect 7830 25292 7855 25348
rect 7911 25292 7936 25348
rect 7992 25292 8017 25348
rect 8073 25292 8098 25348
rect 8154 25292 8179 25348
rect 8235 25292 8260 25348
rect 8316 25292 8341 25348
rect 8397 25292 8422 25348
rect 8478 25292 8503 25348
rect 8559 25292 8584 25348
rect 8640 25292 8665 25348
rect 8721 25292 8746 25348
rect 8802 25292 8827 25348
rect 8883 25292 8908 25348
rect 8964 25292 8989 25348
rect 9045 25292 9070 25348
rect 9126 25292 9151 25348
rect 9207 25292 9232 25348
rect 9288 25292 9313 25348
rect 9369 25292 9394 25348
rect 9450 25292 9475 25348
rect 9531 25292 9556 25348
rect 9612 25292 9637 25348
rect 9693 25292 9718 25348
rect 9774 25292 9799 25348
rect 9855 25292 9880 25348
rect 9936 25292 9961 25348
rect 10017 25292 10042 25348
rect 10098 25292 10123 25348
rect 10179 25292 10204 25348
rect 10260 25292 10285 25348
rect 10341 25292 10366 25348
rect 10422 25292 10447 25348
rect 10503 25292 10528 25348
rect 10584 25292 10609 25348
rect 10665 25292 10690 25348
rect 10746 25292 10771 25348
rect 10827 25292 10852 25348
rect 10908 25292 10933 25348
rect 10989 25292 11014 25348
rect 11070 25292 11095 25348
rect 11151 25292 11176 25348
rect 11232 25292 11257 25348
rect 11313 25292 11338 25348
rect 11394 25292 11419 25348
rect 11475 25292 11500 25348
rect 2472 25278 11500 25292
rect 1852 25268 11500 25278
rect 1852 25253 5425 25268
rect 1852 25197 2170 25253
rect 2226 25197 2252 25253
rect 2308 25197 2334 25253
rect 2390 25197 2416 25253
rect 2472 25212 5425 25253
rect 5481 25212 5506 25268
rect 5562 25212 5587 25268
rect 5643 25212 5668 25268
rect 5724 25212 5749 25268
rect 5805 25212 5830 25268
rect 5886 25212 5911 25268
rect 5967 25212 5992 25268
rect 6048 25212 6073 25268
rect 6129 25212 6154 25268
rect 6210 25212 6235 25268
rect 6291 25212 6316 25268
rect 6372 25212 6397 25268
rect 6453 25212 6478 25268
rect 6534 25212 6559 25268
rect 6615 25212 6640 25268
rect 6696 25212 6721 25268
rect 6777 25212 6802 25268
rect 6858 25212 6883 25268
rect 6939 25212 6964 25268
rect 7020 25212 7045 25268
rect 7101 25212 7126 25268
rect 7182 25212 7207 25268
rect 7263 25212 7288 25268
rect 7344 25212 7369 25268
rect 7425 25212 7450 25268
rect 7506 25212 7531 25268
rect 7587 25212 7612 25268
rect 7668 25212 7693 25268
rect 7749 25212 7774 25268
rect 7830 25212 7855 25268
rect 7911 25212 7936 25268
rect 7992 25212 8017 25268
rect 8073 25212 8098 25268
rect 8154 25212 8179 25268
rect 8235 25212 8260 25268
rect 8316 25212 8341 25268
rect 8397 25212 8422 25268
rect 8478 25212 8503 25268
rect 8559 25212 8584 25268
rect 8640 25212 8665 25268
rect 8721 25212 8746 25268
rect 8802 25212 8827 25268
rect 8883 25212 8908 25268
rect 8964 25212 8989 25268
rect 9045 25212 9070 25268
rect 9126 25212 9151 25268
rect 9207 25212 9232 25268
rect 9288 25212 9313 25268
rect 9369 25212 9394 25268
rect 9450 25212 9475 25268
rect 9531 25212 9556 25268
rect 9612 25212 9637 25268
rect 9693 25212 9718 25268
rect 9774 25212 9799 25268
rect 9855 25212 9880 25268
rect 9936 25212 9961 25268
rect 10017 25212 10042 25268
rect 10098 25212 10123 25268
rect 10179 25212 10204 25268
rect 10260 25212 10285 25268
rect 10341 25212 10366 25268
rect 10422 25212 10447 25268
rect 10503 25212 10528 25268
rect 10584 25212 10609 25268
rect 10665 25212 10690 25268
rect 10746 25212 10771 25268
rect 10827 25212 10852 25268
rect 10908 25212 10933 25268
rect 10989 25212 11014 25268
rect 11070 25212 11095 25268
rect 11151 25212 11176 25268
rect 11232 25212 11257 25268
rect 11313 25212 11338 25268
rect 11394 25212 11419 25268
rect 11475 25212 11500 25268
rect 2472 25197 11500 25212
rect 1852 25188 11500 25197
rect 1852 25172 5425 25188
rect 1852 25116 2170 25172
rect 2226 25116 2252 25172
rect 2308 25116 2334 25172
rect 2390 25116 2416 25172
rect 2472 25132 5425 25172
rect 5481 25132 5506 25188
rect 5562 25132 5587 25188
rect 5643 25132 5668 25188
rect 5724 25132 5749 25188
rect 5805 25132 5830 25188
rect 5886 25132 5911 25188
rect 5967 25132 5992 25188
rect 6048 25132 6073 25188
rect 6129 25132 6154 25188
rect 6210 25132 6235 25188
rect 6291 25132 6316 25188
rect 6372 25132 6397 25188
rect 6453 25132 6478 25188
rect 6534 25132 6559 25188
rect 6615 25132 6640 25188
rect 6696 25132 6721 25188
rect 6777 25132 6802 25188
rect 6858 25132 6883 25188
rect 6939 25132 6964 25188
rect 7020 25132 7045 25188
rect 7101 25132 7126 25188
rect 7182 25132 7207 25188
rect 7263 25132 7288 25188
rect 7344 25132 7369 25188
rect 7425 25132 7450 25188
rect 7506 25132 7531 25188
rect 7587 25132 7612 25188
rect 7668 25132 7693 25188
rect 7749 25132 7774 25188
rect 7830 25132 7855 25188
rect 7911 25132 7936 25188
rect 7992 25132 8017 25188
rect 8073 25132 8098 25188
rect 8154 25132 8179 25188
rect 8235 25132 8260 25188
rect 8316 25132 8341 25188
rect 8397 25132 8422 25188
rect 8478 25132 8503 25188
rect 8559 25132 8584 25188
rect 8640 25132 8665 25188
rect 8721 25132 8746 25188
rect 8802 25132 8827 25188
rect 8883 25132 8908 25188
rect 8964 25132 8989 25188
rect 9045 25132 9070 25188
rect 9126 25132 9151 25188
rect 9207 25132 9232 25188
rect 9288 25132 9313 25188
rect 9369 25132 9394 25188
rect 9450 25132 9475 25188
rect 9531 25132 9556 25188
rect 9612 25132 9637 25188
rect 9693 25132 9718 25188
rect 9774 25132 9799 25188
rect 9855 25132 9880 25188
rect 9936 25132 9961 25188
rect 10017 25132 10042 25188
rect 10098 25132 10123 25188
rect 10179 25132 10204 25188
rect 10260 25132 10285 25188
rect 10341 25132 10366 25188
rect 10422 25132 10447 25188
rect 10503 25132 10528 25188
rect 10584 25132 10609 25188
rect 10665 25132 10690 25188
rect 10746 25132 10771 25188
rect 10827 25132 10852 25188
rect 10908 25132 10933 25188
rect 10989 25132 11014 25188
rect 11070 25132 11095 25188
rect 11151 25132 11176 25188
rect 11232 25132 11257 25188
rect 11313 25132 11338 25188
rect 11394 25132 11419 25188
rect 11475 25132 11500 25188
rect 2472 25116 11500 25132
rect 1852 25108 11500 25116
rect 1852 25091 5425 25108
rect 1852 25035 2170 25091
rect 2226 25035 2252 25091
rect 2308 25035 2334 25091
rect 2390 25035 2416 25091
rect 2472 25052 5425 25091
rect 5481 25052 5506 25108
rect 5562 25052 5587 25108
rect 5643 25052 5668 25108
rect 5724 25052 5749 25108
rect 5805 25052 5830 25108
rect 5886 25052 5911 25108
rect 5967 25052 5992 25108
rect 6048 25052 6073 25108
rect 6129 25052 6154 25108
rect 6210 25052 6235 25108
rect 6291 25052 6316 25108
rect 6372 25052 6397 25108
rect 6453 25052 6478 25108
rect 6534 25052 6559 25108
rect 6615 25052 6640 25108
rect 6696 25052 6721 25108
rect 6777 25052 6802 25108
rect 6858 25052 6883 25108
rect 6939 25052 6964 25108
rect 7020 25052 7045 25108
rect 7101 25052 7126 25108
rect 7182 25052 7207 25108
rect 7263 25052 7288 25108
rect 7344 25052 7369 25108
rect 7425 25052 7450 25108
rect 7506 25052 7531 25108
rect 7587 25052 7612 25108
rect 7668 25052 7693 25108
rect 7749 25052 7774 25108
rect 7830 25052 7855 25108
rect 7911 25052 7936 25108
rect 7992 25052 8017 25108
rect 8073 25052 8098 25108
rect 8154 25052 8179 25108
rect 8235 25052 8260 25108
rect 8316 25052 8341 25108
rect 8397 25052 8422 25108
rect 8478 25052 8503 25108
rect 8559 25052 8584 25108
rect 8640 25052 8665 25108
rect 8721 25052 8746 25108
rect 8802 25052 8827 25108
rect 8883 25052 8908 25108
rect 8964 25052 8989 25108
rect 9045 25052 9070 25108
rect 9126 25052 9151 25108
rect 9207 25052 9232 25108
rect 9288 25052 9313 25108
rect 9369 25052 9394 25108
rect 9450 25052 9475 25108
rect 9531 25052 9556 25108
rect 9612 25052 9637 25108
rect 9693 25052 9718 25108
rect 9774 25052 9799 25108
rect 9855 25052 9880 25108
rect 9936 25052 9961 25108
rect 10017 25052 10042 25108
rect 10098 25052 10123 25108
rect 10179 25052 10204 25108
rect 10260 25052 10285 25108
rect 10341 25052 10366 25108
rect 10422 25052 10447 25108
rect 10503 25052 10528 25108
rect 10584 25052 10609 25108
rect 10665 25052 10690 25108
rect 10746 25052 10771 25108
rect 10827 25052 10852 25108
rect 10908 25052 10933 25108
rect 10989 25052 11014 25108
rect 11070 25052 11095 25108
rect 11151 25052 11176 25108
rect 11232 25052 11257 25108
rect 11313 25052 11338 25108
rect 11394 25052 11419 25108
rect 11475 25052 11500 25108
rect 2472 25035 11500 25052
rect 1852 25028 11500 25035
rect 1852 25010 5425 25028
rect 1852 24954 2170 25010
rect 2226 24954 2252 25010
rect 2308 24954 2334 25010
rect 2390 24954 2416 25010
rect 2472 24972 5425 25010
rect 5481 24972 5506 25028
rect 5562 24972 5587 25028
rect 5643 24972 5668 25028
rect 5724 24972 5749 25028
rect 5805 24972 5830 25028
rect 5886 24972 5911 25028
rect 5967 24972 5992 25028
rect 6048 24972 6073 25028
rect 6129 24972 6154 25028
rect 6210 24972 6235 25028
rect 6291 24972 6316 25028
rect 6372 24972 6397 25028
rect 6453 24972 6478 25028
rect 6534 24972 6559 25028
rect 6615 24972 6640 25028
rect 6696 24972 6721 25028
rect 6777 24972 6802 25028
rect 6858 24972 6883 25028
rect 6939 24972 6964 25028
rect 7020 24972 7045 25028
rect 7101 24972 7126 25028
rect 7182 24972 7207 25028
rect 7263 24972 7288 25028
rect 7344 24972 7369 25028
rect 7425 24972 7450 25028
rect 7506 24972 7531 25028
rect 7587 24972 7612 25028
rect 7668 24972 7693 25028
rect 7749 24972 7774 25028
rect 7830 24972 7855 25028
rect 7911 24972 7936 25028
rect 7992 24972 8017 25028
rect 8073 24972 8098 25028
rect 8154 24972 8179 25028
rect 8235 24972 8260 25028
rect 8316 24972 8341 25028
rect 8397 24972 8422 25028
rect 8478 24972 8503 25028
rect 8559 24972 8584 25028
rect 8640 24972 8665 25028
rect 8721 24972 8746 25028
rect 8802 24972 8827 25028
rect 8883 24972 8908 25028
rect 8964 24972 8989 25028
rect 9045 24972 9070 25028
rect 9126 24972 9151 25028
rect 9207 24972 9232 25028
rect 9288 24972 9313 25028
rect 9369 24972 9394 25028
rect 9450 24972 9475 25028
rect 9531 24972 9556 25028
rect 9612 24972 9637 25028
rect 9693 24972 9718 25028
rect 9774 24972 9799 25028
rect 9855 24972 9880 25028
rect 9936 24972 9961 25028
rect 10017 24972 10042 25028
rect 10098 24972 10123 25028
rect 10179 24972 10204 25028
rect 10260 24972 10285 25028
rect 10341 24972 10366 25028
rect 10422 24972 10447 25028
rect 10503 24972 10528 25028
rect 10584 24972 10609 25028
rect 10665 24972 10690 25028
rect 10746 24972 10771 25028
rect 10827 24972 10852 25028
rect 10908 24972 10933 25028
rect 10989 24972 11014 25028
rect 11070 24972 11095 25028
rect 11151 24972 11176 25028
rect 11232 24972 11257 25028
rect 11313 24972 11338 25028
rect 11394 24972 11419 25028
rect 11475 24972 11500 25028
rect 2472 24954 11500 24972
rect 1852 24948 11500 24954
rect 1852 24929 5425 24948
rect 1852 24873 2170 24929
rect 2226 24873 2252 24929
rect 2308 24873 2334 24929
rect 2390 24873 2416 24929
rect 2472 24892 5425 24929
rect 5481 24892 5506 24948
rect 5562 24892 5587 24948
rect 5643 24892 5668 24948
rect 5724 24892 5749 24948
rect 5805 24892 5830 24948
rect 5886 24892 5911 24948
rect 5967 24892 5992 24948
rect 6048 24892 6073 24948
rect 6129 24892 6154 24948
rect 6210 24892 6235 24948
rect 6291 24892 6316 24948
rect 6372 24892 6397 24948
rect 6453 24892 6478 24948
rect 6534 24892 6559 24948
rect 6615 24892 6640 24948
rect 6696 24892 6721 24948
rect 6777 24892 6802 24948
rect 6858 24892 6883 24948
rect 6939 24892 6964 24948
rect 7020 24892 7045 24948
rect 7101 24892 7126 24948
rect 7182 24892 7207 24948
rect 7263 24892 7288 24948
rect 7344 24892 7369 24948
rect 7425 24892 7450 24948
rect 7506 24892 7531 24948
rect 7587 24892 7612 24948
rect 7668 24892 7693 24948
rect 7749 24892 7774 24948
rect 7830 24892 7855 24948
rect 7911 24892 7936 24948
rect 7992 24892 8017 24948
rect 8073 24892 8098 24948
rect 8154 24892 8179 24948
rect 8235 24892 8260 24948
rect 8316 24892 8341 24948
rect 8397 24892 8422 24948
rect 8478 24892 8503 24948
rect 8559 24892 8584 24948
rect 8640 24892 8665 24948
rect 8721 24892 8746 24948
rect 8802 24892 8827 24948
rect 8883 24892 8908 24948
rect 8964 24892 8989 24948
rect 9045 24892 9070 24948
rect 9126 24892 9151 24948
rect 9207 24892 9232 24948
rect 9288 24892 9313 24948
rect 9369 24892 9394 24948
rect 9450 24892 9475 24948
rect 9531 24892 9556 24948
rect 9612 24892 9637 24948
rect 9693 24892 9718 24948
rect 9774 24892 9799 24948
rect 9855 24892 9880 24948
rect 9936 24892 9961 24948
rect 10017 24892 10042 24948
rect 10098 24892 10123 24948
rect 10179 24892 10204 24948
rect 10260 24892 10285 24948
rect 10341 24892 10366 24948
rect 10422 24892 10447 24948
rect 10503 24892 10528 24948
rect 10584 24892 10609 24948
rect 10665 24892 10690 24948
rect 10746 24892 10771 24948
rect 10827 24892 10852 24948
rect 10908 24892 10933 24948
rect 10989 24892 11014 24948
rect 11070 24892 11095 24948
rect 11151 24892 11176 24948
rect 11232 24892 11257 24948
rect 11313 24892 11338 24948
rect 11394 24892 11419 24948
rect 11475 24892 11500 24948
rect 2472 24873 11500 24892
rect 1852 24868 11500 24873
rect 1852 24848 5425 24868
rect 1852 24792 2170 24848
rect 2226 24792 2252 24848
rect 2308 24792 2334 24848
rect 2390 24792 2416 24848
rect 2472 24812 5425 24848
rect 5481 24812 5506 24868
rect 5562 24812 5587 24868
rect 5643 24812 5668 24868
rect 5724 24812 5749 24868
rect 5805 24812 5830 24868
rect 5886 24812 5911 24868
rect 5967 24812 5992 24868
rect 6048 24812 6073 24868
rect 6129 24812 6154 24868
rect 6210 24812 6235 24868
rect 6291 24812 6316 24868
rect 6372 24812 6397 24868
rect 6453 24812 6478 24868
rect 6534 24812 6559 24868
rect 6615 24812 6640 24868
rect 6696 24812 6721 24868
rect 6777 24812 6802 24868
rect 6858 24812 6883 24868
rect 6939 24812 6964 24868
rect 7020 24812 7045 24868
rect 7101 24812 7126 24868
rect 7182 24812 7207 24868
rect 7263 24812 7288 24868
rect 7344 24812 7369 24868
rect 7425 24812 7450 24868
rect 7506 24812 7531 24868
rect 7587 24812 7612 24868
rect 7668 24812 7693 24868
rect 7749 24812 7774 24868
rect 7830 24812 7855 24868
rect 7911 24812 7936 24868
rect 7992 24812 8017 24868
rect 8073 24812 8098 24868
rect 8154 24812 8179 24868
rect 8235 24812 8260 24868
rect 8316 24812 8341 24868
rect 8397 24812 8422 24868
rect 8478 24812 8503 24868
rect 8559 24812 8584 24868
rect 8640 24812 8665 24868
rect 8721 24812 8746 24868
rect 8802 24812 8827 24868
rect 8883 24812 8908 24868
rect 8964 24812 8989 24868
rect 9045 24812 9070 24868
rect 9126 24812 9151 24868
rect 9207 24812 9232 24868
rect 9288 24812 9313 24868
rect 9369 24812 9394 24868
rect 9450 24812 9475 24868
rect 9531 24812 9556 24868
rect 9612 24812 9637 24868
rect 9693 24812 9718 24868
rect 9774 24812 9799 24868
rect 9855 24812 9880 24868
rect 9936 24812 9961 24868
rect 10017 24812 10042 24868
rect 10098 24812 10123 24868
rect 10179 24812 10204 24868
rect 10260 24812 10285 24868
rect 10341 24812 10366 24868
rect 10422 24812 10447 24868
rect 10503 24812 10528 24868
rect 10584 24812 10609 24868
rect 10665 24812 10690 24868
rect 10746 24812 10771 24868
rect 10827 24812 10852 24868
rect 10908 24812 10933 24868
rect 10989 24812 11014 24868
rect 11070 24812 11095 24868
rect 11151 24812 11176 24868
rect 11232 24812 11257 24868
rect 11313 24812 11338 24868
rect 11394 24812 11419 24868
rect 11475 24812 11500 24868
rect 2472 24792 11500 24812
rect 1852 24788 11500 24792
rect 1852 24767 5425 24788
rect 1852 24711 2170 24767
rect 2226 24711 2252 24767
rect 2308 24711 2334 24767
rect 2390 24711 2416 24767
rect 2472 24732 5425 24767
rect 5481 24732 5506 24788
rect 5562 24732 5587 24788
rect 5643 24732 5668 24788
rect 5724 24732 5749 24788
rect 5805 24732 5830 24788
rect 5886 24732 5911 24788
rect 5967 24732 5992 24788
rect 6048 24732 6073 24788
rect 6129 24732 6154 24788
rect 6210 24732 6235 24788
rect 6291 24732 6316 24788
rect 6372 24732 6397 24788
rect 6453 24732 6478 24788
rect 6534 24732 6559 24788
rect 6615 24732 6640 24788
rect 6696 24732 6721 24788
rect 6777 24732 6802 24788
rect 6858 24732 6883 24788
rect 6939 24732 6964 24788
rect 7020 24732 7045 24788
rect 7101 24732 7126 24788
rect 7182 24732 7207 24788
rect 7263 24732 7288 24788
rect 7344 24732 7369 24788
rect 7425 24732 7450 24788
rect 7506 24732 7531 24788
rect 7587 24732 7612 24788
rect 7668 24732 7693 24788
rect 7749 24732 7774 24788
rect 7830 24732 7855 24788
rect 7911 24732 7936 24788
rect 7992 24732 8017 24788
rect 8073 24732 8098 24788
rect 8154 24732 8179 24788
rect 8235 24732 8260 24788
rect 8316 24732 8341 24788
rect 8397 24732 8422 24788
rect 8478 24732 8503 24788
rect 8559 24732 8584 24788
rect 8640 24732 8665 24788
rect 8721 24732 8746 24788
rect 8802 24732 8827 24788
rect 8883 24732 8908 24788
rect 8964 24732 8989 24788
rect 9045 24732 9070 24788
rect 9126 24732 9151 24788
rect 9207 24732 9232 24788
rect 9288 24732 9313 24788
rect 9369 24732 9394 24788
rect 9450 24732 9475 24788
rect 9531 24732 9556 24788
rect 9612 24732 9637 24788
rect 9693 24732 9718 24788
rect 9774 24732 9799 24788
rect 9855 24732 9880 24788
rect 9936 24732 9961 24788
rect 10017 24732 10042 24788
rect 10098 24732 10123 24788
rect 10179 24732 10204 24788
rect 10260 24732 10285 24788
rect 10341 24732 10366 24788
rect 10422 24732 10447 24788
rect 10503 24732 10528 24788
rect 10584 24732 10609 24788
rect 10665 24732 10690 24788
rect 10746 24732 10771 24788
rect 10827 24732 10852 24788
rect 10908 24732 10933 24788
rect 10989 24732 11014 24788
rect 11070 24732 11095 24788
rect 11151 24732 11176 24788
rect 11232 24732 11257 24788
rect 11313 24732 11338 24788
rect 11394 24732 11419 24788
rect 11475 24732 11500 24788
rect 2472 24711 11500 24732
rect 1852 24708 11500 24711
rect 1852 24686 5425 24708
rect 1852 24630 2170 24686
rect 2226 24630 2252 24686
rect 2308 24630 2334 24686
rect 2390 24630 2416 24686
rect 2472 24652 5425 24686
rect 5481 24652 5506 24708
rect 5562 24652 5587 24708
rect 5643 24652 5668 24708
rect 5724 24652 5749 24708
rect 5805 24652 5830 24708
rect 5886 24652 5911 24708
rect 5967 24652 5992 24708
rect 6048 24652 6073 24708
rect 6129 24652 6154 24708
rect 6210 24652 6235 24708
rect 6291 24652 6316 24708
rect 6372 24652 6397 24708
rect 6453 24652 6478 24708
rect 6534 24652 6559 24708
rect 6615 24652 6640 24708
rect 6696 24652 6721 24708
rect 6777 24652 6802 24708
rect 6858 24652 6883 24708
rect 6939 24652 6964 24708
rect 7020 24652 7045 24708
rect 7101 24652 7126 24708
rect 7182 24652 7207 24708
rect 7263 24652 7288 24708
rect 7344 24652 7369 24708
rect 7425 24652 7450 24708
rect 7506 24652 7531 24708
rect 7587 24652 7612 24708
rect 7668 24652 7693 24708
rect 7749 24652 7774 24708
rect 7830 24652 7855 24708
rect 7911 24652 7936 24708
rect 7992 24652 8017 24708
rect 8073 24652 8098 24708
rect 8154 24652 8179 24708
rect 8235 24652 8260 24708
rect 8316 24652 8341 24708
rect 8397 24652 8422 24708
rect 8478 24652 8503 24708
rect 8559 24652 8584 24708
rect 8640 24652 8665 24708
rect 8721 24652 8746 24708
rect 8802 24652 8827 24708
rect 8883 24652 8908 24708
rect 8964 24652 8989 24708
rect 9045 24652 9070 24708
rect 9126 24652 9151 24708
rect 9207 24652 9232 24708
rect 9288 24652 9313 24708
rect 9369 24652 9394 24708
rect 9450 24652 9475 24708
rect 9531 24652 9556 24708
rect 9612 24652 9637 24708
rect 9693 24652 9718 24708
rect 9774 24652 9799 24708
rect 9855 24652 9880 24708
rect 9936 24652 9961 24708
rect 10017 24652 10042 24708
rect 10098 24652 10123 24708
rect 10179 24652 10204 24708
rect 10260 24652 10285 24708
rect 10341 24652 10366 24708
rect 10422 24652 10447 24708
rect 10503 24652 10528 24708
rect 10584 24652 10609 24708
rect 10665 24652 10690 24708
rect 10746 24652 10771 24708
rect 10827 24652 10852 24708
rect 10908 24652 10933 24708
rect 10989 24652 11014 24708
rect 11070 24652 11095 24708
rect 11151 24652 11176 24708
rect 11232 24652 11257 24708
rect 11313 24652 11338 24708
rect 11394 24652 11419 24708
rect 11475 24652 11500 24708
rect 13076 25822 15047 25828
rect 13076 25766 14509 25822
rect 14565 25766 14603 25822
rect 14659 25766 14697 25822
rect 14753 25766 14791 25822
rect 14847 25766 14885 25822
rect 14941 25766 14979 25822
rect 15035 25766 15047 25822
rect 13076 25741 15047 25766
rect 13076 25685 14509 25741
rect 14565 25685 14603 25741
rect 14659 25685 14697 25741
rect 14753 25685 14791 25741
rect 14847 25685 14885 25741
rect 14941 25685 14979 25741
rect 15035 25685 15047 25741
rect 13076 25660 15047 25685
rect 13076 25604 14509 25660
rect 14565 25604 14603 25660
rect 14659 25604 14697 25660
rect 14753 25604 14791 25660
rect 14847 25604 14885 25660
rect 14941 25604 14979 25660
rect 15035 25604 15047 25660
rect 13076 25579 15047 25604
rect 13076 25523 14509 25579
rect 14565 25523 14603 25579
rect 14659 25523 14697 25579
rect 14753 25523 14791 25579
rect 14847 25523 14885 25579
rect 14941 25523 14979 25579
rect 15035 25523 15047 25579
rect 13076 25498 15047 25523
rect 13076 25442 14509 25498
rect 14565 25442 14603 25498
rect 14659 25442 14697 25498
rect 14753 25442 14791 25498
rect 14847 25442 14885 25498
rect 14941 25442 14979 25498
rect 15035 25442 15047 25498
rect 13076 25417 15047 25442
rect 13076 25361 14509 25417
rect 14565 25361 14603 25417
rect 14659 25361 14697 25417
rect 14753 25361 14791 25417
rect 14847 25361 14885 25417
rect 14941 25361 14979 25417
rect 15035 25361 15047 25417
rect 13076 25336 15047 25361
rect 13076 25280 14509 25336
rect 14565 25280 14603 25336
rect 14659 25280 14697 25336
rect 14753 25280 14791 25336
rect 14847 25280 14885 25336
rect 14941 25280 14979 25336
rect 15035 25280 15047 25336
rect 13076 25255 15047 25280
rect 13076 25199 14509 25255
rect 14565 25199 14603 25255
rect 14659 25199 14697 25255
rect 14753 25199 14791 25255
rect 14847 25199 14885 25255
rect 14941 25199 14979 25255
rect 15035 25199 15047 25255
rect 13076 25174 15047 25199
rect 13076 25118 14509 25174
rect 14565 25118 14603 25174
rect 14659 25118 14697 25174
rect 14753 25118 14791 25174
rect 14847 25118 14885 25174
rect 14941 25118 14979 25174
rect 15035 25118 15047 25174
rect 13076 25093 15047 25118
rect 13076 25037 14509 25093
rect 14565 25037 14603 25093
rect 14659 25037 14697 25093
rect 14753 25037 14791 25093
rect 14847 25037 14885 25093
rect 14941 25037 14979 25093
rect 15035 25037 15047 25093
rect 13076 25011 15047 25037
rect 13076 24955 14509 25011
rect 14565 24955 14603 25011
rect 14659 24955 14697 25011
rect 14753 24955 14791 25011
rect 14847 24955 14885 25011
rect 14941 24955 14979 25011
rect 15035 24955 15047 25011
rect 13076 24929 15047 24955
rect 13076 24873 14509 24929
rect 14565 24873 14603 24929
rect 14659 24873 14697 24929
rect 14753 24873 14791 24929
rect 14847 24873 14885 24929
rect 14941 24873 14979 24929
rect 15035 24873 15047 24929
rect 13076 24847 15047 24873
rect 13076 24791 14509 24847
rect 14565 24791 14603 24847
rect 14659 24791 14697 24847
rect 14753 24791 14791 24847
rect 14847 24791 14885 24847
rect 14941 24791 14979 24847
rect 15035 24791 15047 24847
rect 13076 24765 15047 24791
rect 13076 24709 14509 24765
rect 14565 24709 14603 24765
rect 14659 24709 14697 24765
rect 14753 24709 14791 24765
rect 14847 24709 14885 24765
rect 14941 24709 14979 24765
rect 15035 24709 15047 24765
rect 13076 24683 15047 24709
rect 13076 24652 14509 24683
rect 2472 24630 14509 24652
rect 1852 24627 14509 24630
rect 14565 24627 14603 24683
rect 14659 24627 14697 24683
rect 14753 24627 14791 24683
rect 14847 24627 14885 24683
rect 14941 24627 14979 24683
rect 15035 24627 15047 24683
rect 1852 24604 15047 24627
rect 1852 24548 2170 24604
rect 2226 24548 2252 24604
rect 2308 24548 2334 24604
rect 2390 24548 2416 24604
rect 2472 24601 15047 24604
rect 2472 24548 14509 24601
rect 1852 24545 14509 24548
rect 14565 24545 14603 24601
rect 14659 24545 14697 24601
rect 14753 24545 14791 24601
rect 14847 24545 14885 24601
rect 14941 24545 14979 24601
rect 15035 24545 15047 24601
rect 1852 24522 15047 24545
rect 1852 24466 2170 24522
rect 2226 24466 2252 24522
rect 2308 24466 2334 24522
rect 2390 24466 2416 24522
rect 2472 24519 15047 24522
rect 2472 24466 14509 24519
rect 1852 24463 14509 24466
rect 14565 24463 14603 24519
rect 14659 24463 14697 24519
rect 14753 24463 14791 24519
rect 14847 24463 14885 24519
rect 14941 24463 14979 24519
rect 15035 24463 15047 24519
rect 1852 24440 15047 24463
rect 1852 24384 2170 24440
rect 2226 24384 2252 24440
rect 2308 24384 2334 24440
rect 2390 24384 2416 24440
rect 2472 24437 15047 24440
rect 2472 24384 14509 24437
rect 1852 24381 14509 24384
rect 14565 24381 14603 24437
rect 14659 24381 14697 24437
rect 14753 24381 14791 24437
rect 14847 24381 14885 24437
rect 14941 24381 14979 24437
rect 15035 24381 15047 24437
rect 1852 24358 15047 24381
rect 1852 24302 2170 24358
rect 2226 24302 2252 24358
rect 2308 24302 2334 24358
rect 2390 24302 2416 24358
rect 2472 24355 15047 24358
rect 2472 24323 14509 24355
rect 2472 24302 5425 24323
rect 1852 24276 5425 24302
rect 1852 24220 2170 24276
rect 2226 24220 2252 24276
rect 2308 24220 2334 24276
rect 2390 24220 2416 24276
rect 2472 24267 5425 24276
rect 5481 24267 5506 24323
rect 5562 24267 5587 24323
rect 5643 24267 5668 24323
rect 5724 24267 5749 24323
rect 5805 24267 5830 24323
rect 5886 24267 5911 24323
rect 5967 24267 5992 24323
rect 6048 24267 6073 24323
rect 6129 24267 6154 24323
rect 6210 24267 6235 24323
rect 6291 24267 6316 24323
rect 6372 24267 6397 24323
rect 6453 24267 6478 24323
rect 6534 24267 6559 24323
rect 6615 24267 6640 24323
rect 6696 24267 6721 24323
rect 6777 24267 6802 24323
rect 6858 24267 6883 24323
rect 6939 24267 6964 24323
rect 7020 24267 7045 24323
rect 7101 24267 7126 24323
rect 7182 24267 7207 24323
rect 7263 24267 7288 24323
rect 7344 24267 7369 24323
rect 7425 24267 7450 24323
rect 7506 24267 7531 24323
rect 7587 24267 7612 24323
rect 7668 24267 7693 24323
rect 7749 24267 7774 24323
rect 7830 24267 7855 24323
rect 7911 24267 7936 24323
rect 7992 24267 8017 24323
rect 8073 24267 8098 24323
rect 8154 24267 8179 24323
rect 8235 24267 8260 24323
rect 8316 24267 8341 24323
rect 8397 24267 8422 24323
rect 8478 24267 8503 24323
rect 8559 24267 8584 24323
rect 8640 24267 8665 24323
rect 8721 24267 8746 24323
rect 8802 24267 8827 24323
rect 8883 24267 8908 24323
rect 8964 24267 8989 24323
rect 9045 24267 9070 24323
rect 9126 24267 9151 24323
rect 9207 24267 9232 24323
rect 9288 24267 9313 24323
rect 9369 24267 9394 24323
rect 9450 24267 9475 24323
rect 9531 24267 9556 24323
rect 9612 24267 9637 24323
rect 9693 24267 9718 24323
rect 9774 24267 9799 24323
rect 9855 24267 9880 24323
rect 9936 24267 9961 24323
rect 10017 24267 10042 24323
rect 10098 24267 10123 24323
rect 10179 24267 10204 24323
rect 10260 24267 10285 24323
rect 10341 24267 10366 24323
rect 10422 24267 10447 24323
rect 10503 24267 10528 24323
rect 10584 24267 10609 24323
rect 10665 24267 10690 24323
rect 10746 24267 10771 24323
rect 10827 24267 10852 24323
rect 10908 24267 10933 24323
rect 10989 24267 11014 24323
rect 11070 24267 11095 24323
rect 11151 24267 11176 24323
rect 11232 24267 11257 24323
rect 11313 24267 11338 24323
rect 11394 24267 11419 24323
rect 11475 24267 11500 24323
rect 2472 24243 11500 24267
rect 2472 24220 5425 24243
rect 1852 24194 5425 24220
rect 1852 24138 2170 24194
rect 2226 24138 2252 24194
rect 2308 24138 2334 24194
rect 2390 24138 2416 24194
rect 2472 24187 5425 24194
rect 5481 24187 5506 24243
rect 5562 24187 5587 24243
rect 5643 24187 5668 24243
rect 5724 24187 5749 24243
rect 5805 24187 5830 24243
rect 5886 24187 5911 24243
rect 5967 24187 5992 24243
rect 6048 24187 6073 24243
rect 6129 24187 6154 24243
rect 6210 24187 6235 24243
rect 6291 24187 6316 24243
rect 6372 24187 6397 24243
rect 6453 24187 6478 24243
rect 6534 24187 6559 24243
rect 6615 24187 6640 24243
rect 6696 24187 6721 24243
rect 6777 24187 6802 24243
rect 6858 24187 6883 24243
rect 6939 24187 6964 24243
rect 7020 24187 7045 24243
rect 7101 24187 7126 24243
rect 7182 24187 7207 24243
rect 7263 24187 7288 24243
rect 7344 24187 7369 24243
rect 7425 24187 7450 24243
rect 7506 24187 7531 24243
rect 7587 24187 7612 24243
rect 7668 24187 7693 24243
rect 7749 24187 7774 24243
rect 7830 24187 7855 24243
rect 7911 24187 7936 24243
rect 7992 24187 8017 24243
rect 8073 24187 8098 24243
rect 8154 24187 8179 24243
rect 8235 24187 8260 24243
rect 8316 24187 8341 24243
rect 8397 24187 8422 24243
rect 8478 24187 8503 24243
rect 8559 24187 8584 24243
rect 8640 24187 8665 24243
rect 8721 24187 8746 24243
rect 8802 24187 8827 24243
rect 8883 24187 8908 24243
rect 8964 24187 8989 24243
rect 9045 24187 9070 24243
rect 9126 24187 9151 24243
rect 9207 24187 9232 24243
rect 9288 24187 9313 24243
rect 9369 24187 9394 24243
rect 9450 24187 9475 24243
rect 9531 24187 9556 24243
rect 9612 24187 9637 24243
rect 9693 24187 9718 24243
rect 9774 24187 9799 24243
rect 9855 24187 9880 24243
rect 9936 24187 9961 24243
rect 10017 24187 10042 24243
rect 10098 24187 10123 24243
rect 10179 24187 10204 24243
rect 10260 24187 10285 24243
rect 10341 24187 10366 24243
rect 10422 24187 10447 24243
rect 10503 24187 10528 24243
rect 10584 24187 10609 24243
rect 10665 24187 10690 24243
rect 10746 24187 10771 24243
rect 10827 24187 10852 24243
rect 10908 24187 10933 24243
rect 10989 24187 11014 24243
rect 11070 24187 11095 24243
rect 11151 24187 11176 24243
rect 11232 24187 11257 24243
rect 11313 24187 11338 24243
rect 11394 24187 11419 24243
rect 11475 24187 11500 24243
rect 2472 24163 11500 24187
rect 2472 24138 5425 24163
rect 1852 24112 5425 24138
rect 1852 24056 2170 24112
rect 2226 24056 2252 24112
rect 2308 24056 2334 24112
rect 2390 24056 2416 24112
rect 2472 24107 5425 24112
rect 5481 24107 5506 24163
rect 5562 24107 5587 24163
rect 5643 24107 5668 24163
rect 5724 24107 5749 24163
rect 5805 24107 5830 24163
rect 5886 24107 5911 24163
rect 5967 24107 5992 24163
rect 6048 24107 6073 24163
rect 6129 24107 6154 24163
rect 6210 24107 6235 24163
rect 6291 24107 6316 24163
rect 6372 24107 6397 24163
rect 6453 24107 6478 24163
rect 6534 24107 6559 24163
rect 6615 24107 6640 24163
rect 6696 24107 6721 24163
rect 6777 24107 6802 24163
rect 6858 24107 6883 24163
rect 6939 24107 6964 24163
rect 7020 24107 7045 24163
rect 7101 24107 7126 24163
rect 7182 24107 7207 24163
rect 7263 24107 7288 24163
rect 7344 24107 7369 24163
rect 7425 24107 7450 24163
rect 7506 24107 7531 24163
rect 7587 24107 7612 24163
rect 7668 24107 7693 24163
rect 7749 24107 7774 24163
rect 7830 24107 7855 24163
rect 7911 24107 7936 24163
rect 7992 24107 8017 24163
rect 8073 24107 8098 24163
rect 8154 24107 8179 24163
rect 8235 24107 8260 24163
rect 8316 24107 8341 24163
rect 8397 24107 8422 24163
rect 8478 24107 8503 24163
rect 8559 24107 8584 24163
rect 8640 24107 8665 24163
rect 8721 24107 8746 24163
rect 8802 24107 8827 24163
rect 8883 24107 8908 24163
rect 8964 24107 8989 24163
rect 9045 24107 9070 24163
rect 9126 24107 9151 24163
rect 9207 24107 9232 24163
rect 9288 24107 9313 24163
rect 9369 24107 9394 24163
rect 9450 24107 9475 24163
rect 9531 24107 9556 24163
rect 9612 24107 9637 24163
rect 9693 24107 9718 24163
rect 9774 24107 9799 24163
rect 9855 24107 9880 24163
rect 9936 24107 9961 24163
rect 10017 24107 10042 24163
rect 10098 24107 10123 24163
rect 10179 24107 10204 24163
rect 10260 24107 10285 24163
rect 10341 24107 10366 24163
rect 10422 24107 10447 24163
rect 10503 24107 10528 24163
rect 10584 24107 10609 24163
rect 10665 24107 10690 24163
rect 10746 24107 10771 24163
rect 10827 24107 10852 24163
rect 10908 24107 10933 24163
rect 10989 24107 11014 24163
rect 11070 24107 11095 24163
rect 11151 24107 11176 24163
rect 11232 24107 11257 24163
rect 11313 24107 11338 24163
rect 11394 24107 11419 24163
rect 11475 24107 11500 24163
rect 2472 24083 11500 24107
rect 2472 24056 5425 24083
rect 1852 24030 5425 24056
rect 1852 23974 2170 24030
rect 2226 23974 2252 24030
rect 2308 23974 2334 24030
rect 2390 23974 2416 24030
rect 2472 24027 5425 24030
rect 5481 24027 5506 24083
rect 5562 24027 5587 24083
rect 5643 24027 5668 24083
rect 5724 24027 5749 24083
rect 5805 24027 5830 24083
rect 5886 24027 5911 24083
rect 5967 24027 5992 24083
rect 6048 24027 6073 24083
rect 6129 24027 6154 24083
rect 6210 24027 6235 24083
rect 6291 24027 6316 24083
rect 6372 24027 6397 24083
rect 6453 24027 6478 24083
rect 6534 24027 6559 24083
rect 6615 24027 6640 24083
rect 6696 24027 6721 24083
rect 6777 24027 6802 24083
rect 6858 24027 6883 24083
rect 6939 24027 6964 24083
rect 7020 24027 7045 24083
rect 7101 24027 7126 24083
rect 7182 24027 7207 24083
rect 7263 24027 7288 24083
rect 7344 24027 7369 24083
rect 7425 24027 7450 24083
rect 7506 24027 7531 24083
rect 7587 24027 7612 24083
rect 7668 24027 7693 24083
rect 7749 24027 7774 24083
rect 7830 24027 7855 24083
rect 7911 24027 7936 24083
rect 7992 24027 8017 24083
rect 8073 24027 8098 24083
rect 8154 24027 8179 24083
rect 8235 24027 8260 24083
rect 8316 24027 8341 24083
rect 8397 24027 8422 24083
rect 8478 24027 8503 24083
rect 8559 24027 8584 24083
rect 8640 24027 8665 24083
rect 8721 24027 8746 24083
rect 8802 24027 8827 24083
rect 8883 24027 8908 24083
rect 8964 24027 8989 24083
rect 9045 24027 9070 24083
rect 9126 24027 9151 24083
rect 9207 24027 9232 24083
rect 9288 24027 9313 24083
rect 9369 24027 9394 24083
rect 9450 24027 9475 24083
rect 9531 24027 9556 24083
rect 9612 24027 9637 24083
rect 9693 24027 9718 24083
rect 9774 24027 9799 24083
rect 9855 24027 9880 24083
rect 9936 24027 9961 24083
rect 10017 24027 10042 24083
rect 10098 24027 10123 24083
rect 10179 24027 10204 24083
rect 10260 24027 10285 24083
rect 10341 24027 10366 24083
rect 10422 24027 10447 24083
rect 10503 24027 10528 24083
rect 10584 24027 10609 24083
rect 10665 24027 10690 24083
rect 10746 24027 10771 24083
rect 10827 24027 10852 24083
rect 10908 24027 10933 24083
rect 10989 24027 11014 24083
rect 11070 24027 11095 24083
rect 11151 24027 11176 24083
rect 11232 24027 11257 24083
rect 11313 24027 11338 24083
rect 11394 24027 11419 24083
rect 11475 24027 11500 24083
rect 2472 24003 11500 24027
rect 2472 23974 5425 24003
rect 1852 23948 5425 23974
rect 1852 23892 2170 23948
rect 2226 23892 2252 23948
rect 2308 23892 2334 23948
rect 2390 23892 2416 23948
rect 2472 23947 5425 23948
rect 5481 23947 5506 24003
rect 5562 23947 5587 24003
rect 5643 23947 5668 24003
rect 5724 23947 5749 24003
rect 5805 23947 5830 24003
rect 5886 23947 5911 24003
rect 5967 23947 5992 24003
rect 6048 23947 6073 24003
rect 6129 23947 6154 24003
rect 6210 23947 6235 24003
rect 6291 23947 6316 24003
rect 6372 23947 6397 24003
rect 6453 23947 6478 24003
rect 6534 23947 6559 24003
rect 6615 23947 6640 24003
rect 6696 23947 6721 24003
rect 6777 23947 6802 24003
rect 6858 23947 6883 24003
rect 6939 23947 6964 24003
rect 7020 23947 7045 24003
rect 7101 23947 7126 24003
rect 7182 23947 7207 24003
rect 7263 23947 7288 24003
rect 7344 23947 7369 24003
rect 7425 23947 7450 24003
rect 7506 23947 7531 24003
rect 7587 23947 7612 24003
rect 7668 23947 7693 24003
rect 7749 23947 7774 24003
rect 7830 23947 7855 24003
rect 7911 23947 7936 24003
rect 7992 23947 8017 24003
rect 8073 23947 8098 24003
rect 8154 23947 8179 24003
rect 8235 23947 8260 24003
rect 8316 23947 8341 24003
rect 8397 23947 8422 24003
rect 8478 23947 8503 24003
rect 8559 23947 8584 24003
rect 8640 23947 8665 24003
rect 8721 23947 8746 24003
rect 8802 23947 8827 24003
rect 8883 23947 8908 24003
rect 8964 23947 8989 24003
rect 9045 23947 9070 24003
rect 9126 23947 9151 24003
rect 9207 23947 9232 24003
rect 9288 23947 9313 24003
rect 9369 23947 9394 24003
rect 9450 23947 9475 24003
rect 9531 23947 9556 24003
rect 9612 23947 9637 24003
rect 9693 23947 9718 24003
rect 9774 23947 9799 24003
rect 9855 23947 9880 24003
rect 9936 23947 9961 24003
rect 10017 23947 10042 24003
rect 10098 23947 10123 24003
rect 10179 23947 10204 24003
rect 10260 23947 10285 24003
rect 10341 23947 10366 24003
rect 10422 23947 10447 24003
rect 10503 23947 10528 24003
rect 10584 23947 10609 24003
rect 10665 23947 10690 24003
rect 10746 23947 10771 24003
rect 10827 23947 10852 24003
rect 10908 23947 10933 24003
rect 10989 23947 11014 24003
rect 11070 23947 11095 24003
rect 11151 23947 11176 24003
rect 11232 23947 11257 24003
rect 11313 23947 11338 24003
rect 11394 23947 11419 24003
rect 11475 23947 11500 24003
rect 2472 23923 11500 23947
rect 2472 23892 5425 23923
rect 1852 23867 5425 23892
rect 5481 23867 5506 23923
rect 5562 23867 5587 23923
rect 5643 23867 5668 23923
rect 5724 23867 5749 23923
rect 5805 23867 5830 23923
rect 5886 23867 5911 23923
rect 5967 23867 5992 23923
rect 6048 23867 6073 23923
rect 6129 23867 6154 23923
rect 6210 23867 6235 23923
rect 6291 23867 6316 23923
rect 6372 23867 6397 23923
rect 6453 23867 6478 23923
rect 6534 23867 6559 23923
rect 6615 23867 6640 23923
rect 6696 23867 6721 23923
rect 6777 23867 6802 23923
rect 6858 23867 6883 23923
rect 6939 23867 6964 23923
rect 7020 23867 7045 23923
rect 7101 23867 7126 23923
rect 7182 23867 7207 23923
rect 7263 23867 7288 23923
rect 7344 23867 7369 23923
rect 7425 23867 7450 23923
rect 7506 23867 7531 23923
rect 7587 23867 7612 23923
rect 7668 23867 7693 23923
rect 7749 23867 7774 23923
rect 7830 23867 7855 23923
rect 7911 23867 7936 23923
rect 7992 23867 8017 23923
rect 8073 23867 8098 23923
rect 8154 23867 8179 23923
rect 8235 23867 8260 23923
rect 8316 23867 8341 23923
rect 8397 23867 8422 23923
rect 8478 23867 8503 23923
rect 8559 23867 8584 23923
rect 8640 23867 8665 23923
rect 8721 23867 8746 23923
rect 8802 23867 8827 23923
rect 8883 23867 8908 23923
rect 8964 23867 8989 23923
rect 9045 23867 9070 23923
rect 9126 23867 9151 23923
rect 9207 23867 9232 23923
rect 9288 23867 9313 23923
rect 9369 23867 9394 23923
rect 9450 23867 9475 23923
rect 9531 23867 9556 23923
rect 9612 23867 9637 23923
rect 9693 23867 9718 23923
rect 9774 23867 9799 23923
rect 9855 23867 9880 23923
rect 9936 23867 9961 23923
rect 10017 23867 10042 23923
rect 10098 23867 10123 23923
rect 10179 23867 10204 23923
rect 10260 23867 10285 23923
rect 10341 23867 10366 23923
rect 10422 23867 10447 23923
rect 10503 23867 10528 23923
rect 10584 23867 10609 23923
rect 10665 23867 10690 23923
rect 10746 23867 10771 23923
rect 10827 23867 10852 23923
rect 10908 23867 10933 23923
rect 10989 23867 11014 23923
rect 11070 23867 11095 23923
rect 11151 23867 11176 23923
rect 11232 23867 11257 23923
rect 11313 23867 11338 23923
rect 11394 23867 11419 23923
rect 11475 23867 11500 23923
rect 1852 23866 11500 23867
rect 1852 23810 2170 23866
rect 2226 23810 2252 23866
rect 2308 23810 2334 23866
rect 2390 23810 2416 23866
rect 2472 23843 11500 23866
rect 2472 23810 5425 23843
rect 1852 23787 5425 23810
rect 5481 23787 5506 23843
rect 5562 23787 5587 23843
rect 5643 23787 5668 23843
rect 5724 23787 5749 23843
rect 5805 23787 5830 23843
rect 5886 23787 5911 23843
rect 5967 23787 5992 23843
rect 6048 23787 6073 23843
rect 6129 23787 6154 23843
rect 6210 23787 6235 23843
rect 6291 23787 6316 23843
rect 6372 23787 6397 23843
rect 6453 23787 6478 23843
rect 6534 23787 6559 23843
rect 6615 23787 6640 23843
rect 6696 23787 6721 23843
rect 6777 23787 6802 23843
rect 6858 23787 6883 23843
rect 6939 23787 6964 23843
rect 7020 23787 7045 23843
rect 7101 23787 7126 23843
rect 7182 23787 7207 23843
rect 7263 23787 7288 23843
rect 7344 23787 7369 23843
rect 7425 23787 7450 23843
rect 7506 23787 7531 23843
rect 7587 23787 7612 23843
rect 7668 23787 7693 23843
rect 7749 23787 7774 23843
rect 7830 23787 7855 23843
rect 7911 23787 7936 23843
rect 7992 23787 8017 23843
rect 8073 23787 8098 23843
rect 8154 23787 8179 23843
rect 8235 23787 8260 23843
rect 8316 23787 8341 23843
rect 8397 23787 8422 23843
rect 8478 23787 8503 23843
rect 8559 23787 8584 23843
rect 8640 23787 8665 23843
rect 8721 23787 8746 23843
rect 8802 23787 8827 23843
rect 8883 23787 8908 23843
rect 8964 23787 8989 23843
rect 9045 23787 9070 23843
rect 9126 23787 9151 23843
rect 9207 23787 9232 23843
rect 9288 23787 9313 23843
rect 9369 23787 9394 23843
rect 9450 23787 9475 23843
rect 9531 23787 9556 23843
rect 9612 23787 9637 23843
rect 9693 23787 9718 23843
rect 9774 23787 9799 23843
rect 9855 23787 9880 23843
rect 9936 23787 9961 23843
rect 10017 23787 10042 23843
rect 10098 23787 10123 23843
rect 10179 23787 10204 23843
rect 10260 23787 10285 23843
rect 10341 23787 10366 23843
rect 10422 23787 10447 23843
rect 10503 23787 10528 23843
rect 10584 23787 10609 23843
rect 10665 23787 10690 23843
rect 10746 23787 10771 23843
rect 10827 23787 10852 23843
rect 10908 23787 10933 23843
rect 10989 23787 11014 23843
rect 11070 23787 11095 23843
rect 11151 23787 11176 23843
rect 11232 23787 11257 23843
rect 11313 23787 11338 23843
rect 11394 23787 11419 23843
rect 11475 23787 11500 23843
rect 1852 23784 11500 23787
rect 1852 23728 2170 23784
rect 2226 23728 2252 23784
rect 2308 23728 2334 23784
rect 2390 23728 2416 23784
rect 2472 23763 11500 23784
rect 2472 23728 5425 23763
rect 1852 23707 5425 23728
rect 5481 23707 5506 23763
rect 5562 23707 5587 23763
rect 5643 23707 5668 23763
rect 5724 23707 5749 23763
rect 5805 23707 5830 23763
rect 5886 23707 5911 23763
rect 5967 23707 5992 23763
rect 6048 23707 6073 23763
rect 6129 23707 6154 23763
rect 6210 23707 6235 23763
rect 6291 23707 6316 23763
rect 6372 23707 6397 23763
rect 6453 23707 6478 23763
rect 6534 23707 6559 23763
rect 6615 23707 6640 23763
rect 6696 23707 6721 23763
rect 6777 23707 6802 23763
rect 6858 23707 6883 23763
rect 6939 23707 6964 23763
rect 7020 23707 7045 23763
rect 7101 23707 7126 23763
rect 7182 23707 7207 23763
rect 7263 23707 7288 23763
rect 7344 23707 7369 23763
rect 7425 23707 7450 23763
rect 7506 23707 7531 23763
rect 7587 23707 7612 23763
rect 7668 23707 7693 23763
rect 7749 23707 7774 23763
rect 7830 23707 7855 23763
rect 7911 23707 7936 23763
rect 7992 23707 8017 23763
rect 8073 23707 8098 23763
rect 8154 23707 8179 23763
rect 8235 23707 8260 23763
rect 8316 23707 8341 23763
rect 8397 23707 8422 23763
rect 8478 23707 8503 23763
rect 8559 23707 8584 23763
rect 8640 23707 8665 23763
rect 8721 23707 8746 23763
rect 8802 23707 8827 23763
rect 8883 23707 8908 23763
rect 8964 23707 8989 23763
rect 9045 23707 9070 23763
rect 9126 23707 9151 23763
rect 9207 23707 9232 23763
rect 9288 23707 9313 23763
rect 9369 23707 9394 23763
rect 9450 23707 9475 23763
rect 9531 23707 9556 23763
rect 9612 23707 9637 23763
rect 9693 23707 9718 23763
rect 9774 23707 9799 23763
rect 9855 23707 9880 23763
rect 9936 23707 9961 23763
rect 10017 23707 10042 23763
rect 10098 23707 10123 23763
rect 10179 23707 10204 23763
rect 10260 23707 10285 23763
rect 10341 23707 10366 23763
rect 10422 23707 10447 23763
rect 10503 23707 10528 23763
rect 10584 23707 10609 23763
rect 10665 23707 10690 23763
rect 10746 23707 10771 23763
rect 10827 23707 10852 23763
rect 10908 23707 10933 23763
rect 10989 23707 11014 23763
rect 11070 23707 11095 23763
rect 11151 23707 11176 23763
rect 11232 23707 11257 23763
rect 11313 23707 11338 23763
rect 11394 23707 11419 23763
rect 11475 23707 11500 23763
rect 1852 23702 11500 23707
rect 1852 23646 2170 23702
rect 2226 23646 2252 23702
rect 2308 23646 2334 23702
rect 2390 23646 2416 23702
rect 2472 23683 11500 23702
rect 2472 23646 5425 23683
rect 1852 23627 5425 23646
rect 5481 23627 5506 23683
rect 5562 23627 5587 23683
rect 5643 23627 5668 23683
rect 5724 23627 5749 23683
rect 5805 23627 5830 23683
rect 5886 23627 5911 23683
rect 5967 23627 5992 23683
rect 6048 23627 6073 23683
rect 6129 23627 6154 23683
rect 6210 23627 6235 23683
rect 6291 23627 6316 23683
rect 6372 23627 6397 23683
rect 6453 23627 6478 23683
rect 6534 23627 6559 23683
rect 6615 23627 6640 23683
rect 6696 23627 6721 23683
rect 6777 23627 6802 23683
rect 6858 23627 6883 23683
rect 6939 23627 6964 23683
rect 7020 23627 7045 23683
rect 7101 23627 7126 23683
rect 7182 23627 7207 23683
rect 7263 23627 7288 23683
rect 7344 23627 7369 23683
rect 7425 23627 7450 23683
rect 7506 23627 7531 23683
rect 7587 23627 7612 23683
rect 7668 23627 7693 23683
rect 7749 23627 7774 23683
rect 7830 23627 7855 23683
rect 7911 23627 7936 23683
rect 7992 23627 8017 23683
rect 8073 23627 8098 23683
rect 8154 23627 8179 23683
rect 8235 23627 8260 23683
rect 8316 23627 8341 23683
rect 8397 23627 8422 23683
rect 8478 23627 8503 23683
rect 8559 23627 8584 23683
rect 8640 23627 8665 23683
rect 8721 23627 8746 23683
rect 8802 23627 8827 23683
rect 8883 23627 8908 23683
rect 8964 23627 8989 23683
rect 9045 23627 9070 23683
rect 9126 23627 9151 23683
rect 9207 23627 9232 23683
rect 9288 23627 9313 23683
rect 9369 23627 9394 23683
rect 9450 23627 9475 23683
rect 9531 23627 9556 23683
rect 9612 23627 9637 23683
rect 9693 23627 9718 23683
rect 9774 23627 9799 23683
rect 9855 23627 9880 23683
rect 9936 23627 9961 23683
rect 10017 23627 10042 23683
rect 10098 23627 10123 23683
rect 10179 23627 10204 23683
rect 10260 23627 10285 23683
rect 10341 23627 10366 23683
rect 10422 23627 10447 23683
rect 10503 23627 10528 23683
rect 10584 23627 10609 23683
rect 10665 23627 10690 23683
rect 10746 23627 10771 23683
rect 10827 23627 10852 23683
rect 10908 23627 10933 23683
rect 10989 23627 11014 23683
rect 11070 23627 11095 23683
rect 11151 23627 11176 23683
rect 11232 23627 11257 23683
rect 11313 23627 11338 23683
rect 11394 23627 11419 23683
rect 11475 23627 11500 23683
rect 1852 23620 11500 23627
rect 1852 23564 2170 23620
rect 2226 23564 2252 23620
rect 2308 23564 2334 23620
rect 2390 23564 2416 23620
rect 2472 23603 11500 23620
rect 2472 23564 5425 23603
rect 1852 23547 5425 23564
rect 5481 23547 5506 23603
rect 5562 23547 5587 23603
rect 5643 23547 5668 23603
rect 5724 23547 5749 23603
rect 5805 23547 5830 23603
rect 5886 23547 5911 23603
rect 5967 23547 5992 23603
rect 6048 23547 6073 23603
rect 6129 23547 6154 23603
rect 6210 23547 6235 23603
rect 6291 23547 6316 23603
rect 6372 23547 6397 23603
rect 6453 23547 6478 23603
rect 6534 23547 6559 23603
rect 6615 23547 6640 23603
rect 6696 23547 6721 23603
rect 6777 23547 6802 23603
rect 6858 23547 6883 23603
rect 6939 23547 6964 23603
rect 7020 23547 7045 23603
rect 7101 23547 7126 23603
rect 7182 23547 7207 23603
rect 7263 23547 7288 23603
rect 7344 23547 7369 23603
rect 7425 23547 7450 23603
rect 7506 23547 7531 23603
rect 7587 23547 7612 23603
rect 7668 23547 7693 23603
rect 7749 23547 7774 23603
rect 7830 23547 7855 23603
rect 7911 23547 7936 23603
rect 7992 23547 8017 23603
rect 8073 23547 8098 23603
rect 8154 23547 8179 23603
rect 8235 23547 8260 23603
rect 8316 23547 8341 23603
rect 8397 23547 8422 23603
rect 8478 23547 8503 23603
rect 8559 23547 8584 23603
rect 8640 23547 8665 23603
rect 8721 23547 8746 23603
rect 8802 23547 8827 23603
rect 8883 23547 8908 23603
rect 8964 23547 8989 23603
rect 9045 23547 9070 23603
rect 9126 23547 9151 23603
rect 9207 23547 9232 23603
rect 9288 23547 9313 23603
rect 9369 23547 9394 23603
rect 9450 23547 9475 23603
rect 9531 23547 9556 23603
rect 9612 23547 9637 23603
rect 9693 23547 9718 23603
rect 9774 23547 9799 23603
rect 9855 23547 9880 23603
rect 9936 23547 9961 23603
rect 10017 23547 10042 23603
rect 10098 23547 10123 23603
rect 10179 23547 10204 23603
rect 10260 23547 10285 23603
rect 10341 23547 10366 23603
rect 10422 23547 10447 23603
rect 10503 23547 10528 23603
rect 10584 23547 10609 23603
rect 10665 23547 10690 23603
rect 10746 23547 10771 23603
rect 10827 23547 10852 23603
rect 10908 23547 10933 23603
rect 10989 23547 11014 23603
rect 11070 23547 11095 23603
rect 11151 23547 11176 23603
rect 11232 23547 11257 23603
rect 11313 23547 11338 23603
rect 11394 23547 11419 23603
rect 11475 23547 11500 23603
rect 1852 23538 11500 23547
rect 1852 23482 2170 23538
rect 2226 23482 2252 23538
rect 2308 23482 2334 23538
rect 2390 23482 2416 23538
rect 2472 23523 11500 23538
rect 2472 23482 5425 23523
rect 1852 23467 5425 23482
rect 5481 23467 5506 23523
rect 5562 23467 5587 23523
rect 5643 23467 5668 23523
rect 5724 23467 5749 23523
rect 5805 23467 5830 23523
rect 5886 23467 5911 23523
rect 5967 23467 5992 23523
rect 6048 23467 6073 23523
rect 6129 23467 6154 23523
rect 6210 23467 6235 23523
rect 6291 23467 6316 23523
rect 6372 23467 6397 23523
rect 6453 23467 6478 23523
rect 6534 23467 6559 23523
rect 6615 23467 6640 23523
rect 6696 23467 6721 23523
rect 6777 23467 6802 23523
rect 6858 23467 6883 23523
rect 6939 23467 6964 23523
rect 7020 23467 7045 23523
rect 7101 23467 7126 23523
rect 7182 23467 7207 23523
rect 7263 23467 7288 23523
rect 7344 23467 7369 23523
rect 7425 23467 7450 23523
rect 7506 23467 7531 23523
rect 7587 23467 7612 23523
rect 7668 23467 7693 23523
rect 7749 23467 7774 23523
rect 7830 23467 7855 23523
rect 7911 23467 7936 23523
rect 7992 23467 8017 23523
rect 8073 23467 8098 23523
rect 8154 23467 8179 23523
rect 8235 23467 8260 23523
rect 8316 23467 8341 23523
rect 8397 23467 8422 23523
rect 8478 23467 8503 23523
rect 8559 23467 8584 23523
rect 8640 23467 8665 23523
rect 8721 23467 8746 23523
rect 8802 23467 8827 23523
rect 8883 23467 8908 23523
rect 8964 23467 8989 23523
rect 9045 23467 9070 23523
rect 9126 23467 9151 23523
rect 9207 23467 9232 23523
rect 9288 23467 9313 23523
rect 9369 23467 9394 23523
rect 9450 23467 9475 23523
rect 9531 23467 9556 23523
rect 9612 23467 9637 23523
rect 9693 23467 9718 23523
rect 9774 23467 9799 23523
rect 9855 23467 9880 23523
rect 9936 23467 9961 23523
rect 10017 23467 10042 23523
rect 10098 23467 10123 23523
rect 10179 23467 10204 23523
rect 10260 23467 10285 23523
rect 10341 23467 10366 23523
rect 10422 23467 10447 23523
rect 10503 23467 10528 23523
rect 10584 23467 10609 23523
rect 10665 23467 10690 23523
rect 10746 23467 10771 23523
rect 10827 23467 10852 23523
rect 10908 23467 10933 23523
rect 10989 23467 11014 23523
rect 11070 23467 11095 23523
rect 11151 23467 11176 23523
rect 11232 23467 11257 23523
rect 11313 23467 11338 23523
rect 11394 23467 11419 23523
rect 11475 23467 11500 23523
rect 1852 23456 11500 23467
rect 1852 23400 2170 23456
rect 2226 23400 2252 23456
rect 2308 23400 2334 23456
rect 2390 23400 2416 23456
rect 2472 23443 11500 23456
rect 2472 23400 5425 23443
rect 1852 23387 5425 23400
rect 5481 23387 5506 23443
rect 5562 23387 5587 23443
rect 5643 23387 5668 23443
rect 5724 23387 5749 23443
rect 5805 23387 5830 23443
rect 5886 23387 5911 23443
rect 5967 23387 5992 23443
rect 6048 23387 6073 23443
rect 6129 23387 6154 23443
rect 6210 23387 6235 23443
rect 6291 23387 6316 23443
rect 6372 23387 6397 23443
rect 6453 23387 6478 23443
rect 6534 23387 6559 23443
rect 6615 23387 6640 23443
rect 6696 23387 6721 23443
rect 6777 23387 6802 23443
rect 6858 23387 6883 23443
rect 6939 23387 6964 23443
rect 7020 23387 7045 23443
rect 7101 23387 7126 23443
rect 7182 23387 7207 23443
rect 7263 23387 7288 23443
rect 7344 23387 7369 23443
rect 7425 23387 7450 23443
rect 7506 23387 7531 23443
rect 7587 23387 7612 23443
rect 7668 23387 7693 23443
rect 7749 23387 7774 23443
rect 7830 23387 7855 23443
rect 7911 23387 7936 23443
rect 7992 23387 8017 23443
rect 8073 23387 8098 23443
rect 8154 23387 8179 23443
rect 8235 23387 8260 23443
rect 8316 23387 8341 23443
rect 8397 23387 8422 23443
rect 8478 23387 8503 23443
rect 8559 23387 8584 23443
rect 8640 23387 8665 23443
rect 8721 23387 8746 23443
rect 8802 23387 8827 23443
rect 8883 23387 8908 23443
rect 8964 23387 8989 23443
rect 9045 23387 9070 23443
rect 9126 23387 9151 23443
rect 9207 23387 9232 23443
rect 9288 23387 9313 23443
rect 9369 23387 9394 23443
rect 9450 23387 9475 23443
rect 9531 23387 9556 23443
rect 9612 23387 9637 23443
rect 9693 23387 9718 23443
rect 9774 23387 9799 23443
rect 9855 23387 9880 23443
rect 9936 23387 9961 23443
rect 10017 23387 10042 23443
rect 10098 23387 10123 23443
rect 10179 23387 10204 23443
rect 10260 23387 10285 23443
rect 10341 23387 10366 23443
rect 10422 23387 10447 23443
rect 10503 23387 10528 23443
rect 10584 23387 10609 23443
rect 10665 23387 10690 23443
rect 10746 23387 10771 23443
rect 10827 23387 10852 23443
rect 10908 23387 10933 23443
rect 10989 23387 11014 23443
rect 11070 23387 11095 23443
rect 11151 23387 11176 23443
rect 11232 23387 11257 23443
rect 11313 23387 11338 23443
rect 11394 23387 11419 23443
rect 11475 23387 11500 23443
rect 1852 23374 11500 23387
rect 1852 23318 2170 23374
rect 2226 23318 2252 23374
rect 2308 23318 2334 23374
rect 2390 23318 2416 23374
rect 2472 23363 11500 23374
rect 2472 23318 5425 23363
rect 1852 23307 5425 23318
rect 5481 23307 5506 23363
rect 5562 23307 5587 23363
rect 5643 23307 5668 23363
rect 5724 23307 5749 23363
rect 5805 23307 5830 23363
rect 5886 23307 5911 23363
rect 5967 23307 5992 23363
rect 6048 23307 6073 23363
rect 6129 23307 6154 23363
rect 6210 23307 6235 23363
rect 6291 23307 6316 23363
rect 6372 23307 6397 23363
rect 6453 23307 6478 23363
rect 6534 23307 6559 23363
rect 6615 23307 6640 23363
rect 6696 23307 6721 23363
rect 6777 23307 6802 23363
rect 6858 23307 6883 23363
rect 6939 23307 6964 23363
rect 7020 23307 7045 23363
rect 7101 23307 7126 23363
rect 7182 23307 7207 23363
rect 7263 23307 7288 23363
rect 7344 23307 7369 23363
rect 7425 23307 7450 23363
rect 7506 23307 7531 23363
rect 7587 23307 7612 23363
rect 7668 23307 7693 23363
rect 7749 23307 7774 23363
rect 7830 23307 7855 23363
rect 7911 23307 7936 23363
rect 7992 23307 8017 23363
rect 8073 23307 8098 23363
rect 8154 23307 8179 23363
rect 8235 23307 8260 23363
rect 8316 23307 8341 23363
rect 8397 23307 8422 23363
rect 8478 23307 8503 23363
rect 8559 23307 8584 23363
rect 8640 23307 8665 23363
rect 8721 23307 8746 23363
rect 8802 23307 8827 23363
rect 8883 23307 8908 23363
rect 8964 23307 8989 23363
rect 9045 23307 9070 23363
rect 9126 23307 9151 23363
rect 9207 23307 9232 23363
rect 9288 23307 9313 23363
rect 9369 23307 9394 23363
rect 9450 23307 9475 23363
rect 9531 23307 9556 23363
rect 9612 23307 9637 23363
rect 9693 23307 9718 23363
rect 9774 23307 9799 23363
rect 9855 23307 9880 23363
rect 9936 23307 9961 23363
rect 10017 23307 10042 23363
rect 10098 23307 10123 23363
rect 10179 23307 10204 23363
rect 10260 23307 10285 23363
rect 10341 23307 10366 23363
rect 10422 23307 10447 23363
rect 10503 23307 10528 23363
rect 10584 23307 10609 23363
rect 10665 23307 10690 23363
rect 10746 23307 10771 23363
rect 10827 23307 10852 23363
rect 10908 23307 10933 23363
rect 10989 23307 11014 23363
rect 11070 23307 11095 23363
rect 11151 23307 11176 23363
rect 11232 23307 11257 23363
rect 11313 23307 11338 23363
rect 11394 23307 11419 23363
rect 11475 23307 11500 23363
rect 1852 23292 11500 23307
rect 1852 23236 2170 23292
rect 2226 23236 2252 23292
rect 2308 23236 2334 23292
rect 2390 23236 2416 23292
rect 2472 23283 11500 23292
rect 2472 23236 5425 23283
rect 1852 23227 5425 23236
rect 5481 23227 5506 23283
rect 5562 23227 5587 23283
rect 5643 23227 5668 23283
rect 5724 23227 5749 23283
rect 5805 23227 5830 23283
rect 5886 23227 5911 23283
rect 5967 23227 5992 23283
rect 6048 23227 6073 23283
rect 6129 23227 6154 23283
rect 6210 23227 6235 23283
rect 6291 23227 6316 23283
rect 6372 23227 6397 23283
rect 6453 23227 6478 23283
rect 6534 23227 6559 23283
rect 6615 23227 6640 23283
rect 6696 23227 6721 23283
rect 6777 23227 6802 23283
rect 6858 23227 6883 23283
rect 6939 23227 6964 23283
rect 7020 23227 7045 23283
rect 7101 23227 7126 23283
rect 7182 23227 7207 23283
rect 7263 23227 7288 23283
rect 7344 23227 7369 23283
rect 7425 23227 7450 23283
rect 7506 23227 7531 23283
rect 7587 23227 7612 23283
rect 7668 23227 7693 23283
rect 7749 23227 7774 23283
rect 7830 23227 7855 23283
rect 7911 23227 7936 23283
rect 7992 23227 8017 23283
rect 8073 23227 8098 23283
rect 8154 23227 8179 23283
rect 8235 23227 8260 23283
rect 8316 23227 8341 23283
rect 8397 23227 8422 23283
rect 8478 23227 8503 23283
rect 8559 23227 8584 23283
rect 8640 23227 8665 23283
rect 8721 23227 8746 23283
rect 8802 23227 8827 23283
rect 8883 23227 8908 23283
rect 8964 23227 8989 23283
rect 9045 23227 9070 23283
rect 9126 23227 9151 23283
rect 9207 23227 9232 23283
rect 9288 23227 9313 23283
rect 9369 23227 9394 23283
rect 9450 23227 9475 23283
rect 9531 23227 9556 23283
rect 9612 23227 9637 23283
rect 9693 23227 9718 23283
rect 9774 23227 9799 23283
rect 9855 23227 9880 23283
rect 9936 23227 9961 23283
rect 10017 23227 10042 23283
rect 10098 23227 10123 23283
rect 10179 23227 10204 23283
rect 10260 23227 10285 23283
rect 10341 23227 10366 23283
rect 10422 23227 10447 23283
rect 10503 23227 10528 23283
rect 10584 23227 10609 23283
rect 10665 23227 10690 23283
rect 10746 23227 10771 23283
rect 10827 23227 10852 23283
rect 10908 23227 10933 23283
rect 10989 23227 11014 23283
rect 11070 23227 11095 23283
rect 11151 23227 11176 23283
rect 11232 23227 11257 23283
rect 11313 23227 11338 23283
rect 11394 23227 11419 23283
rect 11475 23227 11500 23283
rect 1852 23210 11500 23227
rect 1852 23154 2170 23210
rect 2226 23154 2252 23210
rect 2308 23154 2334 23210
rect 2390 23154 2416 23210
rect 2472 23203 11500 23210
rect 2472 23154 5425 23203
rect 1852 23147 5425 23154
rect 5481 23147 5506 23203
rect 5562 23147 5587 23203
rect 5643 23147 5668 23203
rect 5724 23147 5749 23203
rect 5805 23147 5830 23203
rect 5886 23147 5911 23203
rect 5967 23147 5992 23203
rect 6048 23147 6073 23203
rect 6129 23147 6154 23203
rect 6210 23147 6235 23203
rect 6291 23147 6316 23203
rect 6372 23147 6397 23203
rect 6453 23147 6478 23203
rect 6534 23147 6559 23203
rect 6615 23147 6640 23203
rect 6696 23147 6721 23203
rect 6777 23147 6802 23203
rect 6858 23147 6883 23203
rect 6939 23147 6964 23203
rect 7020 23147 7045 23203
rect 7101 23147 7126 23203
rect 7182 23147 7207 23203
rect 7263 23147 7288 23203
rect 7344 23147 7369 23203
rect 7425 23147 7450 23203
rect 7506 23147 7531 23203
rect 7587 23147 7612 23203
rect 7668 23147 7693 23203
rect 7749 23147 7774 23203
rect 7830 23147 7855 23203
rect 7911 23147 7936 23203
rect 7992 23147 8017 23203
rect 8073 23147 8098 23203
rect 8154 23147 8179 23203
rect 8235 23147 8260 23203
rect 8316 23147 8341 23203
rect 8397 23147 8422 23203
rect 8478 23147 8503 23203
rect 8559 23147 8584 23203
rect 8640 23147 8665 23203
rect 8721 23147 8746 23203
rect 8802 23147 8827 23203
rect 8883 23147 8908 23203
rect 8964 23147 8989 23203
rect 9045 23147 9070 23203
rect 9126 23147 9151 23203
rect 9207 23147 9232 23203
rect 9288 23147 9313 23203
rect 9369 23147 9394 23203
rect 9450 23147 9475 23203
rect 9531 23147 9556 23203
rect 9612 23147 9637 23203
rect 9693 23147 9718 23203
rect 9774 23147 9799 23203
rect 9855 23147 9880 23203
rect 9936 23147 9961 23203
rect 10017 23147 10042 23203
rect 10098 23147 10123 23203
rect 10179 23147 10204 23203
rect 10260 23147 10285 23203
rect 10341 23147 10366 23203
rect 10422 23147 10447 23203
rect 10503 23147 10528 23203
rect 10584 23147 10609 23203
rect 10665 23147 10690 23203
rect 10746 23147 10771 23203
rect 10827 23147 10852 23203
rect 10908 23147 10933 23203
rect 10989 23147 11014 23203
rect 11070 23147 11095 23203
rect 11151 23147 11176 23203
rect 11232 23147 11257 23203
rect 11313 23147 11338 23203
rect 11394 23147 11419 23203
rect 11475 23147 11500 23203
rect 13076 24299 14509 24323
rect 14565 24299 14603 24355
rect 14659 24299 14697 24355
rect 14753 24299 14791 24355
rect 14847 24299 14885 24355
rect 14941 24299 14979 24355
rect 15035 24299 15047 24355
rect 13076 24273 15047 24299
rect 13076 24217 14509 24273
rect 14565 24217 14603 24273
rect 14659 24217 14697 24273
rect 14753 24217 14791 24273
rect 14847 24217 14885 24273
rect 14941 24217 14979 24273
rect 15035 24217 15047 24273
rect 13076 24191 15047 24217
rect 13076 24135 14509 24191
rect 14565 24135 14603 24191
rect 14659 24135 14697 24191
rect 14753 24135 14791 24191
rect 14847 24135 14885 24191
rect 14941 24135 14979 24191
rect 15035 24135 15047 24191
rect 13076 24109 15047 24135
rect 13076 24053 14509 24109
rect 14565 24053 14603 24109
rect 14659 24053 14697 24109
rect 14753 24053 14791 24109
rect 14847 24053 14885 24109
rect 14941 24053 14979 24109
rect 15035 24053 15047 24109
rect 13076 24027 15047 24053
rect 13076 23971 14509 24027
rect 14565 23971 14603 24027
rect 14659 23971 14697 24027
rect 14753 23971 14791 24027
rect 14847 23971 14885 24027
rect 14941 23971 14979 24027
rect 15035 23971 15047 24027
rect 13076 23945 15047 23971
rect 13076 23889 14509 23945
rect 14565 23889 14603 23945
rect 14659 23889 14697 23945
rect 14753 23889 14791 23945
rect 14847 23889 14885 23945
rect 14941 23889 14979 23945
rect 15035 23889 15047 23945
rect 13076 23863 15047 23889
rect 13076 23807 14509 23863
rect 14565 23807 14603 23863
rect 14659 23807 14697 23863
rect 14753 23807 14791 23863
rect 14847 23807 14885 23863
rect 14941 23807 14979 23863
rect 15035 23807 15047 23863
rect 13076 23781 15047 23807
rect 13076 23725 14509 23781
rect 14565 23725 14603 23781
rect 14659 23725 14697 23781
rect 14753 23725 14791 23781
rect 14847 23725 14885 23781
rect 14941 23725 14979 23781
rect 15035 23725 15047 23781
rect 13076 23699 15047 23725
rect 13076 23643 14509 23699
rect 14565 23643 14603 23699
rect 14659 23643 14697 23699
rect 14753 23643 14791 23699
rect 14847 23643 14885 23699
rect 14941 23643 14979 23699
rect 15035 23643 15047 23699
rect 13076 23617 15047 23643
rect 13076 23561 14509 23617
rect 14565 23561 14603 23617
rect 14659 23561 14697 23617
rect 14753 23561 14791 23617
rect 14847 23561 14885 23617
rect 14941 23561 14979 23617
rect 15035 23561 15047 23617
rect 13076 23535 15047 23561
rect 13076 23479 14509 23535
rect 14565 23479 14603 23535
rect 14659 23479 14697 23535
rect 14753 23479 14791 23535
rect 14847 23479 14885 23535
rect 14941 23479 14979 23535
rect 15035 23479 15047 23535
rect 13076 23453 15047 23479
rect 13076 23397 14509 23453
rect 14565 23397 14603 23453
rect 14659 23397 14697 23453
rect 14753 23397 14791 23453
rect 14847 23397 14885 23453
rect 14941 23397 14979 23453
rect 15035 23397 15047 23453
rect 13076 23371 15047 23397
rect 13076 23315 14509 23371
rect 14565 23315 14603 23371
rect 14659 23315 14697 23371
rect 14753 23315 14791 23371
rect 14847 23315 14885 23371
rect 14941 23315 14979 23371
rect 15035 23315 15047 23371
rect 13076 23289 15047 23315
rect 13076 23233 14509 23289
rect 14565 23233 14603 23289
rect 14659 23233 14697 23289
rect 14753 23233 14791 23289
rect 14847 23233 14885 23289
rect 14941 23233 14979 23289
rect 15035 23233 15047 23289
rect 13076 23207 15047 23233
rect 13076 23151 14509 23207
rect 14565 23151 14603 23207
rect 14659 23151 14697 23207
rect 14753 23151 14791 23207
rect 14847 23151 14885 23207
rect 14941 23151 14979 23207
rect 15035 23151 15047 23207
rect 13076 23147 15047 23151
rect 1852 23136 15047 23147
rect 148 23094 850 23106
rect 148 23042 149 23094
rect 201 23042 247 23094
rect 299 23042 456 23094
rect 508 23042 524 23094
rect 576 23042 592 23094
rect 644 23042 660 23094
rect 712 23042 728 23094
rect 780 23042 796 23094
rect 848 23042 850 23094
rect 148 23030 850 23042
rect 148 22978 149 23030
rect 201 22978 247 23030
rect 299 22978 456 23030
rect 508 22978 524 23030
rect 576 22978 592 23030
rect 644 22978 660 23030
rect 712 22978 728 23030
rect 780 22978 796 23030
rect 848 22978 850 23030
rect 148 22966 850 22978
rect 148 22914 149 22966
rect 201 22914 247 22966
rect 299 22914 456 22966
rect 508 22914 524 22966
rect 576 22914 592 22966
rect 644 22914 660 22966
rect 712 22914 728 22966
rect 780 22914 796 22966
rect 848 22914 850 22966
rect 148 22902 850 22914
rect 148 22850 149 22902
rect 201 22850 247 22902
rect 299 22850 456 22902
rect 508 22850 524 22902
rect 576 22850 592 22902
rect 644 22850 660 22902
rect 712 22850 728 22902
rect 780 22850 796 22902
rect 848 22850 850 22902
rect 148 22838 850 22850
rect 148 22786 149 22838
rect 201 22786 247 22838
rect 299 22786 456 22838
rect 508 22786 524 22838
rect 576 22786 592 22838
rect 644 22786 660 22838
rect 712 22786 728 22838
rect 780 22786 796 22838
rect 848 22786 850 22838
rect 148 22774 850 22786
rect 148 22722 149 22774
rect 201 22722 247 22774
rect 299 22722 456 22774
rect 508 22722 524 22774
rect 576 22722 592 22774
rect 644 22722 660 22774
rect 712 22722 728 22774
rect 780 22722 796 22774
rect 848 22722 850 22774
rect 148 22710 850 22722
rect 148 22658 149 22710
rect 201 22658 247 22710
rect 299 22658 456 22710
rect 508 22658 524 22710
rect 576 22658 592 22710
rect 644 22658 660 22710
rect 712 22658 728 22710
rect 780 22658 796 22710
rect 848 22658 850 22710
rect 148 22646 850 22658
rect 148 22594 149 22646
rect 201 22594 247 22646
rect 299 22594 456 22646
rect 508 22594 524 22646
rect 576 22594 592 22646
rect 644 22594 660 22646
rect 712 22594 728 22646
rect 780 22594 796 22646
rect 848 22594 850 22646
rect 148 22582 850 22594
rect 148 22530 149 22582
rect 201 22530 247 22582
rect 299 22530 456 22582
rect 508 22530 524 22582
rect 576 22530 592 22582
rect 644 22530 660 22582
rect 712 22530 728 22582
rect 780 22530 796 22582
rect 848 22530 850 22582
rect 148 22518 850 22530
rect 148 22466 149 22518
rect 201 22466 247 22518
rect 299 22466 456 22518
rect 508 22466 524 22518
rect 576 22466 592 22518
rect 644 22466 660 22518
rect 712 22466 728 22518
rect 780 22466 796 22518
rect 848 22466 850 22518
rect 148 22454 850 22466
rect 148 22402 149 22454
rect 201 22402 247 22454
rect 299 22402 456 22454
rect 508 22402 524 22454
rect 576 22402 592 22454
rect 644 22402 660 22454
rect 712 22402 728 22454
rect 780 22402 796 22454
rect 848 22402 850 22454
rect 148 22390 850 22402
rect 148 22338 149 22390
rect 201 22338 247 22390
rect 299 22338 456 22390
rect 508 22338 524 22390
rect 576 22338 592 22390
rect 644 22338 660 22390
rect 712 22338 728 22390
rect 780 22338 796 22390
rect 848 22338 850 22390
rect 148 22326 850 22338
rect 148 22274 149 22326
rect 201 22274 247 22326
rect 299 22274 456 22326
rect 508 22274 524 22326
rect 576 22274 592 22326
rect 644 22274 660 22326
rect 712 22274 728 22326
rect 780 22274 796 22326
rect 848 22274 850 22326
rect 148 22262 850 22274
rect 148 22210 149 22262
rect 201 22210 247 22262
rect 299 22210 456 22262
rect 508 22210 524 22262
rect 576 22210 592 22262
rect 644 22210 660 22262
rect 712 22210 728 22262
rect 780 22210 796 22262
rect 848 22210 850 22262
rect 148 22198 850 22210
rect 148 22146 149 22198
rect 201 22146 247 22198
rect 299 22146 456 22198
rect 508 22146 524 22198
rect 576 22146 592 22198
rect 644 22146 660 22198
rect 712 22146 728 22198
rect 780 22146 796 22198
rect 848 22146 850 22198
rect 148 22134 850 22146
rect 148 22082 149 22134
rect 201 22082 247 22134
rect 299 22082 456 22134
rect 508 22082 524 22134
rect 576 22082 592 22134
rect 644 22082 660 22134
rect 712 22082 728 22134
rect 780 22082 796 22134
rect 848 22082 850 22134
rect 148 22070 850 22082
rect 148 22018 149 22070
rect 201 22018 247 22070
rect 299 22018 456 22070
rect 508 22018 524 22070
rect 576 22018 592 22070
rect 644 22018 660 22070
rect 712 22018 728 22070
rect 780 22018 796 22070
rect 848 22018 850 22070
rect 148 22006 850 22018
rect 148 21954 149 22006
rect 201 21954 247 22006
rect 299 21954 456 22006
rect 508 21954 524 22006
rect 576 21954 592 22006
rect 644 21954 660 22006
rect 712 21954 728 22006
rect 780 21954 796 22006
rect 848 21954 850 22006
rect 148 21942 850 21954
rect 148 21890 149 21942
rect 201 21890 247 21942
rect 299 21890 456 21942
rect 508 21890 524 21942
rect 576 21890 592 21942
rect 644 21890 660 21942
rect 712 21890 728 21942
rect 780 21890 796 21942
rect 848 21890 850 21942
rect 148 21878 850 21890
rect 148 21826 149 21878
rect 201 21826 247 21878
rect 299 21826 456 21878
rect 508 21826 524 21878
rect 576 21826 592 21878
rect 644 21826 660 21878
rect 712 21826 728 21878
rect 780 21826 796 21878
rect 848 21826 850 21878
rect 148 21814 850 21826
rect 148 21762 149 21814
rect 201 21762 247 21814
rect 299 21762 456 21814
rect 508 21762 524 21814
rect 576 21762 592 21814
rect 644 21762 660 21814
rect 712 21762 728 21814
rect 780 21762 796 21814
rect 848 21762 850 21814
rect 148 21750 850 21762
rect 148 21698 149 21750
rect 201 21698 247 21750
rect 299 21698 456 21750
rect 508 21698 524 21750
rect 576 21698 592 21750
rect 644 21698 660 21750
rect 712 21698 728 21750
rect 780 21698 796 21750
rect 848 21698 850 21750
rect 148 21686 850 21698
rect 148 21634 149 21686
rect 201 21634 247 21686
rect 299 21634 456 21686
rect 508 21634 524 21686
rect 576 21634 592 21686
rect 644 21634 660 21686
rect 712 21634 728 21686
rect 780 21634 796 21686
rect 848 21634 850 21686
rect 148 21622 850 21634
rect 148 21570 149 21622
rect 201 21570 247 21622
rect 299 21570 456 21622
rect 508 21570 524 21622
rect 576 21570 592 21622
rect 644 21570 660 21622
rect 712 21570 728 21622
rect 780 21570 796 21622
rect 848 21570 850 21622
rect 148 21558 850 21570
rect 148 21506 149 21558
rect 201 21506 247 21558
rect 299 21506 456 21558
rect 508 21506 524 21558
rect 576 21506 592 21558
rect 644 21506 660 21558
rect 712 21506 728 21558
rect 780 21506 796 21558
rect 848 21506 850 21558
rect 148 21494 850 21506
rect 148 21442 149 21494
rect 201 21442 247 21494
rect 299 21442 456 21494
rect 508 21442 524 21494
rect 576 21442 592 21494
rect 644 21442 660 21494
rect 712 21442 728 21494
rect 780 21442 796 21494
rect 848 21442 850 21494
rect 148 21430 850 21442
rect 148 21378 149 21430
rect 201 21378 247 21430
rect 299 21378 456 21430
rect 508 21378 524 21430
rect 576 21378 592 21430
rect 644 21378 660 21430
rect 712 21378 728 21430
rect 780 21378 796 21430
rect 848 21378 850 21430
rect 148 21366 850 21378
rect 148 21314 149 21366
rect 201 21314 247 21366
rect 299 21314 456 21366
rect 508 21314 524 21366
rect 576 21314 592 21366
rect 644 21314 660 21366
rect 712 21314 728 21366
rect 780 21314 796 21366
rect 848 21314 850 21366
rect 148 21302 850 21314
rect 148 21250 149 21302
rect 201 21250 247 21302
rect 299 21250 456 21302
rect 508 21250 524 21302
rect 576 21250 592 21302
rect 644 21250 660 21302
rect 712 21250 728 21302
rect 780 21250 796 21302
rect 848 21250 850 21302
rect 148 21238 850 21250
rect 148 21186 149 21238
rect 201 21186 247 21238
rect 299 21186 456 21238
rect 508 21186 524 21238
rect 576 21186 592 21238
rect 644 21186 660 21238
rect 712 21186 728 21238
rect 780 21186 796 21238
rect 848 21186 850 21238
rect 148 21174 850 21186
rect 148 21122 149 21174
rect 201 21122 247 21174
rect 299 21122 456 21174
rect 508 21122 524 21174
rect 576 21122 592 21174
rect 644 21122 660 21174
rect 712 21122 728 21174
rect 780 21122 796 21174
rect 848 21122 850 21174
rect 148 21110 850 21122
rect 148 21058 149 21110
rect 201 21058 247 21110
rect 299 21058 456 21110
rect 508 21058 524 21110
rect 576 21058 592 21110
rect 644 21058 660 21110
rect 712 21058 728 21110
rect 780 21058 796 21110
rect 848 21058 850 21110
rect 148 21046 850 21058
rect 148 20994 149 21046
rect 201 20994 247 21046
rect 299 20994 456 21046
rect 508 20994 524 21046
rect 576 20994 592 21046
rect 644 20994 660 21046
rect 712 20994 728 21046
rect 780 20994 796 21046
rect 848 20994 850 21046
rect 148 20982 850 20994
rect 148 20930 149 20982
rect 201 20930 247 20982
rect 299 20930 456 20982
rect 508 20930 524 20982
rect 576 20930 592 20982
rect 644 20930 660 20982
rect 712 20930 728 20982
rect 780 20930 796 20982
rect 848 20930 850 20982
rect 148 20923 850 20930
rect 148 20918 670 20923
rect 726 20918 794 20923
rect 148 20866 149 20918
rect 201 20866 247 20918
rect 299 20866 456 20918
rect 508 20866 524 20918
rect 576 20866 592 20918
rect 644 20866 660 20918
rect 726 20867 728 20918
rect 712 20866 728 20867
rect 780 20867 794 20918
rect 780 20866 796 20867
rect 848 20866 850 20867
rect 148 20854 850 20866
rect 148 20802 149 20854
rect 201 20802 247 20854
rect 299 20802 456 20854
rect 508 20802 524 20854
rect 576 20802 592 20854
rect 644 20802 660 20854
rect 712 20832 728 20854
rect 726 20802 728 20832
rect 780 20832 796 20854
rect 848 20832 850 20854
rect 780 20802 794 20832
rect 148 20790 670 20802
rect 726 20790 794 20802
rect 148 20738 149 20790
rect 201 20738 247 20790
rect 299 20738 456 20790
rect 508 20738 524 20790
rect 576 20738 592 20790
rect 644 20738 660 20790
rect 726 20776 728 20790
rect 712 20741 728 20776
rect 726 20738 728 20741
rect 780 20776 794 20790
rect 780 20741 796 20776
rect 848 20741 850 20776
rect 780 20738 794 20741
rect 148 20726 670 20738
rect 726 20726 794 20738
rect 148 20674 149 20726
rect 201 20674 247 20726
rect 299 20674 456 20726
rect 508 20674 524 20726
rect 576 20674 592 20726
rect 644 20674 660 20726
rect 726 20685 728 20726
rect 712 20674 728 20685
rect 780 20685 794 20726
rect 780 20674 796 20685
rect 848 20674 850 20685
rect 148 20662 850 20674
rect 148 20610 149 20662
rect 201 20610 247 20662
rect 299 20610 456 20662
rect 508 20610 524 20662
rect 576 20610 592 20662
rect 644 20610 660 20662
rect 712 20650 728 20662
rect 726 20610 728 20650
rect 780 20650 796 20662
rect 848 20650 850 20662
rect 780 20610 794 20650
rect 148 20598 670 20610
rect 726 20598 794 20610
rect 148 20546 149 20598
rect 201 20546 247 20598
rect 299 20546 456 20598
rect 508 20546 524 20598
rect 576 20546 592 20598
rect 644 20546 660 20598
rect 726 20594 728 20598
rect 712 20559 728 20594
rect 726 20546 728 20559
rect 780 20594 794 20598
rect 780 20559 796 20594
rect 848 20559 850 20594
rect 780 20546 794 20559
rect 148 20534 670 20546
rect 726 20534 794 20546
rect 148 20482 149 20534
rect 201 20482 247 20534
rect 299 20482 456 20534
rect 508 20482 524 20534
rect 576 20482 592 20534
rect 644 20482 660 20534
rect 726 20503 728 20534
rect 712 20482 728 20503
rect 780 20503 794 20534
rect 780 20482 796 20503
rect 848 20482 850 20503
rect 148 20470 850 20482
rect 148 20418 149 20470
rect 201 20418 247 20470
rect 299 20418 456 20470
rect 508 20418 524 20470
rect 576 20418 592 20470
rect 644 20418 660 20470
rect 712 20468 728 20470
rect 726 20418 728 20468
rect 780 20468 796 20470
rect 848 20468 850 20470
rect 780 20418 794 20468
rect 148 20412 670 20418
rect 726 20412 794 20418
rect 148 20406 850 20412
rect 148 20354 149 20406
rect 201 20354 247 20406
rect 299 20354 456 20406
rect 508 20354 524 20406
rect 576 20354 592 20406
rect 644 20354 660 20406
rect 712 20354 728 20406
rect 780 20354 796 20406
rect 848 20354 850 20406
rect 1625 20931 3768 20932
rect 1625 20923 2790 20931
rect 1625 20867 1627 20923
rect 1683 20867 1715 20923
rect 1771 20867 1803 20923
rect 1859 20867 1891 20923
rect 1947 20867 1979 20923
rect 2035 20867 2067 20923
rect 2123 20875 2790 20923
rect 2846 20875 2873 20931
rect 2929 20875 2956 20931
rect 3012 20875 3039 20931
rect 3095 20875 3122 20931
rect 3178 20875 3205 20931
rect 3261 20875 3288 20931
rect 3344 20875 3371 20931
rect 3427 20875 3454 20931
rect 3510 20875 3537 20931
rect 3593 20875 3620 20931
rect 3676 20875 3703 20931
rect 3759 20875 3768 20931
rect 2123 20867 3768 20875
rect 1625 20837 3768 20867
rect 1625 20832 2790 20837
rect 1625 20776 1627 20832
rect 1683 20776 1715 20832
rect 1771 20776 1803 20832
rect 1859 20776 1891 20832
rect 1947 20776 1979 20832
rect 2035 20776 2067 20832
rect 2123 20781 2790 20832
rect 2846 20781 2873 20837
rect 2929 20781 2956 20837
rect 3012 20781 3039 20837
rect 3095 20781 3122 20837
rect 3178 20781 3205 20837
rect 3261 20781 3288 20837
rect 3344 20781 3371 20837
rect 3427 20781 3454 20837
rect 3510 20781 3537 20837
rect 3593 20781 3620 20837
rect 3676 20781 3703 20837
rect 3759 20781 3768 20837
rect 2123 20776 3768 20781
rect 1625 20743 3768 20776
rect 1625 20741 2790 20743
rect 1625 20685 1627 20741
rect 1683 20685 1715 20741
rect 1771 20685 1803 20741
rect 1859 20685 1891 20741
rect 1947 20685 1979 20741
rect 2035 20685 2067 20741
rect 2123 20687 2790 20741
rect 2846 20687 2873 20743
rect 2929 20687 2956 20743
rect 3012 20687 3039 20743
rect 3095 20687 3122 20743
rect 3178 20687 3205 20743
rect 3261 20687 3288 20743
rect 3344 20687 3371 20743
rect 3427 20687 3454 20743
rect 3510 20687 3537 20743
rect 3593 20687 3620 20743
rect 3676 20687 3703 20743
rect 3759 20687 3768 20743
rect 2123 20685 3768 20687
rect 1625 20650 3768 20685
rect 1625 20594 1627 20650
rect 1683 20594 1715 20650
rect 1771 20594 1803 20650
rect 1859 20594 1891 20650
rect 1947 20594 1979 20650
rect 2035 20594 2067 20650
rect 2123 20649 3768 20650
rect 2123 20594 2790 20649
rect 1625 20593 2790 20594
rect 2846 20593 2873 20649
rect 2929 20593 2956 20649
rect 3012 20593 3039 20649
rect 3095 20593 3122 20649
rect 3178 20593 3205 20649
rect 3261 20593 3288 20649
rect 3344 20593 3371 20649
rect 3427 20593 3454 20649
rect 3510 20593 3537 20649
rect 3593 20593 3620 20649
rect 3676 20593 3703 20649
rect 3759 20593 3768 20649
rect 1625 20571 3768 20593
rect 1625 20559 2784 20571
rect 1625 20503 1627 20559
rect 1683 20503 1715 20559
rect 1771 20503 1803 20559
rect 1859 20503 1891 20559
rect 1947 20503 1979 20559
rect 2035 20503 2067 20559
rect 2123 20519 2784 20559
rect 2836 20555 2853 20571
rect 2905 20555 2922 20571
rect 2974 20555 2991 20571
rect 3043 20555 3060 20571
rect 3112 20555 3128 20571
rect 2846 20519 2853 20555
rect 3112 20519 3122 20555
rect 3180 20519 3196 20571
rect 3248 20555 3264 20571
rect 3316 20555 3332 20571
rect 3384 20555 3400 20571
rect 3452 20555 3468 20571
rect 3261 20519 3264 20555
rect 3452 20519 3454 20555
rect 3520 20519 3536 20571
rect 3588 20555 3604 20571
rect 3656 20555 3672 20571
rect 3724 20555 3768 20571
rect 3593 20519 3604 20555
rect 2123 20503 2790 20519
rect 1625 20499 2790 20503
rect 2846 20499 2873 20519
rect 2929 20499 2956 20519
rect 3012 20499 3039 20519
rect 3095 20499 3122 20519
rect 3178 20499 3205 20519
rect 3261 20499 3288 20519
rect 3344 20499 3371 20519
rect 3427 20499 3454 20519
rect 3510 20499 3537 20519
rect 3593 20499 3620 20519
rect 3676 20499 3703 20519
rect 3759 20499 3768 20555
rect 1625 20468 3768 20499
rect 1625 20412 1627 20468
rect 1683 20412 1715 20468
rect 1771 20412 1803 20468
rect 1859 20412 1891 20468
rect 1947 20412 1979 20468
rect 2035 20412 2067 20468
rect 2123 20461 3768 20468
rect 2123 20459 2790 20461
rect 2846 20459 2873 20461
rect 2929 20459 2956 20461
rect 3012 20459 3039 20461
rect 3095 20459 3122 20461
rect 3178 20459 3205 20461
rect 3261 20459 3288 20461
rect 3344 20459 3371 20461
rect 3427 20459 3454 20461
rect 3510 20459 3537 20461
rect 3593 20459 3620 20461
rect 3676 20459 3703 20461
rect 2123 20412 2784 20459
rect 1625 20407 2784 20412
rect 2846 20407 2853 20459
rect 3112 20407 3122 20459
rect 3180 20407 3196 20459
rect 3261 20407 3264 20459
rect 3452 20407 3454 20459
rect 3520 20407 3536 20459
rect 3593 20407 3604 20459
rect 1625 20405 2790 20407
rect 2846 20405 2873 20407
rect 2929 20405 2956 20407
rect 3012 20405 3039 20407
rect 3095 20405 3122 20407
rect 3178 20405 3205 20407
rect 3261 20405 3288 20407
rect 3344 20405 3371 20407
rect 3427 20405 3454 20407
rect 3510 20405 3537 20407
rect 3593 20405 3620 20407
rect 3676 20405 3703 20407
rect 3759 20405 3768 20461
rect 1625 20403 3768 20405
rect 12199 20566 12251 20572
rect 12199 20496 12251 20514
rect 12199 20425 12251 20444
rect 148 20342 850 20354
rect 148 20290 149 20342
rect 201 20290 247 20342
rect 299 20290 456 20342
rect 508 20290 524 20342
rect 576 20290 592 20342
rect 644 20290 660 20342
rect 712 20290 728 20342
rect 780 20290 796 20342
rect 848 20290 850 20342
rect 148 20277 850 20290
rect 148 20225 149 20277
rect 201 20225 247 20277
rect 299 20225 456 20277
rect 508 20225 524 20277
rect 576 20225 592 20277
rect 644 20225 660 20277
rect 712 20225 728 20277
rect 780 20225 796 20277
rect 848 20225 850 20277
rect 148 20212 850 20225
rect 148 20160 149 20212
rect 201 20160 247 20212
rect 299 20160 456 20212
rect 508 20160 524 20212
rect 576 20160 592 20212
rect 644 20160 660 20212
rect 712 20160 728 20212
rect 780 20160 796 20212
rect 848 20160 850 20212
rect 148 20147 850 20160
rect 148 20095 149 20147
rect 201 20095 247 20147
rect 299 20095 456 20147
rect 508 20095 524 20147
rect 576 20095 592 20147
rect 644 20095 660 20147
rect 712 20095 728 20147
rect 780 20095 796 20147
rect 848 20095 850 20147
rect 148 20082 850 20095
rect 148 20030 149 20082
rect 201 20030 247 20082
rect 299 20030 456 20082
rect 508 20030 524 20082
rect 576 20030 592 20082
rect 644 20030 660 20082
rect 712 20030 728 20082
rect 780 20030 796 20082
rect 848 20030 850 20082
rect 148 20017 850 20030
rect 148 19965 149 20017
rect 201 19965 247 20017
rect 299 19965 456 20017
rect 508 19965 524 20017
rect 576 19965 592 20017
rect 644 19965 660 20017
rect 712 19965 728 20017
rect 780 19965 796 20017
rect 848 19965 850 20017
rect 148 19952 850 19965
rect 148 19900 149 19952
rect 201 19900 247 19952
rect 299 19900 456 19952
rect 508 19900 524 19952
rect 576 19900 592 19952
rect 644 19900 660 19952
rect 712 19900 728 19952
rect 780 19900 796 19952
rect 848 19900 850 19952
rect 148 19887 850 19900
rect 148 19835 149 19887
rect 201 19835 247 19887
rect 299 19835 456 19887
rect 508 19835 524 19887
rect 576 19835 592 19887
rect 644 19835 660 19887
rect 712 19835 728 19887
rect 780 19835 796 19887
rect 848 19835 850 19887
rect 148 19822 850 19835
rect 148 19770 149 19822
rect 201 19770 247 19822
rect 299 19770 456 19822
rect 508 19770 524 19822
rect 576 19770 592 19822
rect 644 19770 660 19822
rect 712 19770 728 19822
rect 780 19770 796 19822
rect 848 19770 850 19822
rect 148 19757 850 19770
rect 148 19705 149 19757
rect 201 19705 247 19757
rect 299 19705 456 19757
rect 508 19705 524 19757
rect 576 19705 592 19757
rect 644 19705 660 19757
rect 712 19705 728 19757
rect 780 19705 796 19757
rect 848 19705 850 19757
rect 148 19692 850 19705
rect 148 19640 149 19692
rect 201 19640 247 19692
rect 299 19640 456 19692
rect 508 19640 524 19692
rect 576 19640 592 19692
rect 644 19640 660 19692
rect 712 19640 728 19692
rect 780 19640 796 19692
rect 848 19640 850 19692
rect 12199 20354 12251 20373
rect 12199 20283 12251 20302
rect 12199 20110 12251 20231
rect 12199 20046 12251 20058
rect 12199 19982 12251 19994
rect 12199 19918 12251 19930
rect 12199 19854 12251 19866
rect 12199 19790 12251 19802
rect 12199 19725 12251 19738
rect 12199 19667 12251 19673
rect 148 19627 850 19640
rect 148 19575 149 19627
rect 201 19575 247 19627
rect 299 19575 456 19627
rect 508 19575 524 19627
rect 576 19575 592 19627
rect 644 19575 660 19627
rect 712 19575 728 19627
rect 780 19575 796 19627
rect 848 19575 850 19627
rect 148 19562 850 19575
rect 148 19510 149 19562
rect 201 19510 247 19562
rect 299 19510 456 19562
rect 508 19510 524 19562
rect 576 19510 592 19562
rect 644 19510 660 19562
rect 712 19510 728 19562
rect 780 19510 796 19562
rect 848 19510 850 19562
rect 148 19497 850 19510
rect 148 19445 149 19497
rect 201 19445 247 19497
rect 299 19445 456 19497
rect 508 19445 524 19497
rect 576 19445 592 19497
rect 644 19445 660 19497
rect 712 19445 728 19497
rect 780 19445 796 19497
rect 848 19445 850 19497
rect 148 19432 850 19445
rect 148 19380 149 19432
rect 201 19380 247 19432
rect 299 19380 456 19432
rect 508 19380 524 19432
rect 576 19380 592 19432
rect 644 19380 660 19432
rect 712 19380 728 19432
rect 780 19380 796 19432
rect 848 19380 850 19432
rect 148 19367 850 19380
rect 148 19315 149 19367
rect 201 19315 247 19367
rect 299 19315 456 19367
rect 508 19315 524 19367
rect 576 19315 592 19367
rect 644 19315 660 19367
rect 712 19315 728 19367
rect 780 19315 796 19367
rect 848 19315 850 19367
rect 148 19302 850 19315
rect 148 19250 149 19302
rect 201 19250 247 19302
rect 299 19250 456 19302
rect 508 19250 524 19302
rect 576 19250 592 19302
rect 644 19250 660 19302
rect 712 19250 728 19302
rect 780 19250 796 19302
rect 848 19250 850 19302
rect 148 19237 850 19250
tri 15377 19243 15379 19245 ne
rect 15379 19243 15423 19245
rect 148 19185 149 19237
rect 201 19185 247 19237
rect 299 19185 456 19237
rect 508 19185 524 19237
rect 576 19185 592 19237
rect 644 19185 660 19237
rect 712 19185 728 19237
rect 780 19185 796 19237
rect 848 19185 850 19237
rect 2781 19191 2787 19243
rect 2846 19191 2854 19243
rect 3040 19191 3042 19243
rect 3107 19191 3122 19243
rect 3182 19191 3189 19243
rect 3375 19191 3378 19243
rect 3442 19191 3456 19243
rect 3518 19191 3522 19243
rect 3706 19191 3713 19243
rect 3772 19191 3778 19243
tri 15379 19239 15383 19243 ne
rect 2781 19187 2790 19191
rect 2846 19187 2874 19191
rect 2930 19187 2958 19191
rect 3014 19187 3042 19191
rect 3098 19187 3126 19191
rect 3182 19187 3210 19191
rect 3266 19187 3294 19191
rect 3350 19187 3378 19191
rect 3434 19187 3462 19191
rect 3518 19187 3546 19191
rect 3602 19187 3630 19191
rect 3686 19187 3713 19191
rect 3769 19187 3778 19191
rect 148 19179 850 19185
rect 3016 19069 3025 19073
rect 3081 19069 3111 19073
rect 3167 19069 3197 19073
rect 3253 19069 3283 19073
rect 3339 19069 3369 19073
rect 3425 19069 3455 19073
rect 3511 19069 3541 19073
rect 3597 19069 3627 19073
rect 3683 19069 3713 19073
rect 3769 19069 3778 19073
rect 3016 19017 3022 19069
rect 3081 19017 3092 19069
rect 3354 19017 3369 19069
rect 3425 19017 3442 19069
rect 3511 19017 3512 19069
rect 3703 19017 3713 19069
rect 3772 19017 3778 19069
rect 269 18824 276 18876
rect 328 18824 341 18876
rect 393 18824 406 18876
rect 458 18824 471 18876
rect 523 18824 536 18876
rect 588 18824 601 18876
rect 653 18824 666 18876
rect 718 18824 725 18876
rect 269 18794 725 18824
rect 269 18742 276 18794
rect 328 18742 341 18794
rect 393 18742 406 18794
rect 458 18742 471 18794
rect 523 18742 536 18794
rect 588 18742 601 18794
rect 653 18742 666 18794
rect 718 18742 725 18794
rect 269 18712 725 18742
rect 269 18660 276 18712
rect 328 18660 341 18712
rect 393 18660 406 18712
rect 458 18660 471 18712
rect 523 18660 536 18712
rect 588 18660 601 18712
rect 653 18660 666 18712
rect 718 18660 725 18712
rect 1251 18824 1257 18876
rect 1309 18824 1325 18876
rect 1377 18824 1393 18876
rect 1445 18824 1461 18876
rect 1513 18824 1528 18876
rect 1580 18824 1595 18876
rect 1647 18824 1730 18876
rect 1251 18794 1730 18824
rect 1251 18742 1257 18794
rect 1309 18742 1325 18794
rect 1377 18742 1393 18794
rect 1445 18742 1461 18794
rect 1513 18742 1528 18794
rect 1580 18742 1595 18794
rect 1647 18742 1730 18794
rect 1251 18712 1730 18742
rect 1251 18660 1257 18712
rect 1309 18660 1325 18712
rect 1377 18660 1393 18712
rect 1445 18660 1461 18712
rect 1513 18660 1528 18712
rect 1580 18660 1595 18712
rect 1647 18678 1730 18712
tri 1730 18678 1928 18876 sw
rect 1647 18660 1928 18678
rect 269 18294 725 18660
tri 1578 18517 1721 18660 ne
rect 1721 16857 1928 18660
rect 3198 17349 3207 17353
rect 3198 17297 3204 17349
rect 3263 17297 3289 17353
rect 3345 17349 3354 17353
rect 3348 17297 3354 17349
rect 8445 17283 8941 17285
rect 8445 17227 8454 17283
rect 8510 17227 8604 17283
rect 8660 17227 8754 17283
rect 8810 17227 8903 17283
rect 8959 17227 9052 17283
rect 9108 17227 9117 17283
rect 8445 17195 9117 17227
rect 8445 17139 8454 17195
rect 8510 17139 8604 17195
rect 8660 17139 8754 17195
rect 8810 17139 8903 17195
rect 8959 17139 9052 17195
rect 9108 17139 9117 17195
rect 8445 17107 9117 17139
rect 8445 17051 8454 17107
rect 8510 17051 8604 17107
rect 8660 17051 8754 17107
rect 8810 17051 8903 17107
rect 8959 17051 9052 17107
rect 9108 17051 9117 17107
tri 1721 16777 1801 16857 ne
rect 1801 16777 1928 16857
tri 1928 16777 2107 16956 sw
rect 5731 16795 9142 16802
rect 5731 16777 7041 16795
rect 7097 16777 7121 16795
rect 7177 16777 9142 16795
tri 1801 16725 1853 16777 ne
rect 1853 16725 2107 16777
tri 2107 16725 2159 16777 sw
rect 5731 16725 5737 16777
rect 5789 16725 5802 16777
rect 5854 16725 5867 16777
rect 5919 16725 5932 16777
rect 5984 16725 5997 16777
rect 6049 16725 6062 16777
rect 6114 16725 6127 16777
rect 6179 16725 6192 16777
rect 6244 16725 6257 16777
rect 6309 16725 6322 16777
rect 6374 16725 6387 16777
rect 6439 16725 6452 16777
rect 6504 16725 6517 16777
rect 6569 16725 6582 16777
rect 6634 16725 6647 16777
rect 6699 16725 6712 16777
rect 6764 16725 6777 16777
rect 6829 16725 6842 16777
rect 6894 16725 6907 16777
rect 6959 16725 6972 16777
rect 7024 16725 7036 16777
rect 7097 16739 7100 16777
rect 7088 16725 7100 16739
rect 7152 16725 7164 16739
rect 7216 16725 7228 16777
rect 7280 16725 7292 16777
rect 7344 16725 7356 16777
rect 7408 16725 7420 16777
rect 7472 16725 7484 16777
rect 7536 16725 7548 16777
rect 7600 16725 7612 16777
rect 7664 16725 7676 16777
rect 7728 16725 7740 16777
rect 7792 16725 7804 16777
rect 7856 16725 7868 16777
rect 7920 16725 7932 16777
rect 7984 16725 7996 16777
rect 8048 16725 8060 16777
rect 8112 16725 8124 16777
rect 8176 16725 8188 16777
rect 8240 16725 8252 16777
rect 8304 16725 8316 16777
rect 8368 16725 8380 16777
rect 8432 16725 8444 16777
rect 8496 16725 8508 16777
rect 8560 16725 8572 16777
rect 8624 16725 8636 16777
rect 8688 16725 8700 16777
rect 8752 16725 8764 16777
rect 8816 16725 8828 16777
rect 8880 16725 8892 16777
rect 8944 16725 8956 16777
rect 9008 16725 9020 16777
rect 9072 16725 9084 16777
rect 9136 16725 9142 16777
tri 1853 16689 1889 16725 ne
rect 1889 16689 2159 16725
tri 2159 16689 2195 16725 sw
rect 5731 16700 9142 16725
tri 1889 16650 1928 16689 ne
rect 1928 16650 2195 16689
tri 1928 16383 2195 16650 ne
tri 2195 16383 2501 16689 sw
rect 8445 16395 8454 16451
rect 8510 16395 8604 16451
rect 8660 16395 8754 16451
rect 8810 16395 8903 16451
rect 8959 16395 9052 16451
rect 9108 16395 9117 16451
tri 2195 16167 2411 16383 ne
rect 2411 16327 3894 16383
rect 3950 16327 4019 16383
rect 4075 16327 4144 16383
rect 4200 16327 4269 16383
rect 4325 16327 4334 16383
rect 2411 16303 4334 16327
rect 2411 16247 3894 16303
rect 3950 16247 4019 16303
rect 4075 16247 4144 16303
rect 4200 16247 4269 16303
rect 4325 16247 4334 16303
rect 2411 16223 4334 16247
rect 2411 16167 3894 16223
rect 3950 16167 4019 16223
rect 4075 16167 4144 16223
rect 4200 16167 4269 16223
rect 4325 16167 4334 16223
rect 8445 16363 9117 16395
rect 8445 16307 8454 16363
rect 8510 16307 8604 16363
rect 8660 16307 8754 16363
rect 8810 16307 8903 16363
rect 8959 16307 9052 16363
rect 9108 16307 9117 16363
rect 8445 16275 9117 16307
rect 8445 16219 8454 16275
rect 8510 16219 8604 16275
rect 8660 16219 8754 16275
rect 8810 16219 8903 16275
rect 8959 16219 9052 16275
rect 9108 16219 9117 16275
rect 8445 16217 8941 16219
rect 7396 16154 9292 16155
rect 7396 16102 7402 16154
rect 7454 16102 7469 16154
rect 7521 16102 7536 16154
rect 7588 16102 7602 16154
rect 7654 16102 9196 16154
rect 9248 16102 9292 16154
rect 7396 16082 9292 16102
rect 7396 16030 7402 16082
rect 7454 16030 7469 16082
rect 7521 16030 7536 16082
rect 7588 16030 7602 16082
rect 7654 16030 9196 16082
rect 9248 16030 9292 16082
rect 7396 16010 9292 16030
rect 7396 15958 7402 16010
rect 7454 15958 7469 16010
rect 7521 15958 7536 16010
rect 7588 15958 7602 16010
rect 7654 15958 9196 16010
rect 9248 15958 9292 16010
rect 7396 15957 9292 15958
rect 1584 15457 1590 15509
rect 1642 15457 1654 15509
rect 1706 15457 1712 15509
tri 1608 15423 1642 15457 ne
tri 1620 15017 1642 15039 se
rect 1642 15017 1694 15457
tri 1694 15439 1712 15457 nw
tri 1613 15010 1620 15017 se
rect 1620 15010 1687 15017
tri 1687 15010 1694 15017 nw
tri 1561 14958 1613 15010 se
tri 1539 14821 1561 14843 se
rect 1561 14821 1613 14958
tri 1613 14936 1687 15010 nw
tri 1515 14797 1539 14821 se
rect 1539 14797 1589 14821
tri 1589 14797 1613 14821 nw
tri 1463 14745 1515 14797 se
rect 1463 11292 1515 14745
tri 1515 14723 1589 14797 nw
rect 11002 13900 11276 13930
rect 5816 13865 5868 13871
rect 11002 13844 11011 13900
rect 11067 13844 11111 13900
rect 11167 13844 11211 13900
rect 11267 13844 11276 13900
rect 11002 13814 11276 13844
rect 5816 13801 5868 13813
rect 5816 13562 5868 13749
rect 9470 13574 9536 13580
rect 5816 13498 5868 13510
rect 5816 12910 5868 13446
tri 5812 12846 5816 12850 se
rect 5816 12846 5868 12858
tri 5760 12794 5812 12846 se
rect 5812 12794 5816 12846
tri 5754 12788 5760 12794 se
rect 5760 12788 5868 12794
rect 6025 13554 6077 13560
rect 6025 13490 6077 13502
tri 5742 12776 5754 12788 se
rect 5754 12776 5816 12788
tri 5816 12776 5828 12788 nw
tri 5705 12739 5742 12776 se
rect 5742 12739 5779 12776
tri 5779 12739 5816 12776 nw
rect 4715 12272 5215 12278
rect 4767 12220 5163 12272
rect 4715 12208 5215 12220
rect 4767 12156 5163 12208
rect 4715 12150 5215 12156
rect 5705 11904 5757 12739
tri 5757 12717 5779 12739 nw
rect 5705 11834 5757 11852
rect 5705 11764 5757 11782
rect 5705 11694 5757 11712
rect 2839 11610 2845 11662
rect 2897 11610 2909 11662
rect 2961 11610 2967 11662
tri 2839 11579 2870 11610 ne
rect 2870 11572 2929 11610
tri 2929 11572 2967 11610 nw
rect 5705 11624 5757 11642
tri 1463 11256 1499 11292 ne
rect 1499 11256 1515 11292
tri 1515 11256 1573 11314 sw
tri 1499 11240 1515 11256 ne
rect 1515 11240 1573 11256
tri 1515 11182 1573 11240 ne
tri 1573 11182 1647 11256 sw
tri 1573 11160 1595 11182 ne
rect 1595 10792 1647 11182
tri 1595 10770 1617 10792 ne
rect 1617 10770 1647 10792
tri 1647 10770 1691 10814 sw
tri 1617 10748 1639 10770 ne
rect 266 9413 562 9414
rect 266 9361 272 9413
rect 324 9361 348 9413
rect 400 9361 424 9413
rect 476 9361 500 9413
rect 552 9361 562 9413
rect 266 9339 562 9361
rect 266 9287 272 9339
rect 324 9287 348 9339
rect 400 9287 424 9339
rect 476 9287 500 9339
rect 552 9287 562 9339
rect 266 9265 562 9287
tri 238 9213 266 9241 se
rect 266 9213 272 9265
rect 324 9213 348 9265
rect 400 9213 424 9265
rect 476 9213 500 9265
rect 552 9213 562 9265
tri 232 9207 238 9213 se
rect 238 9207 562 9213
tri 227 9202 232 9207 se
rect 232 9202 562 9207
tri 216 9191 227 9202 se
rect 227 9191 562 9202
tri 164 9139 216 9191 se
rect 216 9139 272 9191
rect 324 9139 348 9191
rect 400 9139 424 9191
rect 476 9139 500 9191
rect 552 9139 562 9191
tri 163 9138 164 9139 se
rect 164 9138 562 9139
tri 158 9133 163 9138 se
rect 163 9133 557 9138
tri 557 9133 562 9138 nw
tri 141 9116 158 9133 se
rect 158 9116 540 9133
tri 540 9116 557 9133 nw
tri 139 9114 141 9116 se
rect 141 9114 535 9116
tri 87 9062 139 9114 se
rect 139 9062 277 9114
rect 329 9111 535 9114
tri 535 9111 540 9116 nw
rect 329 9062 483 9111
tri 84 9059 87 9062 se
rect 87 9059 483 9062
tri 483 9059 535 9111 nw
tri 75 9050 84 9059 se
rect 84 9050 444 9059
tri 67 9042 75 9050 se
rect 75 9042 277 9050
rect 67 8998 277 9042
rect 329 9020 444 9050
tri 444 9020 483 9059 nw
rect 329 8998 392 9020
rect 67 8985 392 8998
rect 67 8933 277 8985
rect 329 8968 392 8985
tri 392 8968 444 9020 nw
rect 1444 8968 1450 9020
rect 1502 8968 1514 9020
rect 1566 8968 1572 9020
rect 329 8933 354 8968
rect 67 8930 354 8933
tri 354 8930 392 8968 nw
tri 1444 8930 1482 8968 ne
rect 67 8927 351 8930
tri 351 8927 354 8930 nw
rect 67 7323 219 8927
tri 219 8795 351 8927 nw
rect 1193 8719 1245 8725
rect 1193 8655 1245 8667
tri 1444 8675 1482 8713 se
rect 1482 8675 1534 8968
tri 1534 8930 1572 8968 nw
rect 1639 8815 1691 10770
rect 2225 9999 2231 10051
rect 2283 10044 2299 10051
rect 2351 10044 2367 10051
rect 2419 10044 2435 10051
rect 2290 9999 2299 10044
rect 2419 9999 2431 10044
rect 2487 9999 2503 10051
rect 2555 10044 2571 10051
rect 2623 10044 2638 10051
rect 2623 9999 2627 10044
rect 2690 9999 2696 10051
rect 2225 9988 2234 9999
rect 2290 9988 2333 9999
rect 2389 9988 2431 9999
rect 2487 9988 2529 9999
rect 2585 9988 2627 9999
rect 2683 9988 2696 9999
rect 2225 9977 2696 9988
rect 2225 9925 2231 9977
rect 2283 9950 2299 9977
rect 2351 9950 2367 9977
rect 2419 9950 2435 9977
rect 2290 9925 2299 9950
rect 2419 9925 2431 9950
rect 2487 9925 2503 9977
rect 2555 9950 2571 9977
rect 2623 9950 2638 9977
rect 2623 9925 2627 9950
rect 2690 9925 2696 9977
rect 2225 9903 2234 9925
rect 2290 9903 2333 9925
rect 2389 9903 2431 9925
rect 2487 9903 2529 9925
rect 2585 9903 2627 9925
rect 2683 9903 2696 9925
rect 2225 9851 2231 9903
rect 2290 9894 2299 9903
rect 2419 9894 2431 9903
rect 2283 9856 2299 9894
rect 2351 9856 2367 9894
rect 2419 9856 2435 9894
rect 2290 9851 2299 9856
rect 2419 9851 2431 9856
rect 2487 9851 2503 9903
rect 2623 9894 2627 9903
rect 2555 9856 2571 9894
rect 2623 9856 2638 9894
rect 2623 9851 2627 9856
rect 2690 9851 2696 9903
rect 2225 9829 2234 9851
rect 2290 9829 2333 9851
rect 2389 9829 2431 9851
rect 2487 9829 2529 9851
rect 2585 9829 2627 9851
rect 2683 9829 2696 9851
rect 2225 9777 2231 9829
rect 2290 9800 2299 9829
rect 2419 9800 2431 9829
rect 2283 9777 2299 9800
rect 2351 9777 2367 9800
rect 2419 9777 2435 9800
rect 2487 9777 2503 9829
rect 2623 9800 2627 9829
rect 2555 9777 2571 9800
rect 2623 9777 2638 9800
rect 2690 9777 2696 9829
rect 2225 9762 2696 9777
rect 2225 9755 2234 9762
rect 2290 9755 2333 9762
rect 2389 9755 2431 9762
rect 2487 9755 2529 9762
rect 2585 9755 2627 9762
rect 2683 9755 2696 9762
rect 2225 9703 2231 9755
rect 2290 9706 2299 9755
rect 2419 9706 2431 9755
rect 2283 9703 2299 9706
rect 2351 9703 2367 9706
rect 2419 9703 2435 9706
rect 2487 9703 2503 9755
rect 2623 9706 2627 9755
rect 2555 9703 2571 9706
rect 2623 9703 2638 9706
rect 2690 9703 2696 9755
tri 2848 9715 2870 9737 se
rect 2870 9715 2922 11572
tri 2922 11565 2929 11572 nw
rect 5705 11553 5757 11572
rect 6025 11630 6077 13438
rect 9470 13522 9477 13574
rect 9529 13522 9536 13574
rect 9470 13510 9536 13522
rect 9470 13458 9477 13510
rect 9529 13458 9536 13510
rect 9346 13077 9411 13086
rect 9402 13059 9411 13077
rect 9346 13007 9359 13021
rect 9346 12997 9411 13007
rect 9402 12995 9411 12997
rect 7533 12945 7585 12951
rect 9402 12941 9411 12943
rect 9346 12932 9411 12941
rect 9470 13080 9536 13458
rect 9470 13024 9475 13080
rect 9531 13024 9536 13080
rect 9470 13000 9536 13024
rect 9470 12944 9475 13000
rect 9531 12944 9536 13000
rect 9470 12935 9536 12944
rect 7533 12881 7585 12893
rect 7533 11755 7585 12829
rect 8023 11840 8079 11849
tri 8020 11777 8023 11780 se
rect 8023 11777 8079 11784
tri 7533 11747 7541 11755 ne
rect 7541 11747 7585 11755
tri 7585 11747 7615 11777 sw
tri 7990 11747 8020 11777 se
rect 8020 11760 8079 11777
rect 8020 11747 8023 11760
tri 7541 11703 7585 11747 ne
rect 7585 11703 7663 11747
tri 7585 11695 7593 11703 ne
rect 7593 11695 7663 11703
rect 7715 11695 7727 11747
rect 7779 11695 7785 11747
rect 7946 11695 7952 11747
rect 8004 11695 8016 11747
rect 8068 11695 8079 11704
tri 6077 11630 6096 11649 sw
rect 6025 11627 6096 11630
tri 6025 11556 6096 11627 ne
tri 6096 11595 6131 11630 sw
rect 6096 11556 6131 11595
tri 6131 11556 6170 11595 sw
tri 6665 11556 6704 11595 se
rect 6704 11586 6760 11595
rect 4616 11472 4625 11528
rect 4681 11472 4715 11528
rect 4771 11501 4876 11528
tri 4876 11501 4903 11528 sw
tri 6096 11504 6148 11556 ne
rect 6148 11530 6704 11556
rect 6148 11506 6760 11530
rect 6148 11504 6704 11506
rect 4771 11491 4903 11501
tri 4903 11491 4913 11501 sw
rect 4771 11482 4913 11491
tri 4913 11482 4922 11491 sw
rect 5705 11482 5757 11501
rect 4771 11472 4922 11482
tri 4854 11430 4896 11472 ne
rect 4896 11430 4922 11472
tri 4922 11430 4974 11482 sw
tri 6641 11441 6704 11504 ne
rect 6704 11441 6760 11450
tri 4896 11413 4913 11430 ne
rect 4913 11424 4974 11430
tri 4974 11424 4980 11430 sw
rect 5705 11424 5757 11430
rect 4913 11413 4980 11424
tri 4980 11413 4991 11424 sw
tri 4913 11391 4935 11413 ne
rect 4935 10651 4991 11413
tri 4935 10598 4988 10651 ne
rect 4988 10640 4991 10651
tri 4991 10640 5024 10673 sw
rect 4988 10622 5024 10640
tri 5024 10622 5042 10640 sw
tri 15365 10622 15383 10640 se
rect 15383 10622 15423 19243
tri 15423 19239 15429 19245 nw
rect 4988 10601 5042 10622
tri 5042 10601 5063 10622 sw
tri 15344 10601 15365 10622 se
rect 15365 10601 15402 10622
tri 15402 10601 15423 10622 nw
rect 4988 10598 5063 10601
tri 5063 10598 5066 10601 sw
tri 15341 10598 15344 10601 se
tri 4988 10595 4991 10598 ne
rect 4991 10595 5066 10598
tri 4991 10520 5066 10595 ne
tri 5066 10543 5121 10598 sw
tri 15286 10543 15341 10598 se
rect 15341 10543 15344 10598
tri 15344 10543 15402 10601 nw
rect 5066 10520 5121 10543
tri 5121 10520 5144 10543 sw
tri 15263 10520 15286 10543 se
tri 5066 10442 5144 10520 ne
tri 5144 10442 5222 10520 sw
tri 15246 10503 15263 10520 se
rect 15263 10503 15286 10520
tri 5144 10398 5188 10442 ne
rect 5188 10398 5947 10442
tri 5947 10398 5991 10442 sw
rect 2990 10342 2999 10398
rect 3055 10385 3088 10398
rect 3144 10385 3177 10398
rect 3233 10385 3265 10398
rect 3321 10385 3353 10398
rect 3409 10385 3441 10398
rect 3497 10385 3529 10398
rect 3585 10385 3617 10398
rect 3673 10385 3705 10398
rect 3055 10342 3065 10385
rect 2990 10333 3000 10342
rect 3052 10333 3065 10342
rect 3117 10333 3130 10342
rect 3182 10333 3194 10342
rect 3246 10333 3258 10385
rect 3321 10342 3322 10385
rect 3438 10342 3441 10385
rect 3310 10333 3322 10342
rect 3374 10333 3386 10342
rect 3438 10333 3450 10342
rect 3502 10333 3514 10385
rect 3694 10342 3705 10385
rect 3761 10342 3770 10398
tri 5188 10390 5196 10398 ne
rect 5196 10390 5991 10398
tri 5991 10390 5999 10398 sw
tri 5196 10386 5200 10390 ne
rect 5200 10386 5999 10390
rect 3566 10333 3578 10342
rect 3630 10333 3642 10342
rect 3694 10333 3706 10342
rect 3758 10333 3770 10342
tri 5925 10333 5978 10386 ne
rect 5978 10333 5999 10386
tri 5999 10333 6056 10390 sw
rect 2990 10318 3770 10333
rect 2990 10262 2999 10318
rect 3055 10309 3088 10318
rect 3144 10309 3177 10318
rect 3233 10309 3265 10318
rect 3321 10309 3353 10318
rect 3409 10309 3441 10318
rect 3497 10309 3529 10318
rect 3585 10309 3617 10318
rect 3673 10309 3705 10318
rect 3055 10262 3065 10309
rect 2990 10257 3000 10262
rect 3052 10257 3065 10262
rect 3117 10257 3130 10262
rect 3182 10257 3194 10262
rect 3246 10257 3258 10309
rect 3321 10262 3322 10309
rect 3438 10262 3441 10309
rect 3310 10257 3322 10262
rect 3374 10257 3386 10262
rect 3438 10257 3450 10262
rect 3502 10257 3514 10309
rect 3694 10262 3705 10309
rect 3761 10262 3770 10318
tri 5978 10312 5999 10333 ne
rect 5999 10312 6056 10333
tri 6056 10312 6077 10333 sw
tri 5999 10286 6025 10312 ne
rect 3566 10257 3578 10262
rect 3630 10257 3642 10262
rect 3694 10257 3706 10262
rect 3758 10257 3770 10262
rect 3987 10079 3993 10131
rect 4045 10079 4057 10131
rect 4109 10079 4115 10131
rect 4540 10079 4546 10131
rect 4598 10079 4610 10131
rect 4662 10079 4668 10131
tri 2844 9711 2848 9715 se
rect 2848 9711 2918 9715
tri 2918 9711 2922 9715 nw
tri 2836 9703 2844 9711 se
rect 2844 9703 2910 9711
tri 2910 9703 2918 9711 nw
tri 2770 9637 2836 9703 se
rect 2836 9637 2844 9703
tri 2844 9637 2910 9703 nw
tri 2768 9635 2770 9637 se
rect 2770 9635 2842 9637
tri 2842 9635 2844 9637 nw
tri 2748 9615 2768 9635 se
rect 2768 9615 2790 9635
tri 2356 9583 2388 9615 se
rect 2388 9583 2790 9615
tri 2790 9583 2842 9635 nw
tri 2336 9563 2356 9583 se
rect 2356 9563 2770 9583
tri 2770 9563 2790 9583 nw
tri 2316 9543 2336 9563 se
rect 2336 9543 2390 9563
tri 2390 9543 2410 9563 nw
tri 2302 9529 2316 9543 se
rect 2316 9529 2376 9543
tri 2376 9529 2390 9543 nw
tri 2264 9491 2302 9529 se
rect 2302 9491 2338 9529
tri 2338 9491 2376 9529 nw
tri 2250 9477 2264 9491 se
rect 2264 9477 2314 9491
rect 2250 9467 2314 9477
tri 2314 9467 2338 9491 nw
tri 1639 8814 1640 8815 ne
rect 1640 8814 1691 8815
tri 1691 8814 1714 8837 sw
tri 1640 8763 1691 8814 ne
rect 1691 8763 1714 8814
tri 1691 8740 1714 8763 ne
tri 1714 8759 1769 8814 sw
rect 2250 8767 2302 9467
tri 2302 9455 2314 9467 nw
rect 2778 9259 2789 9260
rect 2845 9259 2921 9260
rect 2977 9259 3053 9260
rect 3109 9259 3185 9260
rect 3241 9259 3317 9260
rect 3373 9259 3449 9260
rect 3505 9259 3581 9260
rect 3637 9259 3713 9260
rect 3769 9259 3778 9260
rect 2778 9207 2784 9259
rect 2845 9207 2851 9259
rect 2903 9207 2918 9259
rect 2977 9207 2985 9259
rect 3037 9207 3052 9259
rect 3109 9207 3119 9259
rect 3171 9207 3185 9259
rect 3241 9207 3253 9259
rect 3305 9207 3317 9259
rect 3373 9207 3387 9259
rect 3439 9207 3449 9259
rect 3506 9207 3521 9259
rect 3573 9207 3581 9259
rect 3640 9207 3654 9259
rect 3706 9207 3713 9259
rect 3772 9207 3778 9259
rect 2778 9204 2789 9207
rect 2845 9204 2921 9207
rect 2977 9204 3053 9207
rect 3109 9204 3185 9207
rect 3241 9204 3317 9207
rect 3373 9204 3449 9207
rect 3505 9204 3581 9207
rect 3637 9204 3713 9207
rect 3769 9204 3778 9207
rect 2778 9185 3778 9204
rect 2778 9133 2784 9185
rect 2836 9133 2851 9185
rect 2903 9133 2918 9185
rect 2970 9133 2985 9185
rect 3037 9133 3052 9185
rect 3104 9133 3119 9185
rect 3171 9133 3186 9185
rect 3238 9133 3253 9185
rect 3305 9133 3320 9185
rect 3372 9133 3387 9185
rect 3439 9133 3454 9185
rect 3506 9133 3521 9185
rect 3573 9133 3588 9185
rect 3640 9133 3654 9185
rect 3706 9133 3720 9185
rect 3772 9133 3778 9185
rect 2778 9120 3778 9133
rect 2778 9111 2789 9120
rect 2845 9111 2921 9120
rect 2977 9111 3053 9120
rect 3109 9111 3185 9120
rect 3241 9111 3317 9120
rect 3373 9111 3449 9120
rect 3505 9111 3581 9120
rect 3637 9111 3713 9120
rect 3769 9111 3778 9120
rect 2778 9059 2784 9111
rect 2845 9064 2851 9111
rect 2836 9059 2851 9064
rect 2903 9059 2918 9111
rect 2977 9064 2985 9111
rect 2970 9059 2985 9064
rect 3037 9059 3052 9111
rect 3109 9064 3119 9111
rect 3104 9059 3119 9064
rect 3171 9064 3185 9111
rect 3241 9064 3253 9111
rect 3171 9059 3186 9064
rect 3238 9059 3253 9064
rect 3305 9064 3317 9111
rect 3373 9064 3387 9111
rect 3305 9059 3320 9064
rect 3372 9059 3387 9064
rect 3439 9064 3449 9111
rect 3439 9059 3454 9064
rect 3506 9059 3521 9111
rect 3573 9064 3581 9111
rect 3573 9059 3588 9064
rect 3640 9059 3654 9111
rect 3706 9064 3713 9111
rect 3706 9059 3720 9064
rect 3772 9059 3778 9111
rect 2778 9058 3778 9059
tri 2250 8759 2258 8767 ne
rect 2258 8759 2302 8767
tri 2302 8759 2332 8789 sw
rect 1714 8740 1769 8759
tri 1769 8740 1788 8759 sw
tri 2258 8740 2277 8759 ne
rect 2277 8740 2332 8759
tri 1714 8713 1741 8740 ne
rect 1741 8715 1788 8740
tri 1788 8715 1813 8740 sw
tri 2277 8715 2302 8740 ne
rect 2302 8715 2332 8740
rect 1741 8713 1813 8715
tri 1813 8713 1815 8715 sw
tri 2302 8713 2304 8715 ne
rect 2304 8713 2332 8715
tri 2332 8713 2378 8759 sw
tri 1534 8675 1572 8713 sw
rect 1444 8623 1450 8675
rect 1502 8623 1514 8675
rect 1566 8623 1572 8675
tri 1741 8666 1788 8713 ne
rect 1788 8685 1815 8713
tri 1815 8685 1843 8713 sw
tri 2304 8685 2332 8713 ne
rect 2332 8685 2378 8713
tri 2378 8685 2406 8713 sw
rect 1788 8666 1843 8685
tri 1843 8666 1862 8685 sw
tri 2332 8666 2351 8685 ne
rect 2351 8666 2406 8685
tri 1788 8623 1831 8666 ne
rect 1831 8623 1862 8666
tri 1862 8623 1905 8666 sw
tri 2351 8623 2394 8666 ne
rect 2394 8623 2406 8666
tri 2406 8623 2468 8685 sw
rect 1193 8597 1245 8603
tri 1193 8595 1195 8597 ne
rect 1195 7884 1241 8597
tri 1241 8593 1245 8597 nw
tri 1831 8593 1861 8623 ne
rect 1861 8611 1905 8623
tri 1905 8611 1917 8623 sw
tri 2394 8611 2406 8623 ne
rect 2406 8611 2468 8623
tri 2468 8611 2480 8623 sw
rect 1861 8593 1917 8611
tri 1861 8592 1862 8593 ne
rect 1862 8592 1917 8593
tri 1917 8592 1936 8611 sw
tri 2406 8592 2425 8611 ne
rect 2425 8592 2480 8611
tri 1862 8591 1863 8592 ne
rect 1863 8591 1936 8592
tri 1936 8591 1937 8592 sw
tri 2425 8591 2426 8592 ne
rect 2426 8591 2480 8592
tri 2480 8591 2500 8611 sw
tri 1863 8585 1869 8591 ne
rect 1869 8585 1937 8591
tri 1937 8585 1943 8591 sw
tri 2426 8585 2432 8591 ne
rect 2432 8585 2500 8591
tri 2500 8585 2506 8591 sw
tri 1869 8533 1921 8585 ne
rect 1921 8537 1943 8585
tri 1943 8537 1991 8585 sw
tri 2432 8537 2480 8585 ne
rect 2480 8537 2506 8585
tri 2506 8537 2554 8585 sw
rect 1921 8533 1991 8537
tri 1991 8533 1995 8537 sw
tri 2480 8533 2484 8537 ne
rect 2484 8533 2554 8537
tri 2554 8533 2558 8537 sw
tri 1921 8521 1933 8533 ne
rect 1933 8521 1995 8533
tri 1995 8521 2007 8533 sw
tri 2484 8521 2496 8533 ne
rect 2496 8521 2558 8533
tri 2558 8521 2570 8533 sw
tri 1933 8518 1936 8521 ne
rect 1936 8518 2007 8521
tri 2007 8518 2010 8521 sw
tri 2496 8518 2499 8521 ne
rect 2499 8518 2570 8521
tri 1936 8469 1985 8518 ne
rect 1985 8469 2010 8518
tri 2010 8469 2059 8518 sw
tri 2499 8469 2548 8518 ne
rect 2548 8469 2570 8518
tri 2570 8469 2622 8521 sw
tri 1985 8444 2010 8469 ne
rect 2010 8463 2059 8469
tri 2059 8463 2065 8469 sw
tri 2548 8463 2554 8469 ne
rect 2554 8463 2622 8469
tri 2622 8463 2628 8469 sw
rect 2010 8444 2065 8463
tri 2065 8444 2084 8463 sw
tri 2554 8444 2573 8463 ne
rect 2573 8444 2628 8463
tri 2010 8370 2084 8444 ne
tri 2084 8389 2139 8444 sw
tri 2573 8389 2628 8444 ne
tri 2628 8389 2702 8463 sw
rect 2084 8370 2139 8389
tri 2139 8370 2158 8389 sw
tri 2628 8370 2647 8389 ne
rect 2647 8370 2702 8389
tri 2084 8350 2104 8370 ne
rect 2104 8350 2158 8370
tri 2158 8350 2178 8370 sw
tri 2647 8350 2667 8370 ne
rect 2667 8350 2702 8370
tri 2702 8350 2741 8389 sw
tri 2104 8349 2105 8350 ne
rect 2105 8349 2178 8350
tri 2178 8349 2179 8350 sw
tri 2667 8349 2668 8350 ne
rect 2668 8349 2741 8350
tri 2741 8349 2742 8350 sw
tri 2105 8297 2157 8349 ne
rect 2157 8315 2179 8349
tri 2179 8315 2213 8349 sw
tri 2668 8315 2702 8349 ne
rect 2702 8315 2742 8349
tri 2742 8315 2776 8349 sw
rect 2157 8297 2213 8315
tri 2213 8297 2231 8315 sw
tri 2702 8297 2720 8315 ne
rect 2720 8297 2776 8315
tri 2157 8296 2158 8297 ne
rect 2158 8296 2231 8297
tri 2231 8296 2232 8297 sw
tri 2720 8296 2721 8297 ne
rect 2721 8296 2776 8297
tri 2158 8272 2182 8296 ne
rect 2182 8293 2232 8296
tri 2232 8293 2235 8296 sw
tri 2721 8293 2724 8296 ne
rect 2182 8272 2235 8293
tri 2235 8272 2256 8293 sw
tri 2182 8269 2185 8272 ne
rect 2185 8269 2256 8272
tri 2256 8269 2259 8272 sw
tri 2185 8222 2232 8269 ne
rect 2232 8222 2259 8269
tri 2259 8222 2306 8269 sw
tri 2232 8217 2237 8222 ne
rect 2237 8217 2306 8222
tri 2306 8217 2311 8222 sw
tri 2237 8191 2263 8217 ne
rect 2263 8191 2311 8217
tri 2311 8191 2337 8217 sw
tri 2263 8148 2306 8191 ne
rect 2306 8148 2337 8191
tri 2337 8148 2380 8191 sw
tri 2306 8139 2315 8148 ne
rect 2315 8139 2380 8148
tri 2380 8139 2389 8148 sw
tri 2315 8086 2368 8139 ne
rect 2368 8086 2389 8139
tri 2389 8086 2442 8139 sw
rect 2724 8086 2776 8296
rect 2839 8217 2845 8269
rect 2897 8232 2913 8269
rect 2906 8217 2913 8232
rect 2965 8232 2981 8269
rect 2965 8217 2974 8232
rect 3033 8217 3049 8269
rect 3101 8232 3117 8269
rect 3169 8217 3184 8269
rect 3236 8232 3251 8269
rect 3303 8217 3318 8269
rect 3370 8232 3385 8269
rect 3437 8217 3452 8269
rect 3504 8232 3519 8269
rect 3571 8217 3586 8269
rect 3638 8232 3653 8269
rect 3646 8217 3653 8232
rect 3705 8232 3720 8269
rect 3705 8217 3713 8232
rect 3772 8217 3778 8269
rect 2839 8191 2850 8217
rect 2906 8191 2974 8217
rect 3030 8191 3098 8217
rect 3154 8191 3221 8217
rect 3277 8191 3344 8217
rect 3400 8191 3467 8217
rect 3523 8191 3590 8217
rect 3646 8191 3713 8217
rect 3769 8191 3778 8217
rect 2839 8139 2845 8191
rect 2906 8176 2913 8191
rect 2897 8139 2913 8176
rect 2965 8176 2974 8191
rect 2965 8139 2981 8176
rect 3033 8139 3049 8191
rect 3101 8139 3117 8176
rect 3169 8139 3184 8191
rect 3236 8139 3251 8176
rect 3303 8139 3318 8191
rect 3370 8139 3385 8176
rect 3437 8139 3452 8191
rect 3504 8139 3519 8176
rect 3571 8139 3586 8191
rect 3646 8176 3653 8191
rect 3638 8139 3653 8176
rect 3705 8176 3713 8191
rect 3705 8139 3720 8176
rect 3772 8139 3778 8191
tri 2776 8086 2798 8108 sw
rect 1535 8077 2133 8086
rect 1535 8021 1536 8077
rect 1592 8021 1626 8077
rect 1682 8021 1716 8077
rect 1772 8021 1806 8077
rect 1862 8021 1896 8077
rect 1952 8021 1986 8077
rect 2042 8021 2076 8077
rect 2132 8021 2133 8077
tri 2368 8074 2380 8086 ne
rect 2380 8074 2442 8086
tri 2442 8074 2454 8086 sw
tri 2724 8074 2736 8086 ne
rect 2736 8074 2798 8086
rect 1535 7993 2133 8021
tri 2380 8000 2454 8074 ne
tri 2454 8058 2470 8074 sw
tri 2736 8058 2752 8074 ne
rect 2752 8058 2798 8074
tri 2798 8058 2826 8086 sw
rect 2454 8034 2470 8058
tri 2470 8034 2494 8058 sw
tri 2752 8034 2776 8058 ne
rect 2776 8034 2826 8058
rect 2454 8000 2494 8034
tri 2494 8000 2528 8034 sw
tri 2776 8000 2810 8034 ne
rect 2810 8000 2826 8034
rect 1535 7937 1536 7993
rect 1592 7937 1626 7993
rect 1682 7937 1716 7993
rect 1772 7937 1806 7993
rect 1862 7937 1896 7993
rect 1952 7937 1986 7993
rect 2042 7937 2076 7993
rect 2132 7937 2133 7993
rect 1535 7909 2133 7937
tri 2454 7926 2528 8000 ne
tri 2528 7984 2544 8000 sw
tri 2810 7984 2826 8000 ne
tri 2826 7984 2900 8058 sw
rect 2528 7945 2544 7984
tri 2544 7945 2583 7984 sw
tri 2826 7945 2865 7984 ne
rect 2865 7945 3084 7984
tri 3084 7945 3123 7984 sw
rect 2528 7932 2583 7945
tri 2583 7932 2596 7945 sw
tri 2865 7932 2878 7945 ne
rect 2878 7932 3123 7945
rect 2528 7926 2596 7932
tri 2596 7926 2602 7932 sw
tri 3062 7926 3068 7932 ne
rect 3068 7926 3123 7932
tri 1195 7850 1229 7884 ne
rect 1229 7850 1241 7884
tri 1241 7850 1295 7904 sw
rect 1535 7853 1536 7909
rect 1592 7853 1626 7909
rect 1682 7853 1716 7909
rect 1772 7853 1806 7909
rect 1862 7853 1896 7909
rect 1952 7853 1986 7909
rect 2042 7853 2076 7909
rect 2132 7853 2133 7909
tri 1229 7838 1241 7850 ne
rect 1241 7838 1295 7850
tri 1241 7796 1283 7838 ne
rect 1283 7796 1295 7838
tri 1295 7796 1349 7850 sw
rect 1535 7825 2133 7853
tri 2528 7852 2602 7926 ne
tri 2602 7871 2657 7926 sw
tri 3068 7871 3123 7926 ne
tri 3123 7871 3197 7945 sw
rect 2602 7852 2657 7871
tri 2657 7852 2676 7871 sw
tri 3123 7852 3142 7871 ne
rect 3142 7852 3197 7871
tri 1283 7791 1288 7796 ne
rect 1288 7791 1349 7796
tri 1349 7791 1354 7796 sw
tri 1288 7784 1295 7791 ne
rect 1295 7784 1354 7791
tri 1354 7784 1361 7791 sw
tri 1295 7764 1315 7784 ne
tri 1060 4172 1106 4218 sw
rect 1054 4166 1106 4172
rect 1054 4102 1106 4114
rect 1054 4044 1106 4050
rect 941 2813 997 2822
rect 42 2802 94 2808
rect 42 2738 94 2750
rect 42 2680 94 2686
rect 941 2733 997 2757
tri 923 2652 941 2670 se
rect 941 2652 997 2677
tri 920 2649 923 2652 se
rect 923 2649 994 2652
tri 994 2649 997 2652 nw
tri 918 2647 920 2649 se
rect 920 2647 992 2649
tri 992 2647 994 2649 nw
tri 917 2646 918 2647 se
rect 918 2646 991 2647
tri 991 2646 992 2647 nw
tri 868 2597 917 2646 se
rect 917 2597 939 2646
rect 868 2594 939 2597
tri 939 2594 991 2646 nw
tri 818 2188 868 2238 se
rect 868 2188 920 2594
tri 920 2575 939 2594 nw
tri 805 2175 818 2188 se
rect 818 2175 920 2188
tri 920 2175 933 2188 sw
rect 324 2123 330 2175
rect 382 2123 394 2175
rect 446 2123 452 2175
rect 805 2123 811 2175
rect 863 2123 875 2175
rect 927 2123 933 2175
tri 1250 1840 1315 1905 se
rect 1315 1885 1361 7784
rect 1535 7769 1536 7825
rect 1592 7769 1626 7825
rect 1682 7769 1716 7825
rect 1772 7769 1806 7825
rect 1862 7769 1896 7825
rect 1952 7769 1986 7825
rect 2042 7769 2076 7825
rect 2132 7769 2133 7825
tri 2602 7796 2658 7852 ne
rect 2658 7797 2676 7852
tri 2676 7797 2731 7852 sw
tri 3142 7797 3197 7852 ne
tri 3197 7826 3242 7871 sw
rect 3197 7797 3242 7826
tri 3242 7797 3271 7826 sw
rect 2658 7796 2731 7797
tri 2731 7796 2732 7797 sw
tri 3197 7796 3198 7797 ne
rect 3198 7796 3271 7797
tri 3271 7796 3272 7797 sw
tri 2658 7791 2663 7796 ne
rect 2663 7791 2732 7796
tri 2732 7791 2737 7796 sw
tri 3198 7791 3203 7796 ne
rect 3203 7791 3272 7796
tri 3272 7791 3277 7796 sw
tri 2663 7778 2676 7791 ne
rect 2676 7778 2737 7791
tri 2737 7778 2750 7791 sw
tri 3203 7778 3216 7791 ne
rect 3216 7778 3277 7791
rect 1535 7741 2133 7769
rect 1535 7685 1536 7741
rect 1592 7685 1626 7741
rect 1682 7685 1716 7741
rect 1772 7685 1806 7741
rect 1862 7685 1896 7741
rect 1952 7685 1986 7741
rect 2042 7685 2076 7741
rect 2132 7685 2133 7741
tri 2676 7739 2715 7778 ne
rect 2715 7739 2750 7778
tri 2750 7739 2789 7778 sw
tri 3216 7739 3255 7778 ne
rect 3255 7739 3277 7778
tri 3277 7739 3329 7791 sw
rect 4619 7739 4625 7791
rect 4677 7739 4689 7791
rect 4741 7739 4747 7791
tri 2715 7704 2750 7739 ne
rect 2750 7723 2789 7739
tri 2789 7723 2805 7739 sw
tri 3255 7723 3271 7739 ne
rect 3271 7723 3329 7739
tri 3329 7723 3345 7739 sw
tri 4639 7723 4655 7739 ne
rect 4655 7723 4747 7739
rect 2750 7704 2805 7723
tri 2805 7704 2824 7723 sw
tri 3271 7704 3290 7723 ne
rect 3290 7709 3345 7723
tri 3345 7709 3359 7723 sw
tri 4655 7709 4669 7723 ne
rect 4669 7709 4747 7723
rect 3290 7704 3359 7709
rect 1535 7657 2133 7685
rect 1535 7601 1536 7657
rect 1592 7601 1626 7657
rect 1682 7601 1716 7657
rect 1772 7601 1806 7657
rect 1862 7601 1896 7657
rect 1952 7601 1986 7657
rect 2042 7601 2076 7657
rect 2132 7601 2133 7657
tri 2750 7630 2824 7704 ne
tri 2824 7649 2879 7704 sw
tri 3290 7649 3345 7704 ne
rect 3345 7683 3359 7704
tri 3359 7683 3385 7709 sw
tri 4669 7683 4695 7709 ne
rect 3345 7649 3385 7683
tri 3385 7649 3419 7683 sw
rect 2824 7630 2879 7649
tri 2879 7630 2898 7649 sw
tri 3345 7630 3364 7649 ne
rect 3364 7630 3419 7649
rect 1535 7573 2133 7601
rect 1535 7517 1536 7573
rect 1592 7517 1626 7573
rect 1682 7517 1716 7573
rect 1772 7517 1806 7573
rect 1862 7517 1896 7573
rect 1952 7517 1986 7573
rect 2042 7517 2076 7573
rect 2132 7517 2133 7573
tri 2824 7556 2898 7630 ne
tri 2898 7575 2953 7630 sw
tri 3364 7575 3419 7630 ne
tri 3419 7575 3493 7649 sw
rect 2898 7556 2953 7575
tri 2953 7556 2972 7575 sw
tri 3419 7556 3438 7575 ne
rect 3438 7556 3493 7575
rect 1535 7489 2133 7517
rect 1535 7433 1536 7489
rect 1592 7433 1626 7489
rect 1682 7433 1716 7489
rect 1772 7433 1806 7489
rect 1862 7433 1896 7489
rect 1952 7433 1986 7489
rect 2042 7433 2076 7489
rect 2132 7433 2133 7489
tri 2898 7482 2972 7556 ne
tri 2972 7501 3027 7556 sw
tri 3438 7501 3493 7556 ne
tri 3493 7501 3567 7575 sw
rect 2972 7482 3027 7501
tri 3027 7482 3046 7501 sw
tri 2972 7479 2975 7482 ne
rect 2975 7479 3046 7482
tri 3493 7479 3515 7501 ne
tri 2975 7460 2994 7479 ne
rect 1535 7405 2133 7433
rect 1535 7349 1536 7405
rect 1592 7349 1626 7405
rect 1682 7349 1716 7405
rect 1772 7349 1806 7405
rect 1862 7349 1896 7405
rect 1952 7349 1986 7405
rect 2042 7349 2076 7405
rect 2132 7349 2133 7405
rect 1535 7321 2133 7349
rect 1535 7265 1536 7321
rect 1592 7265 1626 7321
rect 1682 7265 1716 7321
rect 1772 7265 1806 7321
rect 1862 7265 1896 7321
rect 1952 7265 1986 7321
rect 2042 7265 2076 7321
rect 2132 7265 2133 7321
rect 1535 7237 2133 7265
rect 1535 7181 1536 7237
rect 1592 7181 1626 7237
rect 1682 7181 1716 7237
rect 1772 7181 1806 7237
rect 1862 7181 1896 7237
rect 1952 7181 1986 7237
rect 2042 7181 2076 7237
rect 2132 7181 2133 7237
rect 1535 7152 2133 7181
rect 1535 7096 1536 7152
rect 1592 7096 1626 7152
rect 1682 7096 1716 7152
rect 1772 7096 1806 7152
rect 1862 7096 1896 7152
rect 1952 7096 1986 7152
rect 2042 7096 2076 7152
rect 2132 7096 2133 7152
rect 1535 7067 2133 7096
rect 1535 7011 1536 7067
rect 1592 7011 1626 7067
rect 1682 7011 1716 7067
rect 1772 7011 1806 7067
rect 1862 7011 1896 7067
rect 1952 7011 1986 7067
rect 2042 7011 2076 7067
rect 2132 7011 2133 7067
rect 1535 6982 2133 7011
rect 1535 6926 1536 6982
rect 1592 6926 1626 6982
rect 1682 6926 1716 6982
rect 1772 6926 1806 6982
rect 1862 6926 1896 6982
rect 1952 6926 1986 6982
rect 2042 6926 2076 6982
rect 2132 6926 2133 6982
rect 1535 6897 2133 6926
rect 1535 6841 1536 6897
rect 1592 6841 1626 6897
rect 1682 6841 1716 6897
rect 1772 6841 1806 6897
rect 1862 6841 1896 6897
rect 1952 6841 1986 6897
rect 2042 6841 2076 6897
rect 2132 6841 2133 6897
rect 1535 6812 2133 6841
rect 1535 6756 1536 6812
rect 1592 6756 1626 6812
rect 1682 6756 1716 6812
rect 1772 6756 1806 6812
rect 1862 6756 1896 6812
rect 1952 6756 1986 6812
rect 2042 6756 2076 6812
rect 2132 6756 2133 6812
rect 1535 6727 2133 6756
rect 1535 6671 1536 6727
rect 1592 6671 1626 6727
rect 1682 6671 1716 6727
rect 1772 6671 1806 6727
rect 1862 6671 1896 6727
rect 1952 6671 1986 6727
rect 2042 6671 2076 6727
rect 2132 6671 2133 6727
rect 1535 6662 2133 6671
rect 1709 6635 2117 6644
rect 1765 6579 1797 6635
rect 1853 6579 1885 6635
rect 1941 6579 1973 6635
rect 2029 6579 2061 6635
rect 1709 6551 2117 6579
rect 1765 6495 1797 6551
rect 1853 6495 1885 6551
rect 1941 6495 1973 6551
rect 2029 6495 2061 6551
rect 1709 6467 2117 6495
rect 1765 6411 1797 6467
rect 1853 6411 1885 6467
rect 1941 6411 1973 6467
rect 2029 6411 2061 6467
rect 1709 6383 2117 6411
rect 1765 6327 1797 6383
rect 1853 6327 1885 6383
rect 1941 6327 1973 6383
rect 2029 6327 2061 6383
rect 2994 6405 3046 7479
tri 3441 7032 3515 7106 se
rect 3515 7084 3567 7501
tri 3515 7032 3567 7084 nw
tri 3367 6958 3441 7032 se
tri 3441 6958 3515 7032 nw
tri 3293 6884 3367 6958 se
tri 3367 6884 3441 6958 nw
tri 3273 6864 3293 6884 se
rect 3293 6864 3347 6884
tri 3347 6864 3367 6884 nw
tri 3046 6405 3055 6414 sw
rect 2994 6392 3055 6405
tri 2994 6356 3030 6392 ne
rect 3030 6356 3055 6392
tri 3055 6356 3104 6405 sw
tri 3030 6331 3055 6356 ne
rect 3055 6331 3104 6356
tri 3104 6331 3129 6356 sw
rect 1709 6299 2117 6327
tri 3055 6309 3077 6331 ne
rect 1765 6243 1797 6299
rect 1853 6243 1885 6299
rect 1941 6243 1973 6299
rect 2029 6243 2061 6299
rect 1709 6215 2117 6243
rect 1765 6159 1797 6215
rect 1853 6159 1885 6215
rect 1941 6159 1973 6215
rect 2029 6159 2061 6215
rect 1709 6131 2117 6159
rect 1765 6075 1797 6131
rect 1853 6075 1885 6131
rect 1941 6075 1973 6131
rect 2029 6075 2061 6131
rect 1709 6046 2117 6075
rect 1765 5990 1797 6046
rect 1853 5990 1885 6046
rect 1941 5990 1973 6046
rect 2029 5990 2061 6046
rect 1709 5961 2117 5990
rect 1765 5905 1797 5961
rect 1853 5905 1885 5961
rect 1941 5905 1973 5961
rect 2029 5905 2061 5961
rect 1709 5896 2117 5905
rect 1708 5836 1976 5845
rect 1764 5780 1814 5836
rect 1870 5780 1920 5836
rect 1708 5754 1976 5780
rect 1764 5698 1814 5754
rect 1870 5698 1920 5754
rect 1708 5672 1976 5698
rect 1764 5616 1814 5672
rect 1870 5616 1920 5672
rect 1708 5590 1976 5616
rect 1764 5534 1814 5590
rect 1870 5534 1920 5590
rect 1708 5508 1976 5534
rect 1764 5452 1814 5508
rect 1870 5452 1920 5508
rect 1708 5426 1976 5452
rect 1764 5370 1814 5426
rect 1870 5370 1920 5426
rect 1708 5343 1976 5370
rect 1764 5287 1814 5343
rect 1870 5287 1920 5343
rect 1708 5278 1976 5287
rect 1709 5228 2117 5237
rect 1765 5172 1797 5228
rect 1853 5172 1885 5228
rect 1941 5172 1973 5228
rect 2029 5172 2061 5228
rect 1709 5148 2117 5172
rect 1765 5092 1797 5148
rect 1853 5092 1885 5148
rect 1941 5092 1973 5148
rect 2029 5092 2061 5148
rect 1709 5068 2117 5092
rect 1765 5012 1797 5068
rect 1853 5012 1885 5068
rect 1941 5012 1973 5068
rect 2029 5012 2061 5068
rect 1709 4988 2117 5012
rect 1765 4932 1797 4988
rect 1853 4932 1885 4988
rect 1941 4932 1973 4988
rect 2029 4932 2061 4988
rect 1709 4908 2117 4932
rect 1765 4852 1797 4908
rect 1853 4852 1885 4908
rect 1941 4852 1973 4908
rect 2029 4852 2061 4908
rect 1709 4828 2117 4852
rect 1765 4772 1797 4828
rect 1853 4772 1885 4828
rect 1941 4772 1973 4828
rect 2029 4772 2061 4828
rect 1709 4747 2117 4772
rect 1765 4691 1797 4747
rect 1853 4691 1885 4747
rect 1941 4691 1973 4747
rect 2029 4691 2061 4747
rect 1709 4666 2117 4691
rect 1765 4610 1797 4666
rect 1853 4610 1885 4666
rect 1941 4610 1973 4666
rect 2029 4610 2061 4666
rect 1709 4585 2117 4610
rect 1765 4529 1797 4585
rect 1853 4529 1885 4585
rect 1941 4529 1973 4585
rect 2029 4529 2061 4585
rect 1709 4504 2117 4529
rect 1765 4448 1797 4504
rect 1853 4448 1885 4504
rect 1941 4448 1973 4504
rect 2029 4448 2061 4504
rect 1709 4423 2117 4448
rect 1765 4367 1797 4423
rect 1853 4367 1885 4423
rect 1941 4367 1973 4423
rect 2029 4367 2061 4423
rect 1709 4342 2117 4367
rect 1765 4286 1797 4342
rect 1853 4286 1885 4342
rect 1941 4286 1973 4342
rect 2029 4286 2061 4342
rect 1709 4261 2117 4286
rect 1765 4205 1797 4261
rect 1853 4205 1885 4261
rect 1941 4205 1973 4261
rect 2029 4205 2061 4261
rect 1709 4180 2117 4205
rect 1765 4124 1797 4180
rect 1853 4124 1885 4180
rect 1941 4124 1973 4180
rect 2029 4124 2061 4180
rect 1451 4071 1457 4123
rect 1509 4071 1521 4123
rect 1573 4071 1633 4123
tri 1506 3996 1581 4071 ne
rect 1581 3791 1633 4071
rect 1709 4099 2117 4124
rect 1765 4043 1797 4099
rect 1853 4043 1885 4099
rect 1941 4043 1973 4099
rect 2029 4043 2061 4099
rect 1709 4018 2117 4043
rect 1765 3962 1797 4018
rect 1853 3962 1885 4018
rect 1941 3962 1973 4018
rect 2029 3962 2061 4018
rect 1709 3937 2117 3962
rect 1765 3881 1797 3937
rect 1853 3881 1885 3937
rect 1941 3881 1973 3937
rect 2029 3881 2061 3937
rect 1709 3872 2117 3881
tri 3021 3872 3077 3928 se
rect 3077 3906 3129 6331
rect 3273 6312 3325 6864
tri 3325 6842 3347 6864 nw
tri 3325 6312 3347 6334 sw
tri 3273 6304 3281 6312 ne
rect 3281 6304 3347 6312
tri 3347 6304 3355 6312 sw
tri 3281 6263 3322 6304 ne
rect 3322 6285 3355 6304
tri 3355 6285 3374 6304 sw
tri 3003 3854 3021 3872 se
rect 3021 3854 3077 3872
tri 3077 3854 3129 3906 nw
tri 2962 3813 3003 3854 se
tri 1581 3770 1602 3791 ne
rect 1602 3770 1633 3791
tri 1633 3770 1676 3813 sw
tri 2929 3780 2962 3813 se
rect 2962 3780 3003 3813
tri 3003 3780 3077 3854 nw
tri 2919 3770 2929 3780 se
tri 1602 3739 1633 3770 ne
rect 1633 3739 2297 3770
tri 1633 3718 1654 3739 ne
rect 1654 3718 2297 3739
tri 2275 3697 2296 3718 ne
rect 2296 3697 2297 3718
tri 2297 3697 2370 3770 sw
tri 2855 3706 2919 3770 se
rect 2919 3706 2929 3770
tri 2929 3706 3003 3780 nw
tri 2296 3696 2297 3697 ne
rect 2297 3696 2370 3697
tri 2297 3675 2318 3696 ne
rect 1960 3622 1966 3674
rect 2018 3622 2030 3674
rect 2082 3622 2088 3674
tri 1996 3582 2036 3622 ne
rect 2036 3526 2088 3622
tri 2036 3511 2051 3526 ne
rect 2051 3511 2088 3526
tri 2088 3511 2125 3548 sw
tri 2051 3474 2088 3511 ne
rect 2088 3474 2125 3511
tri 2088 3437 2125 3474 ne
tri 2125 3437 2199 3511 sw
tri 2125 3415 2147 3437 ne
rect 1315 1840 1316 1885
tri 1316 1840 1361 1885 nw
tri 1249 1839 1250 1840 se
rect 1250 1839 1315 1840
tri 1315 1839 1316 1840 nw
tri 1220 1810 1249 1839 se
rect 1249 1810 1286 1839
tri 1286 1810 1315 1839 nw
tri 1214 1804 1220 1810 se
rect 1220 1804 1280 1810
tri 1280 1804 1286 1810 nw
rect 1497 1804 1625 1840
tri 1183 1773 1214 1804 se
rect 1214 1773 1249 1804
tri 1249 1773 1280 1804 nw
tri 1162 1752 1183 1773 se
rect 1183 1752 1228 1773
tri 1228 1752 1249 1773 nw
rect 1549 1752 1573 1804
tri 1148 1738 1162 1752 se
rect 1162 1738 1214 1752
tri 1214 1738 1228 1752 nw
rect 1497 1738 1625 1752
tri 1117 1707 1148 1738 se
rect 1148 1707 1183 1738
tri 1183 1707 1214 1738 nw
tri 1096 1686 1117 1707 se
rect 1117 1686 1162 1707
tri 1162 1686 1183 1707 nw
rect 1549 1686 1573 1738
tri 1090 1680 1096 1686 se
rect 1096 1680 1156 1686
tri 1156 1680 1162 1686 nw
rect 1497 1680 1625 1686
tri 1080 1670 1090 1680 se
rect 1090 1670 1146 1680
tri 1146 1670 1156 1680 nw
rect 1080 1653 1129 1670
tri 1129 1653 1146 1670 nw
rect 1080 1652 1128 1653
tri 1128 1652 1129 1653 nw
rect 1080 1651 1127 1652
tri 1127 1651 1128 1652 nw
tri 1039 1034 1080 1075 se
rect 1080 1055 1126 1651
tri 1126 1650 1127 1651 nw
rect 1498 1646 1507 1652
rect 1498 1594 1499 1646
rect 1563 1596 1590 1652
rect 1646 1646 1655 1652
rect 1551 1594 1603 1596
rect 1498 1577 1655 1594
rect 1498 1525 1499 1577
rect 1551 1525 1603 1577
rect 1498 1508 1655 1525
rect 1498 1456 1499 1508
rect 1551 1506 1603 1508
rect 1498 1450 1507 1456
rect 1563 1450 1590 1506
rect 1646 1450 1655 1456
rect 1780 1651 1789 1653
rect 1780 1599 1786 1651
rect 1780 1597 1789 1599
rect 1845 1597 1858 1653
rect 1780 1577 1858 1597
rect 1780 1525 1786 1577
rect 1838 1525 1858 1577
rect 1780 1507 1858 1525
rect 1780 1503 1789 1507
rect 1780 1451 1786 1503
rect 1845 1451 1858 1507
rect 1780 1450 1858 1451
rect 1182 1285 1188 1337
rect 1240 1285 1252 1337
rect 1304 1285 1310 1337
tri 1229 1250 1264 1285 ne
rect 1080 1034 1105 1055
tri 1105 1034 1126 1055 nw
tri 1223 1034 1264 1075 se
rect 1264 1055 1310 1285
rect 1264 1034 1289 1055
tri 1289 1034 1310 1055 nw
tri 1031 1026 1039 1034 se
rect 1039 1026 1097 1034
tri 1097 1026 1105 1034 nw
tri 1215 1026 1223 1034 se
rect 1223 1026 1281 1034
tri 1281 1026 1289 1034 nw
tri 1025 1020 1031 1026 se
rect 1031 1020 1091 1026
tri 1091 1020 1097 1026 nw
tri 1209 1020 1215 1026 se
rect 1215 1020 1269 1026
tri 794 1014 800 1020 se
rect 800 1014 1085 1020
tri 1085 1014 1091 1020 nw
tri 1203 1014 1209 1020 se
rect 1209 1014 1269 1020
tri 1269 1014 1281 1026 nw
tri 790 1010 794 1014 se
rect 794 1010 1081 1014
tri 1081 1010 1085 1014 nw
tri 1199 1010 1203 1014 se
rect 1203 1010 1265 1014
tri 1265 1010 1269 1014 nw
tri 789 1009 790 1010 se
rect 790 1009 1080 1010
tri 1080 1009 1081 1010 nw
tri 1198 1009 1199 1010 se
rect 1199 1009 1264 1010
tri 1264 1009 1265 1010 nw
tri 738 958 789 1009 se
rect 789 974 1045 1009
tri 1045 974 1080 1009 nw
tri 1163 974 1198 1009 se
rect 1198 974 1213 1009
rect 789 958 804 974
tri 804 958 820 974 nw
tri 1147 958 1163 974 se
rect 1163 958 1213 974
tri 1213 958 1264 1009 nw
tri 734 954 738 958 se
rect 738 954 800 958
tri 800 954 804 958 nw
tri 1143 954 1147 958 se
rect 1147 954 1198 958
tri 723 943 734 954 se
rect 734 943 789 954
tri 789 943 800 954 nw
tri 1132 943 1143 954 se
rect 1143 943 1198 954
tri 1198 943 1213 958 nw
tri 714 934 723 943 se
rect 723 934 780 943
tri 780 934 789 943 nw
tri 1123 934 1132 943 se
rect 1132 934 1189 943
tri 1189 934 1198 943 nw
tri 675 895 714 934 se
rect 714 895 741 934
tri 741 895 780 934 nw
tri 1084 895 1123 934 se
rect 1123 895 1150 934
tri 1150 895 1189 934 nw
rect 675 882 728 895
tri 728 882 741 895 nw
rect 1084 882 1137 895
tri 1137 882 1150 895 nw
rect 675 878 724 882
tri 724 878 728 882 nw
rect 1084 878 1133 882
tri 1133 878 1137 882 nw
rect 288 330 344 339
rect 288 250 344 274
rect 288 185 344 194
rect 675 0 721 878
tri 721 875 724 878 nw
rect 1084 0 1130 878
tri 1130 875 1133 878 nw
tri 1651 735 1689 773 se
rect 1689 751 1741 1356
rect 2147 1026 2199 3437
tri 2296 3223 2318 3245 se
rect 2318 3223 2370 3696
tri 2823 3674 2855 3706 se
rect 2855 3674 2897 3706
tri 2897 3674 2929 3706 nw
tri 2293 3220 2296 3223 se
rect 2296 3220 2367 3223
tri 2367 3220 2370 3223 nw
tri 2794 3645 2823 3674 se
rect 2823 3645 2868 3674
tri 2868 3645 2897 3674 nw
tri 2292 3219 2293 3220 se
rect 2293 3219 2366 3220
tri 2366 3219 2367 3220 nw
tri 2273 3200 2292 3219 se
rect 2292 3200 2347 3219
tri 2347 3200 2366 3219 nw
tri 2244 3171 2273 3200 se
rect 2273 3171 2296 3200
rect 2244 1208 2296 3171
tri 2296 3149 2347 3200 nw
rect 2440 2646 2761 2647
rect 2440 2594 2446 2646
rect 2498 2594 2511 2646
rect 2563 2594 2575 2646
rect 2627 2594 2639 2646
rect 2691 2594 2703 2646
rect 2755 2594 2761 2646
rect 2440 2574 2761 2594
rect 2440 2522 2446 2574
rect 2498 2522 2511 2574
rect 2563 2522 2575 2574
rect 2627 2522 2639 2574
rect 2691 2522 2703 2574
rect 2755 2522 2761 2574
rect 2440 2502 2761 2522
rect 2440 2450 2446 2502
rect 2498 2450 2511 2502
rect 2563 2450 2575 2502
rect 2627 2450 2639 2502
rect 2691 2450 2703 2502
rect 2755 2450 2761 2502
rect 2440 2449 2761 2450
tri 2720 1239 2794 1313 se
rect 2794 1291 2846 3645
tri 2846 3623 2868 3645 nw
rect 3322 2495 3374 6285
rect 4695 5036 4747 7709
rect 6025 7602 6077 10312
rect 11001 10281 11007 10333
rect 11059 10326 11081 10333
rect 11133 10326 11155 10333
rect 11207 10326 11229 10333
rect 11071 10281 11081 10326
rect 11207 10281 11216 10326
rect 11281 10281 11287 10333
rect 11001 10270 11015 10281
rect 11071 10270 11116 10281
rect 11172 10270 11216 10281
rect 11272 10270 11287 10281
rect 11001 10269 11287 10270
rect 7399 10244 7625 10257
rect 7399 10192 7406 10244
rect 7458 10192 7487 10244
rect 7539 10192 7567 10244
rect 7619 10192 7625 10244
rect 6891 10079 6897 10131
rect 6949 10079 6961 10131
rect 7013 10079 7019 10131
tri 6891 10051 6919 10079 ne
rect 6919 10051 6995 10079
tri 6995 10055 7019 10079 nw
tri 6919 10028 6942 10051 ne
rect 6942 10028 6995 10051
tri 6942 10027 6943 10028 ne
rect 6943 9977 6995 10028
rect 6943 9913 6995 9925
tri 6913 7796 6943 7826 se
rect 6943 7796 6995 9861
rect 7214 9976 7220 10028
rect 7272 9976 7284 10028
rect 7336 9976 7342 10028
tri 6908 7791 6913 7796 se
rect 6913 7791 6995 7796
rect 6867 7739 6873 7791
rect 6925 7739 6937 7791
rect 6989 7739 6995 7791
tri 7181 7796 7214 7829 se
rect 7214 7796 7266 9976
tri 7266 9942 7300 9976 nw
rect 7399 9635 7625 10192
rect 11001 10217 11007 10269
rect 11059 10217 11081 10269
rect 11133 10217 11155 10269
rect 11207 10217 11229 10269
rect 11281 10217 11287 10269
rect 11001 10216 11287 10217
rect 11001 10205 11015 10216
rect 11071 10205 11116 10216
rect 11172 10205 11216 10216
rect 11272 10205 11287 10216
rect 11001 10153 11007 10205
rect 11071 10160 11081 10205
rect 11207 10160 11216 10205
rect 11059 10153 11081 10160
rect 11133 10153 11155 10160
rect 11207 10153 11229 10160
rect 11281 10153 11287 10205
rect 15246 10152 15286 10503
tri 15286 10485 15344 10543 nw
tri 15246 10134 15264 10152 ne
rect 15264 10134 15286 10152
tri 15286 10134 15322 10170 sw
tri 15264 10131 15267 10134 ne
rect 15267 10131 15322 10134
tri 15322 10131 15325 10134 sw
tri 15267 10112 15286 10131 ne
rect 15286 10112 15325 10131
tri 15286 10076 15322 10112 ne
rect 15322 10076 15325 10112
tri 15325 10076 15380 10131 sw
tri 15322 10055 15343 10076 ne
rect 15343 10055 15380 10076
tri 15380 10055 15401 10076 sw
tri 15343 10039 15359 10055 ne
rect 15359 10039 15401 10055
rect 7816 10030 7947 10039
rect 7816 10028 7872 10030
rect 7928 10028 7947 10030
tri 15359 10028 15370 10039 ne
rect 15370 10028 15401 10039
tri 15401 10028 15428 10055 sw
rect 7816 9976 7822 10028
rect 7938 9976 7947 10028
tri 15370 10018 15380 10028 ne
rect 15380 10018 15428 10028
tri 15428 10018 15438 10028 sw
tri 15380 9997 15401 10018 ne
rect 15401 9997 15438 10018
rect 7816 9974 7872 9976
rect 7928 9974 7947 9976
rect 7816 9950 7947 9974
rect 7816 9894 7872 9950
rect 7928 9894 7947 9950
rect 7816 9885 7947 9894
rect 9645 9988 9776 9997
rect 9645 9932 9682 9988
rect 9738 9932 9776 9988
tri 15401 9960 15438 9997 ne
tri 15438 9960 15496 10018 sw
rect 9645 9908 9776 9932
rect 9645 9907 9682 9908
rect 9738 9907 9776 9908
rect 9645 9855 9654 9907
rect 9770 9855 9776 9907
tri 15438 9902 15496 9960 ne
tri 15496 9902 15554 9960 sw
rect 9645 9852 9682 9855
rect 9738 9852 9776 9855
rect 9645 9843 9776 9852
tri 15496 9844 15554 9902 ne
tri 15554 9844 15612 9902 sw
tri 15554 9843 15555 9844 ne
rect 15555 9843 15612 9844
tri 15555 9786 15612 9843 ne
tri 15612 9786 15670 9844 sw
tri 15612 9728 15670 9786 ne
tri 15670 9728 15728 9786 sw
tri 15670 9670 15728 9728 ne
tri 15728 9670 15786 9728 sw
rect 7399 9583 7409 9635
rect 7461 9583 7488 9635
rect 7540 9583 7567 9635
rect 7619 9583 7625 9635
tri 15728 9612 15786 9670 ne
tri 15786 9612 15844 9670 sw
rect 7399 9543 7625 9583
tri 15786 9554 15844 9612 ne
tri 15844 9554 15902 9612 sw
rect 7399 9491 7434 9543
rect 7486 9491 7625 9543
tri 15844 9534 15864 9554 ne
rect 7399 9467 7625 9491
rect 7399 9415 7434 9467
rect 7486 9415 7625 9467
rect 7399 9254 7625 9415
rect 10896 9500 11287 9501
rect 10896 9448 10902 9500
rect 10954 9471 10968 9500
rect 10954 9448 10956 9471
rect 11020 9448 11034 9500
rect 11086 9471 11099 9500
rect 11151 9471 11164 9500
rect 11095 9448 11099 9471
rect 11216 9448 11229 9500
rect 11281 9448 11287 9500
rect 10896 9426 10956 9448
rect 11012 9426 11039 9448
rect 11095 9426 11122 9448
rect 11178 9426 11287 9448
rect 10896 9374 10902 9426
rect 10954 9415 10956 9426
rect 10954 9387 10968 9415
rect 10954 9374 10956 9387
rect 11020 9374 11034 9426
rect 11095 9415 11099 9426
rect 11086 9387 11099 9415
rect 11151 9387 11164 9415
rect 11095 9374 11099 9387
rect 11216 9374 11229 9426
rect 11281 9374 11287 9426
rect 10896 9352 10956 9374
rect 11012 9352 11039 9374
rect 11095 9352 11122 9374
rect 11178 9352 11287 9374
rect 10896 9300 10902 9352
rect 10954 9331 10956 9352
rect 10954 9300 10968 9331
rect 11020 9300 11034 9352
rect 11095 9331 11099 9352
rect 11086 9300 11099 9331
rect 11151 9300 11164 9331
rect 11216 9300 11229 9352
rect 11281 9300 11287 9352
rect 10896 9299 11287 9300
rect 7451 9202 7519 9254
rect 7571 9202 7625 9254
rect 7399 9185 7625 9202
rect 7451 9133 7519 9185
rect 7571 9133 7625 9185
rect 7399 9116 7625 9133
rect 7451 9064 7519 9116
rect 7571 9064 7625 9116
rect 7399 9058 7625 9064
rect 9118 9265 9564 9274
rect 9118 9209 9121 9265
rect 9177 9209 9217 9265
rect 9273 9209 9313 9265
rect 9369 9209 9409 9265
rect 9465 9209 9505 9265
rect 9561 9209 9564 9265
rect 9118 9178 9564 9209
rect 9118 9122 9121 9178
rect 9177 9122 9217 9178
rect 9273 9122 9313 9178
rect 9369 9122 9409 9178
rect 9465 9122 9505 9178
rect 9561 9122 9564 9178
rect 9118 9091 9564 9122
rect 9118 9035 9121 9091
rect 9177 9035 9217 9091
rect 9273 9035 9313 9091
rect 9369 9035 9409 9091
rect 9465 9035 9505 9091
rect 9561 9035 9564 9091
rect 9118 9004 9564 9035
rect 9118 8948 9121 9004
rect 9177 8948 9217 9004
rect 9273 8948 9313 9004
rect 9369 8948 9409 9004
rect 9465 8948 9505 9004
rect 9561 8948 9564 9004
rect 9118 8917 9564 8948
rect 9118 8861 9121 8917
rect 9177 8861 9217 8917
rect 9273 8861 9313 8917
rect 9369 8861 9409 8917
rect 9465 8861 9505 8917
rect 9561 8861 9564 8917
rect 9118 8830 9564 8861
rect 9118 8774 9121 8830
rect 9177 8774 9217 8830
rect 9273 8774 9313 8830
rect 9369 8774 9409 8830
rect 9465 8774 9505 8830
rect 9561 8774 9564 8830
rect 9118 8742 9564 8774
rect 9118 8686 9121 8742
rect 9177 8686 9217 8742
rect 9273 8686 9313 8742
rect 9369 8686 9409 8742
rect 9465 8686 9505 8742
rect 9561 8686 9564 8742
rect 9118 8654 9564 8686
rect 9118 8598 9121 8654
rect 9177 8598 9217 8654
rect 9273 8598 9313 8654
rect 9369 8598 9409 8654
rect 9465 8598 9505 8654
rect 9561 8598 9564 8654
rect 9118 8566 9564 8598
rect 9118 8510 9121 8566
rect 9177 8510 9217 8566
rect 9273 8510 9313 8566
rect 9369 8510 9409 8566
rect 9465 8510 9505 8566
rect 9561 8510 9564 8566
rect 9118 8478 9564 8510
rect 9118 8422 9121 8478
rect 9177 8422 9217 8478
rect 9273 8422 9313 8478
rect 9369 8422 9409 8478
rect 9465 8422 9505 8478
rect 9561 8422 9564 8478
rect 9118 8390 9564 8422
rect 9118 8334 9121 8390
rect 9177 8334 9217 8390
rect 9273 8334 9313 8390
rect 9369 8334 9409 8390
rect 9465 8334 9505 8390
rect 9561 8334 9564 8390
rect 15783 8585 15835 8591
rect 15783 8521 15835 8533
rect 9118 8325 9564 8334
rect 9782 8297 9788 8349
rect 9840 8297 9852 8349
rect 9904 8297 9910 8349
rect 11591 8297 11597 8349
rect 11649 8297 11661 8349
rect 11713 8297 11719 8349
rect 9782 8272 9863 8297
tri 9863 8272 9888 8297 nw
tri 11591 8272 11616 8297 ne
rect 11616 8272 11694 8297
tri 11694 8272 11719 8297 nw
rect 13568 8313 13820 8350
rect 13872 8313 13892 8350
rect 13944 8313 13964 8350
rect 14016 8313 14036 8350
rect 9782 8269 9860 8272
tri 9860 8269 9863 8272 nw
tri 11616 8269 11619 8272 ne
rect 11619 8269 11681 8272
rect 9782 8259 9850 8269
tri 9850 8259 9860 8269 nw
tri 9768 8139 9782 8153 se
rect 9782 8139 9834 8259
tri 9834 8243 9850 8259 nw
rect 10496 8217 10502 8269
rect 10554 8235 10591 8269
rect 10643 8235 10680 8269
rect 10496 8191 10506 8217
rect 10496 8139 10502 8191
rect 10562 8179 10587 8235
rect 10643 8179 10668 8235
rect 10732 8217 10738 8269
tri 11619 8259 11629 8269 ne
rect 10724 8191 10738 8217
rect 10554 8139 10591 8179
rect 10643 8139 10680 8179
rect 10732 8139 10738 8191
tri 9708 8079 9768 8139 se
rect 9768 8131 9834 8139
rect 9768 8079 9782 8131
tri 9782 8079 9834 8131 nw
tri 9634 8005 9708 8079 se
tri 9708 8005 9782 8079 nw
tri 9560 7931 9634 8005 se
tri 9634 7931 9708 8005 nw
tri 9486 7857 9560 7931 se
tri 9560 7857 9634 7931 nw
tri 9468 7839 9486 7857 se
rect 9486 7839 9499 7857
tri 7266 7796 7309 7839 sw
tri 9425 7796 9468 7839 se
rect 9468 7796 9499 7839
tri 9499 7796 9560 7857 nw
rect 7181 7744 7187 7796
rect 7239 7744 7251 7796
rect 7303 7744 7309 7796
tri 9412 7783 9425 7796 se
rect 9425 7783 9486 7796
tri 9486 7783 9499 7796 nw
tri 9373 7744 9412 7783 se
rect 9412 7744 9447 7783
tri 9447 7744 9486 7783 nw
rect 10325 7744 10331 7796
rect 10383 7744 10395 7796
rect 10447 7744 10453 7796
tri 9368 7739 9373 7744 se
rect 9373 7739 9412 7744
tri 9338 7709 9368 7739 se
rect 9368 7709 9412 7739
tri 9412 7709 9447 7744 nw
tri 9287 7658 9338 7709 se
rect 9338 7658 9361 7709
tri 9361 7658 9412 7709 nw
rect 10325 7698 10453 7744
tri 10325 7658 10365 7698 ne
rect 10365 7658 10453 7698
tri 6025 7571 6056 7602 ne
rect 6056 7571 6077 7602
tri 6077 7571 6130 7624 sw
tri 6056 7550 6077 7571 ne
rect 6077 7550 6130 7571
tri 6077 7549 6078 7550 ne
tri 6056 7322 6078 7344 se
rect 6078 7322 6130 7550
tri 6025 7291 6056 7322 se
rect 6056 7291 6077 7322
tri 4695 5022 4709 5036 ne
rect 4709 5022 4747 5036
tri 4747 5022 4783 5058 sw
tri 4709 5000 4731 5022 ne
tri 4657 3001 4731 3075 se
rect 4731 3053 4783 5022
tri 5591 3674 5641 3724 sw
rect 5515 3622 5521 3674
rect 5573 3622 5585 3674
rect 5637 3622 5643 3674
rect 6025 3531 6077 7291
tri 6077 7269 6130 7322 nw
rect 6852 4231 6858 4283
rect 6910 4231 6922 4283
rect 6974 4231 6980 4283
rect 8631 4239 8637 4291
rect 8689 4239 8701 4291
rect 8753 4239 8759 4291
tri 8759 4239 8811 4291 sw
tri 8737 4232 8744 4239 ne
rect 8744 4232 8811 4239
tri 8811 4232 8818 4239 sw
tri 8744 4231 8745 4232 ne
rect 8745 4231 8818 4232
tri 8818 4231 8819 4232 sw
tri 6852 4195 6888 4231 ne
rect 6888 4217 6966 4231
tri 6966 4217 6980 4231 nw
tri 8745 4217 8759 4231 ne
rect 8759 4217 8819 4231
rect 6888 4195 6944 4217
tri 6944 4195 6966 4217 nw
tri 8759 4195 8781 4217 ne
rect 8781 4199 8819 4217
tri 8819 4199 8851 4231 sw
rect 8781 4195 8851 4199
tri 6888 4191 6892 4195 ne
rect 6892 3585 6944 4195
tri 8781 4158 8818 4195 ne
rect 8818 4158 8851 4195
tri 8851 4158 8892 4199 sw
tri 9246 4158 9287 4199 se
rect 9287 4177 9339 7658
tri 9339 7636 9361 7658 nw
tri 10365 7656 10367 7658 ne
rect 10367 7656 10453 7658
tri 10367 7636 10387 7656 ne
rect 10387 7636 10453 7656
tri 10453 7636 10473 7656 sw
tri 10387 7597 10426 7636 ne
rect 10426 7597 10473 7636
tri 10473 7597 10512 7636 sw
tri 10426 7570 10453 7597 ne
rect 10453 7570 10512 7597
tri 10453 7511 10512 7570 ne
tri 10512 7511 10598 7597 sw
tri 10512 7425 10598 7511 ne
tri 10598 7425 10684 7511 sw
tri 10598 7391 10632 7425 ne
rect 10632 6991 10684 7425
tri 10632 6946 10677 6991 ne
rect 10677 6946 10684 6991
tri 10684 6946 10751 7013 sw
tri 10677 6939 10684 6946 ne
rect 10684 6939 10751 6946
tri 10684 6872 10751 6939 ne
tri 10751 6872 10825 6946 sw
tri 10751 6850 10773 6872 ne
rect 10773 6356 10825 6872
tri 10825 6356 10901 6432 sw
rect 10773 6304 10779 6356
rect 10831 6304 10843 6356
rect 10895 6304 10901 6356
rect 11629 5824 11681 8269
tri 11681 8259 11694 8272 nw
rect 13568 8257 13577 8313
rect 13633 8257 13661 8313
rect 13717 8257 13745 8313
rect 13801 8298 13820 8313
rect 13885 8298 13892 8313
rect 14088 8298 14107 8350
rect 14159 8298 14178 8350
rect 14230 8298 14249 8350
rect 14301 8298 14307 8350
rect 13801 8272 13829 8298
rect 13885 8272 13912 8298
rect 13968 8272 13995 8298
rect 14051 8272 14307 8298
rect 13801 8257 13820 8272
rect 13885 8257 13892 8272
rect 13568 8220 13820 8257
rect 13872 8220 13892 8257
rect 13944 8220 13964 8257
rect 14016 8220 14036 8257
rect 14088 8220 14107 8272
rect 14159 8220 14178 8272
rect 14230 8220 14249 8272
rect 14301 8220 14307 8272
rect 14141 8183 14341 8192
rect 14197 8127 14285 8183
rect 14141 8102 14341 8127
rect 14197 8046 14285 8102
rect 14141 8021 14341 8046
rect 14197 7965 14285 8021
rect 14141 7940 14341 7965
rect 14197 7884 14285 7940
rect 14141 7859 14341 7884
rect 14197 7803 14285 7859
rect 14141 7778 14341 7803
rect 14197 7722 14285 7778
rect 14141 7697 14341 7722
rect 14197 7641 14285 7697
rect 14141 7616 14341 7641
rect 14197 7560 14285 7616
rect 14141 7535 14341 7560
rect 14197 7479 14285 7535
rect 14141 7454 14341 7479
rect 14197 7398 14285 7454
rect 14141 7373 14341 7398
rect 14197 7317 14285 7373
rect 14141 7291 14341 7317
rect 14197 7235 14285 7291
rect 14141 7209 14341 7235
rect 14197 7153 14285 7209
rect 14141 7127 14341 7153
rect 14197 7071 14285 7127
rect 14141 7045 14341 7071
rect 14197 6989 14285 7045
rect 14141 6963 14341 6989
rect 14197 6907 14285 6963
rect 14141 6881 14341 6907
rect 14197 6825 14285 6881
rect 14141 6799 14341 6825
rect 14197 6743 14285 6799
rect 14141 6717 14341 6743
rect 14197 6661 14285 6717
rect 14141 6635 14341 6661
rect 14197 6579 14285 6635
rect 14141 6553 14341 6579
rect 14197 6497 14285 6553
rect 14141 6471 14341 6497
rect 14197 6415 14285 6471
rect 14141 6389 14341 6415
rect 12030 6304 12036 6356
rect 12088 6304 12100 6356
rect 12152 6304 12158 6356
rect 14197 6333 14285 6389
rect 14141 6324 14341 6333
tri 12030 6266 12068 6304 ne
rect 12068 6242 12158 6304
tri 12068 6226 12084 6242 ne
rect 12084 6226 12158 6242
tri 12084 6216 12094 6226 ne
rect 12094 6216 12158 6226
tri 12158 6216 12168 6226 sw
tri 12094 6152 12158 6216 ne
rect 12158 6152 12168 6216
tri 12158 6142 12168 6152 ne
tri 12168 6142 12242 6216 sw
tri 12168 6068 12242 6142 ne
tri 12242 6068 12316 6142 sw
tri 12242 6046 12264 6068 ne
rect 11808 5975 11814 6027
rect 11866 5975 11878 6027
rect 11930 5975 11936 6027
tri 11842 5933 11884 5975 ne
rect 11884 5597 11936 5975
tri 11884 5559 11922 5597 ne
rect 11922 5559 11936 5597
tri 11936 5559 11996 5619 sw
tri 11922 5545 11936 5559 ne
rect 11936 5545 11996 5559
tri 11936 5537 11944 5545 ne
rect 9287 4158 9320 4177
tri 9320 4158 9339 4177 nw
tri 11891 4984 11944 5037 se
rect 11944 5015 11996 5545
rect 12264 5091 12316 6068
tri 12513 6027 12543 6057 sw
rect 12461 5975 12467 6027
rect 12519 5975 12531 6027
rect 12583 5975 12589 6027
tri 12513 5945 12543 5975 nw
tri 12264 5051 12304 5091 ne
rect 12304 5051 12316 5091
tri 12316 5051 12378 5113 sw
tri 12304 5039 12316 5051 ne
rect 12316 5039 12378 5051
rect 11944 4984 11965 5015
tri 11965 4984 11996 5015 nw
tri 12316 4984 12371 5039 ne
rect 12371 4984 12378 5039
tri 12378 4984 12445 5051 sw
tri 8818 4106 8870 4158 ne
rect 8870 4106 9268 4158
tri 9268 4106 9320 4158 nw
tri 6944 3585 6948 3589 sw
rect 6892 3567 6948 3585
tri 6892 3548 6911 3567 ne
rect 6911 3548 6948 3567
tri 6077 3531 6094 3548 sw
tri 6911 3531 6928 3548 ne
rect 6928 3531 6948 3548
rect 6025 3526 6094 3531
tri 6025 3457 6094 3526 ne
tri 6094 3511 6114 3531 sw
tri 6928 3511 6948 3531 ne
tri 6948 3511 7022 3585 sw
rect 6094 3457 6114 3511
tri 6114 3457 6168 3511 sw
tri 6948 3457 7002 3511 ne
rect 7002 3457 7022 3511
tri 6094 3399 6152 3457 ne
rect 6152 3437 6168 3457
tri 6168 3437 6188 3457 sw
tri 7002 3437 7022 3457 ne
tri 7022 3437 7096 3511 sw
rect 6152 3399 6188 3437
tri 6188 3399 6226 3437 sw
tri 7022 3399 7060 3437 ne
rect 7060 3399 7096 3437
tri 7096 3399 7134 3437 sw
tri 6152 3383 6168 3399 ne
rect 6168 3383 6226 3399
tri 6226 3383 6242 3399 sw
tri 7060 3383 7076 3399 ne
rect 7076 3383 7134 3399
tri 6168 3347 6204 3383 ne
rect 6204 3363 6242 3383
tri 6242 3363 6262 3383 sw
tri 7076 3363 7096 3383 ne
rect 7096 3363 7134 3383
tri 7134 3363 7170 3399 sw
rect 6204 3358 6262 3363
tri 6262 3358 6267 3363 sw
tri 7096 3358 7101 3363 ne
rect 7101 3358 7170 3363
rect 6204 3347 6267 3358
tri 6267 3347 6278 3358 sw
tri 7101 3347 7112 3358 ne
rect 7112 3347 7170 3358
tri 11880 3347 11891 3358 se
rect 11891 3347 11936 4984
tri 11936 4955 11965 4984 nw
tri 12371 4977 12378 4984 ne
rect 12378 4977 12445 4984
tri 12445 4977 12452 4984 sw
tri 12378 4955 12400 4977 ne
tri 6204 3345 6206 3347 ne
rect 6206 3345 6278 3347
tri 6278 3345 6280 3347 sw
tri 7112 3345 7114 3347 ne
rect 7114 3345 7170 3347
tri 11878 3345 11880 3347 se
rect 11880 3345 11936 3347
tri 6206 3344 6207 3345 ne
rect 6207 3344 6280 3345
tri 6280 3344 6281 3345 sw
rect 6847 3344 7071 3345
tri 6207 3309 6242 3344 ne
rect 6242 3309 6281 3344
tri 6281 3309 6316 3344 sw
tri 6242 3292 6259 3309 ne
rect 6259 3292 6316 3309
tri 6316 3292 6333 3309 sw
rect 6847 3292 6854 3344
rect 6906 3292 6934 3344
rect 6986 3292 7013 3344
rect 7065 3292 7071 3344
tri 7114 3341 7118 3345 ne
tri 6259 3272 6279 3292 ne
rect 6279 3272 6333 3292
tri 6333 3272 6353 3292 sw
rect 6847 3272 7071 3292
tri 6279 3235 6316 3272 ne
rect 6316 3235 6353 3272
tri 6353 3235 6390 3272 sw
tri 6316 3220 6331 3235 ne
rect 6331 3220 6390 3235
tri 6331 3219 6332 3220 ne
rect 6332 3219 6390 3220
tri 6332 3213 6338 3219 ne
tri 4731 3001 4783 3053 nw
tri 4583 2927 4657 3001 se
tri 4657 2927 4731 3001 nw
tri 4553 2897 4583 2927 se
rect 4583 2897 4627 2927
tri 4627 2897 4657 2927 nw
tri 3322 2476 3341 2495 ne
tri 3322 2308 3341 2327 se
rect 3341 2308 3374 2495
rect 3627 2646 4312 2647
rect 3627 2594 3633 2646
rect 3685 2639 3702 2646
rect 3754 2639 3771 2646
rect 3823 2639 3840 2646
rect 3892 2639 3909 2646
rect 3961 2639 3978 2646
rect 4030 2639 4047 2646
rect 4099 2639 4116 2646
rect 4168 2639 4185 2646
rect 4237 2639 4254 2646
rect 3754 2594 3756 2639
rect 3823 2594 3837 2639
rect 3893 2594 3909 2639
rect 3974 2594 3978 2639
rect 4237 2594 4242 2639
rect 4306 2594 4312 2646
rect 3627 2583 3674 2594
rect 3730 2583 3756 2594
rect 3812 2583 3837 2594
rect 3893 2583 3918 2594
rect 3974 2583 3999 2594
rect 4055 2583 4080 2594
rect 4136 2583 4161 2594
rect 4217 2583 4242 2594
rect 4298 2583 4312 2594
rect 3627 2574 4312 2583
rect 3627 2522 3633 2574
rect 3685 2522 3702 2574
rect 3754 2522 3771 2574
rect 3823 2522 3840 2574
rect 3892 2522 3909 2574
rect 3961 2522 3978 2574
rect 4030 2522 4047 2574
rect 4099 2522 4116 2574
rect 4168 2522 4185 2574
rect 4237 2522 4254 2574
rect 4306 2522 4312 2574
rect 3627 2509 4312 2522
rect 3627 2502 3674 2509
rect 3730 2502 3756 2509
rect 3812 2502 3837 2509
rect 3893 2502 3918 2509
rect 3974 2502 3999 2509
rect 4055 2502 4080 2509
rect 4136 2502 4161 2509
rect 4217 2502 4242 2509
rect 4298 2502 4312 2509
rect 3627 2450 3633 2502
rect 3754 2453 3756 2502
rect 3823 2453 3837 2502
rect 3893 2453 3909 2502
rect 3974 2453 3978 2502
rect 4237 2453 4242 2502
rect 3685 2450 3702 2453
rect 3754 2450 3771 2453
rect 3823 2450 3840 2453
rect 3892 2450 3909 2453
rect 3961 2450 3978 2453
rect 4030 2450 4047 2453
rect 4099 2450 4116 2453
rect 4168 2450 4185 2453
rect 4237 2450 4254 2453
rect 4306 2450 4312 2502
rect 3627 2449 4312 2450
tri 2972 2207 3048 2283 ne
rect 3048 2135 3100 2283
tri 3100 2135 3112 2147 sw
rect 3048 2125 3112 2135
tri 3048 2105 3068 2125 ne
rect 3068 2105 3112 2125
tri 3112 2105 3142 2135 sw
tri 3068 2061 3112 2105 ne
rect 3112 2061 3142 2105
tri 3142 2061 3186 2105 sw
tri 3112 2053 3120 2061 ne
rect 3120 2053 3186 2061
tri 3186 2053 3194 2061 sw
tri 3120 2047 3126 2053 ne
rect 3126 2047 3194 2053
tri 3194 2047 3200 2053 sw
tri 3126 2033 3140 2047 ne
rect 3140 2033 3200 2047
tri 3200 2033 3214 2047 sw
tri 3140 1987 3186 2033 ne
rect 3186 1987 3214 2033
tri 3214 1987 3260 2033 sw
tri 3186 1981 3192 1987 ne
rect 3192 1981 3260 1987
tri 3192 1967 3206 1981 ne
rect 3206 1967 3260 1981
tri 3206 1965 3208 1967 ne
tri 2794 1239 2846 1291 nw
tri 2711 1230 2720 1239 se
rect 2720 1230 2731 1239
tri 2244 1176 2276 1208 ne
rect 2276 1176 2296 1208
tri 2296 1176 2350 1230 sw
tri 2657 1176 2711 1230 se
rect 2711 1176 2731 1230
tri 2731 1176 2794 1239 nw
rect 3208 1176 3260 1967
rect 3322 1451 3374 2308
rect 3847 1651 4275 1652
rect 3847 1599 3853 1651
rect 3905 1599 3926 1651
rect 3978 1599 3999 1651
rect 4051 1599 4072 1651
rect 4124 1599 4145 1651
rect 4197 1599 4217 1651
rect 4269 1599 4275 1651
rect 3847 1577 4275 1599
rect 3847 1525 3853 1577
rect 3905 1525 3926 1577
rect 3978 1525 3999 1577
rect 4051 1525 4072 1577
rect 4124 1525 4145 1577
rect 4197 1525 4217 1577
rect 4269 1525 4275 1577
rect 3847 1503 4275 1525
tri 3374 1451 3377 1454 sw
rect 3847 1451 3853 1503
rect 3905 1451 3926 1503
rect 3978 1451 3999 1503
rect 4051 1451 4072 1503
rect 4124 1451 4145 1503
rect 4197 1451 4217 1503
rect 4269 1451 4275 1503
rect 3322 1432 3377 1451
tri 3377 1432 3396 1451 sw
tri 3322 1358 3396 1432 ne
tri 3396 1409 3419 1432 sw
rect 3396 1358 3419 1409
tri 3419 1358 3470 1409 sw
tri 3396 1335 3419 1358 ne
rect 3419 1357 3470 1358
tri 3470 1357 3471 1358 sw
tri 3260 1176 3336 1252 sw
tri 2276 1164 2288 1176 ne
rect 2288 1164 2350 1176
tri 2350 1164 2362 1176 sw
tri 2646 1165 2657 1176 se
rect 2657 1165 2720 1176
tri 2720 1165 2731 1176 nw
tri 2645 1164 2646 1165 se
rect 2646 1164 2679 1165
tri 2288 1156 2296 1164 ne
rect 2296 1156 2362 1164
tri 2296 1124 2328 1156 ne
rect 2328 1124 2362 1156
tri 2362 1124 2402 1164 sw
tri 2605 1124 2645 1164 se
rect 2645 1124 2679 1164
tri 2679 1124 2720 1165 nw
rect 3208 1124 3214 1176
rect 3266 1124 3278 1176
rect 3330 1124 3336 1176
tri 2328 1109 2343 1124 ne
rect 2343 1109 2402 1124
tri 2402 1109 2417 1124 sw
tri 2590 1109 2605 1124 se
rect 2605 1109 2664 1124
tri 2664 1109 2679 1124 nw
tri 2343 1090 2362 1109 ne
rect 2362 1090 2417 1109
tri 2417 1090 2436 1109 sw
tri 2572 1091 2590 1109 se
rect 2590 1091 2646 1109
tri 2646 1091 2664 1109 nw
tri 2571 1090 2572 1091 se
rect 2572 1090 2645 1091
tri 2645 1090 2646 1091 nw
tri 2362 1087 2365 1090 ne
rect 2365 1087 2436 1090
tri 2568 1087 2571 1090 se
rect 2571 1087 2642 1090
tri 2642 1087 2645 1090 nw
tri 2365 1086 2366 1087 ne
rect 2366 1086 2436 1087
tri 2567 1086 2568 1087 se
rect 2568 1086 2641 1087
tri 2641 1086 2642 1087 nw
rect 2779 1086 2788 1087
rect 2844 1086 2889 1087
rect 2945 1086 2990 1087
rect 3046 1086 3091 1087
rect 3147 1086 3192 1087
rect 3248 1086 3293 1087
tri 2366 1068 2384 1086 ne
tri 2199 1026 2204 1031 sw
rect 2147 1014 2204 1026
tri 2204 1014 2216 1026 sw
rect 2147 1010 2216 1014
tri 2216 1010 2220 1014 sw
rect 2147 1009 2220 1010
tri 2147 972 2184 1009 ne
rect 2184 972 2220 1009
tri 2220 972 2258 1010 sw
tri 2184 958 2198 972 ne
rect 2198 958 2258 972
tri 2198 957 2199 958 ne
rect 2199 957 2258 958
tri 2199 950 2206 957 ne
rect 1689 735 1725 751
tri 1725 735 1741 751 nw
tri 1636 720 1651 735 se
rect 1651 720 1710 735
tri 1710 720 1725 735 nw
tri 1615 699 1636 720 se
rect 1636 699 1689 720
tri 1689 699 1710 720 nw
tri 1592 676 1615 699 se
rect 1615 676 1658 699
tri 1201 551 1213 563 se
rect 1213 551 1265 676
tri 1584 668 1592 676 se
rect 1592 668 1658 676
tri 1658 668 1689 699 nw
tri 1571 655 1584 668 se
rect 1584 655 1645 668
tri 1645 655 1658 668 nw
tri 1561 645 1571 655 se
rect 1571 645 1635 655
tri 1635 645 1645 655 nw
tri 1556 640 1561 645 se
rect 1561 640 1630 645
tri 1630 640 1635 645 nw
tri 1541 625 1556 640 se
rect 1556 625 1615 640
tri 1615 625 1630 640 nw
tri 1525 609 1541 625 se
rect 1541 609 1599 625
tri 1599 609 1615 625 nw
tri 1510 594 1525 609 se
rect 1525 594 1584 609
tri 1584 594 1599 609 nw
tri 2191 594 2206 609 se
rect 2206 594 2258 957
tri 2383 621 2384 622 se
rect 2384 621 2436 1086
tri 2356 594 2383 621 se
rect 2383 594 2436 621
tri 1492 576 1510 594 se
rect 1510 576 1566 594
tri 1566 576 1584 594 nw
tri 2173 576 2191 594 se
rect 2191 587 2258 594
rect 2191 576 2247 587
tri 2247 576 2258 587 nw
tri 2338 576 2356 594 se
rect 2356 576 2436 594
tri 1491 575 1492 576 se
rect 1492 575 1565 576
tri 1565 575 1566 576 nw
tri 2172 575 2173 576 se
rect 2173 575 2246 576
tri 2246 575 2247 576 nw
tri 2337 575 2338 576 se
rect 2338 575 2436 576
tri 1467 551 1491 575 se
rect 1491 551 1541 575
tri 1541 551 1565 575 nw
tri 2148 551 2172 575 se
rect 2172 551 2206 575
tri 1173 523 1201 551 se
rect 1201 523 1265 551
tri 1265 523 1293 551 sw
tri 1451 535 1467 551 se
rect 1467 535 1525 551
tri 1525 535 1541 551 nw
tri 2132 535 2148 551 se
rect 2148 535 2206 551
tri 2206 535 2246 575 nw
tri 1439 523 1451 535 se
rect 1451 523 1513 535
tri 1513 523 1525 535 nw
tri 2120 523 2132 535 se
rect 2132 523 2194 535
tri 2194 523 2206 535 nw
rect 2308 523 2314 575
rect 2366 523 2378 575
rect 2430 523 2436 575
tri 2551 1070 2567 1086 se
rect 2567 1070 2625 1086
tri 2625 1070 2641 1086 nw
tri 1169 519 1173 523 se
rect 1173 519 1293 523
tri 1293 519 1297 523 sw
tri 1435 519 1439 523 se
rect 1439 519 1509 523
tri 1509 519 1513 523 nw
tri 2116 519 2120 523 se
rect 2120 519 2190 523
tri 2190 519 2194 523 nw
rect 1169 467 1175 519
rect 1227 467 1239 519
rect 1291 467 1297 519
tri 1393 477 1435 519 se
rect 1435 477 1467 519
tri 1467 477 1509 519 nw
tri 1383 467 1393 477 se
rect 1393 467 1457 477
tri 1457 467 1467 477 nw
rect 1896 467 1902 519
rect 1954 467 1966 519
rect 2018 512 2183 519
tri 2183 512 2190 519 nw
rect 2018 506 2177 512
tri 2177 506 2183 512 nw
rect 2018 498 2169 506
tri 2169 498 2177 506 nw
rect 2018 483 2154 498
tri 2154 483 2169 498 nw
rect 2018 467 2138 483
tri 2138 467 2154 483 nw
tri 1347 431 1383 467 se
rect 1383 431 1421 467
tri 1421 431 1457 467 nw
tri 1319 403 1347 431 se
rect 1347 403 1393 431
tri 1393 403 1421 431 nw
tri 1293 377 1319 403 se
rect 1319 377 1367 403
tri 1367 377 1393 403 nw
tri 1253 337 1293 377 se
rect 1293 337 1327 377
tri 1327 337 1367 377 nw
tri 1245 329 1253 337 se
rect 1253 329 1319 337
tri 1319 329 1327 337 nw
tri 1226 310 1245 329 se
rect 1245 310 1300 329
tri 1300 310 1319 329 nw
rect 1226 0 1278 310
tri 1278 288 1300 310 nw
rect 1379 200 1388 256
rect 1444 255 1475 256
rect 1531 255 1562 256
rect 1531 203 1548 255
rect 1444 200 1475 203
rect 1531 200 1562 203
rect 1618 200 1648 256
rect 1704 255 1734 256
rect 1790 255 1820 256
rect 1876 255 1906 256
rect 1962 255 1992 256
rect 1708 203 1734 255
rect 1816 203 1820 255
rect 1962 203 1978 255
rect 1704 200 1734 203
rect 1790 200 1820 203
rect 1876 200 1906 203
rect 1962 200 1992 203
rect 2048 200 2078 256
rect 2134 255 2143 256
rect 2137 203 2143 255
rect 2134 200 2143 203
rect 1379 181 2143 200
rect 1379 129 1440 181
rect 1492 129 1548 181
rect 1600 129 1656 181
rect 1708 129 1764 181
rect 1816 129 1871 181
rect 1923 129 1978 181
rect 2030 129 2085 181
rect 2137 129 2143 181
rect 1379 110 2143 129
rect 1379 54 1388 110
rect 1444 107 1475 110
rect 1531 107 1562 110
rect 1531 55 1548 107
rect 1444 54 1475 55
rect 1531 54 1562 55
rect 1618 54 1648 110
rect 1704 107 1734 110
rect 1790 107 1820 110
rect 1876 107 1906 110
rect 1962 107 1992 110
rect 1708 55 1734 107
rect 1816 55 1820 107
rect 1962 55 1978 107
rect 1704 54 1734 55
rect 1790 54 1820 55
rect 1876 54 1906 55
rect 1962 54 1992 55
rect 2048 54 2078 110
rect 2134 107 2143 110
rect 2137 55 2143 107
rect 2134 54 2143 55
rect 2551 0 2603 1070
tri 2603 1048 2625 1070 nw
rect 2779 1034 2785 1086
rect 2844 1034 2857 1086
rect 2980 1034 2990 1086
rect 3051 1034 3070 1086
rect 3264 1034 3283 1086
rect 2779 1031 2788 1034
rect 2844 1031 2889 1034
rect 2945 1031 2990 1034
rect 3046 1031 3091 1034
rect 3147 1031 3192 1034
rect 3248 1031 3293 1034
rect 3349 1031 3358 1087
rect 2779 1010 3358 1031
rect 2779 958 2785 1010
rect 2837 958 2857 1010
rect 2909 958 2928 1010
rect 2980 958 2999 1010
rect 3051 958 3070 1010
rect 3122 958 3141 1010
rect 3193 958 3212 1010
rect 3264 958 3283 1010
rect 3335 958 3358 1010
rect 2779 937 3358 958
rect 2779 934 2788 937
rect 2844 934 2889 937
rect 2945 934 2990 937
rect 3046 934 3091 937
rect 3147 934 3192 937
rect 3248 934 3293 937
rect 2779 882 2785 934
rect 2844 882 2857 934
rect 2980 882 2990 934
rect 3051 882 3070 934
rect 3264 882 3283 934
rect 2779 881 2788 882
rect 2844 881 2889 882
rect 2945 881 2990 882
rect 3046 881 3091 882
rect 3147 881 3192 882
rect 3248 881 3293 882
rect 3349 881 3358 937
tri 3392 594 3419 621 se
rect 3419 599 3471 1357
rect 3419 594 3466 599
tri 3466 594 3471 599 nw
tri 3374 576 3392 594 se
rect 3392 576 3448 594
tri 3448 576 3466 594 nw
tri 3362 564 3374 576 se
rect 3374 564 3436 576
tri 3436 564 3448 576 nw
tri 3345 547 3362 564 se
rect 3362 547 3419 564
tri 3419 547 3436 564 nw
tri 3333 535 3345 547 se
rect 3345 535 3384 547
tri 3317 519 3333 535 se
rect 3333 519 3384 535
tri 3310 512 3317 519 se
rect 3317 512 3384 519
tri 3384 512 3419 547 nw
tri 3304 506 3310 512 se
rect 3310 506 3378 512
tri 3378 506 3384 512 nw
tri 3296 498 3304 506 se
rect 3304 498 3370 506
tri 3370 498 3378 506 nw
tri 3281 483 3296 498 se
rect 3296 483 3355 498
tri 3355 483 3370 498 nw
tri 3271 473 3281 483 se
rect 3281 473 3345 483
tri 3345 473 3355 483 nw
tri 3265 467 3271 473 se
rect 3271 467 3336 473
tri 3262 464 3265 467 se
rect 3265 464 3336 467
tri 3336 464 3345 473 nw
rect 3262 0 3314 464
tri 3314 442 3336 464 nw
rect 3847 255 4275 1451
tri 4511 1325 4553 1367 se
rect 4553 1345 4605 2897
tri 4605 2875 4627 2897 nw
rect 4553 1325 4585 1345
tri 4585 1325 4605 1345 nw
rect 4848 1651 4857 1653
rect 4913 1651 4940 1653
rect 4996 1651 5023 1653
rect 5079 1651 5106 1653
rect 5162 1651 5188 1653
rect 5244 1651 5253 1653
rect 4848 1599 4854 1651
rect 4913 1599 4923 1651
rect 5179 1599 5188 1651
rect 5247 1599 5253 1651
rect 4848 1597 4857 1599
rect 4913 1597 4940 1599
rect 4996 1597 5023 1599
rect 5079 1597 5106 1599
rect 5162 1597 5188 1599
rect 5244 1597 5253 1599
rect 4848 1577 5253 1597
rect 4848 1525 4854 1577
rect 4906 1525 4923 1577
rect 4975 1525 4991 1577
rect 5043 1525 5059 1577
rect 5111 1525 5127 1577
rect 5179 1525 5195 1577
rect 5247 1525 5253 1577
rect 4848 1507 5253 1525
rect 4848 1503 4857 1507
rect 4913 1503 4940 1507
rect 4996 1503 5023 1507
rect 5079 1503 5106 1507
rect 5162 1503 5188 1507
rect 5244 1503 5253 1507
rect 4848 1451 4854 1503
rect 4913 1451 4923 1503
rect 5179 1451 5188 1503
rect 5247 1451 5253 1503
rect 4848 1409 5253 1451
tri 4479 1293 4511 1325 se
rect 4511 1293 4553 1325
tri 4553 1293 4585 1325 nw
rect 3847 203 3853 255
rect 3905 203 3926 255
rect 3978 203 3999 255
rect 4051 203 4072 255
rect 4124 203 4145 255
rect 4197 203 4217 255
rect 4269 203 4275 255
rect 3847 181 4275 203
rect 3847 129 3853 181
rect 3905 129 3926 181
rect 3978 129 3999 181
rect 4051 129 4072 181
rect 4124 129 4145 181
rect 4197 129 4217 181
rect 4269 129 4275 181
rect 3847 107 4275 129
rect 3847 55 3853 107
rect 3905 55 3926 107
rect 3978 55 3999 107
rect 4051 55 4072 107
rect 4124 55 4145 107
rect 4197 55 4217 107
rect 4269 55 4275 107
rect 3847 54 4275 55
tri 4471 1285 4479 1293 se
rect 4479 1285 4545 1293
tri 4545 1285 4553 1293 nw
rect 4471 0 4523 1285
tri 4523 1263 4545 1285 nw
rect 4848 713 4862 1409
rect 5238 713 5253 1409
tri 5814 930 5842 958 se
rect 5842 936 5894 1356
tri 6330 958 6338 966 se
rect 6338 958 6390 3219
rect 6847 3220 6854 3272
rect 6906 3220 6934 3272
rect 6986 3220 7013 3272
rect 7065 3220 7071 3272
rect 6847 3200 7071 3220
rect 6847 3148 6854 3200
rect 6906 3148 6934 3200
rect 6986 3148 7013 3200
rect 7065 3148 7071 3200
rect 6847 3145 7071 3148
rect 6903 3089 6931 3145
rect 6987 3089 7015 3145
rect 6847 3022 7071 3089
rect 6903 2966 6931 3022
rect 6987 2966 7015 3022
rect 6847 2899 7071 2966
rect 6903 2843 6931 2899
rect 6987 2843 7015 2899
rect 6847 2776 7071 2843
rect 6903 2720 6931 2776
rect 6987 2720 7015 2776
rect 6847 2653 7071 2720
rect 6903 2597 6931 2653
rect 6987 2597 7015 2653
rect 6847 2530 7071 2597
rect 6903 2474 6931 2530
rect 6987 2474 7015 2530
rect 6847 2407 7071 2474
rect 6903 2351 6931 2407
rect 6987 2351 7015 2407
rect 6847 2284 7071 2351
rect 6903 2228 6931 2284
rect 6987 2228 7015 2284
rect 8615 3293 8621 3345
rect 8673 3293 8717 3345
rect 8769 3293 8775 3345
tri 11866 3333 11878 3345 se
rect 11878 3333 11936 3345
rect 8615 3271 8775 3293
tri 11817 3284 11866 3333 se
rect 11866 3329 11936 3333
rect 11866 3284 11891 3329
tri 11891 3284 11936 3329 nw
rect 8615 3219 8621 3271
rect 8673 3219 8717 3271
rect 8769 3219 8775 3271
rect 8615 3197 8775 3219
tri 11743 3210 11817 3284 se
tri 11817 3210 11891 3284 nw
rect 8615 3145 8621 3197
rect 8673 3145 8717 3197
rect 8769 3145 8775 3197
tri 11678 3145 11743 3210 se
rect 8671 3089 8719 3145
tri 11669 3136 11678 3145 se
rect 11678 3136 11743 3145
tri 11743 3136 11817 3210 nw
rect 8615 3023 8775 3089
rect 8671 2967 8719 3023
rect 8615 2901 8775 2967
rect 8671 2845 8719 2901
rect 8615 2779 8775 2845
rect 8671 2723 8719 2779
rect 8615 2657 8775 2723
rect 8671 2601 8719 2657
tri 11657 3124 11669 3136 se
rect 11669 3124 11731 3136
tri 11731 3124 11743 3136 nw
rect 8615 2535 8775 2601
rect 8671 2479 8719 2535
rect 8615 2412 8775 2479
rect 10506 2595 10512 2647
rect 10564 2637 10579 2647
rect 10631 2637 10707 2647
rect 10759 2637 10780 2647
rect 10832 2637 10853 2647
rect 10905 2637 10926 2647
rect 10978 2637 10999 2647
rect 10578 2595 10579 2637
rect 10506 2581 10522 2595
rect 10578 2581 10614 2595
rect 10670 2581 10706 2637
rect 10762 2595 10780 2637
rect 10978 2595 10982 2637
rect 11051 2595 11057 2647
rect 10762 2581 10798 2595
rect 10854 2581 10890 2595
rect 10946 2581 10982 2595
rect 11038 2581 11057 2595
rect 10506 2575 11057 2581
rect 10506 2523 10512 2575
rect 10564 2523 10579 2575
rect 10631 2523 10707 2575
rect 10759 2523 10780 2575
rect 10832 2523 10853 2575
rect 10905 2523 10926 2575
rect 10978 2523 10999 2575
rect 11051 2523 11057 2575
rect 10506 2515 11057 2523
rect 10506 2503 10522 2515
rect 10578 2503 10614 2515
rect 10506 2451 10512 2503
rect 10578 2459 10579 2503
rect 10670 2459 10706 2515
rect 10762 2503 10798 2515
rect 10854 2503 10890 2515
rect 10946 2503 10982 2515
rect 11038 2503 11057 2515
rect 10762 2459 10780 2503
rect 10978 2459 10982 2503
rect 10564 2451 10579 2459
rect 10631 2451 10707 2459
rect 10759 2451 10780 2459
rect 10832 2451 10853 2459
rect 10905 2451 10926 2459
rect 10978 2451 10999 2459
rect 11051 2451 11057 2503
rect 10506 2448 11057 2451
tri 10559 2429 10578 2448 ne
rect 10578 2429 10760 2448
tri 10760 2429 10779 2448 nw
tri 10578 2423 10584 2429 ne
rect 10584 2423 10754 2429
tri 10754 2423 10760 2429 nw
rect 8671 2356 8719 2412
tri 10584 2371 10636 2423 ne
rect 10636 2371 10702 2423
tri 10702 2371 10754 2423 nw
tri 10636 2364 10643 2371 ne
rect 10643 2364 10695 2371
tri 10695 2364 10702 2371 nw
rect 8615 2289 8775 2356
rect 6847 2161 7071 2228
tri 7736 2207 7812 2283 ne
rect 6903 2105 6931 2161
rect 6987 2105 7015 2161
rect 6847 2038 7071 2105
rect 6903 1982 6931 2038
rect 6987 1982 7015 2038
rect 6847 1915 7071 1982
rect 6903 1859 6931 1915
rect 6987 1859 7015 1915
rect 6847 1810 7071 1859
rect 6847 1758 6854 1810
rect 6906 1758 6934 1810
rect 6986 1758 7013 1810
rect 7065 1758 7071 1810
rect 6847 1732 7071 1758
rect 6847 1680 6854 1732
rect 6906 1680 6934 1732
rect 6986 1680 7013 1732
rect 7065 1680 7071 1732
rect 6838 1651 7057 1652
rect 6838 1599 6844 1651
rect 6896 1599 6922 1651
rect 6974 1599 6999 1651
rect 7051 1599 7057 1651
rect 6838 1577 7057 1599
rect 6838 1525 6844 1577
rect 6896 1525 6922 1577
rect 6974 1525 6999 1577
rect 7051 1525 7057 1577
rect 7812 1606 7864 2283
rect 8671 2233 8719 2289
rect 8615 2166 8775 2233
rect 8671 2110 8719 2166
rect 8615 2043 8775 2110
rect 8671 1987 8719 2043
rect 8615 1810 8775 1987
rect 8615 1758 8621 1810
rect 8673 1758 8717 1810
rect 8769 1758 8775 1810
rect 8615 1732 8775 1758
rect 8615 1680 8621 1732
rect 8673 1680 8717 1732
rect 8769 1680 8775 1732
tri 7812 1560 7858 1606 ne
rect 7858 1560 7864 1606
tri 7864 1560 7932 1628 sw
tri 7858 1554 7864 1560 ne
rect 7864 1554 7932 1560
rect 6838 1503 7057 1525
rect 6838 1451 6844 1503
rect 6896 1451 6922 1503
rect 6974 1451 6999 1503
rect 7051 1451 7057 1503
tri 7864 1486 7932 1554 ne
tri 7932 1486 8006 1560 sw
tri 7932 1464 7954 1486 ne
tri 6689 1176 6838 1325 se
rect 6838 1236 7057 1451
rect 6838 1176 6997 1236
tri 6997 1176 7057 1236 nw
rect 5842 930 5888 936
tri 5888 930 5894 936 nw
tri 6302 930 6330 958 se
rect 6330 944 6390 958
rect 6330 930 6376 944
tri 6376 930 6390 944 nw
tri 6680 1167 6689 1176 se
rect 6689 1167 6988 1176
tri 6988 1167 6997 1176 nw
rect 6680 1124 6945 1167
tri 6945 1124 6988 1167 nw
tri 5776 892 5814 930 se
rect 5814 892 5850 930
tri 5850 892 5888 930 nw
tri 6264 892 6302 930 se
rect 6302 892 6338 930
tri 6338 892 6376 930 nw
tri 5768 884 5776 892 se
rect 5776 884 5842 892
tri 5842 884 5850 892 nw
tri 6261 889 6264 892 se
rect 6264 889 6335 892
tri 6335 889 6338 892 nw
tri 5762 878 5768 884 se
rect 5768 878 5836 884
tri 5836 878 5842 884 nw
rect 6261 878 6324 889
tri 6324 878 6335 889 nw
tri 5754 870 5762 878 se
rect 5762 870 5828 878
tri 5828 870 5836 878 nw
rect 6261 870 6316 878
tri 6316 870 6324 878 nw
tri 5723 839 5754 870 se
rect 5754 839 5797 870
tri 5797 839 5828 870 nw
rect 4848 688 5253 713
rect 4848 632 4862 688
rect 4918 632 4942 688
rect 4998 632 5022 688
rect 5078 632 5102 688
rect 5158 632 5182 688
rect 5238 632 5253 688
rect 4848 607 5253 632
rect 4848 551 4862 607
rect 4918 551 4942 607
rect 4998 551 5022 607
rect 5078 551 5102 607
rect 5158 551 5182 607
rect 5238 551 5253 607
rect 4848 526 5253 551
rect 4848 470 4862 526
rect 4918 470 4942 526
rect 4998 470 5022 526
rect 5078 470 5102 526
rect 5158 470 5182 526
rect 5238 470 5253 526
tri 4833 431 4848 446 se
rect 4848 445 5253 470
rect 4848 431 4862 445
tri 4779 377 4833 431 se
rect 4833 389 4862 431
rect 4918 389 4942 445
rect 4998 389 5022 445
rect 5078 389 5102 445
rect 5158 389 5182 445
rect 5238 389 5253 445
rect 4833 377 5253 389
tri 4739 337 4779 377 se
rect 4779 364 5253 377
rect 4779 337 4862 364
tri 4701 299 4739 337 se
rect 4739 308 4862 337
rect 4918 308 4942 364
rect 4998 308 5022 364
rect 5078 308 5102 364
rect 5158 308 5182 364
rect 5238 308 5253 364
tri 5698 814 5723 839 se
rect 5723 814 5772 839
tri 5772 814 5797 839 nw
rect 4739 299 5253 308
tri 4687 285 4701 299 se
rect 4701 285 5253 299
tri 4663 261 4687 285 se
rect 4687 261 5253 285
tri 4659 257 4663 261 se
rect 4663 257 5253 261
rect 4599 201 4608 257
rect 4664 256 4691 257
rect 4747 256 4774 257
rect 4747 204 4767 256
rect 4664 201 4691 204
rect 4747 201 4774 204
rect 4830 201 4857 257
rect 4913 256 4940 257
rect 4996 256 5023 257
rect 5079 256 5106 257
rect 4926 204 4940 256
rect 5079 204 5088 256
rect 4913 201 4940 204
rect 4996 201 5023 204
rect 5079 201 5106 204
rect 5162 201 5188 257
rect 5244 256 5253 257
rect 5247 204 5253 256
rect 5244 201 5253 204
rect 4599 182 5253 201
rect 4599 130 4660 182
rect 4712 130 4767 182
rect 4819 130 4874 182
rect 4926 130 4981 182
rect 5033 130 5088 182
rect 5140 130 5195 182
rect 5247 130 5253 182
rect 4599 111 5253 130
rect 4599 55 4608 111
rect 4664 108 4691 111
rect 4747 108 4774 111
rect 4747 56 4767 108
rect 4664 55 4691 56
rect 4747 55 4774 56
rect 4830 55 4857 111
rect 4913 108 4940 111
rect 4996 108 5023 111
rect 5079 108 5106 111
rect 4926 56 4940 108
rect 5079 56 5088 108
rect 4913 55 4940 56
rect 4996 55 5023 56
rect 5079 55 5106 56
rect 5162 55 5188 111
rect 5244 108 5253 111
rect 5247 56 5253 108
rect 5244 55 5253 56
rect 5320 0 5372 339
rect 5698 0 5750 814
tri 5750 792 5772 814 nw
tri 6248 551 6261 564 se
rect 6261 551 6313 870
tri 6313 867 6316 870 nw
tri 6216 519 6248 551 se
rect 6248 542 6313 551
rect 6248 519 6283 542
tri 6209 512 6216 519 se
rect 6216 512 6283 519
tri 6283 512 6313 542 nw
rect 6363 787 6415 793
rect 6363 720 6415 735
tri 6203 506 6209 512 se
rect 6209 506 6277 512
tri 6277 506 6283 512 nw
tri 6195 498 6203 506 se
rect 6203 498 6269 506
tri 6269 498 6277 506 nw
tri 6187 490 6195 498 se
rect 6195 490 6261 498
tri 6261 490 6269 498 nw
tri 6180 483 6187 490 se
rect 6187 483 6254 490
tri 6254 483 6261 490 nw
tri 6164 467 6180 483 se
rect 6180 467 6224 483
tri 6150 453 6164 467 se
rect 6164 453 6224 467
tri 6224 453 6254 483 nw
rect 6150 0 6202 453
tri 6202 431 6224 453 nw
rect 6363 0 6415 668
rect 6680 255 6934 1124
tri 6934 1113 6945 1124 nw
rect 7027 771 7079 777
rect 7027 707 7079 719
rect 7027 445 7079 655
tri 7027 431 7041 445 ne
rect 7041 431 7079 445
tri 7079 431 7115 467 sw
tri 7041 402 7070 431 ne
rect 7070 402 7115 431
tri 7115 402 7144 431 sw
tri 7070 380 7092 402 ne
rect 6680 203 6686 255
rect 6738 203 6781 255
rect 6833 203 6876 255
rect 6928 203 6934 255
rect 6680 181 6934 203
rect 6680 129 6686 181
rect 6738 129 6781 181
rect 6833 129 6876 181
rect 6928 129 6934 181
rect 6680 107 6934 129
rect 6680 55 6686 107
rect 6738 55 6781 107
rect 6833 55 6876 107
rect 6928 55 6934 107
rect 6680 54 6934 55
rect 7092 0 7144 402
rect 7678 0 7730 743
tri 7925 377 7954 406 se
rect 7954 377 8006 1486
tri 9966 1356 9971 1361 se
rect 8932 1124 8938 1176
rect 8990 1124 9002 1176
rect 9054 1124 9060 1176
tri 8932 1120 8936 1124 ne
rect 8936 1120 9056 1124
tri 9056 1120 9060 1124 nw
tri 9151 1120 9171 1140 se
rect 9171 1120 9223 1356
tri 9949 1339 9966 1356 se
rect 9966 1339 10023 1356
rect 8936 1113 9049 1120
tri 9049 1113 9056 1120 nw
tri 9144 1113 9151 1120 se
rect 9151 1118 9223 1120
rect 9151 1113 9214 1118
rect 8936 1109 9045 1113
tri 9045 1109 9049 1113 nw
tri 9140 1109 9144 1113 se
rect 9144 1109 9214 1113
tri 9214 1109 9223 1118 nw
tri 9925 1315 9949 1339 se
rect 9949 1315 9977 1339
rect 8936 1090 9026 1109
tri 9026 1090 9045 1109 nw
tri 9121 1090 9140 1109 se
rect 9140 1090 9195 1109
tri 9195 1090 9214 1109 nw
rect 8936 839 8988 1090
tri 8988 1052 9026 1090 nw
tri 9097 1066 9121 1090 se
rect 9121 1066 9171 1090
tri 9171 1066 9195 1090 nw
tri 9083 1052 9097 1066 se
rect 9097 1052 9143 1066
tri 9069 1038 9083 1052 se
rect 9083 1038 9143 1052
tri 9143 1038 9171 1066 nw
tri 9057 1026 9069 1038 se
rect 9069 1026 9131 1038
tri 9131 1026 9143 1038 nw
rect 8936 775 8988 787
rect 8936 717 8988 723
tri 9049 1018 9057 1026 se
rect 9057 1018 9123 1026
tri 9123 1018 9131 1026 nw
rect 9049 1014 9119 1018
tri 9119 1014 9123 1018 nw
rect 9049 1010 9115 1014
tri 9115 1010 9119 1014 nw
tri 7885 337 7925 377 se
rect 7925 337 8006 377
rect 7878 285 7884 337
rect 7936 285 7948 337
rect 8000 285 8006 337
rect 9049 0 9101 1010
tri 9101 996 9115 1010 nw
rect 9776 761 9832 767
rect 9828 758 9832 761
rect 9776 697 9832 702
rect 9828 678 9832 697
rect 9776 613 9832 622
rect 9925 483 9977 1315
tri 9977 1293 10023 1339 nw
tri 11354 1092 11366 1104 se
rect 11366 1092 11418 2283
tri 11418 2248 11453 2283 nw
tri 11655 1161 11657 1163 se
rect 11657 1161 11709 3124
tri 11709 3102 11731 3124 nw
rect 12400 2729 12452 4977
tri 15742 3444 15783 3485 se
rect 15783 3463 15835 8469
tri 14211 3347 14263 3399 se
rect 14263 3347 14310 3399
rect 14362 3347 14374 3399
rect 14426 3347 14432 3399
tri 14186 3322 14211 3347 se
rect 14211 3345 14267 3347
tri 14267 3345 14269 3347 nw
rect 14211 3333 14255 3345
tri 14255 3333 14267 3345 nw
rect 14211 3322 14244 3333
tri 14244 3322 14255 3333 nw
tri 14128 3264 14186 3322 se
tri 14186 3264 14244 3322 nw
tri 14110 3246 14128 3264 se
rect 14128 3246 14168 3264
tri 14168 3246 14186 3264 nw
rect 13336 3206 14128 3246
tri 14128 3206 14168 3246 nw
tri 12400 2710 12419 2729 ne
rect 12419 2710 12452 2729
tri 12452 2710 12493 2751 sw
tri 12419 2677 12452 2710 ne
rect 12452 2709 12493 2710
tri 12493 2709 12494 2710 sw
rect 12452 2677 12494 2709
tri 12452 2636 12493 2677 ne
rect 12493 2636 12494 2677
tri 12494 2636 12567 2709 sw
tri 12493 2562 12567 2636 ne
tri 12567 2562 12641 2636 sw
tri 12567 2540 12589 2562 ne
tri 11890 2207 11966 2283 ne
tri 11614 1120 11655 1161 se
rect 11655 1141 11709 1161
rect 11655 1120 11677 1141
tri 11607 1113 11614 1120 se
rect 11614 1113 11677 1120
tri 11603 1109 11607 1113 se
rect 11607 1109 11677 1113
tri 11677 1109 11709 1141 nw
rect 11966 1137 12018 2283
tri 12570 1909 12589 1928 se
rect 12589 1909 12641 2562
rect 14626 2105 14847 3444
tri 15709 3411 15742 3444 se
rect 15742 3411 15783 3444
tri 15783 3411 15835 3463 nw
tri 15704 3406 15709 3411 se
rect 15709 3406 15778 3411
tri 15778 3406 15783 3411 nw
tri 15697 3399 15704 3406 se
rect 15704 3399 15724 3406
rect 15355 3347 15361 3399
rect 15413 3347 15425 3399
rect 15477 3347 15483 3399
tri 15650 3352 15697 3399 se
rect 15697 3352 15724 3399
tri 15724 3352 15778 3406 nw
tri 15810 3352 15864 3406 se
rect 15864 3390 15902 9554
tri 15864 3352 15902 3390 nw
tri 15645 3347 15650 3352 se
rect 15650 3347 15719 3352
tri 15719 3347 15724 3352 nw
tri 15805 3347 15810 3352 se
tri 15355 3345 15357 3347 ne
rect 15357 3345 15469 3347
tri 15357 3333 15369 3345 ne
rect 15369 3333 15469 3345
tri 15469 3333 15483 3347 nw
tri 15635 3337 15645 3347 se
rect 15645 3337 15709 3347
tri 15709 3337 15719 3347 nw
tri 15795 3337 15805 3347 se
rect 15805 3337 15810 3347
tri 15632 3334 15635 3337 se
rect 15635 3334 15706 3337
tri 15706 3334 15709 3337 nw
tri 15792 3334 15795 3337 se
rect 15795 3334 15810 3337
rect 15632 3333 15705 3334
tri 15705 3333 15706 3334 nw
tri 15791 3333 15792 3334 se
rect 15792 3333 15810 3334
rect 15369 2761 15421 3333
tri 15421 3285 15469 3333 nw
tri 15421 2761 15443 2783 sw
tri 15369 2709 15421 2761 ne
rect 15421 2731 15443 2761
tri 15443 2731 15473 2761 sw
rect 15421 2423 15473 2731
rect 15421 2359 15473 2371
rect 15421 2301 15473 2307
rect 14626 2053 14632 2105
rect 14684 2053 14711 2105
rect 14763 2053 14789 2105
rect 14841 2053 14847 2105
rect 14626 2033 14847 2053
rect 14626 1981 14632 2033
rect 14684 1981 14711 2033
rect 14763 1981 14789 2033
rect 14841 1981 14847 2033
rect 14626 1961 14847 1981
rect 14626 1909 14632 1961
rect 14684 1909 14711 1961
rect 14763 1909 14789 1961
rect 14841 1909 14847 1961
rect 15076 2099 15251 2105
rect 15076 2047 15077 2099
rect 15129 2047 15199 2099
rect 15076 2033 15251 2047
rect 15076 1981 15077 2033
rect 15129 1981 15199 2033
rect 15076 1967 15251 1981
rect 15076 1915 15077 1967
rect 15129 1915 15199 1967
rect 15632 1989 15684 3333
tri 15684 3312 15705 3333 nw
tri 15770 3312 15791 3333 se
rect 15791 3312 15810 3333
tri 15756 3298 15770 3312 se
rect 15770 3298 15810 3312
tri 15810 3298 15864 3352 nw
tri 15743 3285 15756 3298 se
rect 15756 3285 15777 3298
tri 15723 3265 15743 3285 se
rect 15743 3265 15777 3285
tri 15777 3265 15810 3298 nw
rect 15723 2068 15761 3265
tri 15761 3249 15777 3265 nw
tri 15761 2068 15782 2089 sw
rect 15723 2053 15782 2068
tri 15723 2034 15742 2053 ne
tri 15684 1989 15706 2011 sw
tri 15632 1960 15661 1989 ne
rect 15661 1982 15706 1989
tri 15706 1982 15713 1989 sw
tri 12515 1854 12570 1909 se
rect 12570 1906 12641 1909
rect 12570 1854 12589 1906
tri 12589 1854 12641 1906 nw
tri 12441 1780 12515 1854 se
tri 12515 1780 12589 1854 nw
tri 12402 1741 12441 1780 se
rect 12441 1741 12476 1780
tri 12476 1741 12515 1780 nw
rect 12402 1363 12454 1741
tri 12454 1719 12476 1741 nw
tri 12454 1363 12476 1385 sw
tri 12402 1289 12476 1363 ne
tri 12476 1301 12538 1363 sw
rect 12476 1289 12538 1301
tri 12476 1279 12486 1289 ne
rect 12486 1161 12538 1289
tri 12538 1161 12614 1237 sw
tri 12018 1137 12026 1145 sw
rect 11966 1123 12026 1137
tri 11966 1109 11980 1123 ne
rect 11980 1109 12026 1123
tri 12026 1109 12054 1137 sw
rect 12486 1109 12492 1161
rect 12544 1109 12556 1161
rect 12608 1109 12614 1161
rect 10505 1090 10831 1092
rect 10505 1038 10511 1090
rect 10563 1076 10577 1090
rect 10629 1076 10643 1090
rect 10695 1076 10708 1090
rect 10760 1076 10773 1090
rect 10575 1038 10577 1076
rect 10760 1038 10763 1076
rect 10825 1038 10831 1090
tri 11351 1089 11354 1092 se
rect 11354 1089 11418 1092
tri 11583 1089 11603 1109 se
rect 11603 1089 11657 1109
tri 11657 1089 11677 1109 nw
tri 11980 1089 12000 1109 ne
rect 12000 1089 12054 1109
tri 12054 1089 12074 1109 sw
tri 11344 1082 11351 1089 se
rect 11351 1082 11418 1089
tri 11340 1078 11344 1082 se
rect 11344 1081 11417 1082
tri 11417 1081 11418 1082 nw
tri 11575 1081 11583 1089 se
rect 11583 1081 11646 1089
rect 11344 1078 11414 1081
tri 11414 1078 11417 1081 nw
tri 11572 1078 11575 1081 se
rect 11575 1078 11646 1081
tri 11646 1078 11657 1089 nw
tri 12000 1078 12011 1089 ne
rect 12011 1078 12074 1089
tri 12074 1078 12085 1089 sw
rect 12486 1078 12583 1109
tri 12583 1078 12614 1109 nw
rect 15076 1078 15251 1915
tri 15594 1628 15661 1695 se
rect 15661 1673 15713 1982
rect 15661 1628 15668 1673
tri 15668 1628 15713 1673 nw
rect 15594 1486 15650 1628
tri 15650 1610 15668 1628 nw
rect 15594 1404 15650 1430
rect 15594 1322 15650 1348
rect 15594 1257 15650 1266
tri 11316 1054 11340 1078 se
rect 11340 1054 11390 1078
tri 11390 1054 11414 1078 nw
tri 11548 1054 11572 1078 se
rect 11572 1054 11594 1078
rect 10505 1020 10519 1038
rect 10575 1020 10600 1038
rect 10656 1020 10681 1038
rect 10737 1020 10763 1038
rect 10819 1020 10831 1038
tri 11288 1026 11316 1054 se
rect 11316 1026 11362 1054
tri 11362 1026 11390 1054 nw
tri 11520 1026 11548 1054 se
rect 11548 1026 11594 1054
tri 11594 1026 11646 1078 nw
tri 12011 1063 12026 1078 ne
rect 12026 1063 12085 1078
tri 12085 1063 12100 1078 sw
tri 12026 1041 12048 1063 ne
rect 10505 1010 10831 1020
tri 11276 1014 11288 1026 se
rect 11288 1015 11351 1026
tri 11351 1015 11362 1026 nw
tri 11509 1015 11520 1026 se
rect 11520 1015 11583 1026
tri 11583 1015 11594 1026 nw
rect 11288 1014 11350 1015
tri 11350 1014 11351 1015 nw
tri 11508 1014 11509 1015 se
rect 11509 1014 11582 1015
tri 11582 1014 11583 1015 nw
rect 10505 958 10511 1010
rect 10563 994 10577 1010
rect 10629 994 10643 1010
rect 10695 994 10708 1010
rect 10760 994 10773 1010
rect 10575 958 10577 994
rect 10760 958 10763 994
rect 10825 958 10831 1010
tri 11242 980 11276 1014 se
rect 11276 980 11316 1014
tri 11316 980 11350 1014 nw
tri 11474 980 11508 1014 se
rect 11508 980 11545 1014
tri 11224 962 11242 980 se
rect 11242 962 11298 980
tri 11298 962 11316 980 nw
tri 11456 962 11474 980 se
rect 11474 962 11545 980
tri 11545 977 11582 1014 nw
tri 11220 958 11224 962 se
rect 11224 958 11294 962
tri 11294 958 11298 962 nw
tri 11452 958 11456 962 se
rect 11456 958 11545 962
rect 10505 938 10519 958
rect 10575 938 10600 958
rect 10656 938 10681 958
rect 10737 938 10763 958
rect 10819 938 10831 958
rect 10505 930 10831 938
rect 10505 878 10511 930
rect 10563 912 10577 930
rect 10629 912 10643 930
rect 10695 912 10708 930
rect 10760 912 10773 930
rect 10575 878 10577 912
rect 10760 878 10763 912
rect 10825 878 10831 930
rect 10505 856 10519 878
rect 10575 856 10600 878
rect 10656 856 10681 878
rect 10737 856 10763 878
rect 10819 856 10831 878
rect 10505 830 10831 856
rect 10505 774 10519 830
rect 10575 774 10600 830
rect 10656 774 10681 830
rect 10737 774 10763 830
rect 10819 774 10831 830
rect 10216 762 10268 768
rect 10216 692 10268 710
tri 10212 519 10216 523 se
rect 10216 519 10268 640
rect 10320 762 10372 768
rect 10320 692 10372 710
rect 10320 594 10372 640
rect 10505 748 10831 774
rect 10505 692 10519 748
rect 10575 692 10600 748
rect 10656 692 10681 748
rect 10737 692 10763 748
rect 10819 692 10831 748
rect 10505 666 10831 692
tri 10372 594 10389 611 sw
rect 10505 610 10519 666
rect 10575 610 10600 666
rect 10656 610 10681 666
rect 10737 610 10763 666
rect 10819 610 10831 666
rect 10320 589 10389 594
tri 10320 576 10333 589 ne
rect 10333 576 10389 589
tri 10389 576 10407 594 sw
rect 10505 584 10831 610
tri 11190 928 11220 958 se
rect 11220 928 11242 958
rect 11190 619 11242 928
tri 11242 906 11294 958 nw
tri 11410 916 11452 958 se
rect 11452 916 11545 958
rect 11410 776 11545 916
rect 11410 724 11416 776
rect 11468 724 11487 776
rect 11539 724 11545 776
rect 12048 818 12100 1063
tri 12100 818 12128 846 sw
rect 12048 786 12128 818
tri 12128 786 12160 818 sw
rect 12048 770 12160 786
tri 12160 770 12176 786 sw
rect 12048 718 12054 770
rect 12106 718 12118 770
rect 12170 718 12176 770
tri 11190 594 11215 619 ne
rect 11215 594 11242 619
tri 11242 594 11289 641 sw
tri 10333 564 10345 576 ne
rect 10345 564 10407 576
tri 10407 564 10419 576 sw
tri 10345 537 10372 564 ne
rect 10372 537 10419 564
tri 10419 537 10446 564 sw
tri 10372 519 10390 537 ne
rect 10390 519 10446 537
tri 10205 512 10212 519 se
rect 10212 515 10268 519
tri 10268 515 10272 519 sw
tri 10390 515 10394 519 ne
rect 10212 512 10272 515
tri 10272 512 10275 515 sw
tri 10199 506 10205 512 se
rect 10205 506 10275 512
tri 10275 506 10281 512 sw
tri 10191 498 10199 506 se
rect 10199 498 10281 506
tri 10281 498 10289 506 sw
tri 10179 486 10191 498 se
rect 10191 486 10289 498
tri 10289 486 10301 498 sw
tri 9977 483 9980 486 sw
tri 10176 483 10179 486 se
rect 10179 483 10301 486
tri 10301 483 10304 486 sw
tri 9880 431 9925 476 se
rect 9925 431 9980 483
tri 9980 431 10032 483 sw
rect 10176 431 10182 483
rect 10234 431 10246 483
rect 10298 431 10304 483
tri 9879 430 9880 431 se
rect 9880 430 10032 431
tri 10032 430 10033 431 sw
rect 9879 374 9888 430
rect 9944 374 9968 430
rect 10024 374 10033 430
tri 10392 339 10394 341 se
rect 10394 339 10446 519
rect 10505 528 10519 584
rect 10575 528 10600 584
rect 10656 528 10681 584
rect 10737 528 10763 584
rect 10819 528 10831 584
tri 11215 576 11233 594 ne
rect 11233 576 11289 594
tri 11289 576 11307 594 sw
tri 11233 570 11239 576 ne
rect 11239 570 11307 576
tri 11307 570 11313 576 sw
tri 11239 567 11242 570 ne
rect 11242 567 11942 570
tri 11242 564 11245 567 ne
rect 11245 564 11942 567
rect 10505 399 10831 528
tri 11245 518 11291 564 ne
rect 11291 518 11890 564
tri 11756 512 11762 518 ne
rect 11762 512 11890 518
tri 11762 506 11768 512 ne
rect 11768 506 11942 512
tri 11768 498 11776 506 ne
rect 11776 498 11942 506
tri 11776 446 11828 498 ne
rect 11828 446 11890 498
tri 11828 440 11834 446 ne
rect 11834 440 11942 446
tri 10505 383 10521 399 ne
rect 10521 383 10831 399
tri 10521 377 10527 383 ne
rect 10527 377 10831 383
tri 10527 370 10534 377 ne
rect 10534 370 10831 377
rect 12486 377 12538 1078
tri 12538 1033 12583 1078 nw
rect 15076 1026 15092 1078
rect 15144 1026 15193 1078
rect 15245 1026 15251 1078
rect 15076 1014 15251 1026
rect 15076 962 15092 1014
rect 15144 962 15193 1014
rect 15245 962 15251 1014
rect 15430 1046 15578 1047
rect 15430 994 15439 1046
rect 15491 994 15503 1046
rect 15555 994 15578 1046
rect 15430 958 15578 994
rect 15430 906 15439 958
rect 15491 906 15503 958
rect 15555 906 15578 958
rect 15430 870 15578 906
rect 15430 818 15439 870
rect 15491 818 15503 870
rect 15555 818 15578 870
rect 13655 786 13785 792
rect 13707 734 13733 786
rect 13655 716 13785 734
rect 13707 664 13733 716
rect 13655 646 13785 664
rect 13707 594 13733 646
rect 13655 576 13785 594
rect 15430 782 15578 818
rect 15430 730 15439 782
rect 15491 730 15503 782
rect 15555 730 15578 782
rect 13003 483 13012 539
rect 13068 483 13102 539
rect 13158 483 13419 539
rect 13707 524 13733 576
rect 13655 506 13785 524
tri 10534 339 10565 370 ne
rect 10565 339 10831 370
tri 10378 325 10392 339 se
rect 10392 337 10446 339
tri 10446 337 10448 339 sw
tri 10565 337 10567 339 ne
rect 10567 337 10831 339
tri 10831 337 10864 370 sw
rect 10392 325 10448 337
tri 10448 325 10460 337 sw
tri 10567 325 10579 337 ne
rect 10579 325 10864 337
tri 10864 325 10876 337 sw
tri 10366 313 10378 325 se
rect 10378 313 10460 325
tri 10460 313 10472 325 sw
tri 10579 313 10591 325 ne
rect 10591 313 10876 325
tri 10876 313 10888 325 sw
rect 12486 313 12538 325
tri 10346 293 10366 313 se
rect 10366 293 10472 313
tri 10472 293 10492 313 sw
rect 10338 237 10347 293
rect 10403 237 10427 293
rect 10483 237 10492 293
tri 10591 285 10619 313 ne
rect 10619 285 10888 313
tri 10888 285 10916 313 sw
tri 10619 261 10643 285 ne
rect 10643 261 10916 285
tri 10916 261 10940 285 sw
rect 13707 454 13733 506
tri 10643 237 10667 261 ne
rect 10667 255 10940 261
tri 10940 255 10946 261 sw
rect 12486 255 12538 261
rect 10667 237 10946 255
tri 10667 210 10694 237 ne
rect 10694 210 10946 237
tri 10946 210 10991 255 sw
rect 13308 239 13317 295
rect 13373 239 13407 295
rect 13463 239 13472 295
tri 13308 210 13337 239 ne
rect 13337 210 13419 239
tri 10694 180 10724 210 ne
rect 10724 180 13040 210
tri 13337 180 13367 210 ne
tri 10724 165 10739 180 ne
rect 10739 165 12881 180
rect 9918 109 9927 165
rect 9983 109 10007 165
rect 10063 109 10072 165
tri 10739 128 10776 165 ne
rect 10776 128 12881 165
rect 12933 128 12982 180
rect 13034 128 13040 180
tri 9918 104 9923 109 ne
rect 9923 104 10067 109
tri 10067 104 10072 109 nw
tri 10776 104 10800 128 ne
rect 10800 104 13040 128
tri 9923 73 9954 104 ne
rect 9954 73 10036 104
tri 10036 73 10067 104 nw
tri 10800 73 10831 104 ne
rect 10831 73 12881 104
tri 9954 56 9971 73 ne
rect 9971 0 10023 73
tri 10023 60 10036 73 nw
tri 10831 60 10844 73 ne
rect 10844 60 12881 73
tri 10844 52 10852 60 ne
rect 10852 52 12881 60
rect 12933 52 12982 104
rect 13034 52 13040 104
tri 10852 50 10854 52 ne
rect 10854 50 13040 52
rect 13367 0 13419 210
tri 13419 186 13472 239 nw
rect 13655 0 13785 454
tri 15256 411 15430 585 se
rect 15430 519 15578 730
rect 15430 411 15470 519
tri 15470 411 15578 519 nw
rect 15256 0 15384 411
tri 15384 325 15470 411 nw
rect 15478 237 15487 293
rect 15543 237 15577 293
rect 15633 237 15642 293
tri 15741 243 15742 244 se
rect 15742 243 15782 2053
tri 15482 197 15522 237 ne
rect 15522 197 15596 237
tri 15596 197 15636 237 nw
rect 15741 226 15782 243
rect 15522 0 15574 197
tri 15574 175 15596 197 nw
rect 15741 0 15781 226
tri 15781 225 15782 226 nw
rect 15943 0 15983 19200
<< via2 >>
rect 1361 39894 1417 39950
rect 1443 39894 1499 39950
rect 1525 39894 1581 39950
rect 1607 39894 1663 39950
rect 1689 39894 1745 39950
rect 1903 39939 1959 39995
rect 1984 39939 2040 39995
rect 2065 39939 2121 39995
rect 2146 39939 2202 39995
rect 2227 39939 2283 39995
rect 2308 39939 2364 39995
rect 2389 39939 2445 39995
rect 2470 39939 2526 39995
rect 2551 39939 2607 39995
rect 2632 39939 2688 39995
rect 2713 39939 2769 39995
rect 2794 39939 2850 39995
rect 2875 39939 2931 39995
rect 2956 39939 3012 39995
rect 3037 39939 3093 39995
rect 3118 39994 11334 39995
rect 3118 39942 3160 39994
rect 3160 39942 3212 39994
rect 3212 39942 3225 39994
rect 3225 39942 3277 39994
rect 3277 39942 3290 39994
rect 3290 39942 3342 39994
rect 3342 39942 3355 39994
rect 3355 39942 3407 39994
rect 3407 39942 3420 39994
rect 3420 39942 3472 39994
rect 3472 39942 3485 39994
rect 3485 39942 3537 39994
rect 3537 39942 3550 39994
rect 3550 39942 3602 39994
rect 3602 39942 3615 39994
rect 3615 39942 3667 39994
rect 3667 39942 3680 39994
rect 3680 39942 3732 39994
rect 3732 39942 3745 39994
rect 3745 39942 3797 39994
rect 3797 39942 3810 39994
rect 3810 39942 3862 39994
rect 3862 39942 3875 39994
rect 3875 39942 3927 39994
rect 3927 39942 3940 39994
rect 3940 39942 3992 39994
rect 3992 39942 4005 39994
rect 4005 39942 4057 39994
rect 4057 39942 4070 39994
rect 4070 39942 4122 39994
rect 4122 39942 4135 39994
rect 4135 39942 4187 39994
rect 4187 39942 4200 39994
rect 4200 39942 4252 39994
rect 4252 39942 4265 39994
rect 4265 39942 4317 39994
rect 4317 39942 4330 39994
rect 4330 39942 4382 39994
rect 4382 39942 4395 39994
rect 4395 39942 4447 39994
rect 4447 39942 4460 39994
rect 4460 39942 4512 39994
rect 4512 39942 4525 39994
rect 4525 39942 4577 39994
rect 4577 39942 4590 39994
rect 4590 39942 4642 39994
rect 4642 39942 4655 39994
rect 4655 39942 4707 39994
rect 4707 39942 4720 39994
rect 4720 39942 4772 39994
rect 4772 39942 4785 39994
rect 4785 39942 4837 39994
rect 4837 39942 4850 39994
rect 4850 39942 4902 39994
rect 4902 39942 4915 39994
rect 4915 39942 4967 39994
rect 4967 39942 4980 39994
rect 4980 39942 5032 39994
rect 5032 39942 5045 39994
rect 5045 39942 5097 39994
rect 5097 39942 5110 39994
rect 5110 39942 5162 39994
rect 5162 39942 5175 39994
rect 5175 39942 5227 39994
rect 5227 39942 5240 39994
rect 5240 39942 5292 39994
rect 5292 39942 5305 39994
rect 5305 39942 5357 39994
rect 5357 39942 5370 39994
rect 5370 39942 5422 39994
rect 5422 39942 5435 39994
rect 5435 39942 5487 39994
rect 5487 39942 5500 39994
rect 5500 39942 5552 39994
rect 5552 39942 5565 39994
rect 5565 39942 5617 39994
rect 5617 39942 5630 39994
rect 5630 39942 5682 39994
rect 5682 39942 5695 39994
rect 5695 39942 5747 39994
rect 5747 39942 5760 39994
rect 5760 39942 5812 39994
rect 5812 39942 5825 39994
rect 5825 39942 5877 39994
rect 5877 39942 5890 39994
rect 5890 39942 5942 39994
rect 5942 39942 5955 39994
rect 5955 39942 6007 39994
rect 6007 39942 6020 39994
rect 6020 39942 6072 39994
rect 6072 39942 6085 39994
rect 6085 39942 6137 39994
rect 6137 39942 6150 39994
rect 6150 39942 6202 39994
rect 6202 39942 6215 39994
rect 6215 39942 6267 39994
rect 6267 39942 6280 39994
rect 6280 39942 6332 39994
rect 6332 39942 6345 39994
rect 6345 39942 6397 39994
rect 6397 39942 6410 39994
rect 6410 39942 6462 39994
rect 6462 39942 6475 39994
rect 6475 39942 6527 39994
rect 6527 39942 6540 39994
rect 6540 39942 6592 39994
rect 6592 39942 6605 39994
rect 6605 39942 6657 39994
rect 6657 39942 6670 39994
rect 6670 39942 6722 39994
rect 6722 39942 6735 39994
rect 6735 39942 6787 39994
rect 6787 39942 6800 39994
rect 6800 39942 6852 39994
rect 6852 39942 6865 39994
rect 6865 39942 6917 39994
rect 6917 39942 6930 39994
rect 6930 39942 6982 39994
rect 6982 39942 6995 39994
rect 6995 39942 7047 39994
rect 7047 39942 7060 39994
rect 7060 39942 7112 39994
rect 7112 39942 7125 39994
rect 7125 39942 7177 39994
rect 7177 39942 7189 39994
rect 7189 39942 7241 39994
rect 7241 39942 7253 39994
rect 7253 39942 7305 39994
rect 7305 39942 7317 39994
rect 7317 39942 7369 39994
rect 7369 39942 7381 39994
rect 7381 39942 7433 39994
rect 7433 39942 7445 39994
rect 7445 39942 7497 39994
rect 7497 39942 7509 39994
rect 7509 39942 7561 39994
rect 7561 39942 7573 39994
rect 7573 39942 7625 39994
rect 7625 39942 7637 39994
rect 7637 39942 7689 39994
rect 7689 39942 7701 39994
rect 7701 39942 7753 39994
rect 7753 39942 7765 39994
rect 7765 39942 7817 39994
rect 7817 39942 7829 39994
rect 7829 39942 7881 39994
rect 7881 39942 7893 39994
rect 7893 39942 7945 39994
rect 7945 39942 7957 39994
rect 7957 39942 8009 39994
rect 8009 39942 8021 39994
rect 8021 39942 8073 39994
rect 8073 39942 8085 39994
rect 8085 39942 8137 39994
rect 8137 39942 8149 39994
rect 8149 39942 8201 39994
rect 8201 39942 8213 39994
rect 8213 39942 8265 39994
rect 8265 39942 8277 39994
rect 8277 39942 8329 39994
rect 8329 39942 8341 39994
rect 8341 39942 8393 39994
rect 8393 39942 8405 39994
rect 8405 39942 8457 39994
rect 8457 39942 8469 39994
rect 8469 39942 8521 39994
rect 8521 39942 8533 39994
rect 8533 39942 8585 39994
rect 8585 39942 8597 39994
rect 8597 39942 8649 39994
rect 8649 39942 8661 39994
rect 8661 39942 8713 39994
rect 8713 39942 8725 39994
rect 8725 39942 8777 39994
rect 8777 39942 8789 39994
rect 8789 39942 8841 39994
rect 8841 39942 8853 39994
rect 8853 39942 8905 39994
rect 8905 39942 8917 39994
rect 8917 39942 8969 39994
rect 8969 39942 8981 39994
rect 8981 39942 9033 39994
rect 9033 39942 9045 39994
rect 9045 39942 9097 39994
rect 9097 39942 9109 39994
rect 9109 39942 9161 39994
rect 9161 39942 9173 39994
rect 9173 39942 9225 39994
rect 9225 39942 9237 39994
rect 9237 39942 9289 39994
rect 9289 39942 9301 39994
rect 9301 39942 9353 39994
rect 9353 39942 9365 39994
rect 9365 39942 9417 39994
rect 9417 39942 9429 39994
rect 9429 39942 9481 39994
rect 9481 39942 9493 39994
rect 9493 39942 9545 39994
rect 9545 39942 9557 39994
rect 9557 39942 9609 39994
rect 9609 39942 9621 39994
rect 9621 39942 9673 39994
rect 9673 39942 9685 39994
rect 9685 39942 9737 39994
rect 9737 39942 9749 39994
rect 9749 39942 9801 39994
rect 9801 39942 9813 39994
rect 9813 39942 9865 39994
rect 9865 39942 9877 39994
rect 9877 39942 9929 39994
rect 9929 39942 9941 39994
rect 9941 39942 9993 39994
rect 9993 39942 10005 39994
rect 10005 39942 10057 39994
rect 10057 39942 10069 39994
rect 10069 39942 10121 39994
rect 10121 39942 10133 39994
rect 10133 39942 10185 39994
rect 10185 39942 10197 39994
rect 10197 39942 10249 39994
rect 10249 39942 10261 39994
rect 10261 39942 10313 39994
rect 10313 39942 10325 39994
rect 10325 39942 10377 39994
rect 10377 39942 10389 39994
rect 10389 39942 10441 39994
rect 10441 39942 10453 39994
rect 10453 39942 10505 39994
rect 10505 39942 10517 39994
rect 10517 39942 10569 39994
rect 10569 39942 10581 39994
rect 10581 39942 10633 39994
rect 10633 39942 10645 39994
rect 10645 39942 10697 39994
rect 10697 39942 10709 39994
rect 10709 39942 10761 39994
rect 10761 39942 10773 39994
rect 10773 39942 10825 39994
rect 10825 39942 10837 39994
rect 10837 39942 10889 39994
rect 10889 39942 10901 39994
rect 10901 39942 10953 39994
rect 10953 39942 10965 39994
rect 10965 39942 11017 39994
rect 11017 39942 11029 39994
rect 11029 39942 11081 39994
rect 11081 39942 11093 39994
rect 11093 39942 11145 39994
rect 11145 39942 11157 39994
rect 11157 39942 11209 39994
rect 11209 39942 11221 39994
rect 11221 39942 11273 39994
rect 11273 39942 11285 39994
rect 11285 39942 11334 39994
rect 3118 39926 11334 39942
rect 1361 39812 1417 39868
rect 1443 39812 1499 39868
rect 1525 39812 1581 39868
rect 1607 39812 1663 39868
rect 1689 39812 1745 39868
rect 1903 39859 1959 39915
rect 1984 39859 2040 39915
rect 2065 39859 2121 39915
rect 2146 39859 2202 39915
rect 2227 39859 2283 39915
rect 2308 39859 2364 39915
rect 2389 39859 2445 39915
rect 2470 39859 2526 39915
rect 2551 39859 2607 39915
rect 2632 39859 2688 39915
rect 2713 39859 2769 39915
rect 2794 39859 2850 39915
rect 2875 39859 2931 39915
rect 2956 39859 3012 39915
rect 3037 39859 3093 39915
rect 3118 39874 3160 39926
rect 3160 39874 3212 39926
rect 3212 39874 3225 39926
rect 3225 39874 3277 39926
rect 3277 39874 3290 39926
rect 3290 39874 3342 39926
rect 3342 39874 3355 39926
rect 3355 39874 3407 39926
rect 3407 39874 3420 39926
rect 3420 39874 3472 39926
rect 3472 39874 3485 39926
rect 3485 39874 3537 39926
rect 3537 39874 3550 39926
rect 3550 39874 3602 39926
rect 3602 39874 3615 39926
rect 3615 39874 3667 39926
rect 3667 39874 3680 39926
rect 3680 39874 3732 39926
rect 3732 39874 3745 39926
rect 3745 39874 3797 39926
rect 3797 39874 3810 39926
rect 3810 39874 3862 39926
rect 3862 39874 3875 39926
rect 3875 39874 3927 39926
rect 3927 39874 3940 39926
rect 3940 39874 3992 39926
rect 3992 39874 4005 39926
rect 4005 39874 4057 39926
rect 4057 39874 4070 39926
rect 4070 39874 4122 39926
rect 4122 39874 4135 39926
rect 4135 39874 4187 39926
rect 4187 39874 4200 39926
rect 4200 39874 4252 39926
rect 4252 39874 4265 39926
rect 4265 39874 4317 39926
rect 4317 39874 4330 39926
rect 4330 39874 4382 39926
rect 4382 39874 4395 39926
rect 4395 39874 4447 39926
rect 4447 39874 4460 39926
rect 4460 39874 4512 39926
rect 4512 39874 4525 39926
rect 4525 39874 4577 39926
rect 4577 39874 4590 39926
rect 4590 39874 4642 39926
rect 4642 39874 4655 39926
rect 4655 39874 4707 39926
rect 4707 39874 4720 39926
rect 4720 39874 4772 39926
rect 4772 39874 4785 39926
rect 4785 39874 4837 39926
rect 4837 39874 4850 39926
rect 4850 39874 4902 39926
rect 4902 39874 4915 39926
rect 4915 39874 4967 39926
rect 4967 39874 4980 39926
rect 4980 39874 5032 39926
rect 5032 39874 5045 39926
rect 5045 39874 5097 39926
rect 5097 39874 5110 39926
rect 5110 39874 5162 39926
rect 5162 39874 5175 39926
rect 5175 39874 5227 39926
rect 5227 39874 5240 39926
rect 5240 39874 5292 39926
rect 5292 39874 5305 39926
rect 5305 39874 5357 39926
rect 5357 39874 5370 39926
rect 5370 39874 5422 39926
rect 5422 39874 5435 39926
rect 5435 39874 5487 39926
rect 5487 39874 5500 39926
rect 5500 39874 5552 39926
rect 5552 39874 5565 39926
rect 5565 39874 5617 39926
rect 5617 39874 5630 39926
rect 5630 39874 5682 39926
rect 5682 39874 5695 39926
rect 5695 39874 5747 39926
rect 5747 39874 5760 39926
rect 5760 39874 5812 39926
rect 5812 39874 5825 39926
rect 5825 39874 5877 39926
rect 5877 39874 5890 39926
rect 5890 39874 5942 39926
rect 5942 39874 5955 39926
rect 5955 39874 6007 39926
rect 6007 39874 6020 39926
rect 6020 39874 6072 39926
rect 6072 39874 6085 39926
rect 6085 39874 6137 39926
rect 6137 39874 6150 39926
rect 6150 39874 6202 39926
rect 6202 39874 6215 39926
rect 6215 39874 6267 39926
rect 6267 39874 6280 39926
rect 6280 39874 6332 39926
rect 6332 39874 6345 39926
rect 6345 39874 6397 39926
rect 6397 39874 6410 39926
rect 6410 39874 6462 39926
rect 6462 39874 6475 39926
rect 6475 39874 6527 39926
rect 6527 39874 6540 39926
rect 6540 39874 6592 39926
rect 6592 39874 6605 39926
rect 6605 39874 6657 39926
rect 6657 39874 6670 39926
rect 6670 39874 6722 39926
rect 6722 39874 6735 39926
rect 6735 39874 6787 39926
rect 6787 39874 6800 39926
rect 6800 39874 6852 39926
rect 6852 39874 6865 39926
rect 6865 39874 6917 39926
rect 6917 39874 6930 39926
rect 6930 39874 6982 39926
rect 6982 39874 6995 39926
rect 6995 39874 7047 39926
rect 7047 39874 7060 39926
rect 7060 39874 7112 39926
rect 7112 39874 7125 39926
rect 7125 39874 7177 39926
rect 7177 39874 7189 39926
rect 7189 39874 7241 39926
rect 7241 39874 7253 39926
rect 7253 39874 7305 39926
rect 7305 39874 7317 39926
rect 7317 39874 7369 39926
rect 7369 39874 7381 39926
rect 7381 39874 7433 39926
rect 7433 39874 7445 39926
rect 7445 39874 7497 39926
rect 7497 39874 7509 39926
rect 7509 39874 7561 39926
rect 7561 39874 7573 39926
rect 7573 39874 7625 39926
rect 7625 39874 7637 39926
rect 7637 39874 7689 39926
rect 7689 39874 7701 39926
rect 7701 39874 7753 39926
rect 7753 39874 7765 39926
rect 7765 39874 7817 39926
rect 7817 39874 7829 39926
rect 7829 39874 7881 39926
rect 7881 39874 7893 39926
rect 7893 39874 7945 39926
rect 7945 39874 7957 39926
rect 7957 39874 8009 39926
rect 8009 39874 8021 39926
rect 8021 39874 8073 39926
rect 8073 39874 8085 39926
rect 8085 39874 8137 39926
rect 8137 39874 8149 39926
rect 8149 39874 8201 39926
rect 8201 39874 8213 39926
rect 8213 39874 8265 39926
rect 8265 39874 8277 39926
rect 8277 39874 8329 39926
rect 8329 39874 8341 39926
rect 8341 39874 8393 39926
rect 8393 39874 8405 39926
rect 8405 39874 8457 39926
rect 8457 39874 8469 39926
rect 8469 39874 8521 39926
rect 8521 39874 8533 39926
rect 8533 39874 8585 39926
rect 8585 39874 8597 39926
rect 8597 39874 8649 39926
rect 8649 39874 8661 39926
rect 8661 39874 8713 39926
rect 8713 39874 8725 39926
rect 8725 39874 8777 39926
rect 8777 39874 8789 39926
rect 8789 39874 8841 39926
rect 8841 39874 8853 39926
rect 8853 39874 8905 39926
rect 8905 39874 8917 39926
rect 8917 39874 8969 39926
rect 8969 39874 8981 39926
rect 8981 39874 9033 39926
rect 9033 39874 9045 39926
rect 9045 39874 9097 39926
rect 9097 39874 9109 39926
rect 9109 39874 9161 39926
rect 9161 39874 9173 39926
rect 9173 39874 9225 39926
rect 9225 39874 9237 39926
rect 9237 39874 9289 39926
rect 9289 39874 9301 39926
rect 9301 39874 9353 39926
rect 9353 39874 9365 39926
rect 9365 39874 9417 39926
rect 9417 39874 9429 39926
rect 9429 39874 9481 39926
rect 9481 39874 9493 39926
rect 9493 39874 9545 39926
rect 9545 39874 9557 39926
rect 9557 39874 9609 39926
rect 9609 39874 9621 39926
rect 9621 39874 9673 39926
rect 9673 39874 9685 39926
rect 9685 39874 9737 39926
rect 9737 39874 9749 39926
rect 9749 39874 9801 39926
rect 9801 39874 9813 39926
rect 9813 39874 9865 39926
rect 9865 39874 9877 39926
rect 9877 39874 9929 39926
rect 9929 39874 9941 39926
rect 9941 39874 9993 39926
rect 9993 39874 10005 39926
rect 10005 39874 10057 39926
rect 10057 39874 10069 39926
rect 10069 39874 10121 39926
rect 10121 39874 10133 39926
rect 10133 39874 10185 39926
rect 10185 39874 10197 39926
rect 10197 39874 10249 39926
rect 10249 39874 10261 39926
rect 10261 39874 10313 39926
rect 10313 39874 10325 39926
rect 10325 39874 10377 39926
rect 10377 39874 10389 39926
rect 10389 39874 10441 39926
rect 10441 39874 10453 39926
rect 10453 39874 10505 39926
rect 10505 39874 10517 39926
rect 10517 39874 10569 39926
rect 10569 39874 10581 39926
rect 10581 39874 10633 39926
rect 10633 39874 10645 39926
rect 10645 39874 10697 39926
rect 10697 39874 10709 39926
rect 10709 39874 10761 39926
rect 10761 39874 10773 39926
rect 10773 39874 10825 39926
rect 10825 39874 10837 39926
rect 10837 39874 10889 39926
rect 10889 39874 10901 39926
rect 10901 39874 10953 39926
rect 10953 39874 10965 39926
rect 10965 39874 11017 39926
rect 11017 39874 11029 39926
rect 11029 39874 11081 39926
rect 11081 39874 11093 39926
rect 11093 39874 11145 39926
rect 11145 39874 11157 39926
rect 11157 39874 11209 39926
rect 11209 39874 11221 39926
rect 11221 39874 11273 39926
rect 11273 39874 11285 39926
rect 11285 39874 11334 39926
rect 3118 39858 11334 39874
rect 1361 39730 1417 39786
rect 1443 39730 1499 39786
rect 1525 39730 1581 39786
rect 1607 39730 1663 39786
rect 1689 39730 1745 39786
rect 1903 39779 1959 39835
rect 1984 39779 2040 39835
rect 2065 39779 2121 39835
rect 2146 39779 2202 39835
rect 2227 39779 2283 39835
rect 2308 39779 2364 39835
rect 2389 39779 2445 39835
rect 2470 39779 2526 39835
rect 2551 39779 2607 39835
rect 2632 39779 2688 39835
rect 2713 39779 2769 39835
rect 2794 39779 2850 39835
rect 2875 39779 2931 39835
rect 2956 39779 3012 39835
rect 3037 39779 3093 39835
rect 3118 39806 3160 39858
rect 3160 39806 3212 39858
rect 3212 39806 3225 39858
rect 3225 39806 3277 39858
rect 3277 39806 3290 39858
rect 3290 39806 3342 39858
rect 3342 39806 3355 39858
rect 3355 39806 3407 39858
rect 3407 39806 3420 39858
rect 3420 39806 3472 39858
rect 3472 39806 3485 39858
rect 3485 39806 3537 39858
rect 3537 39806 3550 39858
rect 3550 39806 3602 39858
rect 3602 39806 3615 39858
rect 3615 39806 3667 39858
rect 3667 39806 3680 39858
rect 3680 39806 3732 39858
rect 3732 39806 3745 39858
rect 3745 39806 3797 39858
rect 3797 39806 3810 39858
rect 3810 39806 3862 39858
rect 3862 39806 3875 39858
rect 3875 39806 3927 39858
rect 3927 39806 3940 39858
rect 3940 39806 3992 39858
rect 3992 39806 4005 39858
rect 4005 39806 4057 39858
rect 4057 39806 4070 39858
rect 4070 39806 4122 39858
rect 4122 39806 4135 39858
rect 4135 39806 4187 39858
rect 4187 39806 4200 39858
rect 4200 39806 4252 39858
rect 4252 39806 4265 39858
rect 4265 39806 4317 39858
rect 4317 39806 4330 39858
rect 4330 39806 4382 39858
rect 4382 39806 4395 39858
rect 4395 39806 4447 39858
rect 4447 39806 4460 39858
rect 4460 39806 4512 39858
rect 4512 39806 4525 39858
rect 4525 39806 4577 39858
rect 4577 39806 4590 39858
rect 4590 39806 4642 39858
rect 4642 39806 4655 39858
rect 4655 39806 4707 39858
rect 4707 39806 4720 39858
rect 4720 39806 4772 39858
rect 4772 39806 4785 39858
rect 4785 39806 4837 39858
rect 4837 39806 4850 39858
rect 4850 39806 4902 39858
rect 4902 39806 4915 39858
rect 4915 39806 4967 39858
rect 4967 39806 4980 39858
rect 4980 39806 5032 39858
rect 5032 39806 5045 39858
rect 5045 39806 5097 39858
rect 5097 39806 5110 39858
rect 5110 39806 5162 39858
rect 5162 39806 5175 39858
rect 5175 39806 5227 39858
rect 5227 39806 5240 39858
rect 5240 39806 5292 39858
rect 5292 39806 5305 39858
rect 5305 39806 5357 39858
rect 5357 39806 5370 39858
rect 5370 39806 5422 39858
rect 5422 39806 5435 39858
rect 5435 39806 5487 39858
rect 5487 39806 5500 39858
rect 5500 39806 5552 39858
rect 5552 39806 5565 39858
rect 5565 39806 5617 39858
rect 5617 39806 5630 39858
rect 5630 39806 5682 39858
rect 5682 39806 5695 39858
rect 5695 39806 5747 39858
rect 5747 39806 5760 39858
rect 5760 39806 5812 39858
rect 5812 39806 5825 39858
rect 5825 39806 5877 39858
rect 5877 39806 5890 39858
rect 5890 39806 5942 39858
rect 5942 39806 5955 39858
rect 5955 39806 6007 39858
rect 6007 39806 6020 39858
rect 6020 39806 6072 39858
rect 6072 39806 6085 39858
rect 6085 39806 6137 39858
rect 6137 39806 6150 39858
rect 6150 39806 6202 39858
rect 6202 39806 6215 39858
rect 6215 39806 6267 39858
rect 6267 39806 6280 39858
rect 6280 39806 6332 39858
rect 6332 39806 6345 39858
rect 6345 39806 6397 39858
rect 6397 39806 6410 39858
rect 6410 39806 6462 39858
rect 6462 39806 6475 39858
rect 6475 39806 6527 39858
rect 6527 39806 6540 39858
rect 6540 39806 6592 39858
rect 6592 39806 6605 39858
rect 6605 39806 6657 39858
rect 6657 39806 6670 39858
rect 6670 39806 6722 39858
rect 6722 39806 6735 39858
rect 6735 39806 6787 39858
rect 6787 39806 6800 39858
rect 6800 39806 6852 39858
rect 6852 39806 6865 39858
rect 6865 39806 6917 39858
rect 6917 39806 6930 39858
rect 6930 39806 6982 39858
rect 6982 39806 6995 39858
rect 6995 39806 7047 39858
rect 7047 39806 7060 39858
rect 7060 39806 7112 39858
rect 7112 39806 7125 39858
rect 7125 39806 7177 39858
rect 7177 39806 7189 39858
rect 7189 39806 7241 39858
rect 7241 39806 7253 39858
rect 7253 39806 7305 39858
rect 7305 39806 7317 39858
rect 7317 39806 7369 39858
rect 7369 39806 7381 39858
rect 7381 39806 7433 39858
rect 7433 39806 7445 39858
rect 7445 39806 7497 39858
rect 7497 39806 7509 39858
rect 7509 39806 7561 39858
rect 7561 39806 7573 39858
rect 7573 39806 7625 39858
rect 7625 39806 7637 39858
rect 7637 39806 7689 39858
rect 7689 39806 7701 39858
rect 7701 39806 7753 39858
rect 7753 39806 7765 39858
rect 7765 39806 7817 39858
rect 7817 39806 7829 39858
rect 7829 39806 7881 39858
rect 7881 39806 7893 39858
rect 7893 39806 7945 39858
rect 7945 39806 7957 39858
rect 7957 39806 8009 39858
rect 8009 39806 8021 39858
rect 8021 39806 8073 39858
rect 8073 39806 8085 39858
rect 8085 39806 8137 39858
rect 8137 39806 8149 39858
rect 8149 39806 8201 39858
rect 8201 39806 8213 39858
rect 8213 39806 8265 39858
rect 8265 39806 8277 39858
rect 8277 39806 8329 39858
rect 8329 39806 8341 39858
rect 8341 39806 8393 39858
rect 8393 39806 8405 39858
rect 8405 39806 8457 39858
rect 8457 39806 8469 39858
rect 8469 39806 8521 39858
rect 8521 39806 8533 39858
rect 8533 39806 8585 39858
rect 8585 39806 8597 39858
rect 8597 39806 8649 39858
rect 8649 39806 8661 39858
rect 8661 39806 8713 39858
rect 8713 39806 8725 39858
rect 8725 39806 8777 39858
rect 8777 39806 8789 39858
rect 8789 39806 8841 39858
rect 8841 39806 8853 39858
rect 8853 39806 8905 39858
rect 8905 39806 8917 39858
rect 8917 39806 8969 39858
rect 8969 39806 8981 39858
rect 8981 39806 9033 39858
rect 9033 39806 9045 39858
rect 9045 39806 9097 39858
rect 9097 39806 9109 39858
rect 9109 39806 9161 39858
rect 9161 39806 9173 39858
rect 9173 39806 9225 39858
rect 9225 39806 9237 39858
rect 9237 39806 9289 39858
rect 9289 39806 9301 39858
rect 9301 39806 9353 39858
rect 9353 39806 9365 39858
rect 9365 39806 9417 39858
rect 9417 39806 9429 39858
rect 9429 39806 9481 39858
rect 9481 39806 9493 39858
rect 9493 39806 9545 39858
rect 9545 39806 9557 39858
rect 9557 39806 9609 39858
rect 9609 39806 9621 39858
rect 9621 39806 9673 39858
rect 9673 39806 9685 39858
rect 9685 39806 9737 39858
rect 9737 39806 9749 39858
rect 9749 39806 9801 39858
rect 9801 39806 9813 39858
rect 9813 39806 9865 39858
rect 9865 39806 9877 39858
rect 9877 39806 9929 39858
rect 9929 39806 9941 39858
rect 9941 39806 9993 39858
rect 9993 39806 10005 39858
rect 10005 39806 10057 39858
rect 10057 39806 10069 39858
rect 10069 39806 10121 39858
rect 10121 39806 10133 39858
rect 10133 39806 10185 39858
rect 10185 39806 10197 39858
rect 10197 39806 10249 39858
rect 10249 39806 10261 39858
rect 10261 39806 10313 39858
rect 10313 39806 10325 39858
rect 10325 39806 10377 39858
rect 10377 39806 10389 39858
rect 10389 39806 10441 39858
rect 10441 39806 10453 39858
rect 10453 39806 10505 39858
rect 10505 39806 10517 39858
rect 10517 39806 10569 39858
rect 10569 39806 10581 39858
rect 10581 39806 10633 39858
rect 10633 39806 10645 39858
rect 10645 39806 10697 39858
rect 10697 39806 10709 39858
rect 10709 39806 10761 39858
rect 10761 39806 10773 39858
rect 10773 39806 10825 39858
rect 10825 39806 10837 39858
rect 10837 39806 10889 39858
rect 10889 39806 10901 39858
rect 10901 39806 10953 39858
rect 10953 39806 10965 39858
rect 10965 39806 11017 39858
rect 11017 39806 11029 39858
rect 11029 39806 11081 39858
rect 11081 39806 11093 39858
rect 11093 39806 11145 39858
rect 11145 39806 11157 39858
rect 11157 39806 11209 39858
rect 11209 39806 11221 39858
rect 11221 39806 11273 39858
rect 11273 39806 11285 39858
rect 11285 39806 11334 39858
rect 3118 39790 11334 39806
rect 1361 39648 1417 39704
rect 1443 39648 1499 39704
rect 1525 39648 1581 39704
rect 1607 39648 1663 39704
rect 1689 39648 1745 39704
rect 1903 39699 1959 39755
rect 1984 39699 2040 39755
rect 2065 39699 2121 39755
rect 2146 39699 2202 39755
rect 2227 39699 2283 39755
rect 2308 39699 2364 39755
rect 2389 39699 2445 39755
rect 2470 39699 2526 39755
rect 2551 39699 2607 39755
rect 2632 39699 2688 39755
rect 2713 39699 2769 39755
rect 2794 39699 2850 39755
rect 2875 39699 2931 39755
rect 2956 39699 3012 39755
rect 3037 39699 3093 39755
rect 3118 39738 3160 39790
rect 3160 39738 3212 39790
rect 3212 39738 3225 39790
rect 3225 39738 3277 39790
rect 3277 39738 3290 39790
rect 3290 39738 3342 39790
rect 3342 39738 3355 39790
rect 3355 39738 3407 39790
rect 3407 39738 3420 39790
rect 3420 39738 3472 39790
rect 3472 39738 3485 39790
rect 3485 39738 3537 39790
rect 3537 39738 3550 39790
rect 3550 39738 3602 39790
rect 3602 39738 3615 39790
rect 3615 39738 3667 39790
rect 3667 39738 3680 39790
rect 3680 39738 3732 39790
rect 3732 39738 3745 39790
rect 3745 39738 3797 39790
rect 3797 39738 3810 39790
rect 3810 39738 3862 39790
rect 3862 39738 3875 39790
rect 3875 39738 3927 39790
rect 3927 39738 3940 39790
rect 3940 39738 3992 39790
rect 3992 39738 4005 39790
rect 4005 39738 4057 39790
rect 4057 39738 4070 39790
rect 4070 39738 4122 39790
rect 4122 39738 4135 39790
rect 4135 39738 4187 39790
rect 4187 39738 4200 39790
rect 4200 39738 4252 39790
rect 4252 39738 4265 39790
rect 4265 39738 4317 39790
rect 4317 39738 4330 39790
rect 4330 39738 4382 39790
rect 4382 39738 4395 39790
rect 4395 39738 4447 39790
rect 4447 39738 4460 39790
rect 4460 39738 4512 39790
rect 4512 39738 4525 39790
rect 4525 39738 4577 39790
rect 4577 39738 4590 39790
rect 4590 39738 4642 39790
rect 4642 39738 4655 39790
rect 4655 39738 4707 39790
rect 4707 39738 4720 39790
rect 4720 39738 4772 39790
rect 4772 39738 4785 39790
rect 4785 39738 4837 39790
rect 4837 39738 4850 39790
rect 4850 39738 4902 39790
rect 4902 39738 4915 39790
rect 4915 39738 4967 39790
rect 4967 39738 4980 39790
rect 4980 39738 5032 39790
rect 5032 39738 5045 39790
rect 5045 39738 5097 39790
rect 5097 39738 5110 39790
rect 5110 39738 5162 39790
rect 5162 39738 5175 39790
rect 5175 39738 5227 39790
rect 5227 39738 5240 39790
rect 5240 39738 5292 39790
rect 5292 39738 5305 39790
rect 5305 39738 5357 39790
rect 5357 39738 5370 39790
rect 5370 39738 5422 39790
rect 5422 39738 5435 39790
rect 5435 39738 5487 39790
rect 5487 39738 5500 39790
rect 5500 39738 5552 39790
rect 5552 39738 5565 39790
rect 5565 39738 5617 39790
rect 5617 39738 5630 39790
rect 5630 39738 5682 39790
rect 5682 39738 5695 39790
rect 5695 39738 5747 39790
rect 5747 39738 5760 39790
rect 5760 39738 5812 39790
rect 5812 39738 5825 39790
rect 5825 39738 5877 39790
rect 5877 39738 5890 39790
rect 5890 39738 5942 39790
rect 5942 39738 5955 39790
rect 5955 39738 6007 39790
rect 6007 39738 6020 39790
rect 6020 39738 6072 39790
rect 6072 39738 6085 39790
rect 6085 39738 6137 39790
rect 6137 39738 6150 39790
rect 6150 39738 6202 39790
rect 6202 39738 6215 39790
rect 6215 39738 6267 39790
rect 6267 39738 6280 39790
rect 6280 39738 6332 39790
rect 6332 39738 6345 39790
rect 6345 39738 6397 39790
rect 6397 39738 6410 39790
rect 6410 39738 6462 39790
rect 6462 39738 6475 39790
rect 6475 39738 6527 39790
rect 6527 39738 6540 39790
rect 6540 39738 6592 39790
rect 6592 39738 6605 39790
rect 6605 39738 6657 39790
rect 6657 39738 6670 39790
rect 6670 39738 6722 39790
rect 6722 39738 6735 39790
rect 6735 39738 6787 39790
rect 6787 39738 6800 39790
rect 6800 39738 6852 39790
rect 6852 39738 6865 39790
rect 6865 39738 6917 39790
rect 6917 39738 6930 39790
rect 6930 39738 6982 39790
rect 6982 39738 6995 39790
rect 6995 39738 7047 39790
rect 7047 39738 7060 39790
rect 7060 39738 7112 39790
rect 7112 39738 7125 39790
rect 7125 39738 7177 39790
rect 7177 39738 7189 39790
rect 7189 39738 7241 39790
rect 7241 39738 7253 39790
rect 7253 39738 7305 39790
rect 7305 39738 7317 39790
rect 7317 39738 7369 39790
rect 7369 39738 7381 39790
rect 7381 39738 7433 39790
rect 7433 39738 7445 39790
rect 7445 39738 7497 39790
rect 7497 39738 7509 39790
rect 7509 39738 7561 39790
rect 7561 39738 7573 39790
rect 7573 39738 7625 39790
rect 7625 39738 7637 39790
rect 7637 39738 7689 39790
rect 7689 39738 7701 39790
rect 7701 39738 7753 39790
rect 7753 39738 7765 39790
rect 7765 39738 7817 39790
rect 7817 39738 7829 39790
rect 7829 39738 7881 39790
rect 7881 39738 7893 39790
rect 7893 39738 7945 39790
rect 7945 39738 7957 39790
rect 7957 39738 8009 39790
rect 8009 39738 8021 39790
rect 8021 39738 8073 39790
rect 8073 39738 8085 39790
rect 8085 39738 8137 39790
rect 8137 39738 8149 39790
rect 8149 39738 8201 39790
rect 8201 39738 8213 39790
rect 8213 39738 8265 39790
rect 8265 39738 8277 39790
rect 8277 39738 8329 39790
rect 8329 39738 8341 39790
rect 8341 39738 8393 39790
rect 8393 39738 8405 39790
rect 8405 39738 8457 39790
rect 8457 39738 8469 39790
rect 8469 39738 8521 39790
rect 8521 39738 8533 39790
rect 8533 39738 8585 39790
rect 8585 39738 8597 39790
rect 8597 39738 8649 39790
rect 8649 39738 8661 39790
rect 8661 39738 8713 39790
rect 8713 39738 8725 39790
rect 8725 39738 8777 39790
rect 8777 39738 8789 39790
rect 8789 39738 8841 39790
rect 8841 39738 8853 39790
rect 8853 39738 8905 39790
rect 8905 39738 8917 39790
rect 8917 39738 8969 39790
rect 8969 39738 8981 39790
rect 8981 39738 9033 39790
rect 9033 39738 9045 39790
rect 9045 39738 9097 39790
rect 9097 39738 9109 39790
rect 9109 39738 9161 39790
rect 9161 39738 9173 39790
rect 9173 39738 9225 39790
rect 9225 39738 9237 39790
rect 9237 39738 9289 39790
rect 9289 39738 9301 39790
rect 9301 39738 9353 39790
rect 9353 39738 9365 39790
rect 9365 39738 9417 39790
rect 9417 39738 9429 39790
rect 9429 39738 9481 39790
rect 9481 39738 9493 39790
rect 9493 39738 9545 39790
rect 9545 39738 9557 39790
rect 9557 39738 9609 39790
rect 9609 39738 9621 39790
rect 9621 39738 9673 39790
rect 9673 39738 9685 39790
rect 9685 39738 9737 39790
rect 9737 39738 9749 39790
rect 9749 39738 9801 39790
rect 9801 39738 9813 39790
rect 9813 39738 9865 39790
rect 9865 39738 9877 39790
rect 9877 39738 9929 39790
rect 9929 39738 9941 39790
rect 9941 39738 9993 39790
rect 9993 39738 10005 39790
rect 10005 39738 10057 39790
rect 10057 39738 10069 39790
rect 10069 39738 10121 39790
rect 10121 39738 10133 39790
rect 10133 39738 10185 39790
rect 10185 39738 10197 39790
rect 10197 39738 10249 39790
rect 10249 39738 10261 39790
rect 10261 39738 10313 39790
rect 10313 39738 10325 39790
rect 10325 39738 10377 39790
rect 10377 39738 10389 39790
rect 10389 39738 10441 39790
rect 10441 39738 10453 39790
rect 10453 39738 10505 39790
rect 10505 39738 10517 39790
rect 10517 39738 10569 39790
rect 10569 39738 10581 39790
rect 10581 39738 10633 39790
rect 10633 39738 10645 39790
rect 10645 39738 10697 39790
rect 10697 39738 10709 39790
rect 10709 39738 10761 39790
rect 10761 39738 10773 39790
rect 10773 39738 10825 39790
rect 10825 39738 10837 39790
rect 10837 39738 10889 39790
rect 10889 39738 10901 39790
rect 10901 39738 10953 39790
rect 10953 39738 10965 39790
rect 10965 39738 11017 39790
rect 11017 39738 11029 39790
rect 11029 39738 11081 39790
rect 11081 39738 11093 39790
rect 11093 39738 11145 39790
rect 11145 39738 11157 39790
rect 11157 39738 11209 39790
rect 11209 39738 11221 39790
rect 11221 39738 11273 39790
rect 11273 39738 11285 39790
rect 11285 39738 11334 39790
rect 14411 39946 14457 39995
rect 14457 39946 14467 39995
rect 14492 39946 14522 39995
rect 14522 39946 14535 39995
rect 14535 39946 14548 39995
rect 14573 39946 14587 39995
rect 14587 39946 14600 39995
rect 14600 39946 14629 39995
rect 14654 39946 14665 39995
rect 14665 39946 14710 39995
rect 14735 39946 14782 39995
rect 14782 39946 14791 39995
rect 14816 39946 14847 39995
rect 14847 39946 14860 39995
rect 14860 39946 14872 39995
rect 14897 39946 14912 39995
rect 14912 39946 14925 39995
rect 14925 39946 14953 39995
rect 14977 39946 14990 39995
rect 14990 39946 15033 39995
rect 15057 39946 15107 39995
rect 15107 39946 15113 39995
rect 15137 39946 15172 39995
rect 15172 39946 15185 39995
rect 15185 39946 15193 39995
rect 15217 39946 15237 39995
rect 15237 39946 15249 39995
rect 15249 39946 15273 39995
rect 15297 39946 15301 39995
rect 15301 39946 15313 39995
rect 15313 39946 15353 39995
rect 14411 39939 14467 39946
rect 14492 39939 14548 39946
rect 14573 39939 14629 39946
rect 14654 39939 14710 39946
rect 14735 39939 14791 39946
rect 14816 39939 14872 39946
rect 14897 39939 14953 39946
rect 14977 39939 15033 39946
rect 15057 39939 15113 39946
rect 15137 39939 15193 39946
rect 15217 39939 15273 39946
rect 15297 39939 15353 39946
rect 14411 39878 14457 39899
rect 14457 39878 14467 39899
rect 14492 39878 14522 39899
rect 14522 39878 14535 39899
rect 14535 39878 14548 39899
rect 14573 39878 14587 39899
rect 14587 39878 14600 39899
rect 14600 39878 14629 39899
rect 14654 39878 14665 39899
rect 14665 39878 14710 39899
rect 14735 39878 14782 39899
rect 14782 39878 14791 39899
rect 14816 39878 14847 39899
rect 14847 39878 14860 39899
rect 14860 39878 14872 39899
rect 14897 39878 14912 39899
rect 14912 39878 14925 39899
rect 14925 39878 14953 39899
rect 14977 39878 14990 39899
rect 14990 39878 15033 39899
rect 15057 39878 15107 39899
rect 15107 39878 15113 39899
rect 15137 39878 15172 39899
rect 15172 39878 15185 39899
rect 15185 39878 15193 39899
rect 15217 39878 15237 39899
rect 15237 39878 15249 39899
rect 15249 39878 15273 39899
rect 15297 39878 15301 39899
rect 15301 39878 15313 39899
rect 15313 39878 15353 39899
rect 14411 39862 14467 39878
rect 14492 39862 14548 39878
rect 14573 39862 14629 39878
rect 14654 39862 14710 39878
rect 14735 39862 14791 39878
rect 14816 39862 14872 39878
rect 14897 39862 14953 39878
rect 14977 39862 15033 39878
rect 15057 39862 15113 39878
rect 15137 39862 15193 39878
rect 15217 39862 15273 39878
rect 15297 39862 15353 39878
rect 14411 39843 14457 39862
rect 14457 39843 14467 39862
rect 14492 39843 14522 39862
rect 14522 39843 14535 39862
rect 14535 39843 14548 39862
rect 14573 39843 14587 39862
rect 14587 39843 14600 39862
rect 14600 39843 14629 39862
rect 14654 39843 14665 39862
rect 14665 39843 14710 39862
rect 14735 39843 14782 39862
rect 14782 39843 14791 39862
rect 14816 39843 14847 39862
rect 14847 39843 14860 39862
rect 14860 39843 14872 39862
rect 14897 39843 14912 39862
rect 14912 39843 14925 39862
rect 14925 39843 14953 39862
rect 14977 39843 14990 39862
rect 14990 39843 15033 39862
rect 15057 39843 15107 39862
rect 15107 39843 15113 39862
rect 15137 39843 15172 39862
rect 15172 39843 15185 39862
rect 15185 39843 15193 39862
rect 15217 39843 15237 39862
rect 15237 39843 15249 39862
rect 15249 39843 15273 39862
rect 15297 39843 15301 39862
rect 15301 39843 15313 39862
rect 15313 39843 15353 39862
rect 14411 39794 14467 39803
rect 14492 39794 14548 39803
rect 14573 39794 14629 39803
rect 14654 39794 14710 39803
rect 14735 39794 14791 39803
rect 14816 39794 14872 39803
rect 14897 39794 14953 39803
rect 14977 39794 15033 39803
rect 15057 39794 15113 39803
rect 15137 39794 15193 39803
rect 15217 39794 15273 39803
rect 15297 39794 15353 39803
rect 14411 39747 14457 39794
rect 14457 39747 14467 39794
rect 14492 39747 14522 39794
rect 14522 39747 14535 39794
rect 14535 39747 14548 39794
rect 14573 39747 14587 39794
rect 14587 39747 14600 39794
rect 14600 39747 14629 39794
rect 14654 39747 14665 39794
rect 14665 39747 14710 39794
rect 14735 39747 14782 39794
rect 14782 39747 14791 39794
rect 14816 39747 14847 39794
rect 14847 39747 14860 39794
rect 14860 39747 14872 39794
rect 14897 39747 14912 39794
rect 14912 39747 14925 39794
rect 14925 39747 14953 39794
rect 14977 39747 14990 39794
rect 14990 39747 15033 39794
rect 15057 39747 15107 39794
rect 15107 39747 15113 39794
rect 15137 39747 15172 39794
rect 15172 39747 15185 39794
rect 15185 39747 15193 39794
rect 15217 39747 15237 39794
rect 15237 39747 15249 39794
rect 15249 39747 15273 39794
rect 15297 39747 15301 39794
rect 15301 39747 15313 39794
rect 15313 39747 15353 39794
rect 1361 39566 1417 39622
rect 1443 39566 1499 39622
rect 1525 39566 1581 39622
rect 1607 39566 1663 39622
rect 1689 39566 1745 39622
rect 1903 39619 1959 39675
rect 1984 39619 2040 39675
rect 2065 39619 2121 39675
rect 2146 39619 2202 39675
rect 2227 39619 2283 39675
rect 2308 39619 2364 39675
rect 2389 39619 2445 39675
rect 2470 39619 2526 39675
rect 2551 39619 2607 39675
rect 2632 39619 2688 39675
rect 2713 39619 2769 39675
rect 2794 39619 2850 39675
rect 2875 39619 2931 39675
rect 2956 39619 3012 39675
rect 3037 39619 3093 39675
rect 1361 39484 1417 39540
rect 1443 39484 1499 39540
rect 1525 39484 1581 39540
rect 1607 39484 1663 39540
rect 1689 39484 1745 39540
rect 1903 39539 1959 39595
rect 1984 39539 2040 39595
rect 2065 39539 2121 39595
rect 2146 39539 2202 39595
rect 2227 39539 2283 39595
rect 2308 39539 2364 39595
rect 2389 39539 2445 39595
rect 2470 39539 2526 39595
rect 2551 39539 2607 39595
rect 2632 39539 2688 39595
rect 2713 39539 2769 39595
rect 2794 39539 2850 39595
rect 2875 39539 2931 39595
rect 2956 39539 3012 39595
rect 3037 39539 3093 39595
rect 3118 39539 11334 39738
rect 1361 39402 1417 39458
rect 1443 39402 1499 39458
rect 1525 39402 1581 39458
rect 1607 39402 1663 39458
rect 1689 39402 1745 39458
rect 1361 39320 1417 39376
rect 1443 39320 1499 39376
rect 1525 39320 1581 39376
rect 1607 39320 1663 39376
rect 1689 39320 1745 39376
rect 1361 39238 1417 39294
rect 1443 39238 1499 39294
rect 1525 39238 1581 39294
rect 1607 39238 1663 39294
rect 1689 39238 1745 39294
rect 1361 39156 1417 39212
rect 1443 39156 1499 39212
rect 1525 39156 1581 39212
rect 1607 39156 1663 39212
rect 1689 39156 1745 39212
rect 1361 39074 1417 39130
rect 1443 39074 1499 39130
rect 1525 39074 1581 39130
rect 1607 39074 1663 39130
rect 1689 39074 1745 39130
rect 1361 38992 1417 39048
rect 1443 38992 1499 39048
rect 1525 38992 1581 39048
rect 1607 38992 1663 39048
rect 1689 38992 1745 39048
rect 1361 38910 1417 38966
rect 1443 38910 1499 38966
rect 1525 38910 1581 38966
rect 1607 38910 1663 38966
rect 1689 38910 1745 38966
rect 1361 38828 1417 38884
rect 1443 38828 1499 38884
rect 1525 38828 1581 38884
rect 1607 38828 1663 38884
rect 1689 38828 1745 38884
rect 1361 38746 1417 38802
rect 1443 38746 1499 38802
rect 1525 38746 1581 38802
rect 1607 38746 1663 38802
rect 1689 38746 1745 38802
rect 1361 38664 1417 38720
rect 1443 38664 1499 38720
rect 1525 38664 1581 38720
rect 1607 38664 1663 38720
rect 1689 38664 1745 38720
rect 1361 38582 1417 38638
rect 1443 38582 1499 38638
rect 1525 38582 1581 38638
rect 1607 38582 1663 38638
rect 1689 38582 1745 38638
rect 1361 38500 1417 38556
rect 1443 38500 1499 38556
rect 1525 38500 1581 38556
rect 1607 38500 1663 38556
rect 1689 38500 1745 38556
rect 1361 38418 1417 38474
rect 1443 38418 1499 38474
rect 1525 38418 1581 38474
rect 1607 38418 1663 38474
rect 1689 38418 1745 38474
rect 1361 38336 1417 38392
rect 1443 38336 1499 38392
rect 1525 38336 1581 38392
rect 1607 38336 1663 38392
rect 1689 38336 1745 38392
rect 1361 38254 1417 38310
rect 1443 38254 1499 38310
rect 1525 38254 1581 38310
rect 1607 38254 1663 38310
rect 1689 38254 1745 38310
rect 1361 38172 1417 38228
rect 1443 38172 1499 38228
rect 1525 38172 1581 38228
rect 1607 38172 1663 38228
rect 1689 38172 1745 38228
rect 1361 38090 1417 38146
rect 1443 38090 1499 38146
rect 1525 38090 1581 38146
rect 1607 38090 1663 38146
rect 1689 38090 1745 38146
rect 1361 38008 1417 38064
rect 1443 38008 1499 38064
rect 1525 38008 1581 38064
rect 1607 38008 1663 38064
rect 1689 38008 1745 38064
rect 1361 37925 1417 37981
rect 1443 37925 1499 37981
rect 1525 37925 1581 37981
rect 1607 37925 1663 37981
rect 1689 37925 1745 37981
rect 1361 37842 1417 37898
rect 1443 37842 1499 37898
rect 1525 37842 1581 37898
rect 1607 37842 1663 37898
rect 1689 37842 1745 37898
rect 1361 37759 1417 37815
rect 1443 37759 1499 37815
rect 1525 37759 1581 37815
rect 1607 37759 1663 37815
rect 1689 37759 1745 37815
rect 1361 37676 1417 37732
rect 1443 37676 1499 37732
rect 1525 37676 1581 37732
rect 1607 37676 1663 37732
rect 1689 37676 1745 37732
rect 1361 37593 1417 37649
rect 1443 37593 1499 37649
rect 1525 37593 1581 37649
rect 1607 37593 1663 37649
rect 1689 37593 1745 37649
rect 1361 37510 1417 37566
rect 1443 37510 1499 37566
rect 1525 37510 1581 37566
rect 1607 37510 1663 37566
rect 1689 37510 1745 37566
rect 1361 37427 1417 37483
rect 1443 37427 1499 37483
rect 1525 37427 1581 37483
rect 1607 37427 1663 37483
rect 1689 37427 1745 37483
rect 1361 37344 1417 37400
rect 1443 37344 1499 37400
rect 1525 37344 1581 37400
rect 1607 37344 1663 37400
rect 1689 37344 1745 37400
rect 1361 37261 1417 37317
rect 1443 37261 1499 37317
rect 1525 37261 1581 37317
rect 1607 37261 1663 37317
rect 1689 37261 1745 37317
rect 1361 37178 1417 37234
rect 1443 37178 1499 37234
rect 1525 37178 1581 37234
rect 1607 37178 1663 37234
rect 1689 37178 1745 37234
rect 4089 36310 4145 36366
rect 4231 36310 4287 36366
rect 4372 36310 4428 36366
rect 4513 36310 4569 36366
rect 4654 36310 4710 36366
rect 837 36173 893 36229
rect 4089 36210 4145 36266
rect 4231 36210 4287 36266
rect 4372 36210 4428 36266
rect 4513 36210 4569 36266
rect 4654 36210 4710 36266
rect 837 36093 893 36149
rect 2792 36079 2848 36081
rect 2924 36079 2980 36081
rect 3056 36079 3112 36081
rect 3187 36079 3243 36081
rect 3318 36079 3374 36081
rect 3449 36079 3505 36081
rect 3580 36079 3636 36081
rect 3711 36079 3767 36081
rect 2792 36027 2844 36079
rect 2844 36027 2848 36079
rect 2924 36027 2976 36079
rect 2976 36027 2980 36079
rect 3056 36027 3108 36079
rect 3108 36027 3112 36079
rect 3187 36027 3188 36079
rect 3188 36027 3240 36079
rect 3240 36027 3243 36079
rect 3318 36027 3320 36079
rect 3320 36027 3372 36079
rect 3372 36027 3374 36079
rect 3449 36027 3452 36079
rect 3452 36027 3504 36079
rect 3504 36027 3505 36079
rect 3580 36027 3584 36079
rect 3584 36027 3636 36079
rect 3711 36027 3715 36079
rect 3715 36027 3767 36079
rect 2792 36025 2848 36027
rect 2924 36025 2980 36027
rect 3056 36025 3112 36027
rect 3187 36025 3243 36027
rect 3318 36025 3374 36027
rect 3449 36025 3505 36027
rect 3580 36025 3636 36027
rect 3711 36025 3767 36027
rect 2792 35949 2844 35963
rect 2844 35949 2848 35963
rect 2924 35949 2976 35963
rect 2976 35949 2980 35963
rect 3056 35949 3108 35963
rect 3108 35949 3112 35963
rect 3187 35949 3188 35963
rect 3188 35949 3240 35963
rect 3240 35949 3243 35963
rect 3318 35949 3320 35963
rect 3320 35949 3372 35963
rect 3372 35949 3374 35963
rect 3449 35949 3452 35963
rect 3452 35949 3504 35963
rect 3504 35949 3505 35963
rect 3580 35949 3584 35963
rect 3584 35949 3636 35963
rect 3711 35949 3715 35963
rect 3715 35949 3767 35963
rect 2792 35923 2848 35949
rect 2924 35923 2980 35949
rect 3056 35923 3112 35949
rect 3187 35923 3243 35949
rect 3318 35923 3374 35949
rect 3449 35923 3505 35949
rect 3580 35923 3636 35949
rect 3711 35923 3767 35949
rect 2792 35907 2844 35923
rect 2844 35907 2848 35923
rect 2924 35907 2976 35923
rect 2976 35907 2980 35923
rect 3056 35907 3108 35923
rect 3108 35907 3112 35923
rect 3187 35907 3188 35923
rect 3188 35907 3240 35923
rect 3240 35907 3243 35923
rect 3318 35907 3320 35923
rect 3320 35907 3372 35923
rect 3372 35907 3374 35923
rect 3449 35907 3452 35923
rect 3452 35907 3504 35923
rect 3504 35907 3505 35923
rect 3580 35907 3584 35923
rect 3584 35907 3636 35923
rect 3711 35907 3715 35923
rect 3715 35907 3767 35923
rect 2792 35793 2844 35845
rect 2844 35793 2848 35845
rect 2924 35793 2976 35845
rect 2976 35793 2980 35845
rect 3056 35793 3108 35845
rect 3108 35793 3112 35845
rect 3187 35793 3188 35845
rect 3188 35793 3240 35845
rect 3240 35793 3243 35845
rect 3318 35793 3320 35845
rect 3320 35793 3372 35845
rect 3372 35793 3374 35845
rect 3449 35793 3452 35845
rect 3452 35793 3504 35845
rect 3504 35793 3505 35845
rect 3580 35793 3584 35845
rect 3584 35793 3636 35845
rect 3711 35793 3715 35845
rect 3715 35793 3767 35845
rect 2792 35789 2848 35793
rect 2924 35789 2980 35793
rect 3056 35789 3112 35793
rect 3187 35789 3243 35793
rect 3318 35789 3374 35793
rect 3449 35789 3505 35793
rect 3580 35789 3636 35793
rect 3711 35789 3767 35793
rect 298 35562 354 35618
rect 396 35562 452 35618
rect 494 35610 550 35618
rect 592 35610 648 35618
rect 494 35562 506 35610
rect 506 35562 528 35610
rect 528 35562 550 35610
rect 592 35562 602 35610
rect 602 35562 648 35610
rect 298 35482 354 35538
rect 396 35482 452 35538
rect 494 35494 506 35538
rect 506 35494 528 35538
rect 528 35494 550 35538
rect 592 35494 602 35538
rect 602 35494 648 35538
rect 494 35482 550 35494
rect 592 35482 648 35494
rect 298 35402 354 35458
rect 396 35402 452 35458
rect 494 35430 506 35458
rect 506 35430 528 35458
rect 528 35430 550 35458
rect 592 35430 602 35458
rect 602 35430 648 35458
rect 494 35418 550 35430
rect 592 35418 648 35430
rect 494 35402 506 35418
rect 506 35402 528 35418
rect 528 35402 550 35418
rect 592 35402 602 35418
rect 602 35402 648 35418
rect 298 35322 354 35378
rect 396 35322 452 35378
rect 494 35366 506 35378
rect 506 35366 528 35378
rect 528 35366 550 35378
rect 592 35366 602 35378
rect 602 35366 648 35378
rect 494 35354 550 35366
rect 592 35354 648 35366
rect 494 35322 506 35354
rect 506 35322 528 35354
rect 528 35322 550 35354
rect 592 35322 602 35354
rect 602 35322 648 35354
rect 298 35242 354 35298
rect 396 35242 452 35298
rect 494 35290 550 35298
rect 592 35290 648 35298
rect 494 35242 506 35290
rect 506 35242 528 35290
rect 528 35242 550 35290
rect 592 35242 602 35290
rect 602 35242 648 35290
rect 298 35162 354 35218
rect 396 35162 452 35218
rect 494 35174 506 35218
rect 506 35174 528 35218
rect 528 35174 550 35218
rect 592 35174 602 35218
rect 602 35174 648 35218
rect 494 35162 550 35174
rect 592 35162 648 35174
rect 298 35082 354 35138
rect 396 35082 452 35138
rect 494 35110 506 35138
rect 506 35110 528 35138
rect 528 35110 550 35138
rect 592 35110 602 35138
rect 602 35110 648 35138
rect 494 35098 550 35110
rect 592 35098 648 35110
rect 494 35082 506 35098
rect 506 35082 528 35098
rect 528 35082 550 35098
rect 592 35082 602 35098
rect 602 35082 648 35098
rect 298 35002 354 35058
rect 396 35002 452 35058
rect 494 35046 506 35058
rect 506 35046 528 35058
rect 528 35046 550 35058
rect 592 35046 602 35058
rect 602 35046 648 35058
rect 494 35034 550 35046
rect 592 35034 648 35046
rect 494 35002 506 35034
rect 506 35002 528 35034
rect 528 35002 550 35034
rect 592 35002 602 35034
rect 602 35002 648 35034
rect 298 34922 354 34978
rect 396 34922 452 34978
rect 494 34970 550 34978
rect 592 34970 648 34978
rect 494 34922 506 34970
rect 506 34922 528 34970
rect 528 34922 550 34970
rect 592 34922 602 34970
rect 602 34922 648 34970
rect 298 34842 354 34898
rect 396 34842 452 34898
rect 494 34854 506 34898
rect 506 34854 528 34898
rect 528 34854 550 34898
rect 592 34854 602 34898
rect 602 34854 648 34898
rect 494 34842 550 34854
rect 592 34842 648 34854
rect 298 34762 354 34818
rect 396 34762 452 34818
rect 494 34790 506 34818
rect 506 34790 528 34818
rect 528 34790 550 34818
rect 592 34790 602 34818
rect 602 34790 648 34818
rect 494 34778 550 34790
rect 592 34778 648 34790
rect 494 34762 506 34778
rect 506 34762 528 34778
rect 528 34762 550 34778
rect 592 34762 602 34778
rect 602 34762 648 34778
rect 298 34682 354 34738
rect 396 34682 452 34738
rect 494 34726 506 34738
rect 506 34726 528 34738
rect 528 34726 550 34738
rect 592 34726 602 34738
rect 602 34726 648 34738
rect 494 34714 550 34726
rect 592 34714 648 34726
rect 494 34682 506 34714
rect 506 34682 528 34714
rect 528 34682 550 34714
rect 592 34682 602 34714
rect 602 34682 648 34714
rect 298 34602 354 34658
rect 396 34602 452 34658
rect 494 34650 550 34658
rect 592 34650 648 34658
rect 494 34602 506 34650
rect 506 34602 528 34650
rect 528 34602 550 34650
rect 592 34602 602 34650
rect 602 34602 648 34650
rect 298 34522 354 34578
rect 396 34522 452 34578
rect 494 34534 506 34578
rect 506 34534 528 34578
rect 528 34534 550 34578
rect 592 34534 602 34578
rect 602 34534 648 34578
rect 494 34522 550 34534
rect 592 34522 648 34534
rect 298 34442 354 34498
rect 396 34442 452 34498
rect 494 34470 506 34498
rect 506 34470 528 34498
rect 528 34470 550 34498
rect 592 34470 602 34498
rect 602 34470 648 34498
rect 494 34458 550 34470
rect 592 34458 648 34470
rect 494 34442 506 34458
rect 506 34442 528 34458
rect 528 34442 550 34458
rect 592 34442 602 34458
rect 602 34442 648 34458
rect 298 34362 354 34418
rect 396 34362 452 34418
rect 494 34406 506 34418
rect 506 34406 528 34418
rect 528 34406 550 34418
rect 592 34406 602 34418
rect 602 34406 648 34418
rect 494 34394 550 34406
rect 592 34394 648 34406
rect 494 34362 506 34394
rect 506 34362 528 34394
rect 528 34362 550 34394
rect 592 34362 602 34394
rect 602 34362 648 34394
rect 298 34282 354 34338
rect 396 34282 452 34338
rect 494 34330 550 34338
rect 592 34330 648 34338
rect 494 34282 506 34330
rect 506 34282 528 34330
rect 528 34282 550 34330
rect 592 34282 602 34330
rect 602 34282 648 34330
rect 298 34202 354 34258
rect 396 34202 452 34258
rect 494 34214 506 34258
rect 506 34214 528 34258
rect 528 34214 550 34258
rect 592 34214 602 34258
rect 602 34214 648 34258
rect 494 34202 550 34214
rect 592 34202 648 34214
rect 298 34122 354 34178
rect 396 34122 452 34178
rect 494 34150 506 34178
rect 506 34150 528 34178
rect 528 34150 550 34178
rect 592 34150 602 34178
rect 602 34150 648 34178
rect 494 34138 550 34150
rect 592 34138 648 34150
rect 494 34122 506 34138
rect 506 34122 528 34138
rect 528 34122 550 34138
rect 592 34122 602 34138
rect 602 34122 648 34138
rect 298 34042 354 34098
rect 396 34042 452 34098
rect 494 34086 506 34098
rect 506 34086 528 34098
rect 528 34086 550 34098
rect 592 34086 602 34098
rect 602 34086 648 34098
rect 494 34074 550 34086
rect 592 34074 648 34086
rect 494 34042 506 34074
rect 506 34042 528 34074
rect 528 34042 550 34074
rect 592 34042 602 34074
rect 602 34042 648 34074
rect 298 34012 354 34018
rect 298 33962 299 34012
rect 299 33962 354 34012
rect 396 33962 452 34018
rect 494 34010 550 34018
rect 592 34010 648 34018
rect 494 33962 506 34010
rect 506 33962 528 34010
rect 528 33962 550 34010
rect 592 33962 602 34010
rect 602 33962 648 34010
rect 298 33896 299 33938
rect 299 33896 354 33938
rect 298 33884 354 33896
rect 298 33882 299 33884
rect 299 33882 354 33884
rect 396 33882 452 33938
rect 494 33894 506 33938
rect 506 33894 528 33938
rect 528 33894 550 33938
rect 592 33894 602 33938
rect 602 33894 648 33938
rect 494 33882 550 33894
rect 592 33882 648 33894
rect 298 33832 299 33858
rect 299 33832 354 33858
rect 298 33820 354 33832
rect 298 33802 299 33820
rect 299 33802 354 33820
rect 396 33802 452 33858
rect 494 33830 506 33858
rect 506 33830 528 33858
rect 528 33830 550 33858
rect 592 33830 602 33858
rect 602 33830 648 33858
rect 494 33818 550 33830
rect 592 33818 648 33830
rect 494 33802 506 33818
rect 506 33802 528 33818
rect 528 33802 550 33818
rect 592 33802 602 33818
rect 602 33802 648 33818
rect 298 33768 299 33778
rect 299 33768 354 33778
rect 298 33756 354 33768
rect 298 33722 299 33756
rect 299 33722 354 33756
rect 396 33722 452 33778
rect 494 33766 506 33778
rect 506 33766 528 33778
rect 528 33766 550 33778
rect 592 33766 602 33778
rect 602 33766 648 33778
rect 494 33754 550 33766
rect 592 33754 648 33766
rect 494 33722 506 33754
rect 506 33722 528 33754
rect 528 33722 550 33754
rect 592 33722 602 33754
rect 602 33722 648 33754
rect 298 33692 354 33698
rect 298 33642 299 33692
rect 299 33642 354 33692
rect 396 33642 452 33698
rect 494 33690 550 33698
rect 592 33690 648 33698
rect 494 33642 506 33690
rect 506 33642 528 33690
rect 528 33642 550 33690
rect 592 33642 602 33690
rect 602 33642 648 33690
rect 298 33576 299 33618
rect 299 33576 354 33618
rect 298 33564 354 33576
rect 298 33562 299 33564
rect 299 33562 354 33564
rect 396 33562 452 33618
rect 494 33574 506 33618
rect 506 33574 528 33618
rect 528 33574 550 33618
rect 592 33574 602 33618
rect 602 33574 648 33618
rect 494 33562 550 33574
rect 592 33562 648 33574
rect 298 33512 299 33538
rect 299 33512 354 33538
rect 298 33500 354 33512
rect 298 33482 299 33500
rect 299 33482 354 33500
rect 396 33482 452 33538
rect 494 33510 506 33538
rect 506 33510 528 33538
rect 528 33510 550 33538
rect 592 33510 602 33538
rect 602 33510 648 33538
rect 494 33498 550 33510
rect 592 33498 648 33510
rect 494 33482 506 33498
rect 506 33482 528 33498
rect 528 33482 550 33498
rect 592 33482 602 33498
rect 602 33482 648 33498
rect 298 33448 299 33458
rect 299 33448 354 33458
rect 298 33436 354 33448
rect 298 33402 299 33436
rect 299 33402 354 33436
rect 396 33402 452 33458
rect 494 33446 506 33458
rect 506 33446 528 33458
rect 528 33446 550 33458
rect 592 33446 602 33458
rect 602 33446 648 33458
rect 494 33434 550 33446
rect 592 33434 648 33446
rect 494 33402 506 33434
rect 506 33402 528 33434
rect 528 33402 550 33434
rect 592 33402 602 33434
rect 602 33402 648 33434
rect 298 33372 354 33378
rect 298 33322 299 33372
rect 299 33322 354 33372
rect 396 33322 452 33378
rect 494 33370 550 33378
rect 592 33370 648 33378
rect 494 33322 506 33370
rect 506 33322 528 33370
rect 528 33322 550 33370
rect 592 33322 602 33370
rect 602 33322 648 33370
rect 298 33256 299 33298
rect 299 33256 354 33298
rect 298 33244 354 33256
rect 298 33242 299 33244
rect 299 33242 354 33244
rect 396 33242 452 33298
rect 494 33254 506 33298
rect 506 33254 528 33298
rect 528 33254 550 33298
rect 592 33254 602 33298
rect 602 33254 648 33298
rect 494 33242 550 33254
rect 592 33242 648 33254
rect 298 33192 299 33218
rect 299 33192 354 33218
rect 298 33180 354 33192
rect 298 33162 299 33180
rect 299 33162 354 33180
rect 396 33162 452 33218
rect 494 33190 506 33218
rect 506 33190 528 33218
rect 528 33190 550 33218
rect 592 33190 602 33218
rect 602 33190 648 33218
rect 494 33178 550 33190
rect 592 33178 648 33190
rect 494 33162 506 33178
rect 506 33162 528 33178
rect 528 33162 550 33178
rect 592 33162 602 33178
rect 602 33162 648 33178
rect 298 33128 299 33138
rect 299 33128 354 33138
rect 298 33116 354 33128
rect 298 33082 299 33116
rect 299 33082 354 33116
rect 396 33082 452 33138
rect 494 33126 506 33138
rect 506 33126 528 33138
rect 528 33126 550 33138
rect 592 33126 602 33138
rect 602 33126 648 33138
rect 494 33114 550 33126
rect 592 33114 648 33126
rect 494 33082 506 33114
rect 506 33082 528 33114
rect 528 33082 550 33114
rect 592 33082 602 33114
rect 602 33082 648 33114
rect 298 33052 354 33058
rect 298 33002 299 33052
rect 299 33002 354 33052
rect 396 33002 452 33058
rect 494 33050 550 33058
rect 592 33050 648 33058
rect 494 33002 506 33050
rect 506 33002 528 33050
rect 528 33002 550 33050
rect 592 33002 602 33050
rect 602 33002 648 33050
rect 298 32936 299 32978
rect 299 32936 354 32978
rect 298 32924 354 32936
rect 298 32922 299 32924
rect 299 32922 354 32924
rect 396 32922 452 32978
rect 494 32934 506 32978
rect 506 32934 528 32978
rect 528 32934 550 32978
rect 592 32934 602 32978
rect 602 32934 648 32978
rect 494 32922 550 32934
rect 592 32922 648 32934
rect 298 32872 299 32898
rect 299 32872 354 32898
rect 298 32859 354 32872
rect 298 32842 299 32859
rect 299 32842 354 32859
rect 396 32842 452 32898
rect 494 32870 506 32898
rect 506 32870 528 32898
rect 528 32870 550 32898
rect 592 32870 602 32898
rect 602 32870 648 32898
rect 494 32858 550 32870
rect 592 32858 648 32870
rect 494 32842 506 32858
rect 506 32842 528 32858
rect 528 32842 550 32858
rect 592 32842 602 32858
rect 602 32842 648 32858
rect 298 32807 299 32818
rect 299 32807 354 32818
rect 298 32794 354 32807
rect 298 32762 299 32794
rect 299 32762 354 32794
rect 396 32762 452 32818
rect 494 32806 506 32818
rect 506 32806 528 32818
rect 528 32806 550 32818
rect 592 32806 602 32818
rect 602 32806 648 32818
rect 494 32794 550 32806
rect 592 32794 648 32806
rect 494 32762 506 32794
rect 506 32762 528 32794
rect 528 32762 550 32794
rect 592 32762 602 32794
rect 602 32762 648 32794
rect 298 32729 354 32738
rect 298 32682 299 32729
rect 299 32682 354 32729
rect 396 32682 452 32738
rect 494 32729 550 32738
rect 592 32729 648 32738
rect 494 32682 506 32729
rect 506 32682 528 32729
rect 528 32682 550 32729
rect 592 32682 602 32729
rect 602 32682 648 32729
rect 298 32612 299 32658
rect 299 32612 354 32658
rect 298 32602 354 32612
rect 396 32602 452 32658
rect 494 32612 506 32658
rect 506 32612 528 32658
rect 528 32612 550 32658
rect 592 32612 602 32658
rect 602 32612 648 32658
rect 494 32602 550 32612
rect 592 32602 648 32612
rect 298 32547 299 32578
rect 299 32547 354 32578
rect 298 32534 354 32547
rect 298 32522 299 32534
rect 299 32522 354 32534
rect 396 32522 452 32578
rect 494 32547 506 32578
rect 506 32547 528 32578
rect 528 32547 550 32578
rect 592 32547 602 32578
rect 602 32547 648 32578
rect 494 32534 550 32547
rect 592 32534 648 32547
rect 494 32522 506 32534
rect 506 32522 528 32534
rect 528 32522 550 32534
rect 592 32522 602 32534
rect 602 32522 648 32534
rect 298 32482 299 32498
rect 299 32482 354 32498
rect 298 32469 354 32482
rect 298 32442 299 32469
rect 299 32442 354 32469
rect 396 32442 452 32498
rect 494 32482 506 32498
rect 506 32482 528 32498
rect 528 32482 550 32498
rect 592 32482 602 32498
rect 602 32482 648 32498
rect 494 32469 550 32482
rect 592 32469 648 32482
rect 494 32442 506 32469
rect 506 32442 528 32469
rect 528 32442 550 32469
rect 592 32442 602 32469
rect 602 32442 648 32469
rect 298 32417 299 32418
rect 299 32417 354 32418
rect 298 32404 354 32417
rect 298 32362 299 32404
rect 299 32362 354 32404
rect 396 32362 452 32418
rect 494 32417 506 32418
rect 506 32417 528 32418
rect 528 32417 550 32418
rect 592 32417 602 32418
rect 602 32417 648 32418
rect 494 32404 550 32417
rect 592 32404 648 32417
rect 494 32362 506 32404
rect 506 32362 528 32404
rect 528 32362 550 32404
rect 592 32362 602 32404
rect 602 32362 648 32404
rect 298 32287 299 32338
rect 299 32287 354 32338
rect 298 32282 354 32287
rect 396 32282 452 32338
rect 494 32287 506 32338
rect 506 32287 528 32338
rect 528 32287 550 32338
rect 592 32287 602 32338
rect 602 32287 648 32338
rect 494 32282 550 32287
rect 592 32282 648 32287
rect 298 32222 299 32258
rect 299 32222 354 32258
rect 298 32209 354 32222
rect 298 32202 299 32209
rect 299 32202 354 32209
rect 396 32202 452 32258
rect 494 32222 506 32258
rect 506 32222 528 32258
rect 528 32222 550 32258
rect 592 32222 602 32258
rect 602 32222 648 32258
rect 494 32209 550 32222
rect 592 32209 648 32222
rect 494 32202 506 32209
rect 506 32202 528 32209
rect 528 32202 550 32209
rect 592 32202 602 32209
rect 602 32202 648 32209
rect 298 32157 299 32177
rect 299 32157 354 32177
rect 298 32144 354 32157
rect 298 32121 299 32144
rect 299 32121 354 32144
rect 396 32121 452 32177
rect 494 32157 506 32177
rect 506 32157 528 32177
rect 528 32157 550 32177
rect 592 32157 602 32177
rect 602 32157 648 32177
rect 494 32144 550 32157
rect 592 32144 648 32157
rect 494 32121 506 32144
rect 506 32121 528 32144
rect 528 32121 550 32144
rect 592 32121 602 32144
rect 602 32121 648 32144
rect 298 32092 299 32096
rect 299 32092 354 32096
rect 298 32079 354 32092
rect 298 32040 299 32079
rect 299 32040 354 32079
rect 396 32040 452 32096
rect 494 32092 506 32096
rect 506 32092 528 32096
rect 528 32092 550 32096
rect 592 32092 602 32096
rect 602 32092 648 32096
rect 494 32079 550 32092
rect 592 32079 648 32092
rect 494 32040 506 32079
rect 506 32040 528 32079
rect 528 32040 550 32079
rect 592 32040 602 32079
rect 602 32040 648 32079
rect 298 32014 354 32015
rect 298 31962 299 32014
rect 299 31962 354 32014
rect 298 31959 354 31962
rect 396 31959 452 32015
rect 494 32014 550 32015
rect 592 32014 648 32015
rect 494 31962 506 32014
rect 506 31962 528 32014
rect 528 31962 550 32014
rect 592 31962 602 32014
rect 602 31962 648 32014
rect 494 31959 550 31962
rect 592 31959 648 31962
rect 298 31897 299 31934
rect 299 31897 354 31934
rect 298 31884 354 31897
rect 298 31878 299 31884
rect 299 31878 354 31884
rect 396 31878 452 31934
rect 494 31897 506 31934
rect 506 31897 528 31934
rect 528 31897 550 31934
rect 592 31897 602 31934
rect 602 31897 648 31934
rect 494 31884 550 31897
rect 592 31884 648 31897
rect 494 31878 506 31884
rect 506 31878 528 31884
rect 528 31878 550 31884
rect 592 31878 602 31884
rect 602 31878 648 31884
rect 298 31832 299 31853
rect 299 31832 354 31853
rect 298 31819 354 31832
rect 298 31797 299 31819
rect 299 31797 354 31819
rect 396 31797 452 31853
rect 494 31832 506 31853
rect 506 31832 528 31853
rect 528 31832 550 31853
rect 592 31832 602 31853
rect 602 31832 648 31853
rect 494 31819 550 31832
rect 592 31819 648 31832
rect 494 31797 506 31819
rect 506 31797 528 31819
rect 528 31797 550 31819
rect 592 31797 602 31819
rect 602 31797 648 31819
rect 298 31767 299 31772
rect 299 31767 354 31772
rect 298 31754 354 31767
rect 298 31716 299 31754
rect 299 31716 354 31754
rect 396 31716 452 31772
rect 494 31767 506 31772
rect 506 31767 528 31772
rect 528 31767 550 31772
rect 592 31767 602 31772
rect 602 31767 648 31772
rect 494 31754 550 31767
rect 592 31754 648 31767
rect 494 31716 506 31754
rect 506 31716 528 31754
rect 528 31716 550 31754
rect 592 31716 602 31754
rect 602 31716 648 31754
rect 298 31689 354 31691
rect 298 31637 299 31689
rect 299 31637 354 31689
rect 298 31635 354 31637
rect 396 31635 452 31691
rect 494 31689 550 31691
rect 592 31689 648 31691
rect 494 31637 506 31689
rect 506 31637 528 31689
rect 528 31637 550 31689
rect 592 31637 602 31689
rect 602 31637 648 31689
rect 494 31635 550 31637
rect 592 31635 648 31637
rect 298 31572 299 31610
rect 299 31572 354 31610
rect 298 31559 354 31572
rect 298 31554 299 31559
rect 299 31554 354 31559
rect 396 31554 452 31610
rect 494 31572 506 31610
rect 506 31572 528 31610
rect 528 31572 550 31610
rect 592 31572 602 31610
rect 602 31572 648 31610
rect 494 31559 550 31572
rect 592 31559 648 31572
rect 494 31554 506 31559
rect 506 31554 528 31559
rect 528 31554 550 31559
rect 592 31554 602 31559
rect 602 31554 648 31559
rect 298 31507 299 31529
rect 299 31507 354 31529
rect 298 31494 354 31507
rect 298 31473 299 31494
rect 299 31473 354 31494
rect 396 31473 452 31529
rect 494 31507 506 31529
rect 506 31507 528 31529
rect 528 31507 550 31529
rect 592 31507 602 31529
rect 602 31507 648 31529
rect 494 31494 550 31507
rect 592 31494 648 31507
rect 494 31473 506 31494
rect 506 31473 528 31494
rect 528 31473 550 31494
rect 592 31473 602 31494
rect 602 31473 648 31494
rect 5112 32557 5168 32613
rect 5193 32557 5249 32613
rect 5273 32557 5329 32613
rect 5353 32557 5409 32613
rect 5433 32557 5489 32613
rect 5513 32557 5569 32613
rect 5593 32557 5649 32613
rect 5673 32557 5729 32613
rect 5753 32557 5809 32613
rect 5833 32557 5889 32613
rect 5913 32557 5969 32613
rect 5993 32557 6049 32613
rect 6073 32557 6129 32613
rect 6153 32557 6209 32613
rect 6233 32557 6289 32613
rect 5112 32475 5168 32531
rect 5193 32475 5249 32531
rect 5273 32475 5329 32531
rect 5353 32475 5409 32531
rect 5433 32475 5489 32531
rect 5513 32475 5569 32531
rect 5593 32475 5649 32531
rect 5673 32475 5729 32531
rect 5753 32475 5809 32531
rect 5833 32475 5889 32531
rect 5913 32475 5969 32531
rect 5993 32475 6049 32531
rect 6073 32475 6129 32531
rect 6153 32475 6209 32531
rect 6233 32475 6289 32531
rect 5112 32393 5168 32449
rect 5193 32393 5249 32449
rect 5273 32393 5329 32449
rect 5353 32393 5409 32449
rect 5433 32393 5489 32449
rect 5513 32393 5569 32449
rect 5593 32393 5649 32449
rect 5673 32393 5729 32449
rect 5753 32393 5809 32449
rect 5833 32393 5889 32449
rect 5913 32393 5969 32449
rect 5993 32393 6049 32449
rect 6073 32393 6129 32449
rect 6153 32393 6209 32449
rect 6233 32393 6289 32449
rect 5112 32311 5168 32367
rect 5193 32311 5249 32367
rect 5273 32311 5329 32367
rect 5353 32311 5409 32367
rect 5433 32311 5489 32367
rect 5513 32311 5569 32367
rect 5593 32311 5649 32367
rect 5673 32311 5729 32367
rect 5753 32311 5809 32367
rect 5833 32311 5889 32367
rect 5913 32311 5969 32367
rect 5993 32311 6049 32367
rect 6073 32311 6129 32367
rect 6153 32311 6209 32367
rect 6233 32311 6289 32367
rect 5112 32229 5168 32285
rect 5193 32229 5249 32285
rect 5273 32229 5329 32285
rect 5353 32229 5409 32285
rect 5433 32229 5489 32285
rect 5513 32229 5569 32285
rect 5593 32229 5649 32285
rect 5673 32229 5729 32285
rect 5753 32229 5809 32285
rect 5833 32229 5889 32285
rect 5913 32229 5969 32285
rect 5993 32229 6049 32285
rect 6073 32229 6129 32285
rect 6153 32229 6209 32285
rect 6233 32229 6289 32285
rect 5112 32147 5168 32203
rect 5193 32147 5249 32203
rect 5273 32147 5329 32203
rect 5353 32147 5409 32203
rect 5433 32147 5489 32203
rect 5513 32147 5569 32203
rect 5593 32147 5649 32203
rect 5673 32147 5729 32203
rect 5753 32147 5809 32203
rect 5833 32147 5889 32203
rect 5913 32147 5969 32203
rect 5993 32147 6049 32203
rect 6073 32147 6129 32203
rect 6153 32147 6209 32203
rect 6233 32147 6289 32203
rect 5112 32065 5168 32121
rect 5193 32065 5249 32121
rect 5273 32065 5329 32121
rect 5353 32065 5409 32121
rect 5433 32065 5489 32121
rect 5513 32065 5569 32121
rect 5593 32065 5649 32121
rect 5673 32065 5729 32121
rect 5753 32065 5809 32121
rect 5833 32065 5889 32121
rect 5913 32065 5969 32121
rect 5993 32065 6049 32121
rect 6073 32065 6129 32121
rect 6153 32065 6209 32121
rect 6233 32065 6289 32121
rect 5112 31983 5168 32039
rect 5193 31983 5249 32039
rect 5273 31983 5329 32039
rect 5353 31983 5409 32039
rect 5433 31983 5489 32039
rect 5513 31983 5569 32039
rect 5593 31983 5649 32039
rect 5673 31983 5729 32039
rect 5753 31983 5809 32039
rect 5833 31983 5889 32039
rect 5913 31983 5969 32039
rect 5993 31983 6049 32039
rect 6073 31983 6129 32039
rect 6153 31983 6209 32039
rect 6233 31983 6289 32039
rect 5112 31901 5168 31957
rect 5193 31901 5249 31957
rect 5273 31901 5329 31957
rect 5353 31901 5409 31957
rect 5433 31901 5489 31957
rect 5513 31901 5569 31957
rect 5593 31901 5649 31957
rect 5673 31901 5729 31957
rect 5753 31901 5809 31957
rect 5833 31901 5889 31957
rect 5913 31901 5969 31957
rect 5993 31901 6049 31957
rect 6073 31901 6129 31957
rect 6153 31901 6209 31957
rect 6233 31901 6289 31957
rect 5112 31819 5168 31875
rect 5193 31819 5249 31875
rect 5273 31819 5329 31875
rect 5353 31819 5409 31875
rect 5433 31819 5489 31875
rect 5513 31819 5569 31875
rect 5593 31819 5649 31875
rect 5673 31819 5729 31875
rect 5753 31819 5809 31875
rect 5833 31819 5889 31875
rect 5913 31819 5969 31875
rect 5993 31819 6049 31875
rect 6073 31819 6129 31875
rect 6153 31819 6209 31875
rect 6233 31819 6289 31875
rect 5112 31737 5168 31793
rect 5193 31737 5249 31793
rect 5273 31737 5329 31793
rect 5353 31737 5409 31793
rect 5433 31737 5489 31793
rect 5513 31737 5569 31793
rect 5593 31737 5649 31793
rect 5673 31737 5729 31793
rect 5753 31737 5809 31793
rect 5833 31737 5889 31793
rect 5913 31737 5969 31793
rect 5993 31737 6049 31793
rect 6073 31737 6129 31793
rect 6153 31737 6209 31793
rect 6233 31737 6289 31793
rect 5112 31655 5168 31711
rect 5193 31655 5249 31711
rect 5273 31655 5329 31711
rect 5353 31655 5409 31711
rect 5433 31655 5489 31711
rect 5513 31655 5569 31711
rect 5593 31655 5649 31711
rect 5673 31655 5729 31711
rect 5753 31655 5809 31711
rect 5833 31655 5889 31711
rect 5913 31655 5969 31711
rect 5993 31655 6049 31711
rect 6073 31655 6129 31711
rect 6153 31655 6209 31711
rect 6233 31655 6289 31711
rect 5112 31573 5168 31629
rect 5193 31573 5249 31629
rect 5273 31573 5329 31629
rect 5353 31573 5409 31629
rect 5433 31573 5489 31629
rect 5513 31573 5569 31629
rect 5593 31573 5649 31629
rect 5673 31573 5729 31629
rect 5753 31573 5809 31629
rect 5833 31573 5889 31629
rect 5913 31573 5969 31629
rect 5993 31573 6049 31629
rect 6073 31573 6129 31629
rect 6153 31573 6209 31629
rect 6233 31573 6289 31629
rect 5112 31491 5168 31547
rect 5193 31491 5249 31547
rect 5273 31491 5329 31547
rect 5353 31491 5409 31547
rect 5433 31491 5489 31547
rect 5513 31491 5569 31547
rect 5593 31491 5649 31547
rect 5673 31491 5729 31547
rect 5753 31491 5809 31547
rect 5833 31491 5889 31547
rect 5913 31491 5969 31547
rect 5993 31491 6049 31547
rect 6073 31491 6129 31547
rect 6153 31491 6209 31547
rect 6233 31491 6289 31547
rect 6610 32557 6666 32613
rect 6691 32557 6747 32613
rect 6772 32557 6828 32613
rect 6853 32557 6909 32613
rect 6934 32557 6990 32613
rect 7014 32557 7070 32613
rect 7094 32557 7150 32613
rect 7174 32557 7230 32613
rect 7254 32557 7310 32613
rect 7334 32557 7390 32613
rect 7414 32557 7470 32613
rect 7494 32557 7550 32613
rect 7574 32557 7630 32613
rect 7654 32557 7710 32613
rect 7734 32557 7790 32613
rect 6610 32475 6666 32531
rect 6691 32475 6747 32531
rect 6772 32475 6828 32531
rect 6853 32475 6909 32531
rect 6934 32475 6990 32531
rect 7014 32475 7070 32531
rect 7094 32475 7150 32531
rect 7174 32475 7230 32531
rect 7254 32475 7310 32531
rect 7334 32475 7390 32531
rect 7414 32475 7470 32531
rect 7494 32475 7550 32531
rect 7574 32475 7630 32531
rect 7654 32475 7710 32531
rect 7734 32475 7790 32531
rect 6610 32393 6666 32449
rect 6691 32393 6747 32449
rect 6772 32393 6828 32449
rect 6853 32393 6909 32449
rect 6934 32393 6990 32449
rect 7014 32393 7070 32449
rect 7094 32393 7150 32449
rect 7174 32393 7230 32449
rect 7254 32393 7310 32449
rect 7334 32393 7390 32449
rect 7414 32393 7470 32449
rect 7494 32393 7550 32449
rect 7574 32393 7630 32449
rect 7654 32393 7710 32449
rect 7734 32393 7790 32449
rect 6610 32311 6666 32367
rect 6691 32311 6747 32367
rect 6772 32311 6828 32367
rect 6853 32311 6909 32367
rect 6934 32311 6990 32367
rect 7014 32311 7070 32367
rect 7094 32311 7150 32367
rect 7174 32311 7230 32367
rect 7254 32311 7310 32367
rect 7334 32311 7390 32367
rect 7414 32311 7470 32367
rect 7494 32311 7550 32367
rect 7574 32311 7630 32367
rect 7654 32311 7710 32367
rect 7734 32311 7790 32367
rect 6610 32229 6666 32285
rect 6691 32229 6747 32285
rect 6772 32229 6828 32285
rect 6853 32229 6909 32285
rect 6934 32229 6990 32285
rect 7014 32229 7070 32285
rect 7094 32229 7150 32285
rect 7174 32229 7230 32285
rect 7254 32229 7310 32285
rect 7334 32229 7390 32285
rect 7414 32229 7470 32285
rect 7494 32229 7550 32285
rect 7574 32229 7630 32285
rect 7654 32229 7710 32285
rect 7734 32229 7790 32285
rect 6610 32147 6666 32203
rect 6691 32147 6747 32203
rect 6772 32147 6828 32203
rect 6853 32147 6909 32203
rect 6934 32147 6990 32203
rect 7014 32147 7070 32203
rect 7094 32147 7150 32203
rect 7174 32147 7230 32203
rect 7254 32147 7310 32203
rect 7334 32147 7390 32203
rect 7414 32147 7470 32203
rect 7494 32147 7550 32203
rect 7574 32147 7630 32203
rect 7654 32147 7710 32203
rect 7734 32147 7790 32203
rect 6610 32065 6666 32121
rect 6691 32065 6747 32121
rect 6772 32065 6828 32121
rect 6853 32065 6909 32121
rect 6934 32065 6990 32121
rect 7014 32065 7070 32121
rect 7094 32065 7150 32121
rect 7174 32065 7230 32121
rect 7254 32065 7310 32121
rect 7334 32065 7390 32121
rect 7414 32065 7470 32121
rect 7494 32065 7550 32121
rect 7574 32065 7630 32121
rect 7654 32065 7710 32121
rect 7734 32065 7790 32121
rect 6610 31983 6666 32039
rect 6691 31983 6747 32039
rect 6772 31983 6828 32039
rect 6853 31983 6909 32039
rect 6934 31983 6990 32039
rect 7014 31983 7070 32039
rect 7094 31983 7150 32039
rect 7174 31983 7230 32039
rect 7254 31983 7310 32039
rect 7334 31983 7390 32039
rect 7414 31983 7470 32039
rect 7494 31983 7550 32039
rect 7574 31983 7630 32039
rect 7654 31983 7710 32039
rect 7734 31983 7790 32039
rect 6610 31901 6666 31957
rect 6691 31901 6747 31957
rect 6772 31901 6828 31957
rect 6853 31901 6909 31957
rect 6934 31901 6990 31957
rect 7014 31901 7070 31957
rect 7094 31901 7150 31957
rect 7174 31901 7230 31957
rect 7254 31901 7310 31957
rect 7334 31901 7390 31957
rect 7414 31901 7470 31957
rect 7494 31901 7550 31957
rect 7574 31901 7630 31957
rect 7654 31901 7710 31957
rect 7734 31901 7790 31957
rect 6610 31819 6666 31875
rect 6691 31819 6747 31875
rect 6772 31819 6828 31875
rect 6853 31819 6909 31875
rect 6934 31819 6990 31875
rect 7014 31819 7070 31875
rect 7094 31819 7150 31875
rect 7174 31819 7230 31875
rect 7254 31819 7310 31875
rect 7334 31819 7390 31875
rect 7414 31819 7470 31875
rect 7494 31819 7550 31875
rect 7574 31819 7630 31875
rect 7654 31819 7710 31875
rect 7734 31819 7790 31875
rect 6610 31737 6666 31793
rect 6691 31737 6747 31793
rect 6772 31737 6828 31793
rect 6853 31737 6909 31793
rect 6934 31737 6990 31793
rect 7014 31737 7070 31793
rect 7094 31737 7150 31793
rect 7174 31737 7230 31793
rect 7254 31737 7310 31793
rect 7334 31737 7390 31793
rect 7414 31737 7470 31793
rect 7494 31737 7550 31793
rect 7574 31737 7630 31793
rect 7654 31737 7710 31793
rect 7734 31737 7790 31793
rect 6610 31655 6666 31711
rect 6691 31655 6747 31711
rect 6772 31655 6828 31711
rect 6853 31655 6909 31711
rect 6934 31655 6990 31711
rect 7014 31655 7070 31711
rect 7094 31655 7150 31711
rect 7174 31655 7230 31711
rect 7254 31655 7310 31711
rect 7334 31655 7390 31711
rect 7414 31655 7470 31711
rect 7494 31655 7550 31711
rect 7574 31655 7630 31711
rect 7654 31655 7710 31711
rect 7734 31655 7790 31711
rect 6610 31573 6666 31629
rect 6691 31573 6747 31629
rect 6772 31573 6828 31629
rect 6853 31573 6909 31629
rect 6934 31573 6990 31629
rect 7014 31573 7070 31629
rect 7094 31573 7150 31629
rect 7174 31573 7230 31629
rect 7254 31573 7310 31629
rect 7334 31573 7390 31629
rect 7414 31573 7470 31629
rect 7494 31573 7550 31629
rect 7574 31573 7630 31629
rect 7654 31573 7710 31629
rect 7734 31573 7790 31629
rect 6610 31491 6666 31547
rect 6691 31491 6747 31547
rect 6772 31491 6828 31547
rect 6853 31491 6909 31547
rect 6934 31491 6990 31547
rect 7014 31491 7070 31547
rect 7094 31491 7150 31547
rect 7174 31491 7230 31547
rect 7254 31491 7310 31547
rect 7334 31491 7390 31547
rect 7414 31491 7470 31547
rect 7494 31491 7550 31547
rect 7574 31491 7630 31547
rect 7654 31491 7710 31547
rect 7734 31491 7790 31547
rect 8107 32557 8163 32613
rect 8188 32557 8244 32613
rect 8269 32557 8325 32613
rect 8350 32557 8406 32613
rect 8431 32557 8487 32613
rect 8511 32557 8567 32613
rect 8591 32557 8647 32613
rect 8671 32557 8727 32613
rect 8751 32557 8807 32613
rect 8831 32557 8887 32613
rect 8911 32557 8967 32613
rect 8991 32557 9047 32613
rect 9071 32557 9127 32613
rect 9151 32557 9207 32613
rect 9231 32557 9287 32613
rect 8107 32475 8163 32531
rect 8188 32475 8244 32531
rect 8269 32475 8325 32531
rect 8350 32475 8406 32531
rect 8431 32475 8487 32531
rect 8511 32475 8567 32531
rect 8591 32475 8647 32531
rect 8671 32475 8727 32531
rect 8751 32475 8807 32531
rect 8831 32475 8887 32531
rect 8911 32475 8967 32531
rect 8991 32475 9047 32531
rect 9071 32475 9127 32531
rect 9151 32475 9207 32531
rect 9231 32475 9287 32531
rect 8107 32393 8163 32449
rect 8188 32393 8244 32449
rect 8269 32393 8325 32449
rect 8350 32393 8406 32449
rect 8431 32393 8487 32449
rect 8511 32393 8567 32449
rect 8591 32393 8647 32449
rect 8671 32393 8727 32449
rect 8751 32393 8807 32449
rect 8831 32393 8887 32449
rect 8911 32393 8967 32449
rect 8991 32393 9047 32449
rect 9071 32393 9127 32449
rect 9151 32393 9207 32449
rect 9231 32393 9287 32449
rect 8107 32311 8163 32367
rect 8188 32311 8244 32367
rect 8269 32311 8325 32367
rect 8350 32311 8406 32367
rect 8431 32311 8487 32367
rect 8511 32311 8567 32367
rect 8591 32311 8647 32367
rect 8671 32311 8727 32367
rect 8751 32311 8807 32367
rect 8831 32311 8887 32367
rect 8911 32311 8967 32367
rect 8991 32311 9047 32367
rect 9071 32311 9127 32367
rect 9151 32311 9207 32367
rect 9231 32311 9287 32367
rect 8107 32229 8163 32285
rect 8188 32229 8244 32285
rect 8269 32229 8325 32285
rect 8350 32229 8406 32285
rect 8431 32229 8487 32285
rect 8511 32229 8567 32285
rect 8591 32229 8647 32285
rect 8671 32229 8727 32285
rect 8751 32229 8807 32285
rect 8831 32229 8887 32285
rect 8911 32229 8967 32285
rect 8991 32229 9047 32285
rect 9071 32229 9127 32285
rect 9151 32229 9207 32285
rect 9231 32229 9287 32285
rect 8107 32147 8163 32203
rect 8188 32147 8244 32203
rect 8269 32147 8325 32203
rect 8350 32147 8406 32203
rect 8431 32147 8487 32203
rect 8511 32147 8567 32203
rect 8591 32147 8647 32203
rect 8671 32147 8727 32203
rect 8751 32147 8807 32203
rect 8831 32147 8887 32203
rect 8911 32147 8967 32203
rect 8991 32147 9047 32203
rect 9071 32147 9127 32203
rect 9151 32147 9207 32203
rect 9231 32147 9287 32203
rect 8107 32065 8163 32121
rect 8188 32065 8244 32121
rect 8269 32065 8325 32121
rect 8350 32065 8406 32121
rect 8431 32065 8487 32121
rect 8511 32065 8567 32121
rect 8591 32065 8647 32121
rect 8671 32065 8727 32121
rect 8751 32065 8807 32121
rect 8831 32065 8887 32121
rect 8911 32065 8967 32121
rect 8991 32065 9047 32121
rect 9071 32065 9127 32121
rect 9151 32065 9207 32121
rect 9231 32065 9287 32121
rect 8107 31983 8163 32039
rect 8188 31983 8244 32039
rect 8269 31983 8325 32039
rect 8350 31983 8406 32039
rect 8431 31983 8487 32039
rect 8511 31983 8567 32039
rect 8591 31983 8647 32039
rect 8671 31983 8727 32039
rect 8751 31983 8807 32039
rect 8831 31983 8887 32039
rect 8911 31983 8967 32039
rect 8991 31983 9047 32039
rect 9071 31983 9127 32039
rect 9151 31983 9207 32039
rect 9231 31983 9287 32039
rect 8107 31901 8163 31957
rect 8188 31901 8244 31957
rect 8269 31901 8325 31957
rect 8350 31901 8406 31957
rect 8431 31901 8487 31957
rect 8511 31901 8567 31957
rect 8591 31901 8647 31957
rect 8671 31901 8727 31957
rect 8751 31901 8807 31957
rect 8831 31901 8887 31957
rect 8911 31901 8967 31957
rect 8991 31901 9047 31957
rect 9071 31901 9127 31957
rect 9151 31901 9207 31957
rect 9231 31901 9287 31957
rect 8107 31819 8163 31875
rect 8188 31819 8244 31875
rect 8269 31819 8325 31875
rect 8350 31819 8406 31875
rect 8431 31819 8487 31875
rect 8511 31819 8567 31875
rect 8591 31819 8647 31875
rect 8671 31819 8727 31875
rect 8751 31819 8807 31875
rect 8831 31819 8887 31875
rect 8911 31819 8967 31875
rect 8991 31819 9047 31875
rect 9071 31819 9127 31875
rect 9151 31819 9207 31875
rect 9231 31819 9287 31875
rect 8107 31737 8163 31793
rect 8188 31737 8244 31793
rect 8269 31737 8325 31793
rect 8350 31737 8406 31793
rect 8431 31737 8487 31793
rect 8511 31737 8567 31793
rect 8591 31737 8647 31793
rect 8671 31737 8727 31793
rect 8751 31737 8807 31793
rect 8831 31737 8887 31793
rect 8911 31737 8967 31793
rect 8991 31737 9047 31793
rect 9071 31737 9127 31793
rect 9151 31737 9207 31793
rect 9231 31737 9287 31793
rect 8107 31655 8163 31711
rect 8188 31655 8244 31711
rect 8269 31655 8325 31711
rect 8350 31655 8406 31711
rect 8431 31655 8487 31711
rect 8511 31655 8567 31711
rect 8591 31655 8647 31711
rect 8671 31655 8727 31711
rect 8751 31655 8807 31711
rect 8831 31655 8887 31711
rect 8911 31655 8967 31711
rect 8991 31655 9047 31711
rect 9071 31655 9127 31711
rect 9151 31655 9207 31711
rect 9231 31655 9287 31711
rect 8107 31573 8163 31629
rect 8188 31573 8244 31629
rect 8269 31573 8325 31629
rect 8350 31573 8406 31629
rect 8431 31573 8487 31629
rect 8511 31573 8567 31629
rect 8591 31573 8647 31629
rect 8671 31573 8727 31629
rect 8751 31573 8807 31629
rect 8831 31573 8887 31629
rect 8911 31573 8967 31629
rect 8991 31573 9047 31629
rect 9071 31573 9127 31629
rect 9151 31573 9207 31629
rect 9231 31573 9287 31629
rect 8107 31491 8163 31547
rect 8188 31491 8244 31547
rect 8269 31491 8325 31547
rect 8350 31491 8406 31547
rect 8431 31491 8487 31547
rect 8511 31491 8567 31547
rect 8591 31491 8647 31547
rect 8671 31491 8727 31547
rect 8751 31491 8807 31547
rect 8831 31491 8887 31547
rect 8911 31491 8967 31547
rect 8991 31491 9047 31547
rect 9071 31491 9127 31547
rect 9151 31491 9207 31547
rect 9231 31491 9287 31547
rect 9604 32557 9660 32613
rect 9685 32557 9741 32613
rect 9766 32557 9822 32613
rect 9847 32557 9903 32613
rect 9928 32557 9984 32613
rect 10008 32557 10064 32613
rect 10088 32557 10144 32613
rect 10168 32557 10224 32613
rect 10248 32557 10304 32613
rect 10328 32557 10384 32613
rect 10408 32557 10464 32613
rect 10488 32557 10544 32613
rect 10568 32557 10624 32613
rect 10648 32557 10704 32613
rect 10728 32557 10784 32613
rect 9604 32475 9660 32531
rect 9685 32475 9741 32531
rect 9766 32475 9822 32531
rect 9847 32475 9903 32531
rect 9928 32475 9984 32531
rect 10008 32475 10064 32531
rect 10088 32475 10144 32531
rect 10168 32475 10224 32531
rect 10248 32475 10304 32531
rect 10328 32475 10384 32531
rect 10408 32475 10464 32531
rect 10488 32475 10544 32531
rect 10568 32475 10624 32531
rect 10648 32475 10704 32531
rect 10728 32475 10784 32531
rect 9604 32393 9660 32449
rect 9685 32393 9741 32449
rect 9766 32393 9822 32449
rect 9847 32393 9903 32449
rect 9928 32393 9984 32449
rect 10008 32393 10064 32449
rect 10088 32393 10144 32449
rect 10168 32393 10224 32449
rect 10248 32393 10304 32449
rect 10328 32393 10384 32449
rect 10408 32393 10464 32449
rect 10488 32393 10544 32449
rect 10568 32393 10624 32449
rect 10648 32393 10704 32449
rect 10728 32393 10784 32449
rect 9604 32311 9660 32367
rect 9685 32311 9741 32367
rect 9766 32311 9822 32367
rect 9847 32311 9903 32367
rect 9928 32311 9984 32367
rect 10008 32311 10064 32367
rect 10088 32311 10144 32367
rect 10168 32311 10224 32367
rect 10248 32311 10304 32367
rect 10328 32311 10384 32367
rect 10408 32311 10464 32367
rect 10488 32311 10544 32367
rect 10568 32311 10624 32367
rect 10648 32311 10704 32367
rect 10728 32311 10784 32367
rect 9604 32229 9660 32285
rect 9685 32229 9741 32285
rect 9766 32229 9822 32285
rect 9847 32229 9903 32285
rect 9928 32229 9984 32285
rect 10008 32229 10064 32285
rect 10088 32229 10144 32285
rect 10168 32229 10224 32285
rect 10248 32229 10304 32285
rect 10328 32229 10384 32285
rect 10408 32229 10464 32285
rect 10488 32229 10544 32285
rect 10568 32229 10624 32285
rect 10648 32229 10704 32285
rect 10728 32229 10784 32285
rect 9604 32147 9660 32203
rect 9685 32147 9741 32203
rect 9766 32147 9822 32203
rect 9847 32147 9903 32203
rect 9928 32147 9984 32203
rect 10008 32147 10064 32203
rect 10088 32147 10144 32203
rect 10168 32147 10224 32203
rect 10248 32147 10304 32203
rect 10328 32147 10384 32203
rect 10408 32147 10464 32203
rect 10488 32147 10544 32203
rect 10568 32147 10624 32203
rect 10648 32147 10704 32203
rect 10728 32147 10784 32203
rect 9604 32065 9660 32121
rect 9685 32065 9741 32121
rect 9766 32065 9822 32121
rect 9847 32065 9903 32121
rect 9928 32065 9984 32121
rect 10008 32065 10064 32121
rect 10088 32065 10144 32121
rect 10168 32065 10224 32121
rect 10248 32065 10304 32121
rect 10328 32065 10384 32121
rect 10408 32065 10464 32121
rect 10488 32065 10544 32121
rect 10568 32065 10624 32121
rect 10648 32065 10704 32121
rect 10728 32065 10784 32121
rect 9604 31983 9660 32039
rect 9685 31983 9741 32039
rect 9766 31983 9822 32039
rect 9847 31983 9903 32039
rect 9928 31983 9984 32039
rect 10008 31983 10064 32039
rect 10088 31983 10144 32039
rect 10168 31983 10224 32039
rect 10248 31983 10304 32039
rect 10328 31983 10384 32039
rect 10408 31983 10464 32039
rect 10488 31983 10544 32039
rect 10568 31983 10624 32039
rect 10648 31983 10704 32039
rect 10728 31983 10784 32039
rect 9604 31901 9660 31957
rect 9685 31901 9741 31957
rect 9766 31901 9822 31957
rect 9847 31901 9903 31957
rect 9928 31901 9984 31957
rect 10008 31901 10064 31957
rect 10088 31901 10144 31957
rect 10168 31901 10224 31957
rect 10248 31901 10304 31957
rect 10328 31901 10384 31957
rect 10408 31901 10464 31957
rect 10488 31901 10544 31957
rect 10568 31901 10624 31957
rect 10648 31901 10704 31957
rect 10728 31901 10784 31957
rect 9604 31819 9660 31875
rect 9685 31819 9741 31875
rect 9766 31819 9822 31875
rect 9847 31819 9903 31875
rect 9928 31819 9984 31875
rect 10008 31819 10064 31875
rect 10088 31819 10144 31875
rect 10168 31819 10224 31875
rect 10248 31819 10304 31875
rect 10328 31819 10384 31875
rect 10408 31819 10464 31875
rect 10488 31819 10544 31875
rect 10568 31819 10624 31875
rect 10648 31819 10704 31875
rect 10728 31819 10784 31875
rect 9604 31737 9660 31793
rect 9685 31737 9741 31793
rect 9766 31737 9822 31793
rect 9847 31737 9903 31793
rect 9928 31737 9984 31793
rect 10008 31737 10064 31793
rect 10088 31737 10144 31793
rect 10168 31737 10224 31793
rect 10248 31737 10304 31793
rect 10328 31737 10384 31793
rect 10408 31737 10464 31793
rect 10488 31737 10544 31793
rect 10568 31737 10624 31793
rect 10648 31737 10704 31793
rect 10728 31737 10784 31793
rect 9604 31655 9660 31711
rect 9685 31655 9741 31711
rect 9766 31655 9822 31711
rect 9847 31655 9903 31711
rect 9928 31655 9984 31711
rect 10008 31655 10064 31711
rect 10088 31655 10144 31711
rect 10168 31655 10224 31711
rect 10248 31655 10304 31711
rect 10328 31655 10384 31711
rect 10408 31655 10464 31711
rect 10488 31655 10544 31711
rect 10568 31655 10624 31711
rect 10648 31655 10704 31711
rect 10728 31655 10784 31711
rect 9604 31573 9660 31629
rect 9685 31573 9741 31629
rect 9766 31573 9822 31629
rect 9847 31573 9903 31629
rect 9928 31573 9984 31629
rect 10008 31573 10064 31629
rect 10088 31573 10144 31629
rect 10168 31573 10224 31629
rect 10248 31573 10304 31629
rect 10328 31573 10384 31629
rect 10408 31573 10464 31629
rect 10488 31573 10544 31629
rect 10568 31573 10624 31629
rect 10648 31573 10704 31629
rect 10728 31573 10784 31629
rect 9604 31491 9660 31547
rect 9685 31491 9741 31547
rect 9766 31491 9822 31547
rect 9847 31491 9903 31547
rect 9928 31491 9984 31547
rect 10008 31491 10064 31547
rect 10088 31491 10144 31547
rect 10168 31491 10224 31547
rect 10248 31491 10304 31547
rect 10328 31491 10384 31547
rect 10408 31491 10464 31547
rect 10488 31491 10544 31547
rect 10568 31491 10624 31547
rect 10648 31491 10704 31547
rect 10728 31491 10784 31547
rect 11101 32557 11157 32613
rect 11182 32557 11238 32613
rect 11263 32557 11319 32613
rect 11344 32557 11400 32613
rect 11425 32557 11481 32613
rect 11505 32557 11561 32613
rect 11585 32557 11641 32613
rect 11665 32557 11721 32613
rect 11745 32557 11801 32613
rect 11825 32557 11881 32613
rect 11905 32557 11961 32613
rect 11985 32557 12041 32613
rect 12065 32557 12121 32613
rect 12145 32557 12201 32613
rect 12225 32557 12281 32613
rect 11101 32475 11157 32531
rect 11182 32475 11238 32531
rect 11263 32475 11319 32531
rect 11344 32475 11400 32531
rect 11425 32475 11481 32531
rect 11505 32475 11561 32531
rect 11585 32475 11641 32531
rect 11665 32475 11721 32531
rect 11745 32475 11801 32531
rect 11825 32475 11881 32531
rect 11905 32475 11961 32531
rect 11985 32475 12041 32531
rect 12065 32475 12121 32531
rect 12145 32475 12201 32531
rect 12225 32475 12281 32531
rect 11101 32393 11157 32449
rect 11182 32393 11238 32449
rect 11263 32393 11319 32449
rect 11344 32393 11400 32449
rect 11425 32393 11481 32449
rect 11505 32393 11561 32449
rect 11585 32393 11641 32449
rect 11665 32393 11721 32449
rect 11745 32393 11801 32449
rect 11825 32393 11881 32449
rect 11905 32393 11961 32449
rect 11985 32393 12041 32449
rect 12065 32393 12121 32449
rect 12145 32393 12201 32449
rect 12225 32393 12281 32449
rect 11101 32311 11157 32367
rect 11182 32311 11238 32367
rect 11263 32311 11319 32367
rect 11344 32311 11400 32367
rect 11425 32311 11481 32367
rect 11505 32311 11561 32367
rect 11585 32311 11641 32367
rect 11665 32311 11721 32367
rect 11745 32311 11801 32367
rect 11825 32311 11881 32367
rect 11905 32311 11961 32367
rect 11985 32311 12041 32367
rect 12065 32311 12121 32367
rect 12145 32311 12201 32367
rect 12225 32311 12281 32367
rect 11101 32229 11157 32285
rect 11182 32229 11238 32285
rect 11263 32229 11319 32285
rect 11344 32229 11400 32285
rect 11425 32229 11481 32285
rect 11505 32229 11561 32285
rect 11585 32229 11641 32285
rect 11665 32229 11721 32285
rect 11745 32229 11801 32285
rect 11825 32229 11881 32285
rect 11905 32229 11961 32285
rect 11985 32229 12041 32285
rect 12065 32229 12121 32285
rect 12145 32229 12201 32285
rect 12225 32229 12281 32285
rect 11101 32147 11157 32203
rect 11182 32147 11238 32203
rect 11263 32147 11319 32203
rect 11344 32147 11400 32203
rect 11425 32147 11481 32203
rect 11505 32147 11561 32203
rect 11585 32147 11641 32203
rect 11665 32147 11721 32203
rect 11745 32147 11801 32203
rect 11825 32147 11881 32203
rect 11905 32147 11961 32203
rect 11985 32147 12041 32203
rect 12065 32147 12121 32203
rect 12145 32147 12201 32203
rect 12225 32147 12281 32203
rect 11101 32065 11157 32121
rect 11182 32065 11238 32121
rect 11263 32065 11319 32121
rect 11344 32065 11400 32121
rect 11425 32065 11481 32121
rect 11505 32065 11561 32121
rect 11585 32065 11641 32121
rect 11665 32065 11721 32121
rect 11745 32065 11801 32121
rect 11825 32065 11881 32121
rect 11905 32065 11961 32121
rect 11985 32065 12041 32121
rect 12065 32065 12121 32121
rect 12145 32065 12201 32121
rect 12225 32065 12281 32121
rect 11101 31983 11157 32039
rect 11182 31983 11238 32039
rect 11263 31983 11319 32039
rect 11344 31983 11400 32039
rect 11425 31983 11481 32039
rect 11505 31983 11561 32039
rect 11585 31983 11641 32039
rect 11665 31983 11721 32039
rect 11745 31983 11801 32039
rect 11825 31983 11881 32039
rect 11905 31983 11961 32039
rect 11985 31983 12041 32039
rect 12065 31983 12121 32039
rect 12145 31983 12201 32039
rect 12225 31983 12281 32039
rect 11101 31901 11157 31957
rect 11182 31901 11238 31957
rect 11263 31901 11319 31957
rect 11344 31901 11400 31957
rect 11425 31901 11481 31957
rect 11505 31901 11561 31957
rect 11585 31901 11641 31957
rect 11665 31901 11721 31957
rect 11745 31901 11801 31957
rect 11825 31901 11881 31957
rect 11905 31901 11961 31957
rect 11985 31901 12041 31957
rect 12065 31901 12121 31957
rect 12145 31901 12201 31957
rect 12225 31901 12281 31957
rect 11101 31819 11157 31875
rect 11182 31819 11238 31875
rect 11263 31819 11319 31875
rect 11344 31819 11400 31875
rect 11425 31819 11481 31875
rect 11505 31819 11561 31875
rect 11585 31819 11641 31875
rect 11665 31819 11721 31875
rect 11745 31819 11801 31875
rect 11825 31819 11881 31875
rect 11905 31819 11961 31875
rect 11985 31819 12041 31875
rect 12065 31819 12121 31875
rect 12145 31819 12201 31875
rect 12225 31819 12281 31875
rect 11101 31737 11157 31793
rect 11182 31737 11238 31793
rect 11263 31737 11319 31793
rect 11344 31737 11400 31793
rect 11425 31737 11481 31793
rect 11505 31737 11561 31793
rect 11585 31737 11641 31793
rect 11665 31737 11721 31793
rect 11745 31737 11801 31793
rect 11825 31737 11881 31793
rect 11905 31737 11961 31793
rect 11985 31737 12041 31793
rect 12065 31737 12121 31793
rect 12145 31737 12201 31793
rect 12225 31737 12281 31793
rect 11101 31655 11157 31711
rect 11182 31655 11238 31711
rect 11263 31655 11319 31711
rect 11344 31655 11400 31711
rect 11425 31655 11481 31711
rect 11505 31655 11561 31711
rect 11585 31655 11641 31711
rect 11665 31655 11721 31711
rect 11745 31655 11801 31711
rect 11825 31655 11881 31711
rect 11905 31655 11961 31711
rect 11985 31655 12041 31711
rect 12065 31655 12121 31711
rect 12145 31655 12201 31711
rect 12225 31655 12281 31711
rect 11101 31573 11157 31629
rect 11182 31573 11238 31629
rect 11263 31573 11319 31629
rect 11344 31573 11400 31629
rect 11425 31573 11481 31629
rect 11505 31573 11561 31629
rect 11585 31573 11641 31629
rect 11665 31573 11721 31629
rect 11745 31573 11801 31629
rect 11825 31573 11881 31629
rect 11905 31573 11961 31629
rect 11985 31573 12041 31629
rect 12065 31573 12121 31629
rect 12145 31573 12201 31629
rect 12225 31573 12281 31629
rect 11101 31491 11157 31547
rect 11182 31491 11238 31547
rect 11263 31491 11319 31547
rect 11344 31491 11400 31547
rect 11425 31491 11481 31547
rect 11505 31491 11561 31547
rect 11585 31491 11641 31547
rect 11665 31491 11721 31547
rect 11745 31491 11801 31547
rect 11825 31491 11881 31547
rect 11905 31491 11961 31547
rect 11985 31491 12041 31547
rect 12065 31491 12121 31547
rect 12145 31491 12201 31547
rect 12225 31491 12281 31547
rect 12598 32557 12654 32613
rect 12685 32557 12741 32613
rect 12772 32557 12828 32613
rect 12859 32557 12915 32613
rect 12945 32557 13001 32613
rect 13031 32557 13087 32613
rect 13117 32557 13173 32613
rect 13203 32557 13259 32613
rect 12598 32475 12654 32531
rect 12685 32475 12741 32531
rect 12772 32475 12828 32531
rect 12859 32475 12915 32531
rect 12945 32475 13001 32531
rect 13031 32475 13087 32531
rect 13117 32475 13173 32531
rect 13203 32475 13259 32531
rect 12598 32393 12654 32449
rect 12685 32393 12741 32449
rect 12772 32393 12828 32449
rect 12859 32393 12915 32449
rect 12945 32393 13001 32449
rect 13031 32393 13087 32449
rect 13117 32393 13173 32449
rect 13203 32393 13259 32449
rect 12598 32311 12654 32367
rect 12685 32311 12741 32367
rect 12772 32311 12828 32367
rect 12859 32311 12915 32367
rect 12945 32311 13001 32367
rect 13031 32311 13087 32367
rect 13117 32311 13173 32367
rect 13203 32311 13259 32367
rect 12598 32229 12654 32285
rect 12685 32229 12741 32285
rect 12772 32229 12828 32285
rect 12859 32229 12915 32285
rect 12945 32229 13001 32285
rect 13031 32229 13087 32285
rect 13117 32229 13173 32285
rect 13203 32229 13259 32285
rect 12598 32147 12654 32203
rect 12685 32147 12741 32203
rect 12772 32147 12828 32203
rect 12859 32147 12915 32203
rect 12945 32147 13001 32203
rect 13031 32147 13087 32203
rect 13117 32147 13173 32203
rect 13203 32147 13259 32203
rect 12598 32065 12654 32121
rect 12685 32065 12741 32121
rect 12772 32065 12828 32121
rect 12859 32065 12915 32121
rect 12945 32065 13001 32121
rect 13031 32065 13087 32121
rect 13117 32065 13173 32121
rect 13203 32065 13259 32121
rect 12598 31983 12654 32039
rect 12685 31983 12741 32039
rect 12772 31983 12828 32039
rect 12859 31983 12915 32039
rect 12945 31983 13001 32039
rect 13031 31983 13087 32039
rect 13117 31983 13173 32039
rect 13203 31983 13259 32039
rect 12598 31901 12654 31957
rect 12685 31901 12741 31957
rect 12772 31901 12828 31957
rect 12859 31901 12915 31957
rect 12945 31901 13001 31957
rect 13031 31901 13087 31957
rect 13117 31901 13173 31957
rect 13203 31901 13259 31957
rect 12598 31819 12654 31875
rect 12685 31819 12741 31875
rect 12772 31819 12828 31875
rect 12859 31819 12915 31875
rect 12945 31819 13001 31875
rect 13031 31819 13087 31875
rect 13117 31819 13173 31875
rect 13203 31819 13259 31875
rect 12598 31737 12654 31793
rect 12685 31737 12741 31793
rect 12772 31737 12828 31793
rect 12859 31737 12915 31793
rect 12945 31737 13001 31793
rect 13031 31737 13087 31793
rect 13117 31737 13173 31793
rect 13203 31737 13259 31793
rect 12598 31655 12654 31711
rect 12685 31655 12741 31711
rect 12772 31655 12828 31711
rect 12859 31655 12915 31711
rect 12945 31655 13001 31711
rect 13031 31655 13087 31711
rect 13117 31655 13173 31711
rect 13203 31655 13259 31711
rect 12598 31573 12654 31629
rect 12685 31573 12741 31629
rect 12772 31573 12828 31629
rect 12859 31573 12915 31629
rect 12945 31573 13001 31629
rect 13031 31573 13087 31629
rect 13117 31573 13173 31629
rect 13203 31573 13259 31629
rect 12598 31491 12654 31547
rect 12685 31491 12741 31547
rect 12772 31491 12828 31547
rect 12859 31491 12915 31547
rect 12945 31491 13001 31547
rect 13031 31491 13087 31547
rect 13117 31491 13173 31547
rect 13203 31491 13259 31547
rect 298 31442 299 31448
rect 299 31442 354 31448
rect 298 31429 354 31442
rect 298 31392 299 31429
rect 299 31392 354 31429
rect 396 31392 452 31448
rect 494 31442 506 31448
rect 506 31442 528 31448
rect 528 31442 550 31448
rect 592 31442 602 31448
rect 602 31442 648 31448
rect 494 31429 550 31442
rect 592 31429 648 31442
rect 494 31392 506 31429
rect 506 31392 528 31429
rect 528 31392 550 31429
rect 592 31392 602 31429
rect 602 31392 648 31429
rect 298 31364 354 31367
rect 298 31312 299 31364
rect 299 31312 354 31364
rect 298 31311 354 31312
rect 396 31311 452 31367
rect 494 31364 550 31367
rect 592 31364 648 31367
rect 494 31312 506 31364
rect 506 31312 528 31364
rect 528 31312 550 31364
rect 592 31312 602 31364
rect 602 31312 648 31364
rect 494 31311 550 31312
rect 592 31311 648 31312
rect 298 31247 299 31286
rect 299 31247 354 31286
rect 298 31234 354 31247
rect 298 31230 299 31234
rect 299 31230 354 31234
rect 396 31230 452 31286
rect 494 31247 506 31286
rect 506 31247 528 31286
rect 528 31247 550 31286
rect 592 31247 602 31286
rect 602 31247 648 31286
rect 494 31234 550 31247
rect 592 31234 648 31247
rect 494 31230 506 31234
rect 506 31230 528 31234
rect 528 31230 550 31234
rect 592 31230 602 31234
rect 602 31230 648 31234
rect 298 31182 299 31205
rect 299 31182 354 31205
rect 298 31169 354 31182
rect 298 31149 299 31169
rect 299 31149 354 31169
rect 396 31149 452 31205
rect 494 31182 506 31205
rect 506 31182 528 31205
rect 528 31182 550 31205
rect 592 31182 602 31205
rect 602 31182 648 31205
rect 494 31169 550 31182
rect 592 31169 648 31182
rect 494 31149 506 31169
rect 506 31149 528 31169
rect 528 31149 550 31169
rect 592 31149 602 31169
rect 602 31149 648 31169
rect 298 31117 299 31124
rect 299 31117 354 31124
rect 298 31104 354 31117
rect 298 31068 299 31104
rect 299 31068 354 31104
rect 396 31068 452 31124
rect 494 31117 506 31124
rect 506 31117 528 31124
rect 528 31117 550 31124
rect 592 31117 602 31124
rect 602 31117 648 31124
rect 494 31104 550 31117
rect 592 31104 648 31117
rect 494 31068 506 31104
rect 506 31068 528 31104
rect 528 31068 550 31104
rect 592 31068 602 31104
rect 602 31068 648 31104
rect 298 31039 354 31043
rect 298 30987 299 31039
rect 299 30987 354 31039
rect 396 30987 452 31043
rect 494 31039 550 31043
rect 592 31039 648 31043
rect 494 30987 506 31039
rect 506 30987 528 31039
rect 528 30987 550 31039
rect 592 30987 602 31039
rect 602 30987 648 31039
rect 298 30922 299 30962
rect 299 30922 354 30962
rect 298 30909 354 30922
rect 298 30906 299 30909
rect 299 30906 354 30909
rect 396 30906 452 30962
rect 494 30922 506 30962
rect 506 30922 528 30962
rect 528 30922 550 30962
rect 592 30922 602 30962
rect 602 30922 648 30962
rect 494 30909 550 30922
rect 592 30909 648 30922
rect 494 30906 506 30909
rect 506 30906 528 30909
rect 528 30906 550 30909
rect 592 30906 602 30909
rect 602 30906 648 30909
rect 298 30857 299 30881
rect 299 30857 354 30881
rect 298 30844 354 30857
rect 298 30825 299 30844
rect 299 30825 354 30844
rect 396 30825 452 30881
rect 494 30857 506 30881
rect 506 30857 528 30881
rect 528 30857 550 30881
rect 592 30857 602 30881
rect 602 30857 648 30881
rect 494 30844 550 30857
rect 592 30844 648 30857
rect 494 30825 506 30844
rect 506 30825 528 30844
rect 528 30825 550 30844
rect 592 30825 602 30844
rect 602 30825 648 30844
rect 298 30792 299 30800
rect 299 30792 354 30800
rect 298 30779 354 30792
rect 298 30744 299 30779
rect 299 30744 354 30779
rect 396 30744 452 30800
rect 494 30792 506 30800
rect 506 30792 528 30800
rect 528 30792 550 30800
rect 592 30792 602 30800
rect 602 30792 648 30800
rect 494 30779 550 30792
rect 592 30779 648 30792
rect 494 30744 506 30779
rect 506 30744 528 30779
rect 528 30744 550 30779
rect 592 30744 602 30779
rect 602 30744 648 30779
rect 298 30714 354 30719
rect 298 30663 299 30714
rect 299 30663 354 30714
rect 396 30663 452 30719
rect 494 30714 550 30719
rect 592 30714 648 30719
rect 494 30663 506 30714
rect 506 30663 528 30714
rect 528 30663 550 30714
rect 592 30663 602 30714
rect 602 30663 648 30714
rect 298 30597 299 30638
rect 299 30597 354 30638
rect 298 30584 354 30597
rect 298 30582 299 30584
rect 299 30582 354 30584
rect 396 30582 452 30638
rect 494 30597 506 30638
rect 506 30597 528 30638
rect 528 30597 550 30638
rect 592 30597 602 30638
rect 602 30597 648 30638
rect 494 30584 550 30597
rect 592 30584 648 30597
rect 494 30582 506 30584
rect 506 30582 528 30584
rect 528 30582 550 30584
rect 592 30582 602 30584
rect 602 30582 648 30584
rect 298 30532 299 30557
rect 299 30532 354 30557
rect 298 30519 354 30532
rect 298 30501 299 30519
rect 299 30501 354 30519
rect 396 30501 452 30557
rect 494 30532 506 30557
rect 506 30532 528 30557
rect 528 30532 550 30557
rect 592 30532 602 30557
rect 602 30532 648 30557
rect 494 30519 550 30532
rect 592 30519 648 30532
rect 494 30501 506 30519
rect 506 30501 528 30519
rect 528 30501 550 30519
rect 592 30501 602 30519
rect 602 30501 648 30519
rect 298 30467 299 30476
rect 299 30467 354 30476
rect 298 30454 354 30467
rect 298 30420 299 30454
rect 299 30420 354 30454
rect 396 30420 452 30476
rect 494 30467 506 30476
rect 506 30467 528 30476
rect 528 30467 550 30476
rect 592 30467 602 30476
rect 602 30467 648 30476
rect 494 30454 550 30467
rect 592 30454 648 30467
rect 494 30420 506 30454
rect 506 30420 528 30454
rect 528 30420 550 30454
rect 592 30420 602 30454
rect 602 30420 648 30454
rect 298 30389 354 30395
rect 298 30339 299 30389
rect 299 30339 354 30389
rect 396 30339 452 30395
rect 494 30389 550 30395
rect 592 30389 648 30395
rect 494 30339 506 30389
rect 506 30339 528 30389
rect 528 30339 550 30389
rect 592 30339 602 30389
rect 602 30339 648 30389
rect 298 30272 299 30314
rect 299 30272 354 30314
rect 298 30259 354 30272
rect 298 30258 299 30259
rect 299 30258 354 30259
rect 396 30258 452 30314
rect 494 30272 506 30314
rect 506 30272 528 30314
rect 528 30272 550 30314
rect 592 30272 602 30314
rect 602 30272 648 30314
rect 494 30259 550 30272
rect 592 30259 648 30272
rect 494 30258 506 30259
rect 506 30258 528 30259
rect 528 30258 550 30259
rect 592 30258 602 30259
rect 602 30258 648 30259
rect 298 30207 299 30233
rect 299 30207 354 30233
rect 298 30194 354 30207
rect 298 30177 299 30194
rect 299 30177 354 30194
rect 396 30177 452 30233
rect 494 30207 506 30233
rect 506 30207 528 30233
rect 528 30207 550 30233
rect 592 30207 602 30233
rect 602 30207 648 30233
rect 494 30194 550 30207
rect 592 30194 648 30207
rect 494 30177 506 30194
rect 506 30177 528 30194
rect 528 30177 550 30194
rect 592 30177 602 30194
rect 602 30177 648 30194
rect 298 30142 299 30152
rect 299 30142 354 30152
rect 298 30129 354 30142
rect 298 30096 299 30129
rect 299 30096 354 30129
rect 396 30096 452 30152
rect 494 30142 506 30152
rect 506 30142 528 30152
rect 528 30142 550 30152
rect 592 30142 602 30152
rect 602 30142 648 30152
rect 494 30129 550 30142
rect 592 30129 648 30142
rect 494 30096 506 30129
rect 506 30096 528 30129
rect 528 30096 550 30129
rect 592 30096 602 30129
rect 602 30096 648 30129
rect 298 30064 354 30071
rect 298 30015 299 30064
rect 299 30015 354 30064
rect 396 30015 452 30071
rect 494 30064 550 30071
rect 592 30064 648 30071
rect 494 30015 506 30064
rect 506 30015 528 30064
rect 528 30015 550 30064
rect 592 30015 602 30064
rect 602 30015 648 30064
rect 298 29947 299 29990
rect 299 29947 354 29990
rect 298 29934 354 29947
rect 396 29934 452 29990
rect 494 29947 506 29990
rect 506 29947 528 29990
rect 528 29947 550 29990
rect 592 29947 602 29990
rect 602 29947 648 29990
rect 494 29934 550 29947
rect 592 29934 648 29947
rect 298 29882 299 29909
rect 299 29882 354 29909
rect 298 29869 354 29882
rect 298 29853 299 29869
rect 299 29853 354 29869
rect 396 29853 452 29909
rect 494 29882 506 29909
rect 506 29882 528 29909
rect 528 29882 550 29909
rect 592 29882 602 29909
rect 602 29882 648 29909
rect 494 29869 550 29882
rect 592 29869 648 29882
rect 494 29853 506 29869
rect 506 29853 528 29869
rect 528 29853 550 29869
rect 592 29853 602 29869
rect 602 29853 648 29869
rect 298 29817 299 29828
rect 299 29817 354 29828
rect 298 29804 354 29817
rect 298 29772 299 29804
rect 299 29772 354 29804
rect 396 29772 452 29828
rect 494 29817 506 29828
rect 506 29817 528 29828
rect 528 29817 550 29828
rect 592 29817 602 29828
rect 602 29817 648 29828
rect 494 29804 550 29817
rect 592 29804 648 29817
rect 494 29772 506 29804
rect 506 29772 528 29804
rect 528 29772 550 29804
rect 592 29772 602 29804
rect 602 29772 648 29804
rect 298 29739 354 29747
rect 298 29691 299 29739
rect 299 29691 354 29739
rect 396 29691 452 29747
rect 494 29739 550 29747
rect 592 29739 648 29747
rect 494 29691 506 29739
rect 506 29691 528 29739
rect 528 29691 550 29739
rect 592 29691 602 29739
rect 602 29691 648 29739
rect 298 29622 299 29666
rect 299 29622 354 29666
rect 298 29610 354 29622
rect 396 29610 452 29666
rect 494 29622 506 29666
rect 506 29622 528 29666
rect 528 29622 550 29666
rect 592 29622 602 29666
rect 602 29622 648 29666
rect 494 29610 550 29622
rect 592 29610 648 29622
rect 298 29557 299 29585
rect 299 29557 354 29585
rect 298 29544 354 29557
rect 298 29529 299 29544
rect 299 29529 354 29544
rect 396 29529 452 29585
rect 494 29557 506 29585
rect 506 29557 528 29585
rect 528 29557 550 29585
rect 592 29557 602 29585
rect 602 29557 648 29585
rect 494 29544 550 29557
rect 592 29544 648 29557
rect 494 29529 506 29544
rect 506 29529 528 29544
rect 528 29529 550 29544
rect 592 29529 602 29544
rect 602 29529 648 29544
rect 298 29492 299 29504
rect 299 29492 354 29504
rect 298 29479 354 29492
rect 298 29448 299 29479
rect 299 29448 354 29479
rect 396 29448 452 29504
rect 494 29492 506 29504
rect 506 29492 528 29504
rect 528 29492 550 29504
rect 592 29492 602 29504
rect 602 29492 648 29504
rect 494 29479 550 29492
rect 592 29479 648 29492
rect 494 29448 506 29479
rect 506 29448 528 29479
rect 528 29448 550 29479
rect 592 29448 602 29479
rect 602 29448 648 29479
rect 2139 31103 2195 31159
rect 2237 31103 2293 31159
rect 2335 31103 2391 31159
rect 2433 31103 2489 31159
rect 6182 31104 6238 31160
rect 6263 31104 6319 31160
rect 6344 31104 6400 31160
rect 6425 31104 6481 31160
rect 6506 31104 6562 31160
rect 6587 31104 6643 31160
rect 6668 31104 6724 31160
rect 6749 31104 6805 31160
rect 6830 31104 6886 31160
rect 6911 31104 6967 31160
rect 6992 31104 7048 31160
rect 7073 31104 7129 31160
rect 7154 31104 7210 31160
rect 7235 31104 7291 31160
rect 7316 31104 7372 31160
rect 7397 31104 7453 31160
rect 7478 31104 7534 31160
rect 7559 31104 7615 31160
rect 7640 31104 7696 31160
rect 7721 31104 7777 31160
rect 7802 31104 7858 31160
rect 7883 31104 7939 31160
rect 7964 31104 8020 31160
rect 8045 31104 8101 31160
rect 8126 31104 8182 31160
rect 8207 31104 8263 31160
rect 8288 31104 8344 31160
rect 8369 31104 8425 31160
rect 8450 31104 8506 31160
rect 8531 31104 8587 31160
rect 8612 31104 8668 31160
rect 8693 31104 8749 31160
rect 8774 31104 8830 31160
rect 8855 31104 8911 31160
rect 8936 31104 8992 31160
rect 9017 31104 9073 31160
rect 9098 31104 9154 31160
rect 9179 31104 9235 31160
rect 9260 31104 9316 31160
rect 9340 31104 9396 31160
rect 9420 31104 9476 31160
rect 9500 31104 9556 31160
rect 9580 31104 9636 31160
rect 9660 31104 9716 31160
rect 9740 31104 9796 31160
rect 9820 31104 9876 31160
rect 9900 31104 9956 31160
rect 9980 31104 10036 31160
rect 10060 31104 10116 31160
rect 10140 31104 10196 31160
rect 10220 31104 10276 31160
rect 10300 31104 10356 31160
rect 10380 31104 10436 31160
rect 10460 31104 10516 31160
rect 10540 31104 10596 31160
rect 10620 31104 10676 31160
rect 10700 31104 10756 31160
rect 10780 31104 10836 31160
rect 10860 31104 10916 31160
rect 10940 31104 10996 31160
rect 11020 31104 11076 31160
rect 11100 31104 11156 31160
rect 11180 31104 11236 31160
rect 11260 31104 11316 31160
rect 11340 31104 11396 31160
rect 11420 31104 11476 31160
rect 11500 31104 11556 31160
rect 11580 31104 11636 31160
rect 11660 31104 11716 31160
rect 11740 31104 11796 31160
rect 11820 31104 11876 31160
rect 11900 31104 11956 31160
rect 11980 31104 12036 31160
rect 12060 31104 12116 31160
rect 12140 31104 12196 31160
rect 12220 31104 12276 31160
rect 12300 31104 12356 31160
rect 12380 31104 12436 31160
rect 12460 31104 12516 31160
rect 12540 31104 12596 31160
rect 12620 31104 12676 31160
rect 12700 31104 12756 31160
rect 12780 31104 12836 31160
rect 12860 31104 12916 31160
rect 12940 31104 12996 31160
rect 13020 31104 13076 31160
rect 14514 31108 14570 31164
rect 14594 31108 14650 31164
rect 14674 31108 14730 31164
rect 14754 31108 14810 31164
rect 14834 31108 14890 31164
rect 14914 31108 14970 31164
rect 14994 31108 15050 31164
rect 15074 31108 15130 31164
rect 15154 31108 15210 31164
rect 15234 31108 15290 31164
rect 2139 31021 2195 31077
rect 2237 31021 2293 31077
rect 2335 31021 2391 31077
rect 2433 31021 2489 31077
rect 6182 31022 6238 31078
rect 6263 31022 6319 31078
rect 6344 31022 6400 31078
rect 6425 31022 6481 31078
rect 6506 31022 6562 31078
rect 6587 31022 6643 31078
rect 6668 31022 6724 31078
rect 6749 31022 6805 31078
rect 6830 31022 6886 31078
rect 6911 31022 6967 31078
rect 6992 31022 7048 31078
rect 7073 31022 7129 31078
rect 7154 31022 7210 31078
rect 7235 31022 7291 31078
rect 7316 31022 7372 31078
rect 7397 31022 7453 31078
rect 7478 31022 7534 31078
rect 7559 31022 7615 31078
rect 7640 31022 7696 31078
rect 7721 31022 7777 31078
rect 7802 31022 7858 31078
rect 7883 31022 7939 31078
rect 7964 31022 8020 31078
rect 8045 31022 8101 31078
rect 8126 31022 8182 31078
rect 8207 31022 8263 31078
rect 8288 31022 8344 31078
rect 8369 31022 8425 31078
rect 8450 31022 8506 31078
rect 8531 31022 8587 31078
rect 8612 31022 8668 31078
rect 8693 31022 8749 31078
rect 8774 31022 8830 31078
rect 8855 31022 8911 31078
rect 8936 31022 8992 31078
rect 9017 31022 9073 31078
rect 9098 31022 9154 31078
rect 9179 31022 9235 31078
rect 9260 31022 9316 31078
rect 9340 31022 9396 31078
rect 9420 31022 9476 31078
rect 9500 31022 9556 31078
rect 9580 31022 9636 31078
rect 9660 31022 9716 31078
rect 9740 31022 9796 31078
rect 9820 31022 9876 31078
rect 9900 31022 9956 31078
rect 9980 31022 10036 31078
rect 10060 31022 10116 31078
rect 10140 31022 10196 31078
rect 10220 31022 10276 31078
rect 10300 31022 10356 31078
rect 10380 31022 10436 31078
rect 10460 31022 10516 31078
rect 10540 31022 10596 31078
rect 10620 31022 10676 31078
rect 10700 31022 10756 31078
rect 10780 31022 10836 31078
rect 10860 31022 10916 31078
rect 10940 31022 10996 31078
rect 11020 31022 11076 31078
rect 11100 31022 11156 31078
rect 11180 31022 11236 31078
rect 11260 31022 11316 31078
rect 11340 31022 11396 31078
rect 11420 31022 11476 31078
rect 11500 31022 11556 31078
rect 11580 31022 11636 31078
rect 11660 31022 11716 31078
rect 11740 31022 11796 31078
rect 11820 31022 11876 31078
rect 11900 31022 11956 31078
rect 11980 31022 12036 31078
rect 12060 31022 12116 31078
rect 12140 31022 12196 31078
rect 12220 31022 12276 31078
rect 12300 31022 12356 31078
rect 12380 31022 12436 31078
rect 12460 31022 12516 31078
rect 12540 31022 12596 31078
rect 12620 31022 12676 31078
rect 12700 31022 12756 31078
rect 12780 31022 12836 31078
rect 12860 31022 12916 31078
rect 12940 31022 12996 31078
rect 13020 31022 13076 31078
rect 14514 31026 14570 31082
rect 14594 31026 14650 31082
rect 14674 31026 14730 31082
rect 14754 31026 14810 31082
rect 14834 31026 14890 31082
rect 14914 31026 14970 31082
rect 14994 31026 15050 31082
rect 15074 31026 15130 31082
rect 15154 31026 15210 31082
rect 15234 31026 15290 31082
rect 2139 30939 2195 30995
rect 2237 30939 2293 30995
rect 2335 30939 2391 30995
rect 2433 30939 2489 30995
rect 5803 30937 5859 30993
rect 5895 30937 5951 30993
rect 5987 30937 6043 30993
rect 6079 30937 6135 30993
rect 6182 30940 6238 30996
rect 6263 30940 6319 30996
rect 6344 30940 6400 30996
rect 6425 30940 6481 30996
rect 6506 30940 6562 30996
rect 6587 30940 6643 30996
rect 6668 30940 6724 30996
rect 6749 30940 6805 30996
rect 6830 30940 6886 30996
rect 6911 30940 6967 30996
rect 6992 30940 7048 30996
rect 7073 30940 7129 30996
rect 7154 30940 7210 30996
rect 7235 30940 7291 30996
rect 7316 30940 7372 30996
rect 7397 30940 7453 30996
rect 7478 30940 7534 30996
rect 7559 30940 7615 30996
rect 7640 30940 7696 30996
rect 7721 30940 7777 30996
rect 7802 30940 7858 30996
rect 7883 30940 7939 30996
rect 7964 30940 8020 30996
rect 8045 30940 8101 30996
rect 8126 30940 8182 30996
rect 8207 30940 8263 30996
rect 8288 30940 8344 30996
rect 8369 30940 8425 30996
rect 8450 30940 8506 30996
rect 8531 30940 8587 30996
rect 8612 30940 8668 30996
rect 8693 30940 8749 30996
rect 8774 30940 8830 30996
rect 8855 30940 8911 30996
rect 8936 30940 8992 30996
rect 9017 30940 9073 30996
rect 9098 30940 9154 30996
rect 9179 30940 9235 30996
rect 9260 30940 9316 30996
rect 9340 30940 9396 30996
rect 9420 30940 9476 30996
rect 9500 30940 9556 30996
rect 9580 30940 9636 30996
rect 9660 30940 9716 30996
rect 9740 30940 9796 30996
rect 9820 30940 9876 30996
rect 9900 30940 9956 30996
rect 9980 30940 10036 30996
rect 10060 30940 10116 30996
rect 10140 30940 10196 30996
rect 10220 30940 10276 30996
rect 10300 30940 10356 30996
rect 10380 30940 10436 30996
rect 10460 30940 10516 30996
rect 10540 30940 10596 30996
rect 10620 30940 10676 30996
rect 10700 30940 10756 30996
rect 10780 30940 10836 30996
rect 10860 30940 10916 30996
rect 10940 30940 10996 30996
rect 11020 30940 11076 30996
rect 11100 30940 11156 30996
rect 11180 30940 11236 30996
rect 11260 30940 11316 30996
rect 11340 30940 11396 30996
rect 11420 30940 11476 30996
rect 11500 30940 11556 30996
rect 11580 30940 11636 30996
rect 11660 30940 11716 30996
rect 11740 30940 11796 30996
rect 11820 30940 11876 30996
rect 11900 30940 11956 30996
rect 11980 30940 12036 30996
rect 12060 30940 12116 30996
rect 12140 30940 12196 30996
rect 12220 30940 12276 30996
rect 12300 30940 12356 30996
rect 12380 30940 12436 30996
rect 12460 30940 12516 30996
rect 12540 30940 12596 30996
rect 12620 30940 12676 30996
rect 12700 30940 12756 30996
rect 12780 30940 12836 30996
rect 12860 30940 12916 30996
rect 12940 30940 12996 30996
rect 13020 30940 13076 30996
rect 14514 30944 14570 31000
rect 14594 30944 14650 31000
rect 14674 30944 14730 31000
rect 14754 30944 14810 31000
rect 14834 30944 14890 31000
rect 14914 30944 14970 31000
rect 14994 30944 15050 31000
rect 15074 30944 15130 31000
rect 15154 30944 15210 31000
rect 15234 30944 15290 31000
rect 2139 30857 2195 30913
rect 2237 30857 2293 30913
rect 2335 30857 2391 30913
rect 2433 30857 2489 30913
rect 5803 30854 5859 30910
rect 5895 30854 5951 30910
rect 5987 30854 6043 30910
rect 6079 30854 6135 30910
rect 6182 30858 6238 30914
rect 6263 30858 6319 30914
rect 6344 30858 6400 30914
rect 6425 30858 6481 30914
rect 6506 30858 6562 30914
rect 6587 30858 6643 30914
rect 6668 30858 6724 30914
rect 6749 30858 6805 30914
rect 6830 30858 6886 30914
rect 6911 30858 6967 30914
rect 6992 30858 7048 30914
rect 7073 30858 7129 30914
rect 7154 30858 7210 30914
rect 7235 30858 7291 30914
rect 7316 30858 7372 30914
rect 7397 30858 7453 30914
rect 7478 30858 7534 30914
rect 7559 30858 7615 30914
rect 7640 30858 7696 30914
rect 7721 30858 7777 30914
rect 7802 30858 7858 30914
rect 7883 30858 7939 30914
rect 7964 30858 8020 30914
rect 8045 30858 8101 30914
rect 8126 30858 8182 30914
rect 8207 30858 8263 30914
rect 8288 30858 8344 30914
rect 8369 30858 8425 30914
rect 8450 30858 8506 30914
rect 8531 30858 8587 30914
rect 8612 30858 8668 30914
rect 8693 30858 8749 30914
rect 8774 30858 8830 30914
rect 8855 30858 8911 30914
rect 8936 30858 8992 30914
rect 9017 30858 9073 30914
rect 9098 30858 9154 30914
rect 9179 30858 9235 30914
rect 9260 30858 9316 30914
rect 9340 30858 9396 30914
rect 9420 30858 9476 30914
rect 9500 30858 9556 30914
rect 9580 30858 9636 30914
rect 9660 30858 9716 30914
rect 9740 30858 9796 30914
rect 9820 30858 9876 30914
rect 9900 30858 9956 30914
rect 9980 30858 10036 30914
rect 10060 30858 10116 30914
rect 10140 30858 10196 30914
rect 10220 30858 10276 30914
rect 10300 30858 10356 30914
rect 10380 30858 10436 30914
rect 10460 30858 10516 30914
rect 10540 30858 10596 30914
rect 10620 30858 10676 30914
rect 10700 30858 10756 30914
rect 10780 30858 10836 30914
rect 10860 30858 10916 30914
rect 10940 30858 10996 30914
rect 11020 30858 11076 30914
rect 11100 30858 11156 30914
rect 11180 30858 11236 30914
rect 11260 30858 11316 30914
rect 11340 30858 11396 30914
rect 11420 30858 11476 30914
rect 11500 30858 11556 30914
rect 11580 30858 11636 30914
rect 11660 30858 11716 30914
rect 11740 30858 11796 30914
rect 11820 30858 11876 30914
rect 11900 30858 11956 30914
rect 11980 30858 12036 30914
rect 12060 30858 12116 30914
rect 12140 30858 12196 30914
rect 12220 30858 12276 30914
rect 12300 30858 12356 30914
rect 12380 30858 12436 30914
rect 12460 30858 12516 30914
rect 12540 30858 12596 30914
rect 12620 30858 12676 30914
rect 12700 30858 12756 30914
rect 12780 30858 12836 30914
rect 12860 30858 12916 30914
rect 12940 30858 12996 30914
rect 13020 30858 13076 30914
rect 14514 30862 14570 30918
rect 14594 30862 14650 30918
rect 14674 30862 14730 30918
rect 14754 30862 14810 30918
rect 14834 30862 14890 30918
rect 14914 30862 14970 30918
rect 14994 30862 15050 30918
rect 15074 30862 15130 30918
rect 15154 30862 15210 30918
rect 15234 30862 15290 30918
rect 2139 30775 2195 30831
rect 2237 30775 2293 30831
rect 2335 30775 2391 30831
rect 2433 30775 2489 30831
rect 5803 30771 5859 30827
rect 5895 30771 5951 30827
rect 5987 30771 6043 30827
rect 6079 30771 6135 30827
rect 6182 30776 6238 30832
rect 6263 30776 6319 30832
rect 6344 30776 6400 30832
rect 6425 30776 6481 30832
rect 6506 30776 6562 30832
rect 6587 30776 6643 30832
rect 6668 30776 6724 30832
rect 6749 30776 6805 30832
rect 6830 30776 6886 30832
rect 6911 30776 6967 30832
rect 6992 30776 7048 30832
rect 7073 30776 7129 30832
rect 7154 30776 7210 30832
rect 7235 30776 7291 30832
rect 7316 30776 7372 30832
rect 7397 30776 7453 30832
rect 7478 30776 7534 30832
rect 7559 30776 7615 30832
rect 7640 30776 7696 30832
rect 7721 30776 7777 30832
rect 7802 30776 7858 30832
rect 7883 30776 7939 30832
rect 7964 30776 8020 30832
rect 8045 30776 8101 30832
rect 8126 30776 8182 30832
rect 8207 30776 8263 30832
rect 8288 30776 8344 30832
rect 8369 30776 8425 30832
rect 8450 30776 8506 30832
rect 8531 30776 8587 30832
rect 8612 30776 8668 30832
rect 8693 30776 8749 30832
rect 8774 30776 8830 30832
rect 8855 30776 8911 30832
rect 8936 30776 8992 30832
rect 9017 30776 9073 30832
rect 9098 30776 9154 30832
rect 9179 30776 9235 30832
rect 9260 30776 9316 30832
rect 9340 30776 9396 30832
rect 9420 30776 9476 30832
rect 9500 30776 9556 30832
rect 9580 30776 9636 30832
rect 9660 30776 9716 30832
rect 9740 30776 9796 30832
rect 9820 30776 9876 30832
rect 9900 30776 9956 30832
rect 9980 30776 10036 30832
rect 10060 30776 10116 30832
rect 10140 30776 10196 30832
rect 10220 30776 10276 30832
rect 10300 30776 10356 30832
rect 10380 30776 10436 30832
rect 10460 30776 10516 30832
rect 10540 30776 10596 30832
rect 10620 30776 10676 30832
rect 10700 30776 10756 30832
rect 10780 30776 10836 30832
rect 10860 30776 10916 30832
rect 10940 30776 10996 30832
rect 11020 30776 11076 30832
rect 11100 30776 11156 30832
rect 11180 30776 11236 30832
rect 11260 30776 11316 30832
rect 11340 30776 11396 30832
rect 11420 30776 11476 30832
rect 11500 30776 11556 30832
rect 11580 30776 11636 30832
rect 11660 30776 11716 30832
rect 11740 30776 11796 30832
rect 11820 30776 11876 30832
rect 11900 30776 11956 30832
rect 11980 30776 12036 30832
rect 12060 30776 12116 30832
rect 12140 30776 12196 30832
rect 12220 30776 12276 30832
rect 12300 30776 12356 30832
rect 12380 30776 12436 30832
rect 12460 30776 12516 30832
rect 12540 30776 12596 30832
rect 12620 30776 12676 30832
rect 12700 30776 12756 30832
rect 12780 30776 12836 30832
rect 12860 30776 12916 30832
rect 12940 30776 12996 30832
rect 13020 30776 13076 30832
rect 14514 30780 14570 30836
rect 14594 30780 14650 30836
rect 14674 30780 14730 30836
rect 14754 30780 14810 30836
rect 14834 30780 14890 30836
rect 14914 30780 14970 30836
rect 14994 30780 15050 30836
rect 15074 30780 15130 30836
rect 15154 30780 15210 30836
rect 15234 30780 15290 30836
rect 2139 30693 2195 30749
rect 2237 30693 2293 30749
rect 2335 30693 2391 30749
rect 2433 30693 2489 30749
rect 5803 30688 5859 30744
rect 5895 30688 5951 30744
rect 5987 30688 6043 30744
rect 6079 30688 6135 30744
rect 6182 30694 6238 30750
rect 6263 30694 6319 30750
rect 6344 30694 6400 30750
rect 6425 30694 6481 30750
rect 6506 30694 6562 30750
rect 6587 30694 6643 30750
rect 6668 30694 6724 30750
rect 6749 30694 6805 30750
rect 6830 30694 6886 30750
rect 6911 30694 6967 30750
rect 6992 30694 7048 30750
rect 7073 30694 7129 30750
rect 7154 30694 7210 30750
rect 7235 30694 7291 30750
rect 7316 30694 7372 30750
rect 7397 30694 7453 30750
rect 7478 30694 7534 30750
rect 7559 30694 7615 30750
rect 7640 30694 7696 30750
rect 7721 30694 7777 30750
rect 7802 30694 7858 30750
rect 7883 30694 7939 30750
rect 7964 30694 8020 30750
rect 8045 30694 8101 30750
rect 8126 30694 8182 30750
rect 8207 30694 8263 30750
rect 8288 30694 8344 30750
rect 8369 30694 8425 30750
rect 8450 30694 8506 30750
rect 8531 30694 8587 30750
rect 8612 30694 8668 30750
rect 8693 30694 8749 30750
rect 8774 30694 8830 30750
rect 8855 30694 8911 30750
rect 8936 30694 8992 30750
rect 9017 30694 9073 30750
rect 9098 30694 9154 30750
rect 9179 30694 9235 30750
rect 9260 30694 9316 30750
rect 9340 30694 9396 30750
rect 9420 30694 9476 30750
rect 9500 30694 9556 30750
rect 9580 30694 9636 30750
rect 9660 30694 9716 30750
rect 9740 30694 9796 30750
rect 9820 30694 9876 30750
rect 9900 30694 9956 30750
rect 9980 30694 10036 30750
rect 10060 30694 10116 30750
rect 10140 30694 10196 30750
rect 10220 30694 10276 30750
rect 10300 30694 10356 30750
rect 10380 30694 10436 30750
rect 10460 30694 10516 30750
rect 10540 30694 10596 30750
rect 10620 30694 10676 30750
rect 10700 30694 10756 30750
rect 10780 30694 10836 30750
rect 10860 30694 10916 30750
rect 10940 30694 10996 30750
rect 11020 30694 11076 30750
rect 11100 30694 11156 30750
rect 11180 30694 11236 30750
rect 11260 30694 11316 30750
rect 11340 30694 11396 30750
rect 11420 30694 11476 30750
rect 11500 30694 11556 30750
rect 11580 30694 11636 30750
rect 11660 30694 11716 30750
rect 11740 30694 11796 30750
rect 11820 30694 11876 30750
rect 11900 30694 11956 30750
rect 11980 30694 12036 30750
rect 12060 30694 12116 30750
rect 12140 30694 12196 30750
rect 12220 30694 12276 30750
rect 12300 30694 12356 30750
rect 12380 30694 12436 30750
rect 12460 30694 12516 30750
rect 12540 30694 12596 30750
rect 12620 30694 12676 30750
rect 12700 30694 12756 30750
rect 12780 30694 12836 30750
rect 12860 30694 12916 30750
rect 12940 30694 12996 30750
rect 13020 30694 13076 30750
rect 14514 30697 14570 30753
rect 14594 30697 14650 30753
rect 14674 30697 14730 30753
rect 14754 30697 14810 30753
rect 14834 30697 14890 30753
rect 14914 30697 14970 30753
rect 14994 30697 15050 30753
rect 15074 30697 15130 30753
rect 15154 30697 15210 30753
rect 15234 30697 15290 30753
rect 2139 30611 2195 30667
rect 2237 30611 2293 30667
rect 2335 30611 2391 30667
rect 2433 30611 2489 30667
rect 5803 30605 5859 30661
rect 5895 30605 5951 30661
rect 5987 30605 6043 30661
rect 6079 30605 6135 30661
rect 6182 30612 6238 30668
rect 6263 30612 6319 30668
rect 6344 30612 6400 30668
rect 6425 30612 6481 30668
rect 6506 30612 6562 30668
rect 6587 30612 6643 30668
rect 6668 30612 6724 30668
rect 6749 30612 6805 30668
rect 6830 30612 6886 30668
rect 6911 30612 6967 30668
rect 6992 30612 7048 30668
rect 7073 30612 7129 30668
rect 7154 30612 7210 30668
rect 7235 30612 7291 30668
rect 7316 30612 7372 30668
rect 7397 30612 7453 30668
rect 7478 30612 7534 30668
rect 7559 30612 7615 30668
rect 7640 30612 7696 30668
rect 7721 30612 7777 30668
rect 7802 30612 7858 30668
rect 7883 30612 7939 30668
rect 7964 30612 8020 30668
rect 8045 30612 8101 30668
rect 8126 30612 8182 30668
rect 8207 30612 8263 30668
rect 8288 30612 8344 30668
rect 8369 30612 8425 30668
rect 8450 30612 8506 30668
rect 8531 30612 8587 30668
rect 8612 30612 8668 30668
rect 8693 30612 8749 30668
rect 8774 30612 8830 30668
rect 8855 30612 8911 30668
rect 8936 30612 8992 30668
rect 9017 30612 9073 30668
rect 9098 30612 9154 30668
rect 9179 30612 9235 30668
rect 9260 30612 9316 30668
rect 9340 30612 9396 30668
rect 9420 30612 9476 30668
rect 9500 30612 9556 30668
rect 9580 30612 9636 30668
rect 9660 30612 9716 30668
rect 9740 30612 9796 30668
rect 9820 30612 9876 30668
rect 9900 30612 9956 30668
rect 9980 30612 10036 30668
rect 10060 30612 10116 30668
rect 10140 30612 10196 30668
rect 10220 30612 10276 30668
rect 10300 30612 10356 30668
rect 10380 30612 10436 30668
rect 10460 30612 10516 30668
rect 10540 30612 10596 30668
rect 10620 30612 10676 30668
rect 10700 30612 10756 30668
rect 10780 30612 10836 30668
rect 10860 30612 10916 30668
rect 10940 30612 10996 30668
rect 11020 30612 11076 30668
rect 11100 30612 11156 30668
rect 11180 30612 11236 30668
rect 11260 30612 11316 30668
rect 11340 30612 11396 30668
rect 11420 30612 11476 30668
rect 11500 30612 11556 30668
rect 11580 30612 11636 30668
rect 11660 30612 11716 30668
rect 11740 30612 11796 30668
rect 11820 30612 11876 30668
rect 11900 30612 11956 30668
rect 11980 30612 12036 30668
rect 12060 30612 12116 30668
rect 12140 30612 12196 30668
rect 12220 30612 12276 30668
rect 12300 30612 12356 30668
rect 12380 30612 12436 30668
rect 12460 30612 12516 30668
rect 12540 30612 12596 30668
rect 12620 30612 12676 30668
rect 12700 30612 12756 30668
rect 12780 30612 12836 30668
rect 12860 30612 12916 30668
rect 12940 30612 12996 30668
rect 13020 30612 13076 30668
rect 14514 30614 14570 30670
rect 14594 30614 14650 30670
rect 14674 30614 14730 30670
rect 14754 30614 14810 30670
rect 14834 30614 14890 30670
rect 14914 30614 14970 30670
rect 14994 30614 15050 30670
rect 15074 30614 15130 30670
rect 15154 30614 15210 30670
rect 15234 30614 15290 30670
rect 2139 30529 2195 30585
rect 2237 30529 2293 30585
rect 2335 30529 2391 30585
rect 2433 30529 2489 30585
rect 5803 30522 5859 30578
rect 5895 30522 5951 30578
rect 5987 30522 6043 30578
rect 6079 30522 6135 30578
rect 6182 30530 6238 30586
rect 6263 30530 6319 30586
rect 6344 30530 6400 30586
rect 6425 30530 6481 30586
rect 6506 30530 6562 30586
rect 6587 30530 6643 30586
rect 6668 30530 6724 30586
rect 6749 30530 6805 30586
rect 6830 30530 6886 30586
rect 6911 30530 6967 30586
rect 6992 30530 7048 30586
rect 7073 30530 7129 30586
rect 7154 30530 7210 30586
rect 7235 30530 7291 30586
rect 7316 30530 7372 30586
rect 7397 30530 7453 30586
rect 7478 30530 7534 30586
rect 7559 30530 7615 30586
rect 7640 30530 7696 30586
rect 7721 30530 7777 30586
rect 7802 30530 7858 30586
rect 7883 30530 7939 30586
rect 7964 30530 8020 30586
rect 8045 30530 8101 30586
rect 8126 30530 8182 30586
rect 8207 30530 8263 30586
rect 8288 30530 8344 30586
rect 8369 30530 8425 30586
rect 8450 30530 8506 30586
rect 8531 30530 8587 30586
rect 8612 30530 8668 30586
rect 8693 30530 8749 30586
rect 8774 30530 8830 30586
rect 8855 30530 8911 30586
rect 8936 30530 8992 30586
rect 9017 30530 9073 30586
rect 9098 30530 9154 30586
rect 9179 30530 9235 30586
rect 9260 30530 9316 30586
rect 9340 30530 9396 30586
rect 9420 30530 9476 30586
rect 9500 30530 9556 30586
rect 9580 30530 9636 30586
rect 9660 30530 9716 30586
rect 9740 30530 9796 30586
rect 9820 30530 9876 30586
rect 9900 30530 9956 30586
rect 9980 30530 10036 30586
rect 10060 30530 10116 30586
rect 10140 30530 10196 30586
rect 10220 30530 10276 30586
rect 10300 30530 10356 30586
rect 10380 30530 10436 30586
rect 10460 30530 10516 30586
rect 10540 30530 10596 30586
rect 10620 30530 10676 30586
rect 10700 30530 10756 30586
rect 10780 30530 10836 30586
rect 10860 30530 10916 30586
rect 10940 30530 10996 30586
rect 11020 30530 11076 30586
rect 11100 30530 11156 30586
rect 11180 30530 11236 30586
rect 11260 30530 11316 30586
rect 11340 30530 11396 30586
rect 11420 30530 11476 30586
rect 11500 30530 11556 30586
rect 11580 30530 11636 30586
rect 11660 30530 11716 30586
rect 11740 30530 11796 30586
rect 11820 30530 11876 30586
rect 11900 30530 11956 30586
rect 11980 30530 12036 30586
rect 12060 30530 12116 30586
rect 12140 30530 12196 30586
rect 12220 30530 12276 30586
rect 12300 30530 12356 30586
rect 12380 30530 12436 30586
rect 12460 30530 12516 30586
rect 12540 30530 12596 30586
rect 12620 30530 12676 30586
rect 12700 30530 12756 30586
rect 12780 30530 12836 30586
rect 12860 30530 12916 30586
rect 12940 30530 12996 30586
rect 13020 30530 13076 30586
rect 14514 30531 14570 30587
rect 14594 30531 14650 30587
rect 14674 30531 14730 30587
rect 14754 30531 14810 30587
rect 14834 30531 14890 30587
rect 14914 30531 14970 30587
rect 14994 30531 15050 30587
rect 15074 30531 15130 30587
rect 15154 30531 15210 30587
rect 15234 30531 15290 30587
rect 2139 30447 2195 30503
rect 2237 30447 2293 30503
rect 2335 30447 2391 30503
rect 2433 30447 2489 30503
rect 5803 30440 5859 30496
rect 5895 30440 5951 30496
rect 5987 30440 6043 30496
rect 6079 30440 6135 30496
rect 6182 30448 6238 30504
rect 6263 30448 6319 30504
rect 6344 30448 6400 30504
rect 6425 30448 6481 30504
rect 6506 30448 6562 30504
rect 6587 30448 6643 30504
rect 6668 30448 6724 30504
rect 6749 30448 6805 30504
rect 6830 30448 6886 30504
rect 6911 30448 6967 30504
rect 6992 30448 7048 30504
rect 7073 30448 7129 30504
rect 7154 30448 7210 30504
rect 7235 30448 7291 30504
rect 7316 30448 7372 30504
rect 7397 30448 7453 30504
rect 7478 30448 7534 30504
rect 7559 30448 7615 30504
rect 7640 30448 7696 30504
rect 7721 30448 7777 30504
rect 7802 30448 7858 30504
rect 7883 30448 7939 30504
rect 7964 30448 8020 30504
rect 8045 30448 8101 30504
rect 8126 30448 8182 30504
rect 8207 30448 8263 30504
rect 8288 30448 8344 30504
rect 8369 30448 8425 30504
rect 8450 30448 8506 30504
rect 8531 30448 8587 30504
rect 8612 30448 8668 30504
rect 8693 30448 8749 30504
rect 8774 30448 8830 30504
rect 8855 30448 8911 30504
rect 8936 30448 8992 30504
rect 9017 30448 9073 30504
rect 9098 30448 9154 30504
rect 9179 30448 9235 30504
rect 9260 30448 9316 30504
rect 9340 30448 9396 30504
rect 9420 30448 9476 30504
rect 9500 30448 9556 30504
rect 9580 30448 9636 30504
rect 9660 30448 9716 30504
rect 9740 30448 9796 30504
rect 9820 30448 9876 30504
rect 9900 30448 9956 30504
rect 9980 30448 10036 30504
rect 10060 30448 10116 30504
rect 10140 30448 10196 30504
rect 10220 30448 10276 30504
rect 10300 30448 10356 30504
rect 10380 30448 10436 30504
rect 10460 30448 10516 30504
rect 10540 30448 10596 30504
rect 10620 30448 10676 30504
rect 10700 30448 10756 30504
rect 10780 30448 10836 30504
rect 10860 30448 10916 30504
rect 10940 30448 10996 30504
rect 11020 30448 11076 30504
rect 11100 30448 11156 30504
rect 11180 30448 11236 30504
rect 11260 30448 11316 30504
rect 11340 30448 11396 30504
rect 11420 30448 11476 30504
rect 11500 30448 11556 30504
rect 11580 30448 11636 30504
rect 11660 30448 11716 30504
rect 11740 30448 11796 30504
rect 11820 30448 11876 30504
rect 11900 30448 11956 30504
rect 11980 30448 12036 30504
rect 12060 30448 12116 30504
rect 12140 30448 12196 30504
rect 12220 30448 12276 30504
rect 12300 30448 12356 30504
rect 12380 30448 12436 30504
rect 12460 30448 12516 30504
rect 12540 30448 12596 30504
rect 12620 30448 12676 30504
rect 12700 30448 12756 30504
rect 12780 30448 12836 30504
rect 12860 30448 12916 30504
rect 12940 30448 12996 30504
rect 13020 30448 13076 30504
rect 14514 30448 14570 30504
rect 14594 30448 14650 30504
rect 14674 30448 14730 30504
rect 14754 30448 14810 30504
rect 14834 30448 14890 30504
rect 14914 30448 14970 30504
rect 14994 30448 15050 30504
rect 15074 30448 15130 30504
rect 15154 30448 15210 30504
rect 15234 30448 15290 30504
rect 2139 30365 2195 30421
rect 2237 30365 2293 30421
rect 2335 30365 2391 30421
rect 2433 30365 2489 30421
rect 5803 30358 5859 30414
rect 5895 30358 5951 30414
rect 5987 30358 6043 30414
rect 6079 30358 6135 30414
rect 6182 30366 6238 30422
rect 6263 30366 6319 30422
rect 6344 30366 6400 30422
rect 6425 30366 6481 30422
rect 6506 30366 6562 30422
rect 6587 30366 6643 30422
rect 6668 30366 6724 30422
rect 6749 30366 6805 30422
rect 6830 30366 6886 30422
rect 6911 30366 6967 30422
rect 6992 30366 7048 30422
rect 7073 30366 7129 30422
rect 7154 30366 7210 30422
rect 7235 30366 7291 30422
rect 7316 30366 7372 30422
rect 7397 30366 7453 30422
rect 7478 30366 7534 30422
rect 7559 30366 7615 30422
rect 7640 30366 7696 30422
rect 7721 30366 7777 30422
rect 7802 30366 7858 30422
rect 7883 30366 7939 30422
rect 7964 30366 8020 30422
rect 8045 30366 8101 30422
rect 8126 30366 8182 30422
rect 8207 30366 8263 30422
rect 8288 30366 8344 30422
rect 8369 30366 8425 30422
rect 8450 30366 8506 30422
rect 8531 30366 8587 30422
rect 8612 30366 8668 30422
rect 8693 30366 8749 30422
rect 8774 30366 8830 30422
rect 8855 30366 8911 30422
rect 8936 30366 8992 30422
rect 9017 30366 9073 30422
rect 9098 30366 9154 30422
rect 9179 30366 9235 30422
rect 9260 30366 9316 30422
rect 9340 30366 9396 30422
rect 9420 30366 9476 30422
rect 9500 30366 9556 30422
rect 9580 30366 9636 30422
rect 9660 30366 9716 30422
rect 9740 30366 9796 30422
rect 9820 30366 9876 30422
rect 9900 30366 9956 30422
rect 9980 30366 10036 30422
rect 10060 30366 10116 30422
rect 10140 30366 10196 30422
rect 10220 30366 10276 30422
rect 10300 30366 10356 30422
rect 10380 30366 10436 30422
rect 10460 30366 10516 30422
rect 10540 30366 10596 30422
rect 10620 30366 10676 30422
rect 10700 30366 10756 30422
rect 10780 30366 10836 30422
rect 10860 30366 10916 30422
rect 10940 30366 10996 30422
rect 11020 30366 11076 30422
rect 11100 30366 11156 30422
rect 11180 30366 11236 30422
rect 11260 30366 11316 30422
rect 11340 30366 11396 30422
rect 11420 30366 11476 30422
rect 11500 30366 11556 30422
rect 11580 30366 11636 30422
rect 11660 30366 11716 30422
rect 11740 30366 11796 30422
rect 11820 30366 11876 30422
rect 11900 30366 11956 30422
rect 11980 30366 12036 30422
rect 12060 30366 12116 30422
rect 12140 30366 12196 30422
rect 12220 30366 12276 30422
rect 12300 30366 12356 30422
rect 12380 30366 12436 30422
rect 12460 30366 12516 30422
rect 12540 30366 12596 30422
rect 12620 30366 12676 30422
rect 12700 30366 12756 30422
rect 12780 30366 12836 30422
rect 12860 30366 12916 30422
rect 12940 30366 12996 30422
rect 13020 30366 13076 30422
rect 14514 30365 14570 30421
rect 14594 30365 14650 30421
rect 14674 30365 14730 30421
rect 14754 30365 14810 30421
rect 14834 30365 14890 30421
rect 14914 30365 14970 30421
rect 14994 30365 15050 30421
rect 15074 30365 15130 30421
rect 15154 30365 15210 30421
rect 15234 30365 15290 30421
rect 2139 30282 2195 30338
rect 2237 30282 2293 30338
rect 2335 30282 2391 30338
rect 2433 30282 2489 30338
rect 5803 30276 5859 30332
rect 5895 30276 5951 30332
rect 5987 30276 6043 30332
rect 6079 30276 6135 30332
rect 6182 30284 6238 30340
rect 6263 30284 6319 30340
rect 6344 30284 6400 30340
rect 6425 30284 6481 30340
rect 6506 30284 6562 30340
rect 6587 30284 6643 30340
rect 6668 30284 6724 30340
rect 6749 30284 6805 30340
rect 6830 30284 6886 30340
rect 6911 30284 6967 30340
rect 6992 30284 7048 30340
rect 7073 30284 7129 30340
rect 7154 30284 7210 30340
rect 7235 30284 7291 30340
rect 7316 30284 7372 30340
rect 7397 30284 7453 30340
rect 7478 30284 7534 30340
rect 7559 30284 7615 30340
rect 7640 30284 7696 30340
rect 7721 30284 7777 30340
rect 7802 30284 7858 30340
rect 7883 30284 7939 30340
rect 7964 30284 8020 30340
rect 8045 30284 8101 30340
rect 8126 30284 8182 30340
rect 8207 30284 8263 30340
rect 8288 30284 8344 30340
rect 8369 30284 8425 30340
rect 8450 30284 8506 30340
rect 8531 30284 8587 30340
rect 8612 30284 8668 30340
rect 8693 30284 8749 30340
rect 8774 30284 8830 30340
rect 8855 30284 8911 30340
rect 8936 30284 8992 30340
rect 9017 30284 9073 30340
rect 9098 30284 9154 30340
rect 9179 30284 9235 30340
rect 9260 30284 9316 30340
rect 9340 30284 9396 30340
rect 9420 30284 9476 30340
rect 9500 30284 9556 30340
rect 9580 30284 9636 30340
rect 9660 30284 9716 30340
rect 9740 30284 9796 30340
rect 9820 30284 9876 30340
rect 9900 30284 9956 30340
rect 9980 30284 10036 30340
rect 10060 30284 10116 30340
rect 10140 30284 10196 30340
rect 10220 30284 10276 30340
rect 10300 30284 10356 30340
rect 10380 30284 10436 30340
rect 10460 30284 10516 30340
rect 10540 30284 10596 30340
rect 10620 30284 10676 30340
rect 10700 30284 10756 30340
rect 10780 30284 10836 30340
rect 10860 30284 10916 30340
rect 10940 30284 10996 30340
rect 11020 30284 11076 30340
rect 11100 30284 11156 30340
rect 11180 30284 11236 30340
rect 11260 30284 11316 30340
rect 11340 30284 11396 30340
rect 11420 30284 11476 30340
rect 11500 30284 11556 30340
rect 11580 30284 11636 30340
rect 11660 30284 11716 30340
rect 11740 30284 11796 30340
rect 11820 30284 11876 30340
rect 11900 30284 11956 30340
rect 11980 30284 12036 30340
rect 12060 30284 12116 30340
rect 12140 30284 12196 30340
rect 12220 30284 12276 30340
rect 12300 30284 12356 30340
rect 12380 30284 12436 30340
rect 12460 30284 12516 30340
rect 12540 30284 12596 30340
rect 12620 30284 12676 30340
rect 12700 30284 12756 30340
rect 12780 30284 12836 30340
rect 12860 30284 12916 30340
rect 12940 30284 12996 30340
rect 13020 30284 13076 30340
rect 14514 30282 14570 30338
rect 14594 30282 14650 30338
rect 14674 30282 14730 30338
rect 14754 30282 14810 30338
rect 14834 30282 14890 30338
rect 14914 30282 14970 30338
rect 14994 30282 15050 30338
rect 15074 30282 15130 30338
rect 15154 30282 15210 30338
rect 15234 30282 15290 30338
rect 2139 30199 2195 30255
rect 2237 30199 2293 30255
rect 2335 30199 2391 30255
rect 2433 30199 2489 30255
rect 5803 30194 5859 30250
rect 5895 30194 5951 30250
rect 5987 30194 6043 30250
rect 6079 30194 6135 30250
rect 6182 30202 6238 30258
rect 6263 30202 6319 30258
rect 6344 30202 6400 30258
rect 6425 30202 6481 30258
rect 6506 30202 6562 30258
rect 6587 30202 6643 30258
rect 6668 30202 6724 30258
rect 6749 30202 6805 30258
rect 6830 30202 6886 30258
rect 6911 30202 6967 30258
rect 6992 30202 7048 30258
rect 7073 30202 7129 30258
rect 7154 30202 7210 30258
rect 7235 30202 7291 30258
rect 7316 30202 7372 30258
rect 7397 30202 7453 30258
rect 7478 30202 7534 30258
rect 7559 30202 7615 30258
rect 7640 30202 7696 30258
rect 7721 30202 7777 30258
rect 7802 30202 7858 30258
rect 7883 30202 7939 30258
rect 7964 30202 8020 30258
rect 8045 30202 8101 30258
rect 8126 30202 8182 30258
rect 8207 30202 8263 30258
rect 8288 30202 8344 30258
rect 8369 30202 8425 30258
rect 8450 30202 8506 30258
rect 8531 30202 8587 30258
rect 8612 30202 8668 30258
rect 8693 30202 8749 30258
rect 8774 30202 8830 30258
rect 8855 30202 8911 30258
rect 8936 30202 8992 30258
rect 9017 30202 9073 30258
rect 9098 30202 9154 30258
rect 9179 30202 9235 30258
rect 9260 30202 9316 30258
rect 9340 30202 9396 30258
rect 9420 30202 9476 30258
rect 9500 30202 9556 30258
rect 9580 30202 9636 30258
rect 9660 30202 9716 30258
rect 9740 30202 9796 30258
rect 9820 30202 9876 30258
rect 9900 30202 9956 30258
rect 9980 30202 10036 30258
rect 10060 30202 10116 30258
rect 10140 30202 10196 30258
rect 10220 30202 10276 30258
rect 10300 30202 10356 30258
rect 10380 30202 10436 30258
rect 10460 30202 10516 30258
rect 10540 30202 10596 30258
rect 10620 30202 10676 30258
rect 10700 30202 10756 30258
rect 10780 30202 10836 30258
rect 10860 30202 10916 30258
rect 10940 30202 10996 30258
rect 11020 30202 11076 30258
rect 11100 30202 11156 30258
rect 11180 30202 11236 30258
rect 11260 30202 11316 30258
rect 11340 30202 11396 30258
rect 11420 30202 11476 30258
rect 11500 30202 11556 30258
rect 11580 30202 11636 30258
rect 11660 30202 11716 30258
rect 11740 30202 11796 30258
rect 11820 30202 11876 30258
rect 11900 30202 11956 30258
rect 11980 30202 12036 30258
rect 12060 30202 12116 30258
rect 12140 30202 12196 30258
rect 12220 30202 12276 30258
rect 12300 30202 12356 30258
rect 12380 30202 12436 30258
rect 12460 30202 12516 30258
rect 12540 30202 12596 30258
rect 12620 30202 12676 30258
rect 12700 30202 12756 30258
rect 12780 30202 12836 30258
rect 12860 30202 12916 30258
rect 12940 30202 12996 30258
rect 13020 30202 13076 30258
rect 14514 30199 14570 30255
rect 14594 30199 14650 30255
rect 14674 30199 14730 30255
rect 14754 30199 14810 30255
rect 14834 30199 14890 30255
rect 14914 30199 14970 30255
rect 14994 30199 15050 30255
rect 15074 30199 15130 30255
rect 15154 30199 15210 30255
rect 15234 30199 15290 30255
rect 2139 30116 2195 30172
rect 2237 30116 2293 30172
rect 2335 30116 2391 30172
rect 2433 30116 2489 30172
rect 14514 30116 14570 30172
rect 14594 30116 14650 30172
rect 14674 30116 14730 30172
rect 14754 30116 14810 30172
rect 14834 30116 14890 30172
rect 14914 30116 14970 30172
rect 14994 30116 15050 30172
rect 15074 30116 15130 30172
rect 15154 30116 15210 30172
rect 15234 30116 15290 30172
rect 2139 30033 2195 30089
rect 2237 30033 2293 30089
rect 2335 30033 2391 30089
rect 2433 30033 2489 30089
rect 14514 30033 14570 30089
rect 14594 30033 14650 30089
rect 14674 30033 14730 30089
rect 14754 30033 14810 30089
rect 14834 30033 14890 30089
rect 14914 30033 14970 30089
rect 14994 30033 15050 30089
rect 15074 30033 15130 30089
rect 15154 30033 15210 30089
rect 15234 30033 15290 30089
rect 2139 29950 2195 30006
rect 2237 29950 2293 30006
rect 2335 29950 2391 30006
rect 2433 29950 2489 30006
rect 14514 29950 14570 30006
rect 14594 29950 14650 30006
rect 14674 29950 14730 30006
rect 14754 29950 14810 30006
rect 14834 29950 14890 30006
rect 14914 29950 14970 30006
rect 14994 29950 15050 30006
rect 15074 29950 15130 30006
rect 15154 29950 15210 30006
rect 15234 29950 15290 30006
rect 2139 29867 2195 29923
rect 2237 29867 2293 29923
rect 2335 29867 2391 29923
rect 2433 29867 2489 29923
rect 2139 29784 2195 29840
rect 2237 29784 2293 29840
rect 2335 29784 2391 29840
rect 2433 29784 2489 29840
rect 5803 29827 5859 29883
rect 5895 29827 5951 29883
rect 5987 29827 6043 29883
rect 6079 29827 6135 29883
rect 6182 29824 6238 29880
rect 6263 29824 6319 29880
rect 6344 29824 6400 29880
rect 6425 29824 6481 29880
rect 6506 29824 6562 29880
rect 6587 29824 6643 29880
rect 6668 29824 6724 29880
rect 6749 29824 6805 29880
rect 6830 29824 6886 29880
rect 6911 29824 6967 29880
rect 6992 29824 7048 29880
rect 7073 29824 7129 29880
rect 7154 29824 7210 29880
rect 7235 29824 7291 29880
rect 7316 29824 7372 29880
rect 7397 29824 7453 29880
rect 7478 29824 7534 29880
rect 7559 29824 7615 29880
rect 7640 29824 7696 29880
rect 7721 29824 7777 29880
rect 7802 29824 7858 29880
rect 7883 29824 7939 29880
rect 7964 29824 8020 29880
rect 8045 29824 8101 29880
rect 8126 29824 8182 29880
rect 8207 29824 8263 29880
rect 8288 29824 8344 29880
rect 8369 29824 8425 29880
rect 8450 29824 8506 29880
rect 8531 29824 8587 29880
rect 8612 29824 8668 29880
rect 8693 29824 8749 29880
rect 8774 29824 8830 29880
rect 8855 29824 8911 29880
rect 8936 29824 8992 29880
rect 9017 29824 9073 29880
rect 9098 29824 9154 29880
rect 9179 29824 9235 29880
rect 2139 29701 2195 29757
rect 2237 29701 2293 29757
rect 2335 29701 2391 29757
rect 2433 29701 2489 29757
rect 5803 29745 5859 29801
rect 5895 29745 5951 29801
rect 5987 29745 6043 29801
rect 6079 29745 6135 29801
rect 6182 29744 6238 29800
rect 6263 29744 6319 29800
rect 6344 29744 6400 29800
rect 6425 29744 6481 29800
rect 6506 29744 6562 29800
rect 6587 29744 6643 29800
rect 6668 29744 6724 29800
rect 6749 29744 6805 29800
rect 6830 29744 6886 29800
rect 6911 29744 6967 29800
rect 6992 29744 7048 29800
rect 7073 29744 7129 29800
rect 7154 29744 7210 29800
rect 7235 29744 7291 29800
rect 7316 29744 7372 29800
rect 7397 29744 7453 29800
rect 7478 29744 7534 29800
rect 7559 29744 7615 29800
rect 7640 29744 7696 29800
rect 7721 29744 7777 29800
rect 7802 29744 7858 29800
rect 7883 29744 7939 29800
rect 7964 29744 8020 29800
rect 8045 29744 8101 29800
rect 8126 29744 8182 29800
rect 8207 29744 8263 29800
rect 8288 29744 8344 29800
rect 8369 29744 8425 29800
rect 8450 29744 8506 29800
rect 8531 29744 8587 29800
rect 8612 29744 8668 29800
rect 8693 29744 8749 29800
rect 8774 29744 8830 29800
rect 8855 29744 8911 29800
rect 8936 29744 8992 29800
rect 9017 29744 9073 29800
rect 9098 29744 9154 29800
rect 9179 29744 9235 29800
rect 2139 29618 2195 29674
rect 2237 29618 2293 29674
rect 2335 29618 2391 29674
rect 2433 29618 2489 29674
rect 5803 29663 5859 29719
rect 5895 29663 5951 29719
rect 5987 29663 6043 29719
rect 6079 29663 6135 29719
rect 6182 29664 6238 29720
rect 6263 29664 6319 29720
rect 6344 29664 6400 29720
rect 6425 29664 6481 29720
rect 6506 29664 6562 29720
rect 6587 29664 6643 29720
rect 6668 29664 6724 29720
rect 6749 29664 6805 29720
rect 6830 29664 6886 29720
rect 6911 29664 6967 29720
rect 6992 29664 7048 29720
rect 7073 29664 7129 29720
rect 7154 29664 7210 29720
rect 7235 29664 7291 29720
rect 7316 29664 7372 29720
rect 7397 29664 7453 29720
rect 7478 29664 7534 29720
rect 7559 29664 7615 29720
rect 7640 29664 7696 29720
rect 7721 29664 7777 29720
rect 7802 29664 7858 29720
rect 7883 29664 7939 29720
rect 7964 29664 8020 29720
rect 8045 29664 8101 29720
rect 8126 29664 8182 29720
rect 8207 29664 8263 29720
rect 8288 29664 8344 29720
rect 8369 29664 8425 29720
rect 8450 29664 8506 29720
rect 8531 29664 8587 29720
rect 8612 29664 8668 29720
rect 8693 29664 8749 29720
rect 8774 29664 8830 29720
rect 8855 29664 8911 29720
rect 8936 29664 8992 29720
rect 9017 29664 9073 29720
rect 9098 29664 9154 29720
rect 9179 29664 9235 29720
rect 2139 29535 2195 29591
rect 2237 29535 2293 29591
rect 2335 29535 2391 29591
rect 2433 29535 2489 29591
rect 5803 29581 5859 29637
rect 5895 29581 5951 29637
rect 5987 29581 6043 29637
rect 6079 29581 6135 29637
rect 6182 29584 6238 29640
rect 6263 29584 6319 29640
rect 6344 29584 6400 29640
rect 6425 29584 6481 29640
rect 6506 29584 6562 29640
rect 6587 29584 6643 29640
rect 6668 29584 6724 29640
rect 6749 29584 6805 29640
rect 6830 29584 6886 29640
rect 6911 29584 6967 29640
rect 6992 29584 7048 29640
rect 7073 29584 7129 29640
rect 7154 29584 7210 29640
rect 7235 29584 7291 29640
rect 7316 29584 7372 29640
rect 7397 29584 7453 29640
rect 7478 29584 7534 29640
rect 7559 29584 7615 29640
rect 7640 29584 7696 29640
rect 7721 29584 7777 29640
rect 7802 29584 7858 29640
rect 7883 29584 7939 29640
rect 7964 29584 8020 29640
rect 8045 29584 8101 29640
rect 8126 29584 8182 29640
rect 8207 29584 8263 29640
rect 8288 29584 8344 29640
rect 8369 29584 8425 29640
rect 8450 29584 8506 29640
rect 8531 29584 8587 29640
rect 8612 29584 8668 29640
rect 8693 29584 8749 29640
rect 8774 29584 8830 29640
rect 8855 29584 8911 29640
rect 8936 29584 8992 29640
rect 9017 29584 9073 29640
rect 9098 29584 9154 29640
rect 9179 29584 9235 29640
rect 2139 29452 2195 29508
rect 2237 29452 2293 29508
rect 2335 29452 2391 29508
rect 2433 29452 2489 29508
rect 5803 29499 5859 29555
rect 5895 29499 5951 29555
rect 5987 29499 6043 29555
rect 6079 29499 6135 29555
rect 6182 29504 6238 29560
rect 6263 29504 6319 29560
rect 6344 29504 6400 29560
rect 6425 29504 6481 29560
rect 6506 29504 6562 29560
rect 6587 29504 6643 29560
rect 6668 29504 6724 29560
rect 6749 29504 6805 29560
rect 6830 29504 6886 29560
rect 6911 29504 6967 29560
rect 6992 29504 7048 29560
rect 7073 29504 7129 29560
rect 7154 29504 7210 29560
rect 7235 29504 7291 29560
rect 7316 29504 7372 29560
rect 7397 29504 7453 29560
rect 7478 29504 7534 29560
rect 7559 29504 7615 29560
rect 7640 29504 7696 29560
rect 7721 29504 7777 29560
rect 7802 29504 7858 29560
rect 7883 29504 7939 29560
rect 7964 29504 8020 29560
rect 8045 29504 8101 29560
rect 8126 29504 8182 29560
rect 8207 29504 8263 29560
rect 8288 29504 8344 29560
rect 8369 29504 8425 29560
rect 8450 29504 8506 29560
rect 8531 29504 8587 29560
rect 8612 29504 8668 29560
rect 8693 29504 8749 29560
rect 8774 29504 8830 29560
rect 8855 29504 8911 29560
rect 8936 29504 8992 29560
rect 9017 29504 9073 29560
rect 9098 29504 9154 29560
rect 9179 29504 9235 29560
rect 298 29414 354 29423
rect 298 29367 299 29414
rect 299 29367 354 29414
rect 396 29367 452 29423
rect 494 29414 550 29423
rect 592 29414 648 29423
rect 494 29367 506 29414
rect 506 29367 528 29414
rect 528 29367 550 29414
rect 592 29367 602 29414
rect 602 29367 648 29414
rect 298 29297 299 29342
rect 299 29297 354 29342
rect 298 29286 354 29297
rect 396 29286 452 29342
rect 494 29297 506 29342
rect 506 29297 528 29342
rect 528 29297 550 29342
rect 592 29297 602 29342
rect 602 29297 648 29342
rect 494 29286 550 29297
rect 592 29286 648 29297
rect 298 29232 299 29261
rect 299 29232 354 29261
rect 298 29219 354 29232
rect 298 29205 299 29219
rect 299 29205 354 29219
rect 396 29205 452 29261
rect 494 29232 506 29261
rect 506 29232 528 29261
rect 528 29232 550 29261
rect 592 29232 602 29261
rect 602 29232 648 29261
rect 494 29219 550 29232
rect 592 29219 648 29232
rect 494 29205 506 29219
rect 506 29205 528 29219
rect 528 29205 550 29219
rect 592 29205 602 29219
rect 602 29205 648 29219
rect 298 29167 299 29180
rect 299 29167 354 29180
rect 298 29154 354 29167
rect 298 29124 299 29154
rect 299 29124 354 29154
rect 396 29124 452 29180
rect 494 29167 506 29180
rect 506 29167 528 29180
rect 528 29167 550 29180
rect 592 29167 602 29180
rect 602 29167 648 29180
rect 494 29154 550 29167
rect 592 29154 648 29167
rect 494 29124 506 29154
rect 506 29124 528 29154
rect 528 29124 550 29154
rect 592 29124 602 29154
rect 602 29124 648 29154
rect 298 29089 354 29099
rect 298 29043 299 29089
rect 299 29043 354 29089
rect 396 29043 452 29099
rect 494 29089 550 29099
rect 592 29089 648 29099
rect 494 29043 506 29089
rect 506 29043 528 29089
rect 528 29043 550 29089
rect 592 29043 602 29089
rect 602 29043 648 29089
rect 2139 29369 2195 29425
rect 2237 29369 2293 29425
rect 2335 29369 2391 29425
rect 2433 29369 2489 29425
rect 5803 29416 5859 29472
rect 5895 29416 5951 29472
rect 5987 29416 6043 29472
rect 6079 29416 6135 29472
rect 6182 29424 6238 29480
rect 6263 29424 6319 29480
rect 6344 29424 6400 29480
rect 6425 29424 6481 29480
rect 6506 29424 6562 29480
rect 6587 29424 6643 29480
rect 6668 29424 6724 29480
rect 6749 29424 6805 29480
rect 6830 29424 6886 29480
rect 6911 29424 6967 29480
rect 6992 29424 7048 29480
rect 7073 29424 7129 29480
rect 7154 29424 7210 29480
rect 7235 29424 7291 29480
rect 7316 29424 7372 29480
rect 7397 29424 7453 29480
rect 7478 29424 7534 29480
rect 7559 29424 7615 29480
rect 7640 29424 7696 29480
rect 7721 29424 7777 29480
rect 7802 29424 7858 29480
rect 7883 29424 7939 29480
rect 7964 29424 8020 29480
rect 8045 29424 8101 29480
rect 8126 29424 8182 29480
rect 8207 29424 8263 29480
rect 8288 29424 8344 29480
rect 8369 29424 8425 29480
rect 8450 29424 8506 29480
rect 8531 29424 8587 29480
rect 8612 29424 8668 29480
rect 8693 29424 8749 29480
rect 8774 29424 8830 29480
rect 8855 29424 8911 29480
rect 8936 29424 8992 29480
rect 9017 29424 9073 29480
rect 9098 29424 9154 29480
rect 9179 29424 9235 29480
rect 2139 29286 2195 29342
rect 2237 29286 2293 29342
rect 2335 29286 2391 29342
rect 2433 29286 2489 29342
rect 5803 29333 5859 29389
rect 5895 29333 5951 29389
rect 5987 29333 6043 29389
rect 6079 29333 6135 29389
rect 6182 29344 6238 29400
rect 6263 29344 6319 29400
rect 6344 29344 6400 29400
rect 6425 29344 6481 29400
rect 6506 29344 6562 29400
rect 6587 29344 6643 29400
rect 6668 29344 6724 29400
rect 6749 29344 6805 29400
rect 6830 29344 6886 29400
rect 6911 29344 6967 29400
rect 6992 29344 7048 29400
rect 7073 29344 7129 29400
rect 7154 29344 7210 29400
rect 7235 29344 7291 29400
rect 7316 29344 7372 29400
rect 7397 29344 7453 29400
rect 7478 29344 7534 29400
rect 7559 29344 7615 29400
rect 7640 29344 7696 29400
rect 7721 29344 7777 29400
rect 7802 29344 7858 29400
rect 7883 29344 7939 29400
rect 7964 29344 8020 29400
rect 8045 29344 8101 29400
rect 8126 29344 8182 29400
rect 8207 29344 8263 29400
rect 8288 29344 8344 29400
rect 8369 29344 8425 29400
rect 8450 29344 8506 29400
rect 8531 29344 8587 29400
rect 8612 29344 8668 29400
rect 8693 29344 8749 29400
rect 8774 29344 8830 29400
rect 8855 29344 8911 29400
rect 8936 29344 8992 29400
rect 9017 29344 9073 29400
rect 9098 29344 9154 29400
rect 9179 29344 9235 29400
rect 2139 29203 2195 29259
rect 2237 29203 2293 29259
rect 2335 29203 2391 29259
rect 2433 29203 2489 29259
rect 5803 29250 5859 29306
rect 5895 29250 5951 29306
rect 5987 29250 6043 29306
rect 6079 29250 6135 29306
rect 6182 29264 6238 29320
rect 6263 29264 6319 29320
rect 6344 29264 6400 29320
rect 6425 29264 6481 29320
rect 6506 29264 6562 29320
rect 6587 29264 6643 29320
rect 6668 29264 6724 29320
rect 6749 29264 6805 29320
rect 6830 29264 6886 29320
rect 6911 29264 6967 29320
rect 6992 29264 7048 29320
rect 7073 29264 7129 29320
rect 7154 29264 7210 29320
rect 7235 29264 7291 29320
rect 7316 29264 7372 29320
rect 7397 29264 7453 29320
rect 7478 29264 7534 29320
rect 7559 29264 7615 29320
rect 7640 29264 7696 29320
rect 7721 29264 7777 29320
rect 7802 29264 7858 29320
rect 7883 29264 7939 29320
rect 7964 29264 8020 29320
rect 8045 29264 8101 29320
rect 8126 29264 8182 29320
rect 8207 29264 8263 29320
rect 8288 29264 8344 29320
rect 8369 29264 8425 29320
rect 8450 29264 8506 29320
rect 8531 29264 8587 29320
rect 8612 29264 8668 29320
rect 8693 29264 8749 29320
rect 8774 29264 8830 29320
rect 8855 29264 8911 29320
rect 8936 29264 8992 29320
rect 9017 29264 9073 29320
rect 9098 29264 9154 29320
rect 9179 29264 9235 29320
rect 2139 29120 2195 29176
rect 2237 29120 2293 29176
rect 2335 29120 2391 29176
rect 2433 29120 2489 29176
rect 5803 29167 5859 29223
rect 5895 29167 5951 29223
rect 5987 29167 6043 29223
rect 6079 29167 6135 29223
rect 6182 29184 6238 29240
rect 6263 29184 6319 29240
rect 6344 29184 6400 29240
rect 6425 29184 6481 29240
rect 6506 29184 6562 29240
rect 6587 29184 6643 29240
rect 6668 29184 6724 29240
rect 6749 29184 6805 29240
rect 6830 29184 6886 29240
rect 6911 29184 6967 29240
rect 6992 29184 7048 29240
rect 7073 29184 7129 29240
rect 7154 29184 7210 29240
rect 7235 29184 7291 29240
rect 7316 29184 7372 29240
rect 7397 29184 7453 29240
rect 7478 29184 7534 29240
rect 7559 29184 7615 29240
rect 7640 29184 7696 29240
rect 7721 29184 7777 29240
rect 7802 29184 7858 29240
rect 7883 29184 7939 29240
rect 7964 29184 8020 29240
rect 8045 29184 8101 29240
rect 8126 29184 8182 29240
rect 8207 29184 8263 29240
rect 8288 29184 8344 29240
rect 8369 29184 8425 29240
rect 8450 29184 8506 29240
rect 8531 29184 8587 29240
rect 8612 29184 8668 29240
rect 8693 29184 8749 29240
rect 8774 29184 8830 29240
rect 8855 29184 8911 29240
rect 8936 29184 8992 29240
rect 9017 29184 9073 29240
rect 9098 29184 9154 29240
rect 9179 29184 9235 29240
rect 2139 29037 2195 29093
rect 2237 29037 2293 29093
rect 2335 29037 2391 29093
rect 2433 29037 2489 29093
rect 5803 29084 5859 29140
rect 5895 29084 5951 29140
rect 5987 29084 6043 29140
rect 6079 29084 6135 29140
rect 6182 29104 6238 29160
rect 6263 29104 6319 29160
rect 6344 29104 6400 29160
rect 6425 29104 6481 29160
rect 6506 29104 6562 29160
rect 6587 29104 6643 29160
rect 6668 29104 6724 29160
rect 6749 29104 6805 29160
rect 6830 29104 6886 29160
rect 6911 29104 6967 29160
rect 6992 29104 7048 29160
rect 7073 29104 7129 29160
rect 7154 29104 7210 29160
rect 7235 29104 7291 29160
rect 7316 29104 7372 29160
rect 7397 29104 7453 29160
rect 7478 29104 7534 29160
rect 7559 29104 7615 29160
rect 7640 29104 7696 29160
rect 7721 29104 7777 29160
rect 7802 29104 7858 29160
rect 7883 29104 7939 29160
rect 7964 29104 8020 29160
rect 8045 29104 8101 29160
rect 8126 29104 8182 29160
rect 8207 29104 8263 29160
rect 8288 29104 8344 29160
rect 8369 29104 8425 29160
rect 8450 29104 8506 29160
rect 8531 29104 8587 29160
rect 8612 29104 8668 29160
rect 8693 29104 8749 29160
rect 8774 29104 8830 29160
rect 8855 29104 8911 29160
rect 8936 29104 8992 29160
rect 9017 29104 9073 29160
rect 9098 29104 9154 29160
rect 9179 29104 9235 29160
rect 6182 29024 6238 29080
rect 6263 29024 6319 29080
rect 6344 29024 6400 29080
rect 6425 29024 6481 29080
rect 6506 29024 6562 29080
rect 6587 29024 6643 29080
rect 6668 29024 6724 29080
rect 6749 29024 6805 29080
rect 6830 29024 6886 29080
rect 6911 29024 6967 29080
rect 6992 29024 7048 29080
rect 7073 29024 7129 29080
rect 7154 29024 7210 29080
rect 7235 29024 7291 29080
rect 7316 29024 7372 29080
rect 7397 29024 7453 29080
rect 7478 29024 7534 29080
rect 7559 29024 7615 29080
rect 7640 29024 7696 29080
rect 7721 29024 7777 29080
rect 7802 29024 7858 29080
rect 7883 29024 7939 29080
rect 7964 29024 8020 29080
rect 8045 29024 8101 29080
rect 8126 29024 8182 29080
rect 8207 29024 8263 29080
rect 8288 29024 8344 29080
rect 8369 29024 8425 29080
rect 8450 29024 8506 29080
rect 8531 29024 8587 29080
rect 8612 29024 8668 29080
rect 8693 29024 8749 29080
rect 8774 29024 8830 29080
rect 8855 29024 8911 29080
rect 8936 29024 8992 29080
rect 9017 29024 9073 29080
rect 9098 29024 9154 29080
rect 9179 29024 9235 29080
rect 2139 28954 2195 29010
rect 2237 28954 2293 29010
rect 2335 28954 2391 29010
rect 2433 28954 2489 29010
rect 6182 28944 6238 29000
rect 6263 28944 6319 29000
rect 6344 28944 6400 29000
rect 6425 28944 6481 29000
rect 6506 28944 6562 29000
rect 6587 28944 6643 29000
rect 6668 28944 6724 29000
rect 6749 28944 6805 29000
rect 6830 28944 6886 29000
rect 6911 28944 6967 29000
rect 6992 28944 7048 29000
rect 7073 28944 7129 29000
rect 7154 28944 7210 29000
rect 7235 28944 7291 29000
rect 7316 28944 7372 29000
rect 7397 28944 7453 29000
rect 7478 28944 7534 29000
rect 7559 28944 7615 29000
rect 7640 28944 7696 29000
rect 7721 28944 7777 29000
rect 7802 28944 7858 29000
rect 7883 28944 7939 29000
rect 7964 28944 8020 29000
rect 8045 28944 8101 29000
rect 8126 28944 8182 29000
rect 8207 28944 8263 29000
rect 8288 28944 8344 29000
rect 8369 28944 8425 29000
rect 8450 28944 8506 29000
rect 8531 28944 8587 29000
rect 8612 28944 8668 29000
rect 8693 28944 8749 29000
rect 8774 28944 8830 29000
rect 8855 28944 8911 29000
rect 8936 28944 8992 29000
rect 9017 28944 9073 29000
rect 9098 28944 9154 29000
rect 9179 28944 9235 29000
rect 2139 28871 2195 28927
rect 2237 28871 2293 28927
rect 2335 28871 2391 28927
rect 2433 28871 2489 28927
rect 6182 28864 6238 28920
rect 6263 28864 6319 28920
rect 6344 28864 6400 28920
rect 6425 28864 6481 28920
rect 6506 28864 6562 28920
rect 6587 28864 6643 28920
rect 6668 28864 6724 28920
rect 6749 28864 6805 28920
rect 6830 28864 6886 28920
rect 6911 28864 6967 28920
rect 6992 28864 7048 28920
rect 7073 28864 7129 28920
rect 7154 28864 7210 28920
rect 7235 28864 7291 28920
rect 7316 28864 7372 28920
rect 7397 28864 7453 28920
rect 7478 28864 7534 28920
rect 7559 28864 7615 28920
rect 7640 28864 7696 28920
rect 7721 28864 7777 28920
rect 7802 28864 7858 28920
rect 7883 28864 7939 28920
rect 7964 28864 8020 28920
rect 8045 28864 8101 28920
rect 8126 28864 8182 28920
rect 8207 28864 8263 28920
rect 8288 28864 8344 28920
rect 8369 28864 8425 28920
rect 8450 28864 8506 28920
rect 8531 28864 8587 28920
rect 8612 28864 8668 28920
rect 8693 28864 8749 28920
rect 8774 28864 8830 28920
rect 8855 28864 8911 28920
rect 8936 28864 8992 28920
rect 9017 28864 9073 28920
rect 9098 28864 9154 28920
rect 9179 28864 9235 28920
rect 9260 28864 13076 29880
rect 14514 29867 14570 29923
rect 14594 29867 14650 29923
rect 14674 29867 14730 29923
rect 14754 29867 14810 29923
rect 14834 29867 14890 29923
rect 14914 29867 14970 29923
rect 14994 29867 15050 29923
rect 15074 29867 15130 29923
rect 15154 29867 15210 29923
rect 15234 29867 15290 29923
rect 14514 29784 14570 29840
rect 14594 29784 14650 29840
rect 14674 29784 14730 29840
rect 14754 29784 14810 29840
rect 14834 29784 14890 29840
rect 14914 29784 14970 29840
rect 14994 29784 15050 29840
rect 15074 29784 15130 29840
rect 15154 29784 15210 29840
rect 15234 29784 15290 29840
rect 14514 29701 14570 29757
rect 14594 29701 14650 29757
rect 14674 29701 14730 29757
rect 14754 29701 14810 29757
rect 14834 29701 14890 29757
rect 14914 29701 14970 29757
rect 14994 29701 15050 29757
rect 15074 29701 15130 29757
rect 15154 29701 15210 29757
rect 15234 29701 15290 29757
rect 14514 29618 14570 29674
rect 14594 29618 14650 29674
rect 14674 29618 14730 29674
rect 14754 29618 14810 29674
rect 14834 29618 14890 29674
rect 14914 29618 14970 29674
rect 14994 29618 15050 29674
rect 15074 29618 15130 29674
rect 15154 29618 15210 29674
rect 15234 29618 15290 29674
rect 14514 29535 14570 29591
rect 14594 29535 14650 29591
rect 14674 29535 14730 29591
rect 14754 29535 14810 29591
rect 14834 29535 14890 29591
rect 14914 29535 14970 29591
rect 14994 29535 15050 29591
rect 15074 29535 15130 29591
rect 15154 29535 15210 29591
rect 15234 29535 15290 29591
rect 14514 29452 14570 29508
rect 14594 29452 14650 29508
rect 14674 29452 14730 29508
rect 14754 29452 14810 29508
rect 14834 29452 14890 29508
rect 14914 29452 14970 29508
rect 14994 29452 15050 29508
rect 15074 29452 15130 29508
rect 15154 29452 15210 29508
rect 15234 29452 15290 29508
rect 14514 29369 14570 29425
rect 14594 29369 14650 29425
rect 14674 29369 14730 29425
rect 14754 29369 14810 29425
rect 14834 29369 14890 29425
rect 14914 29369 14970 29425
rect 14994 29369 15050 29425
rect 15074 29369 15130 29425
rect 15154 29369 15210 29425
rect 15234 29369 15290 29425
rect 14514 29286 14570 29342
rect 14594 29286 14650 29342
rect 14674 29286 14730 29342
rect 14754 29286 14810 29342
rect 14834 29286 14890 29342
rect 14914 29286 14970 29342
rect 14994 29286 15050 29342
rect 15074 29286 15130 29342
rect 15154 29286 15210 29342
rect 15234 29286 15290 29342
rect 14514 29203 14570 29259
rect 14594 29203 14650 29259
rect 14674 29203 14730 29259
rect 14754 29203 14810 29259
rect 14834 29203 14890 29259
rect 14914 29203 14970 29259
rect 14994 29203 15050 29259
rect 15074 29203 15130 29259
rect 15154 29203 15210 29259
rect 15234 29203 15290 29259
rect 14514 29120 14570 29176
rect 14594 29120 14650 29176
rect 14674 29120 14730 29176
rect 14754 29120 14810 29176
rect 14834 29120 14890 29176
rect 14914 29120 14970 29176
rect 14994 29120 15050 29176
rect 15074 29120 15130 29176
rect 15154 29120 15210 29176
rect 15234 29120 15290 29176
rect 14514 29037 14570 29093
rect 14594 29037 14650 29093
rect 14674 29037 14730 29093
rect 14754 29037 14810 29093
rect 14834 29037 14890 29093
rect 14914 29037 14970 29093
rect 14994 29037 15050 29093
rect 15074 29037 15130 29093
rect 15154 29037 15210 29093
rect 15234 29037 15290 29093
rect 14514 28954 14570 29010
rect 14594 28954 14650 29010
rect 14674 28954 14730 29010
rect 14754 28954 14810 29010
rect 14834 28954 14890 29010
rect 14914 28954 14970 29010
rect 14994 28954 15050 29010
rect 15074 28954 15130 29010
rect 15154 28954 15210 29010
rect 15234 28954 15290 29010
rect 14514 28871 14570 28927
rect 14594 28871 14650 28927
rect 14674 28871 14730 28927
rect 14754 28871 14810 28927
rect 14834 28871 14890 28927
rect 14914 28871 14970 28927
rect 14994 28871 15050 28927
rect 15074 28871 15130 28927
rect 15154 28871 15210 28927
rect 15234 28871 15290 28927
rect 2790 28561 2846 28562
rect 2874 28561 2930 28562
rect 2958 28561 3014 28562
rect 3042 28561 3098 28562
rect 3126 28561 3182 28562
rect 3210 28561 3266 28562
rect 3294 28561 3350 28562
rect 3378 28561 3434 28562
rect 3462 28561 3518 28562
rect 3545 28561 3601 28562
rect 3628 28561 3684 28562
rect 3711 28561 3767 28562
rect 2790 28509 2840 28561
rect 2840 28509 2846 28561
rect 2874 28509 2906 28561
rect 2906 28509 2919 28561
rect 2919 28509 2930 28561
rect 2958 28509 2971 28561
rect 2971 28509 2984 28561
rect 2984 28509 3014 28561
rect 3042 28509 3049 28561
rect 3049 28509 3098 28561
rect 3126 28509 3166 28561
rect 3166 28509 3179 28561
rect 3179 28509 3182 28561
rect 3210 28509 3231 28561
rect 3231 28509 3244 28561
rect 3244 28509 3266 28561
rect 3294 28509 3296 28561
rect 3296 28509 3309 28561
rect 3309 28509 3350 28561
rect 3378 28509 3426 28561
rect 3426 28509 3434 28561
rect 3462 28509 3491 28561
rect 3491 28509 3504 28561
rect 3504 28509 3518 28561
rect 3545 28509 3556 28561
rect 3556 28509 3569 28561
rect 3569 28509 3601 28561
rect 3628 28509 3634 28561
rect 3634 28509 3684 28561
rect 3711 28509 3751 28561
rect 3751 28509 3767 28561
rect 2790 28506 2846 28509
rect 2874 28506 2930 28509
rect 2958 28506 3014 28509
rect 3042 28506 3098 28509
rect 3126 28506 3182 28509
rect 3210 28506 3266 28509
rect 3294 28506 3350 28509
rect 3378 28506 3434 28509
rect 3462 28506 3518 28509
rect 3545 28506 3601 28509
rect 3628 28506 3684 28509
rect 3711 28506 3767 28509
rect 2790 28421 2846 28424
rect 2874 28421 2930 28424
rect 2958 28421 3014 28424
rect 3042 28421 3098 28424
rect 3126 28421 3182 28424
rect 3210 28421 3266 28424
rect 3294 28421 3350 28424
rect 3378 28421 3434 28424
rect 3462 28421 3518 28424
rect 3545 28421 3601 28424
rect 3628 28421 3684 28424
rect 3711 28421 3767 28424
rect 2790 28369 2840 28421
rect 2840 28369 2846 28421
rect 2874 28369 2906 28421
rect 2906 28369 2919 28421
rect 2919 28369 2930 28421
rect 2958 28369 2971 28421
rect 2971 28369 2984 28421
rect 2984 28369 3014 28421
rect 3042 28369 3049 28421
rect 3049 28369 3098 28421
rect 3126 28369 3166 28421
rect 3166 28369 3179 28421
rect 3179 28369 3182 28421
rect 3210 28369 3231 28421
rect 3231 28369 3244 28421
rect 3244 28369 3266 28421
rect 3294 28369 3296 28421
rect 3296 28369 3309 28421
rect 3309 28369 3350 28421
rect 3378 28369 3426 28421
rect 3426 28369 3434 28421
rect 3462 28369 3491 28421
rect 3491 28369 3504 28421
rect 3504 28369 3518 28421
rect 3545 28369 3556 28421
rect 3556 28369 3569 28421
rect 3569 28369 3601 28421
rect 3628 28369 3634 28421
rect 3634 28369 3684 28421
rect 3711 28369 3751 28421
rect 3751 28369 3767 28421
rect 2790 28368 2846 28369
rect 2874 28368 2930 28369
rect 2958 28368 3014 28369
rect 3042 28368 3098 28369
rect 3126 28368 3182 28369
rect 3210 28368 3266 28369
rect 3294 28368 3350 28369
rect 3378 28368 3434 28369
rect 3462 28368 3518 28369
rect 3545 28368 3601 28369
rect 3628 28368 3684 28369
rect 3711 28368 3767 28369
rect 299 27959 355 28015
rect 393 27959 449 28015
rect 487 27972 506 28015
rect 506 27972 528 28015
rect 528 27972 543 28015
rect 581 27972 602 28015
rect 602 27972 637 28015
rect 487 27959 543 27972
rect 581 27959 637 27972
rect 299 27877 355 27933
rect 393 27877 449 27933
rect 487 27906 506 27933
rect 506 27906 528 27933
rect 528 27906 543 27933
rect 581 27906 602 27933
rect 602 27906 637 27933
rect 487 27892 543 27906
rect 581 27892 637 27906
rect 487 27877 506 27892
rect 506 27877 528 27892
rect 528 27877 543 27892
rect 581 27877 602 27892
rect 602 27877 637 27892
rect 299 27795 355 27851
rect 393 27795 449 27851
rect 487 27840 506 27851
rect 506 27840 528 27851
rect 528 27840 543 27851
rect 581 27840 602 27851
rect 602 27840 637 27851
rect 487 27826 543 27840
rect 581 27826 637 27840
rect 487 27795 506 27826
rect 506 27795 528 27826
rect 528 27795 543 27826
rect 581 27795 602 27826
rect 602 27795 637 27826
rect 299 27713 355 27769
rect 393 27713 449 27769
rect 487 27760 543 27769
rect 581 27760 637 27769
rect 487 27713 506 27760
rect 506 27713 528 27760
rect 528 27713 543 27760
rect 581 27713 602 27760
rect 602 27713 637 27760
rect 299 27631 355 27687
rect 393 27631 449 27687
rect 487 27642 506 27687
rect 506 27642 528 27687
rect 528 27642 543 27687
rect 581 27642 602 27687
rect 602 27642 637 27687
rect 487 27631 543 27642
rect 581 27631 637 27642
rect 299 27549 355 27605
rect 393 27549 449 27605
rect 487 27576 506 27605
rect 506 27576 528 27605
rect 528 27576 543 27605
rect 581 27576 602 27605
rect 602 27576 637 27605
rect 487 27562 543 27576
rect 581 27562 637 27576
rect 487 27549 506 27562
rect 506 27549 528 27562
rect 528 27549 543 27562
rect 581 27549 602 27562
rect 602 27549 637 27562
rect 299 27467 355 27523
rect 393 27467 449 27523
rect 487 27510 506 27523
rect 506 27510 528 27523
rect 528 27510 543 27523
rect 581 27510 602 27523
rect 602 27510 637 27523
rect 487 27496 543 27510
rect 581 27496 637 27510
rect 487 27467 506 27496
rect 506 27467 528 27496
rect 528 27467 543 27496
rect 581 27467 602 27496
rect 602 27467 637 27496
rect 299 27385 355 27441
rect 393 27385 449 27441
rect 487 27430 543 27441
rect 581 27430 637 27441
rect 487 27385 506 27430
rect 506 27385 528 27430
rect 528 27385 543 27430
rect 581 27385 602 27430
rect 602 27385 637 27430
rect 299 27303 355 27359
rect 393 27303 449 27359
rect 487 27312 506 27359
rect 506 27312 528 27359
rect 528 27312 543 27359
rect 581 27312 602 27359
rect 602 27312 637 27359
rect 487 27303 543 27312
rect 581 27303 637 27312
rect 299 27221 355 27277
rect 393 27221 449 27277
rect 487 27246 506 27277
rect 506 27246 528 27277
rect 528 27246 543 27277
rect 581 27246 602 27277
rect 602 27246 637 27277
rect 487 27232 543 27246
rect 581 27232 637 27246
rect 487 27221 506 27232
rect 506 27221 528 27232
rect 528 27221 543 27232
rect 581 27221 602 27232
rect 602 27221 637 27232
rect 299 27139 355 27195
rect 393 27139 449 27195
rect 487 27180 506 27195
rect 506 27180 528 27195
rect 528 27180 543 27195
rect 581 27180 602 27195
rect 602 27180 637 27195
rect 487 27167 543 27180
rect 581 27167 637 27180
rect 487 27139 506 27167
rect 506 27139 528 27167
rect 528 27139 543 27167
rect 581 27139 602 27167
rect 602 27139 637 27167
rect 299 27056 355 27112
rect 393 27056 449 27112
rect 487 27102 543 27112
rect 581 27102 637 27112
rect 487 27056 506 27102
rect 506 27056 528 27102
rect 528 27056 543 27102
rect 581 27056 602 27102
rect 602 27056 637 27102
rect 299 26973 355 27029
rect 393 26973 449 27029
rect 487 26985 506 27029
rect 506 26985 528 27029
rect 528 26985 543 27029
rect 581 26985 602 27029
rect 602 26985 637 27029
rect 487 26973 543 26985
rect 581 26973 637 26985
rect 299 26890 355 26946
rect 393 26890 449 26946
rect 487 26920 506 26946
rect 506 26920 528 26946
rect 528 26920 543 26946
rect 581 26920 602 26946
rect 602 26920 637 26946
rect 487 26907 543 26920
rect 581 26907 637 26920
rect 487 26890 506 26907
rect 506 26890 528 26907
rect 528 26890 543 26907
rect 581 26890 602 26907
rect 602 26890 637 26907
rect 299 26807 355 26863
rect 393 26807 449 26863
rect 487 26855 506 26863
rect 506 26855 528 26863
rect 528 26855 543 26863
rect 581 26855 602 26863
rect 602 26855 637 26863
rect 487 26842 543 26855
rect 581 26842 637 26855
rect 487 26807 506 26842
rect 506 26807 528 26842
rect 528 26807 543 26842
rect 581 26807 602 26842
rect 602 26807 637 26842
rect 299 26724 355 26780
rect 393 26724 449 26780
rect 487 26777 543 26780
rect 581 26777 637 26780
rect 487 26725 506 26777
rect 506 26725 528 26777
rect 528 26725 543 26777
rect 581 26725 602 26777
rect 602 26725 637 26777
rect 487 26724 543 26725
rect 581 26724 637 26725
rect 299 26641 355 26697
rect 393 26641 449 26697
rect 487 26660 506 26697
rect 506 26660 528 26697
rect 528 26660 543 26697
rect 581 26660 602 26697
rect 602 26660 637 26697
rect 487 26647 543 26660
rect 581 26647 637 26660
rect 487 26641 506 26647
rect 506 26641 528 26647
rect 528 26641 543 26647
rect 581 26641 602 26647
rect 602 26641 637 26647
rect 299 26558 355 26614
rect 393 26558 449 26614
rect 487 26595 506 26614
rect 506 26595 528 26614
rect 528 26595 543 26614
rect 581 26595 602 26614
rect 602 26595 637 26614
rect 487 26582 543 26595
rect 581 26582 637 26595
rect 487 26558 506 26582
rect 506 26558 528 26582
rect 528 26558 543 26582
rect 581 26558 602 26582
rect 602 26558 637 26582
rect 299 26475 355 26531
rect 393 26475 449 26531
rect 487 26530 506 26531
rect 506 26530 528 26531
rect 528 26530 543 26531
rect 581 26530 602 26531
rect 602 26530 637 26531
rect 487 26517 543 26530
rect 581 26517 637 26530
rect 487 26475 506 26517
rect 506 26475 528 26517
rect 528 26475 543 26517
rect 581 26475 602 26517
rect 602 26475 637 26517
rect 299 26392 355 26448
rect 393 26392 449 26448
rect 487 26400 506 26448
rect 506 26400 528 26448
rect 528 26400 543 26448
rect 581 26400 602 26448
rect 602 26400 637 26448
rect 487 26392 543 26400
rect 581 26392 637 26400
rect 2165 28001 2221 28057
rect 2255 28001 2311 28057
rect 2345 28001 2401 28057
rect 2435 28001 2491 28057
rect 4105 28001 4161 28057
rect 4189 28001 4245 28057
rect 4273 28001 4329 28057
rect 4357 28001 4413 28057
rect 4441 28001 4497 28057
rect 4525 28001 4581 28057
rect 4609 28001 4665 28057
rect 4693 28001 4749 28057
rect 4777 28001 4833 28057
rect 4861 28001 4917 28057
rect 4945 28001 5001 28057
rect 5029 28001 5085 28057
rect 2165 27921 2221 27977
rect 2255 27921 2311 27977
rect 2345 27921 2401 27977
rect 2435 27921 2491 27977
rect 4105 27921 4161 27977
rect 4189 27921 4245 27977
rect 4273 27921 4329 27977
rect 4357 27921 4413 27977
rect 4441 27921 4497 27977
rect 4525 27921 4581 27977
rect 4609 27921 4665 27977
rect 4693 27921 4749 27977
rect 4777 27921 4833 27977
rect 4861 27921 4917 27977
rect 4945 27921 5001 27977
rect 5029 27921 5085 27977
rect 2165 27841 2221 27897
rect 2255 27841 2311 27897
rect 2345 27841 2401 27897
rect 2435 27841 2491 27897
rect 4105 27841 4161 27897
rect 4189 27841 4245 27897
rect 4273 27841 4329 27897
rect 4357 27841 4413 27897
rect 4441 27841 4497 27897
rect 4525 27841 4581 27897
rect 4609 27841 4665 27897
rect 4693 27841 4749 27897
rect 4777 27841 4833 27897
rect 4861 27841 4917 27897
rect 4945 27841 5001 27897
rect 5029 27841 5085 27897
rect 2165 27761 2221 27817
rect 2255 27761 2311 27817
rect 2345 27761 2401 27817
rect 2435 27761 2491 27817
rect 4105 27761 4161 27817
rect 4189 27761 4245 27817
rect 4273 27761 4329 27817
rect 4357 27761 4413 27817
rect 4441 27761 4497 27817
rect 4525 27761 4581 27817
rect 4609 27761 4665 27817
rect 4693 27761 4749 27817
rect 4777 27761 4833 27817
rect 4861 27761 4917 27817
rect 4945 27761 5001 27817
rect 5029 27761 5085 27817
rect 2165 27681 2221 27737
rect 2255 27681 2311 27737
rect 2345 27681 2401 27737
rect 2435 27681 2491 27737
rect 4105 27681 4161 27737
rect 4189 27681 4245 27737
rect 4273 27681 4329 27737
rect 4357 27681 4413 27737
rect 4441 27681 4497 27737
rect 4525 27681 4581 27737
rect 4609 27681 4665 27737
rect 4693 27681 4749 27737
rect 4777 27681 4833 27737
rect 4861 27681 4917 27737
rect 4945 27681 5001 27737
rect 5029 27681 5085 27737
rect 2165 27601 2221 27657
rect 2255 27601 2311 27657
rect 2345 27601 2401 27657
rect 2435 27601 2491 27657
rect 4105 27601 4161 27657
rect 4189 27601 4245 27657
rect 4273 27601 4329 27657
rect 4357 27601 4413 27657
rect 4441 27601 4497 27657
rect 4525 27601 4581 27657
rect 4609 27601 4665 27657
rect 4693 27601 4749 27657
rect 4777 27601 4833 27657
rect 4861 27601 4917 27657
rect 4945 27601 5001 27657
rect 5029 27601 5085 27657
rect 2165 27521 2221 27577
rect 2255 27521 2311 27577
rect 2345 27521 2401 27577
rect 2435 27521 2491 27577
rect 4105 27521 4161 27577
rect 4189 27521 4245 27577
rect 4273 27521 4329 27577
rect 4357 27521 4413 27577
rect 4441 27521 4497 27577
rect 4525 27521 4581 27577
rect 4609 27521 4665 27577
rect 4693 27521 4749 27577
rect 4777 27521 4833 27577
rect 4861 27521 4917 27577
rect 4945 27521 5001 27577
rect 5029 27521 5085 27577
rect 2165 27441 2221 27497
rect 2255 27441 2311 27497
rect 2345 27441 2401 27497
rect 2435 27441 2491 27497
rect 4105 27441 4161 27497
rect 4189 27441 4245 27497
rect 4273 27441 4329 27497
rect 4357 27441 4413 27497
rect 4441 27441 4497 27497
rect 4525 27441 4581 27497
rect 4609 27441 4665 27497
rect 4693 27441 4749 27497
rect 4777 27441 4833 27497
rect 4861 27441 4917 27497
rect 4945 27441 5001 27497
rect 5029 27441 5085 27497
rect 2165 27361 2221 27417
rect 2255 27361 2311 27417
rect 2345 27361 2401 27417
rect 2435 27361 2491 27417
rect 4105 27361 4161 27417
rect 4189 27361 4245 27417
rect 4273 27361 4329 27417
rect 4357 27361 4413 27417
rect 4441 27361 4497 27417
rect 4525 27361 4581 27417
rect 4609 27361 4665 27417
rect 4693 27361 4749 27417
rect 4777 27361 4833 27417
rect 4861 27361 4917 27417
rect 4945 27361 5001 27417
rect 5029 27361 5085 27417
rect 2165 27281 2221 27337
rect 2255 27281 2311 27337
rect 2345 27281 2401 27337
rect 2435 27281 2491 27337
rect 4105 27281 4161 27337
rect 4189 27281 4245 27337
rect 4273 27281 4329 27337
rect 4357 27281 4413 27337
rect 4441 27281 4497 27337
rect 4525 27281 4581 27337
rect 4609 27281 4665 27337
rect 4693 27281 4749 27337
rect 4777 27281 4833 27337
rect 4861 27281 4917 27337
rect 4945 27281 5001 27337
rect 5029 27281 5085 27337
rect 2165 27201 2221 27257
rect 2255 27201 2311 27257
rect 2345 27201 2401 27257
rect 2435 27201 2491 27257
rect 4105 27201 4161 27257
rect 4189 27201 4245 27257
rect 4273 27201 4329 27257
rect 4357 27201 4413 27257
rect 4441 27201 4497 27257
rect 4525 27201 4581 27257
rect 4609 27201 4665 27257
rect 4693 27201 4749 27257
rect 4777 27201 4833 27257
rect 4861 27201 4917 27257
rect 4945 27201 5001 27257
rect 5029 27201 5085 27257
rect 2165 27121 2221 27177
rect 2255 27121 2311 27177
rect 2345 27121 2401 27177
rect 2435 27121 2491 27177
rect 4105 27121 4161 27177
rect 4189 27121 4245 27177
rect 4273 27121 4329 27177
rect 4357 27121 4413 27177
rect 4441 27121 4497 27177
rect 4525 27121 4581 27177
rect 4609 27121 4665 27177
rect 4693 27121 4749 27177
rect 4777 27121 4833 27177
rect 4861 27121 4917 27177
rect 4945 27121 5001 27177
rect 5029 27121 5085 27177
rect 2165 27041 2221 27097
rect 2255 27041 2311 27097
rect 2345 27041 2401 27097
rect 2435 27041 2491 27097
rect 4105 27041 4161 27097
rect 4189 27041 4245 27097
rect 4273 27041 4329 27097
rect 4357 27041 4413 27097
rect 4441 27041 4497 27097
rect 4525 27041 4581 27097
rect 4609 27041 4665 27097
rect 4693 27041 4749 27097
rect 4777 27041 4833 27097
rect 4861 27041 4917 27097
rect 4945 27041 5001 27097
rect 5029 27041 5085 27097
rect 2165 26961 2221 27017
rect 2255 26961 2311 27017
rect 2345 26961 2401 27017
rect 2435 26961 2491 27017
rect 4105 26961 4161 27017
rect 4189 26961 4245 27017
rect 4273 26961 4329 27017
rect 4357 26961 4413 27017
rect 4441 26961 4497 27017
rect 4525 26961 4581 27017
rect 4609 26961 4665 27017
rect 4693 26961 4749 27017
rect 4777 26961 4833 27017
rect 4861 26961 4917 27017
rect 4945 26961 5001 27017
rect 5029 26961 5085 27017
rect 2165 26880 2221 26936
rect 2255 26880 2311 26936
rect 2345 26880 2401 26936
rect 2435 26880 2491 26936
rect 4105 26880 4161 26936
rect 4189 26880 4245 26936
rect 4273 26880 4329 26936
rect 4357 26880 4413 26936
rect 4441 26880 4497 26936
rect 4525 26880 4581 26936
rect 4609 26880 4665 26936
rect 4693 26880 4749 26936
rect 4777 26880 4833 26936
rect 4861 26880 4917 26936
rect 4945 26880 5001 26936
rect 5029 26880 5085 26936
rect 2165 26799 2221 26855
rect 2255 26799 2311 26855
rect 2345 26799 2401 26855
rect 2435 26799 2491 26855
rect 4105 26799 4161 26855
rect 4189 26799 4245 26855
rect 4273 26799 4329 26855
rect 4357 26799 4413 26855
rect 4441 26799 4497 26855
rect 4525 26799 4581 26855
rect 4609 26799 4665 26855
rect 4693 26799 4749 26855
rect 4777 26799 4833 26855
rect 4861 26799 4917 26855
rect 4945 26799 5001 26855
rect 5029 26799 5085 26855
rect 2165 26718 2221 26774
rect 2255 26718 2311 26774
rect 2345 26718 2401 26774
rect 2435 26718 2491 26774
rect 4105 26718 4161 26774
rect 4189 26718 4245 26774
rect 4273 26718 4329 26774
rect 4357 26718 4413 26774
rect 4441 26718 4497 26774
rect 4525 26718 4581 26774
rect 4609 26718 4665 26774
rect 4693 26718 4749 26774
rect 4777 26718 4833 26774
rect 4861 26718 4917 26774
rect 4945 26718 5001 26774
rect 5029 26718 5085 26774
rect 2165 26637 2221 26693
rect 2255 26637 2311 26693
rect 2345 26637 2401 26693
rect 2435 26637 2491 26693
rect 4105 26637 4161 26693
rect 4189 26637 4245 26693
rect 4273 26637 4329 26693
rect 4357 26637 4413 26693
rect 4441 26637 4497 26693
rect 4525 26637 4581 26693
rect 4609 26637 4665 26693
rect 4693 26637 4749 26693
rect 4777 26637 4833 26693
rect 4861 26637 4917 26693
rect 4945 26637 5001 26693
rect 5029 26637 5085 26693
rect 2165 26556 2221 26612
rect 2255 26556 2311 26612
rect 2345 26556 2401 26612
rect 2435 26556 2491 26612
rect 4105 26556 4161 26612
rect 4189 26556 4245 26612
rect 4273 26556 4329 26612
rect 4357 26556 4413 26612
rect 4441 26556 4497 26612
rect 4525 26556 4581 26612
rect 4609 26556 4665 26612
rect 4693 26556 4749 26612
rect 4777 26556 4833 26612
rect 4861 26556 4917 26612
rect 4945 26556 5001 26612
rect 5029 26556 5085 26612
rect 2165 26475 2221 26531
rect 2255 26475 2311 26531
rect 2345 26475 2401 26531
rect 2435 26475 2491 26531
rect 4105 26475 4161 26531
rect 4189 26475 4245 26531
rect 4273 26475 4329 26531
rect 4357 26475 4413 26531
rect 4441 26475 4497 26531
rect 4525 26475 4581 26531
rect 4609 26475 4665 26531
rect 4693 26475 4749 26531
rect 4777 26475 4833 26531
rect 4861 26475 4917 26531
rect 4945 26475 5001 26531
rect 5029 26475 5085 26531
rect 2165 26394 2221 26450
rect 2255 26394 2311 26450
rect 2345 26394 2401 26450
rect 2435 26394 2491 26450
rect 4105 26394 4161 26450
rect 4189 26394 4245 26450
rect 4273 26394 4329 26450
rect 4357 26394 4413 26450
rect 4441 26394 4497 26450
rect 4525 26394 4581 26450
rect 4609 26394 4665 26450
rect 4693 26394 4749 26450
rect 4777 26394 4833 26450
rect 4861 26394 4917 26450
rect 4945 26394 5001 26450
rect 5029 26394 5085 26450
rect 14522 27518 14578 27574
rect 14612 27518 14668 27574
rect 14702 27518 14758 27574
rect 14791 27518 14847 27574
rect 14880 27518 14936 27574
rect 14969 27518 15025 27574
rect 14522 27432 14578 27488
rect 14612 27432 14668 27488
rect 14702 27432 14758 27488
rect 14791 27432 14847 27488
rect 14880 27432 14936 27488
rect 14969 27432 15025 27488
rect 14522 27346 14578 27402
rect 14612 27346 14668 27402
rect 14702 27346 14758 27402
rect 14791 27346 14847 27402
rect 14880 27346 14936 27402
rect 14969 27346 15025 27402
rect 14522 27260 14578 27316
rect 14612 27260 14668 27316
rect 14702 27260 14758 27316
rect 14791 27260 14847 27316
rect 14880 27260 14936 27316
rect 14969 27260 15025 27316
rect 14522 27174 14578 27230
rect 14612 27174 14668 27230
rect 14702 27174 14758 27230
rect 14791 27174 14847 27230
rect 14880 27174 14936 27230
rect 14969 27174 15025 27230
rect 14522 27088 14578 27144
rect 14612 27088 14668 27144
rect 14702 27088 14758 27144
rect 14791 27088 14847 27144
rect 14880 27088 14936 27144
rect 14969 27088 15025 27144
rect 299 26309 355 26365
rect 393 26309 449 26365
rect 487 26335 506 26365
rect 506 26335 528 26365
rect 528 26335 543 26365
rect 581 26335 602 26365
rect 602 26335 637 26365
rect 487 26322 543 26335
rect 581 26322 637 26335
rect 487 26309 506 26322
rect 506 26309 528 26322
rect 528 26309 543 26322
rect 581 26309 602 26322
rect 602 26309 637 26322
rect 299 26226 355 26282
rect 393 26226 449 26282
rect 487 26270 506 26282
rect 506 26270 528 26282
rect 528 26270 543 26282
rect 581 26270 602 26282
rect 602 26270 637 26282
rect 487 26257 543 26270
rect 581 26257 637 26270
rect 487 26226 506 26257
rect 506 26226 528 26257
rect 528 26226 543 26257
rect 581 26226 602 26257
rect 602 26226 637 26257
rect 2170 25764 2226 25820
rect 2252 25764 2308 25820
rect 2334 25764 2390 25820
rect 2416 25764 2472 25820
rect 5425 25772 5481 25828
rect 5506 25772 5562 25828
rect 5587 25772 5643 25828
rect 5668 25772 5724 25828
rect 5749 25772 5805 25828
rect 5830 25772 5886 25828
rect 5911 25772 5967 25828
rect 5992 25772 6048 25828
rect 6073 25772 6129 25828
rect 6154 25772 6210 25828
rect 6235 25772 6291 25828
rect 6316 25772 6372 25828
rect 6397 25772 6453 25828
rect 6478 25772 6534 25828
rect 6559 25772 6615 25828
rect 6640 25772 6696 25828
rect 6721 25772 6777 25828
rect 6802 25772 6858 25828
rect 6883 25772 6939 25828
rect 6964 25772 7020 25828
rect 7045 25772 7101 25828
rect 7126 25772 7182 25828
rect 7207 25772 7263 25828
rect 7288 25772 7344 25828
rect 7369 25772 7425 25828
rect 7450 25772 7506 25828
rect 7531 25772 7587 25828
rect 7612 25772 7668 25828
rect 7693 25772 7749 25828
rect 7774 25772 7830 25828
rect 7855 25772 7911 25828
rect 7936 25772 7992 25828
rect 8017 25772 8073 25828
rect 8098 25772 8154 25828
rect 8179 25772 8235 25828
rect 8260 25772 8316 25828
rect 8341 25772 8397 25828
rect 8422 25772 8478 25828
rect 8503 25772 8559 25828
rect 8584 25772 8640 25828
rect 8665 25772 8721 25828
rect 8746 25772 8802 25828
rect 8827 25772 8883 25828
rect 8908 25772 8964 25828
rect 8989 25772 9045 25828
rect 9070 25772 9126 25828
rect 9151 25772 9207 25828
rect 9232 25772 9288 25828
rect 9313 25772 9369 25828
rect 9394 25772 9450 25828
rect 9475 25772 9531 25828
rect 9556 25772 9612 25828
rect 9637 25772 9693 25828
rect 9718 25772 9774 25828
rect 9799 25772 9855 25828
rect 9880 25772 9936 25828
rect 9961 25772 10017 25828
rect 10042 25772 10098 25828
rect 10123 25772 10179 25828
rect 10204 25772 10260 25828
rect 10285 25772 10341 25828
rect 10366 25772 10422 25828
rect 10447 25772 10503 25828
rect 10528 25772 10584 25828
rect 10609 25772 10665 25828
rect 10690 25772 10746 25828
rect 10771 25772 10827 25828
rect 10852 25772 10908 25828
rect 10933 25772 10989 25828
rect 11014 25772 11070 25828
rect 11095 25772 11151 25828
rect 11176 25772 11232 25828
rect 11257 25772 11313 25828
rect 11338 25772 11394 25828
rect 11419 25772 11475 25828
rect 2170 25683 2226 25739
rect 2252 25683 2308 25739
rect 2334 25683 2390 25739
rect 2416 25683 2472 25739
rect 5425 25692 5481 25748
rect 5506 25692 5562 25748
rect 5587 25692 5643 25748
rect 5668 25692 5724 25748
rect 5749 25692 5805 25748
rect 5830 25692 5886 25748
rect 5911 25692 5967 25748
rect 5992 25692 6048 25748
rect 6073 25692 6129 25748
rect 6154 25692 6210 25748
rect 6235 25692 6291 25748
rect 6316 25692 6372 25748
rect 6397 25692 6453 25748
rect 6478 25692 6534 25748
rect 6559 25692 6615 25748
rect 6640 25692 6696 25748
rect 6721 25692 6777 25748
rect 6802 25692 6858 25748
rect 6883 25692 6939 25748
rect 6964 25692 7020 25748
rect 7045 25692 7101 25748
rect 7126 25692 7182 25748
rect 7207 25692 7263 25748
rect 7288 25692 7344 25748
rect 7369 25692 7425 25748
rect 7450 25692 7506 25748
rect 7531 25692 7587 25748
rect 7612 25692 7668 25748
rect 7693 25692 7749 25748
rect 7774 25692 7830 25748
rect 7855 25692 7911 25748
rect 7936 25692 7992 25748
rect 8017 25692 8073 25748
rect 8098 25692 8154 25748
rect 8179 25692 8235 25748
rect 8260 25692 8316 25748
rect 8341 25692 8397 25748
rect 8422 25692 8478 25748
rect 8503 25692 8559 25748
rect 8584 25692 8640 25748
rect 8665 25692 8721 25748
rect 8746 25692 8802 25748
rect 8827 25692 8883 25748
rect 8908 25692 8964 25748
rect 8989 25692 9045 25748
rect 9070 25692 9126 25748
rect 9151 25692 9207 25748
rect 9232 25692 9288 25748
rect 9313 25692 9369 25748
rect 9394 25692 9450 25748
rect 9475 25692 9531 25748
rect 9556 25692 9612 25748
rect 9637 25692 9693 25748
rect 9718 25692 9774 25748
rect 9799 25692 9855 25748
rect 9880 25692 9936 25748
rect 9961 25692 10017 25748
rect 10042 25692 10098 25748
rect 10123 25692 10179 25748
rect 10204 25692 10260 25748
rect 10285 25692 10341 25748
rect 10366 25692 10422 25748
rect 10447 25692 10503 25748
rect 10528 25692 10584 25748
rect 10609 25692 10665 25748
rect 10690 25692 10746 25748
rect 10771 25692 10827 25748
rect 10852 25692 10908 25748
rect 10933 25692 10989 25748
rect 11014 25692 11070 25748
rect 11095 25692 11151 25748
rect 11176 25692 11232 25748
rect 11257 25692 11313 25748
rect 11338 25692 11394 25748
rect 11419 25692 11475 25748
rect 2170 25602 2226 25658
rect 2252 25602 2308 25658
rect 2334 25602 2390 25658
rect 2416 25602 2472 25658
rect 5425 25612 5481 25668
rect 5506 25612 5562 25668
rect 5587 25612 5643 25668
rect 5668 25612 5724 25668
rect 5749 25612 5805 25668
rect 5830 25612 5886 25668
rect 5911 25612 5967 25668
rect 5992 25612 6048 25668
rect 6073 25612 6129 25668
rect 6154 25612 6210 25668
rect 6235 25612 6291 25668
rect 6316 25612 6372 25668
rect 6397 25612 6453 25668
rect 6478 25612 6534 25668
rect 6559 25612 6615 25668
rect 6640 25612 6696 25668
rect 6721 25612 6777 25668
rect 6802 25612 6858 25668
rect 6883 25612 6939 25668
rect 6964 25612 7020 25668
rect 7045 25612 7101 25668
rect 7126 25612 7182 25668
rect 7207 25612 7263 25668
rect 7288 25612 7344 25668
rect 7369 25612 7425 25668
rect 7450 25612 7506 25668
rect 7531 25612 7587 25668
rect 7612 25612 7668 25668
rect 7693 25612 7749 25668
rect 7774 25612 7830 25668
rect 7855 25612 7911 25668
rect 7936 25612 7992 25668
rect 8017 25612 8073 25668
rect 8098 25612 8154 25668
rect 8179 25612 8235 25668
rect 8260 25612 8316 25668
rect 8341 25612 8397 25668
rect 8422 25612 8478 25668
rect 8503 25612 8559 25668
rect 8584 25612 8640 25668
rect 8665 25612 8721 25668
rect 8746 25612 8802 25668
rect 8827 25612 8883 25668
rect 8908 25612 8964 25668
rect 8989 25612 9045 25668
rect 9070 25612 9126 25668
rect 9151 25612 9207 25668
rect 9232 25612 9288 25668
rect 9313 25612 9369 25668
rect 9394 25612 9450 25668
rect 9475 25612 9531 25668
rect 9556 25612 9612 25668
rect 9637 25612 9693 25668
rect 9718 25612 9774 25668
rect 9799 25612 9855 25668
rect 9880 25612 9936 25668
rect 9961 25612 10017 25668
rect 10042 25612 10098 25668
rect 10123 25612 10179 25668
rect 10204 25612 10260 25668
rect 10285 25612 10341 25668
rect 10366 25612 10422 25668
rect 10447 25612 10503 25668
rect 10528 25612 10584 25668
rect 10609 25612 10665 25668
rect 10690 25612 10746 25668
rect 10771 25612 10827 25668
rect 10852 25612 10908 25668
rect 10933 25612 10989 25668
rect 11014 25612 11070 25668
rect 11095 25612 11151 25668
rect 11176 25612 11232 25668
rect 11257 25612 11313 25668
rect 11338 25612 11394 25668
rect 11419 25612 11475 25668
rect 2170 25521 2226 25577
rect 2252 25521 2308 25577
rect 2334 25521 2390 25577
rect 2416 25521 2472 25577
rect 5425 25532 5481 25588
rect 5506 25532 5562 25588
rect 5587 25532 5643 25588
rect 5668 25532 5724 25588
rect 5749 25532 5805 25588
rect 5830 25532 5886 25588
rect 5911 25532 5967 25588
rect 5992 25532 6048 25588
rect 6073 25532 6129 25588
rect 6154 25532 6210 25588
rect 6235 25532 6291 25588
rect 6316 25532 6372 25588
rect 6397 25532 6453 25588
rect 6478 25532 6534 25588
rect 6559 25532 6615 25588
rect 6640 25532 6696 25588
rect 6721 25532 6777 25588
rect 6802 25532 6858 25588
rect 6883 25532 6939 25588
rect 6964 25532 7020 25588
rect 7045 25532 7101 25588
rect 7126 25532 7182 25588
rect 7207 25532 7263 25588
rect 7288 25532 7344 25588
rect 7369 25532 7425 25588
rect 7450 25532 7506 25588
rect 7531 25532 7587 25588
rect 7612 25532 7668 25588
rect 7693 25532 7749 25588
rect 7774 25532 7830 25588
rect 7855 25532 7911 25588
rect 7936 25532 7992 25588
rect 8017 25532 8073 25588
rect 8098 25532 8154 25588
rect 8179 25532 8235 25588
rect 8260 25532 8316 25588
rect 8341 25532 8397 25588
rect 8422 25532 8478 25588
rect 8503 25532 8559 25588
rect 8584 25532 8640 25588
rect 8665 25532 8721 25588
rect 8746 25532 8802 25588
rect 8827 25532 8883 25588
rect 8908 25532 8964 25588
rect 8989 25532 9045 25588
rect 9070 25532 9126 25588
rect 9151 25532 9207 25588
rect 9232 25532 9288 25588
rect 9313 25532 9369 25588
rect 9394 25532 9450 25588
rect 9475 25532 9531 25588
rect 9556 25532 9612 25588
rect 9637 25532 9693 25588
rect 9718 25532 9774 25588
rect 9799 25532 9855 25588
rect 9880 25532 9936 25588
rect 9961 25532 10017 25588
rect 10042 25532 10098 25588
rect 10123 25532 10179 25588
rect 10204 25532 10260 25588
rect 10285 25532 10341 25588
rect 10366 25532 10422 25588
rect 10447 25532 10503 25588
rect 10528 25532 10584 25588
rect 10609 25532 10665 25588
rect 10690 25532 10746 25588
rect 10771 25532 10827 25588
rect 10852 25532 10908 25588
rect 10933 25532 10989 25588
rect 11014 25532 11070 25588
rect 11095 25532 11151 25588
rect 11176 25532 11232 25588
rect 11257 25532 11313 25588
rect 11338 25532 11394 25588
rect 11419 25532 11475 25588
rect 2170 25440 2226 25496
rect 2252 25440 2308 25496
rect 2334 25440 2390 25496
rect 2416 25440 2472 25496
rect 5425 25452 5481 25508
rect 5506 25452 5562 25508
rect 5587 25452 5643 25508
rect 5668 25452 5724 25508
rect 5749 25452 5805 25508
rect 5830 25452 5886 25508
rect 5911 25452 5967 25508
rect 5992 25452 6048 25508
rect 6073 25452 6129 25508
rect 6154 25452 6210 25508
rect 6235 25452 6291 25508
rect 6316 25452 6372 25508
rect 6397 25452 6453 25508
rect 6478 25452 6534 25508
rect 6559 25452 6615 25508
rect 6640 25452 6696 25508
rect 6721 25452 6777 25508
rect 6802 25452 6858 25508
rect 6883 25452 6939 25508
rect 6964 25452 7020 25508
rect 7045 25452 7101 25508
rect 7126 25452 7182 25508
rect 7207 25452 7263 25508
rect 7288 25452 7344 25508
rect 7369 25452 7425 25508
rect 7450 25452 7506 25508
rect 7531 25452 7587 25508
rect 7612 25452 7668 25508
rect 7693 25452 7749 25508
rect 7774 25452 7830 25508
rect 7855 25452 7911 25508
rect 7936 25452 7992 25508
rect 8017 25452 8073 25508
rect 8098 25452 8154 25508
rect 8179 25452 8235 25508
rect 8260 25452 8316 25508
rect 8341 25452 8397 25508
rect 8422 25452 8478 25508
rect 8503 25452 8559 25508
rect 8584 25452 8640 25508
rect 8665 25452 8721 25508
rect 8746 25452 8802 25508
rect 8827 25452 8883 25508
rect 8908 25452 8964 25508
rect 8989 25452 9045 25508
rect 9070 25452 9126 25508
rect 9151 25452 9207 25508
rect 9232 25452 9288 25508
rect 9313 25452 9369 25508
rect 9394 25452 9450 25508
rect 9475 25452 9531 25508
rect 9556 25452 9612 25508
rect 9637 25452 9693 25508
rect 9718 25452 9774 25508
rect 9799 25452 9855 25508
rect 9880 25452 9936 25508
rect 9961 25452 10017 25508
rect 10042 25452 10098 25508
rect 10123 25452 10179 25508
rect 10204 25452 10260 25508
rect 10285 25452 10341 25508
rect 10366 25452 10422 25508
rect 10447 25452 10503 25508
rect 10528 25452 10584 25508
rect 10609 25452 10665 25508
rect 10690 25452 10746 25508
rect 10771 25452 10827 25508
rect 10852 25452 10908 25508
rect 10933 25452 10989 25508
rect 11014 25452 11070 25508
rect 11095 25452 11151 25508
rect 11176 25452 11232 25508
rect 11257 25452 11313 25508
rect 11338 25452 11394 25508
rect 11419 25452 11475 25508
rect 2170 25359 2226 25415
rect 2252 25359 2308 25415
rect 2334 25359 2390 25415
rect 2416 25359 2472 25415
rect 5425 25372 5481 25428
rect 5506 25372 5562 25428
rect 5587 25372 5643 25428
rect 5668 25372 5724 25428
rect 5749 25372 5805 25428
rect 5830 25372 5886 25428
rect 5911 25372 5967 25428
rect 5992 25372 6048 25428
rect 6073 25372 6129 25428
rect 6154 25372 6210 25428
rect 6235 25372 6291 25428
rect 6316 25372 6372 25428
rect 6397 25372 6453 25428
rect 6478 25372 6534 25428
rect 6559 25372 6615 25428
rect 6640 25372 6696 25428
rect 6721 25372 6777 25428
rect 6802 25372 6858 25428
rect 6883 25372 6939 25428
rect 6964 25372 7020 25428
rect 7045 25372 7101 25428
rect 7126 25372 7182 25428
rect 7207 25372 7263 25428
rect 7288 25372 7344 25428
rect 7369 25372 7425 25428
rect 7450 25372 7506 25428
rect 7531 25372 7587 25428
rect 7612 25372 7668 25428
rect 7693 25372 7749 25428
rect 7774 25372 7830 25428
rect 7855 25372 7911 25428
rect 7936 25372 7992 25428
rect 8017 25372 8073 25428
rect 8098 25372 8154 25428
rect 8179 25372 8235 25428
rect 8260 25372 8316 25428
rect 8341 25372 8397 25428
rect 8422 25372 8478 25428
rect 8503 25372 8559 25428
rect 8584 25372 8640 25428
rect 8665 25372 8721 25428
rect 8746 25372 8802 25428
rect 8827 25372 8883 25428
rect 8908 25372 8964 25428
rect 8989 25372 9045 25428
rect 9070 25372 9126 25428
rect 9151 25372 9207 25428
rect 9232 25372 9288 25428
rect 9313 25372 9369 25428
rect 9394 25372 9450 25428
rect 9475 25372 9531 25428
rect 9556 25372 9612 25428
rect 9637 25372 9693 25428
rect 9718 25372 9774 25428
rect 9799 25372 9855 25428
rect 9880 25372 9936 25428
rect 9961 25372 10017 25428
rect 10042 25372 10098 25428
rect 10123 25372 10179 25428
rect 10204 25372 10260 25428
rect 10285 25372 10341 25428
rect 10366 25372 10422 25428
rect 10447 25372 10503 25428
rect 10528 25372 10584 25428
rect 10609 25372 10665 25428
rect 10690 25372 10746 25428
rect 10771 25372 10827 25428
rect 10852 25372 10908 25428
rect 10933 25372 10989 25428
rect 11014 25372 11070 25428
rect 11095 25372 11151 25428
rect 11176 25372 11232 25428
rect 11257 25372 11313 25428
rect 11338 25372 11394 25428
rect 11419 25372 11475 25428
rect 2170 25278 2226 25334
rect 2252 25278 2308 25334
rect 2334 25278 2390 25334
rect 2416 25278 2472 25334
rect 5425 25292 5481 25348
rect 5506 25292 5562 25348
rect 5587 25292 5643 25348
rect 5668 25292 5724 25348
rect 5749 25292 5805 25348
rect 5830 25292 5886 25348
rect 5911 25292 5967 25348
rect 5992 25292 6048 25348
rect 6073 25292 6129 25348
rect 6154 25292 6210 25348
rect 6235 25292 6291 25348
rect 6316 25292 6372 25348
rect 6397 25292 6453 25348
rect 6478 25292 6534 25348
rect 6559 25292 6615 25348
rect 6640 25292 6696 25348
rect 6721 25292 6777 25348
rect 6802 25292 6858 25348
rect 6883 25292 6939 25348
rect 6964 25292 7020 25348
rect 7045 25292 7101 25348
rect 7126 25292 7182 25348
rect 7207 25292 7263 25348
rect 7288 25292 7344 25348
rect 7369 25292 7425 25348
rect 7450 25292 7506 25348
rect 7531 25292 7587 25348
rect 7612 25292 7668 25348
rect 7693 25292 7749 25348
rect 7774 25292 7830 25348
rect 7855 25292 7911 25348
rect 7936 25292 7992 25348
rect 8017 25292 8073 25348
rect 8098 25292 8154 25348
rect 8179 25292 8235 25348
rect 8260 25292 8316 25348
rect 8341 25292 8397 25348
rect 8422 25292 8478 25348
rect 8503 25292 8559 25348
rect 8584 25292 8640 25348
rect 8665 25292 8721 25348
rect 8746 25292 8802 25348
rect 8827 25292 8883 25348
rect 8908 25292 8964 25348
rect 8989 25292 9045 25348
rect 9070 25292 9126 25348
rect 9151 25292 9207 25348
rect 9232 25292 9288 25348
rect 9313 25292 9369 25348
rect 9394 25292 9450 25348
rect 9475 25292 9531 25348
rect 9556 25292 9612 25348
rect 9637 25292 9693 25348
rect 9718 25292 9774 25348
rect 9799 25292 9855 25348
rect 9880 25292 9936 25348
rect 9961 25292 10017 25348
rect 10042 25292 10098 25348
rect 10123 25292 10179 25348
rect 10204 25292 10260 25348
rect 10285 25292 10341 25348
rect 10366 25292 10422 25348
rect 10447 25292 10503 25348
rect 10528 25292 10584 25348
rect 10609 25292 10665 25348
rect 10690 25292 10746 25348
rect 10771 25292 10827 25348
rect 10852 25292 10908 25348
rect 10933 25292 10989 25348
rect 11014 25292 11070 25348
rect 11095 25292 11151 25348
rect 11176 25292 11232 25348
rect 11257 25292 11313 25348
rect 11338 25292 11394 25348
rect 11419 25292 11475 25348
rect 2170 25197 2226 25253
rect 2252 25197 2308 25253
rect 2334 25197 2390 25253
rect 2416 25197 2472 25253
rect 5425 25212 5481 25268
rect 5506 25212 5562 25268
rect 5587 25212 5643 25268
rect 5668 25212 5724 25268
rect 5749 25212 5805 25268
rect 5830 25212 5886 25268
rect 5911 25212 5967 25268
rect 5992 25212 6048 25268
rect 6073 25212 6129 25268
rect 6154 25212 6210 25268
rect 6235 25212 6291 25268
rect 6316 25212 6372 25268
rect 6397 25212 6453 25268
rect 6478 25212 6534 25268
rect 6559 25212 6615 25268
rect 6640 25212 6696 25268
rect 6721 25212 6777 25268
rect 6802 25212 6858 25268
rect 6883 25212 6939 25268
rect 6964 25212 7020 25268
rect 7045 25212 7101 25268
rect 7126 25212 7182 25268
rect 7207 25212 7263 25268
rect 7288 25212 7344 25268
rect 7369 25212 7425 25268
rect 7450 25212 7506 25268
rect 7531 25212 7587 25268
rect 7612 25212 7668 25268
rect 7693 25212 7749 25268
rect 7774 25212 7830 25268
rect 7855 25212 7911 25268
rect 7936 25212 7992 25268
rect 8017 25212 8073 25268
rect 8098 25212 8154 25268
rect 8179 25212 8235 25268
rect 8260 25212 8316 25268
rect 8341 25212 8397 25268
rect 8422 25212 8478 25268
rect 8503 25212 8559 25268
rect 8584 25212 8640 25268
rect 8665 25212 8721 25268
rect 8746 25212 8802 25268
rect 8827 25212 8883 25268
rect 8908 25212 8964 25268
rect 8989 25212 9045 25268
rect 9070 25212 9126 25268
rect 9151 25212 9207 25268
rect 9232 25212 9288 25268
rect 9313 25212 9369 25268
rect 9394 25212 9450 25268
rect 9475 25212 9531 25268
rect 9556 25212 9612 25268
rect 9637 25212 9693 25268
rect 9718 25212 9774 25268
rect 9799 25212 9855 25268
rect 9880 25212 9936 25268
rect 9961 25212 10017 25268
rect 10042 25212 10098 25268
rect 10123 25212 10179 25268
rect 10204 25212 10260 25268
rect 10285 25212 10341 25268
rect 10366 25212 10422 25268
rect 10447 25212 10503 25268
rect 10528 25212 10584 25268
rect 10609 25212 10665 25268
rect 10690 25212 10746 25268
rect 10771 25212 10827 25268
rect 10852 25212 10908 25268
rect 10933 25212 10989 25268
rect 11014 25212 11070 25268
rect 11095 25212 11151 25268
rect 11176 25212 11232 25268
rect 11257 25212 11313 25268
rect 11338 25212 11394 25268
rect 11419 25212 11475 25268
rect 2170 25116 2226 25172
rect 2252 25116 2308 25172
rect 2334 25116 2390 25172
rect 2416 25116 2472 25172
rect 5425 25132 5481 25188
rect 5506 25132 5562 25188
rect 5587 25132 5643 25188
rect 5668 25132 5724 25188
rect 5749 25132 5805 25188
rect 5830 25132 5886 25188
rect 5911 25132 5967 25188
rect 5992 25132 6048 25188
rect 6073 25132 6129 25188
rect 6154 25132 6210 25188
rect 6235 25132 6291 25188
rect 6316 25132 6372 25188
rect 6397 25132 6453 25188
rect 6478 25132 6534 25188
rect 6559 25132 6615 25188
rect 6640 25132 6696 25188
rect 6721 25132 6777 25188
rect 6802 25132 6858 25188
rect 6883 25132 6939 25188
rect 6964 25132 7020 25188
rect 7045 25132 7101 25188
rect 7126 25132 7182 25188
rect 7207 25132 7263 25188
rect 7288 25132 7344 25188
rect 7369 25132 7425 25188
rect 7450 25132 7506 25188
rect 7531 25132 7587 25188
rect 7612 25132 7668 25188
rect 7693 25132 7749 25188
rect 7774 25132 7830 25188
rect 7855 25132 7911 25188
rect 7936 25132 7992 25188
rect 8017 25132 8073 25188
rect 8098 25132 8154 25188
rect 8179 25132 8235 25188
rect 8260 25132 8316 25188
rect 8341 25132 8397 25188
rect 8422 25132 8478 25188
rect 8503 25132 8559 25188
rect 8584 25132 8640 25188
rect 8665 25132 8721 25188
rect 8746 25132 8802 25188
rect 8827 25132 8883 25188
rect 8908 25132 8964 25188
rect 8989 25132 9045 25188
rect 9070 25132 9126 25188
rect 9151 25132 9207 25188
rect 9232 25132 9288 25188
rect 9313 25132 9369 25188
rect 9394 25132 9450 25188
rect 9475 25132 9531 25188
rect 9556 25132 9612 25188
rect 9637 25132 9693 25188
rect 9718 25132 9774 25188
rect 9799 25132 9855 25188
rect 9880 25132 9936 25188
rect 9961 25132 10017 25188
rect 10042 25132 10098 25188
rect 10123 25132 10179 25188
rect 10204 25132 10260 25188
rect 10285 25132 10341 25188
rect 10366 25132 10422 25188
rect 10447 25132 10503 25188
rect 10528 25132 10584 25188
rect 10609 25132 10665 25188
rect 10690 25132 10746 25188
rect 10771 25132 10827 25188
rect 10852 25132 10908 25188
rect 10933 25132 10989 25188
rect 11014 25132 11070 25188
rect 11095 25132 11151 25188
rect 11176 25132 11232 25188
rect 11257 25132 11313 25188
rect 11338 25132 11394 25188
rect 11419 25132 11475 25188
rect 2170 25035 2226 25091
rect 2252 25035 2308 25091
rect 2334 25035 2390 25091
rect 2416 25035 2472 25091
rect 5425 25052 5481 25108
rect 5506 25052 5562 25108
rect 5587 25052 5643 25108
rect 5668 25052 5724 25108
rect 5749 25052 5805 25108
rect 5830 25052 5886 25108
rect 5911 25052 5967 25108
rect 5992 25052 6048 25108
rect 6073 25052 6129 25108
rect 6154 25052 6210 25108
rect 6235 25052 6291 25108
rect 6316 25052 6372 25108
rect 6397 25052 6453 25108
rect 6478 25052 6534 25108
rect 6559 25052 6615 25108
rect 6640 25052 6696 25108
rect 6721 25052 6777 25108
rect 6802 25052 6858 25108
rect 6883 25052 6939 25108
rect 6964 25052 7020 25108
rect 7045 25052 7101 25108
rect 7126 25052 7182 25108
rect 7207 25052 7263 25108
rect 7288 25052 7344 25108
rect 7369 25052 7425 25108
rect 7450 25052 7506 25108
rect 7531 25052 7587 25108
rect 7612 25052 7668 25108
rect 7693 25052 7749 25108
rect 7774 25052 7830 25108
rect 7855 25052 7911 25108
rect 7936 25052 7992 25108
rect 8017 25052 8073 25108
rect 8098 25052 8154 25108
rect 8179 25052 8235 25108
rect 8260 25052 8316 25108
rect 8341 25052 8397 25108
rect 8422 25052 8478 25108
rect 8503 25052 8559 25108
rect 8584 25052 8640 25108
rect 8665 25052 8721 25108
rect 8746 25052 8802 25108
rect 8827 25052 8883 25108
rect 8908 25052 8964 25108
rect 8989 25052 9045 25108
rect 9070 25052 9126 25108
rect 9151 25052 9207 25108
rect 9232 25052 9288 25108
rect 9313 25052 9369 25108
rect 9394 25052 9450 25108
rect 9475 25052 9531 25108
rect 9556 25052 9612 25108
rect 9637 25052 9693 25108
rect 9718 25052 9774 25108
rect 9799 25052 9855 25108
rect 9880 25052 9936 25108
rect 9961 25052 10017 25108
rect 10042 25052 10098 25108
rect 10123 25052 10179 25108
rect 10204 25052 10260 25108
rect 10285 25052 10341 25108
rect 10366 25052 10422 25108
rect 10447 25052 10503 25108
rect 10528 25052 10584 25108
rect 10609 25052 10665 25108
rect 10690 25052 10746 25108
rect 10771 25052 10827 25108
rect 10852 25052 10908 25108
rect 10933 25052 10989 25108
rect 11014 25052 11070 25108
rect 11095 25052 11151 25108
rect 11176 25052 11232 25108
rect 11257 25052 11313 25108
rect 11338 25052 11394 25108
rect 11419 25052 11475 25108
rect 2170 24954 2226 25010
rect 2252 24954 2308 25010
rect 2334 24954 2390 25010
rect 2416 24954 2472 25010
rect 5425 24972 5481 25028
rect 5506 24972 5562 25028
rect 5587 24972 5643 25028
rect 5668 24972 5724 25028
rect 5749 24972 5805 25028
rect 5830 24972 5886 25028
rect 5911 24972 5967 25028
rect 5992 24972 6048 25028
rect 6073 24972 6129 25028
rect 6154 24972 6210 25028
rect 6235 24972 6291 25028
rect 6316 24972 6372 25028
rect 6397 24972 6453 25028
rect 6478 24972 6534 25028
rect 6559 24972 6615 25028
rect 6640 24972 6696 25028
rect 6721 24972 6777 25028
rect 6802 24972 6858 25028
rect 6883 24972 6939 25028
rect 6964 24972 7020 25028
rect 7045 24972 7101 25028
rect 7126 24972 7182 25028
rect 7207 24972 7263 25028
rect 7288 24972 7344 25028
rect 7369 24972 7425 25028
rect 7450 24972 7506 25028
rect 7531 24972 7587 25028
rect 7612 24972 7668 25028
rect 7693 24972 7749 25028
rect 7774 24972 7830 25028
rect 7855 24972 7911 25028
rect 7936 24972 7992 25028
rect 8017 24972 8073 25028
rect 8098 24972 8154 25028
rect 8179 24972 8235 25028
rect 8260 24972 8316 25028
rect 8341 24972 8397 25028
rect 8422 24972 8478 25028
rect 8503 24972 8559 25028
rect 8584 24972 8640 25028
rect 8665 24972 8721 25028
rect 8746 24972 8802 25028
rect 8827 24972 8883 25028
rect 8908 24972 8964 25028
rect 8989 24972 9045 25028
rect 9070 24972 9126 25028
rect 9151 24972 9207 25028
rect 9232 24972 9288 25028
rect 9313 24972 9369 25028
rect 9394 24972 9450 25028
rect 9475 24972 9531 25028
rect 9556 24972 9612 25028
rect 9637 24972 9693 25028
rect 9718 24972 9774 25028
rect 9799 24972 9855 25028
rect 9880 24972 9936 25028
rect 9961 24972 10017 25028
rect 10042 24972 10098 25028
rect 10123 24972 10179 25028
rect 10204 24972 10260 25028
rect 10285 24972 10341 25028
rect 10366 24972 10422 25028
rect 10447 24972 10503 25028
rect 10528 24972 10584 25028
rect 10609 24972 10665 25028
rect 10690 24972 10746 25028
rect 10771 24972 10827 25028
rect 10852 24972 10908 25028
rect 10933 24972 10989 25028
rect 11014 24972 11070 25028
rect 11095 24972 11151 25028
rect 11176 24972 11232 25028
rect 11257 24972 11313 25028
rect 11338 24972 11394 25028
rect 11419 24972 11475 25028
rect 2170 24873 2226 24929
rect 2252 24873 2308 24929
rect 2334 24873 2390 24929
rect 2416 24873 2472 24929
rect 5425 24892 5481 24948
rect 5506 24892 5562 24948
rect 5587 24892 5643 24948
rect 5668 24892 5724 24948
rect 5749 24892 5805 24948
rect 5830 24892 5886 24948
rect 5911 24892 5967 24948
rect 5992 24892 6048 24948
rect 6073 24892 6129 24948
rect 6154 24892 6210 24948
rect 6235 24892 6291 24948
rect 6316 24892 6372 24948
rect 6397 24892 6453 24948
rect 6478 24892 6534 24948
rect 6559 24892 6615 24948
rect 6640 24892 6696 24948
rect 6721 24892 6777 24948
rect 6802 24892 6858 24948
rect 6883 24892 6939 24948
rect 6964 24892 7020 24948
rect 7045 24892 7101 24948
rect 7126 24892 7182 24948
rect 7207 24892 7263 24948
rect 7288 24892 7344 24948
rect 7369 24892 7425 24948
rect 7450 24892 7506 24948
rect 7531 24892 7587 24948
rect 7612 24892 7668 24948
rect 7693 24892 7749 24948
rect 7774 24892 7830 24948
rect 7855 24892 7911 24948
rect 7936 24892 7992 24948
rect 8017 24892 8073 24948
rect 8098 24892 8154 24948
rect 8179 24892 8235 24948
rect 8260 24892 8316 24948
rect 8341 24892 8397 24948
rect 8422 24892 8478 24948
rect 8503 24892 8559 24948
rect 8584 24892 8640 24948
rect 8665 24892 8721 24948
rect 8746 24892 8802 24948
rect 8827 24892 8883 24948
rect 8908 24892 8964 24948
rect 8989 24892 9045 24948
rect 9070 24892 9126 24948
rect 9151 24892 9207 24948
rect 9232 24892 9288 24948
rect 9313 24892 9369 24948
rect 9394 24892 9450 24948
rect 9475 24892 9531 24948
rect 9556 24892 9612 24948
rect 9637 24892 9693 24948
rect 9718 24892 9774 24948
rect 9799 24892 9855 24948
rect 9880 24892 9936 24948
rect 9961 24892 10017 24948
rect 10042 24892 10098 24948
rect 10123 24892 10179 24948
rect 10204 24892 10260 24948
rect 10285 24892 10341 24948
rect 10366 24892 10422 24948
rect 10447 24892 10503 24948
rect 10528 24892 10584 24948
rect 10609 24892 10665 24948
rect 10690 24892 10746 24948
rect 10771 24892 10827 24948
rect 10852 24892 10908 24948
rect 10933 24892 10989 24948
rect 11014 24892 11070 24948
rect 11095 24892 11151 24948
rect 11176 24892 11232 24948
rect 11257 24892 11313 24948
rect 11338 24892 11394 24948
rect 11419 24892 11475 24948
rect 2170 24792 2226 24848
rect 2252 24792 2308 24848
rect 2334 24792 2390 24848
rect 2416 24792 2472 24848
rect 5425 24812 5481 24868
rect 5506 24812 5562 24868
rect 5587 24812 5643 24868
rect 5668 24812 5724 24868
rect 5749 24812 5805 24868
rect 5830 24812 5886 24868
rect 5911 24812 5967 24868
rect 5992 24812 6048 24868
rect 6073 24812 6129 24868
rect 6154 24812 6210 24868
rect 6235 24812 6291 24868
rect 6316 24812 6372 24868
rect 6397 24812 6453 24868
rect 6478 24812 6534 24868
rect 6559 24812 6615 24868
rect 6640 24812 6696 24868
rect 6721 24812 6777 24868
rect 6802 24812 6858 24868
rect 6883 24812 6939 24868
rect 6964 24812 7020 24868
rect 7045 24812 7101 24868
rect 7126 24812 7182 24868
rect 7207 24812 7263 24868
rect 7288 24812 7344 24868
rect 7369 24812 7425 24868
rect 7450 24812 7506 24868
rect 7531 24812 7587 24868
rect 7612 24812 7668 24868
rect 7693 24812 7749 24868
rect 7774 24812 7830 24868
rect 7855 24812 7911 24868
rect 7936 24812 7992 24868
rect 8017 24812 8073 24868
rect 8098 24812 8154 24868
rect 8179 24812 8235 24868
rect 8260 24812 8316 24868
rect 8341 24812 8397 24868
rect 8422 24812 8478 24868
rect 8503 24812 8559 24868
rect 8584 24812 8640 24868
rect 8665 24812 8721 24868
rect 8746 24812 8802 24868
rect 8827 24812 8883 24868
rect 8908 24812 8964 24868
rect 8989 24812 9045 24868
rect 9070 24812 9126 24868
rect 9151 24812 9207 24868
rect 9232 24812 9288 24868
rect 9313 24812 9369 24868
rect 9394 24812 9450 24868
rect 9475 24812 9531 24868
rect 9556 24812 9612 24868
rect 9637 24812 9693 24868
rect 9718 24812 9774 24868
rect 9799 24812 9855 24868
rect 9880 24812 9936 24868
rect 9961 24812 10017 24868
rect 10042 24812 10098 24868
rect 10123 24812 10179 24868
rect 10204 24812 10260 24868
rect 10285 24812 10341 24868
rect 10366 24812 10422 24868
rect 10447 24812 10503 24868
rect 10528 24812 10584 24868
rect 10609 24812 10665 24868
rect 10690 24812 10746 24868
rect 10771 24812 10827 24868
rect 10852 24812 10908 24868
rect 10933 24812 10989 24868
rect 11014 24812 11070 24868
rect 11095 24812 11151 24868
rect 11176 24812 11232 24868
rect 11257 24812 11313 24868
rect 11338 24812 11394 24868
rect 11419 24812 11475 24868
rect 2170 24711 2226 24767
rect 2252 24711 2308 24767
rect 2334 24711 2390 24767
rect 2416 24711 2472 24767
rect 5425 24732 5481 24788
rect 5506 24732 5562 24788
rect 5587 24732 5643 24788
rect 5668 24732 5724 24788
rect 5749 24732 5805 24788
rect 5830 24732 5886 24788
rect 5911 24732 5967 24788
rect 5992 24732 6048 24788
rect 6073 24732 6129 24788
rect 6154 24732 6210 24788
rect 6235 24732 6291 24788
rect 6316 24732 6372 24788
rect 6397 24732 6453 24788
rect 6478 24732 6534 24788
rect 6559 24732 6615 24788
rect 6640 24732 6696 24788
rect 6721 24732 6777 24788
rect 6802 24732 6858 24788
rect 6883 24732 6939 24788
rect 6964 24732 7020 24788
rect 7045 24732 7101 24788
rect 7126 24732 7182 24788
rect 7207 24732 7263 24788
rect 7288 24732 7344 24788
rect 7369 24732 7425 24788
rect 7450 24732 7506 24788
rect 7531 24732 7587 24788
rect 7612 24732 7668 24788
rect 7693 24732 7749 24788
rect 7774 24732 7830 24788
rect 7855 24732 7911 24788
rect 7936 24732 7992 24788
rect 8017 24732 8073 24788
rect 8098 24732 8154 24788
rect 8179 24732 8235 24788
rect 8260 24732 8316 24788
rect 8341 24732 8397 24788
rect 8422 24732 8478 24788
rect 8503 24732 8559 24788
rect 8584 24732 8640 24788
rect 8665 24732 8721 24788
rect 8746 24732 8802 24788
rect 8827 24732 8883 24788
rect 8908 24732 8964 24788
rect 8989 24732 9045 24788
rect 9070 24732 9126 24788
rect 9151 24732 9207 24788
rect 9232 24732 9288 24788
rect 9313 24732 9369 24788
rect 9394 24732 9450 24788
rect 9475 24732 9531 24788
rect 9556 24732 9612 24788
rect 9637 24732 9693 24788
rect 9718 24732 9774 24788
rect 9799 24732 9855 24788
rect 9880 24732 9936 24788
rect 9961 24732 10017 24788
rect 10042 24732 10098 24788
rect 10123 24732 10179 24788
rect 10204 24732 10260 24788
rect 10285 24732 10341 24788
rect 10366 24732 10422 24788
rect 10447 24732 10503 24788
rect 10528 24732 10584 24788
rect 10609 24732 10665 24788
rect 10690 24732 10746 24788
rect 10771 24732 10827 24788
rect 10852 24732 10908 24788
rect 10933 24732 10989 24788
rect 11014 24732 11070 24788
rect 11095 24732 11151 24788
rect 11176 24732 11232 24788
rect 11257 24732 11313 24788
rect 11338 24732 11394 24788
rect 11419 24732 11475 24788
rect 2170 24630 2226 24686
rect 2252 24630 2308 24686
rect 2334 24630 2390 24686
rect 2416 24630 2472 24686
rect 5425 24652 5481 24708
rect 5506 24652 5562 24708
rect 5587 24652 5643 24708
rect 5668 24652 5724 24708
rect 5749 24652 5805 24708
rect 5830 24652 5886 24708
rect 5911 24652 5967 24708
rect 5992 24652 6048 24708
rect 6073 24652 6129 24708
rect 6154 24652 6210 24708
rect 6235 24652 6291 24708
rect 6316 24652 6372 24708
rect 6397 24652 6453 24708
rect 6478 24652 6534 24708
rect 6559 24652 6615 24708
rect 6640 24652 6696 24708
rect 6721 24652 6777 24708
rect 6802 24652 6858 24708
rect 6883 24652 6939 24708
rect 6964 24652 7020 24708
rect 7045 24652 7101 24708
rect 7126 24652 7182 24708
rect 7207 24652 7263 24708
rect 7288 24652 7344 24708
rect 7369 24652 7425 24708
rect 7450 24652 7506 24708
rect 7531 24652 7587 24708
rect 7612 24652 7668 24708
rect 7693 24652 7749 24708
rect 7774 24652 7830 24708
rect 7855 24652 7911 24708
rect 7936 24652 7992 24708
rect 8017 24652 8073 24708
rect 8098 24652 8154 24708
rect 8179 24652 8235 24708
rect 8260 24652 8316 24708
rect 8341 24652 8397 24708
rect 8422 24652 8478 24708
rect 8503 24652 8559 24708
rect 8584 24652 8640 24708
rect 8665 24652 8721 24708
rect 8746 24652 8802 24708
rect 8827 24652 8883 24708
rect 8908 24652 8964 24708
rect 8989 24652 9045 24708
rect 9070 24652 9126 24708
rect 9151 24652 9207 24708
rect 9232 24652 9288 24708
rect 9313 24652 9369 24708
rect 9394 24652 9450 24708
rect 9475 24652 9531 24708
rect 9556 24652 9612 24708
rect 9637 24652 9693 24708
rect 9718 24652 9774 24708
rect 9799 24652 9855 24708
rect 9880 24652 9936 24708
rect 9961 24652 10017 24708
rect 10042 24652 10098 24708
rect 10123 24652 10179 24708
rect 10204 24652 10260 24708
rect 10285 24652 10341 24708
rect 10366 24652 10422 24708
rect 10447 24652 10503 24708
rect 10528 24652 10584 24708
rect 10609 24652 10665 24708
rect 10690 24652 10746 24708
rect 10771 24652 10827 24708
rect 10852 24652 10908 24708
rect 10933 24652 10989 24708
rect 11014 24652 11070 24708
rect 11095 24652 11151 24708
rect 11176 24652 11232 24708
rect 11257 24652 11313 24708
rect 11338 24652 11394 24708
rect 11419 24652 11475 24708
rect 11500 24652 13076 25828
rect 14509 25766 14565 25822
rect 14603 25766 14659 25822
rect 14697 25766 14753 25822
rect 14791 25766 14847 25822
rect 14885 25766 14941 25822
rect 14979 25766 15035 25822
rect 14509 25685 14565 25741
rect 14603 25685 14659 25741
rect 14697 25685 14753 25741
rect 14791 25685 14847 25741
rect 14885 25685 14941 25741
rect 14979 25685 15035 25741
rect 14509 25604 14565 25660
rect 14603 25604 14659 25660
rect 14697 25604 14753 25660
rect 14791 25604 14847 25660
rect 14885 25604 14941 25660
rect 14979 25604 15035 25660
rect 14509 25523 14565 25579
rect 14603 25523 14659 25579
rect 14697 25523 14753 25579
rect 14791 25523 14847 25579
rect 14885 25523 14941 25579
rect 14979 25523 15035 25579
rect 14509 25442 14565 25498
rect 14603 25442 14659 25498
rect 14697 25442 14753 25498
rect 14791 25442 14847 25498
rect 14885 25442 14941 25498
rect 14979 25442 15035 25498
rect 14509 25361 14565 25417
rect 14603 25361 14659 25417
rect 14697 25361 14753 25417
rect 14791 25361 14847 25417
rect 14885 25361 14941 25417
rect 14979 25361 15035 25417
rect 14509 25280 14565 25336
rect 14603 25280 14659 25336
rect 14697 25280 14753 25336
rect 14791 25280 14847 25336
rect 14885 25280 14941 25336
rect 14979 25280 15035 25336
rect 14509 25199 14565 25255
rect 14603 25199 14659 25255
rect 14697 25199 14753 25255
rect 14791 25199 14847 25255
rect 14885 25199 14941 25255
rect 14979 25199 15035 25255
rect 14509 25118 14565 25174
rect 14603 25118 14659 25174
rect 14697 25118 14753 25174
rect 14791 25118 14847 25174
rect 14885 25118 14941 25174
rect 14979 25118 15035 25174
rect 14509 25037 14565 25093
rect 14603 25037 14659 25093
rect 14697 25037 14753 25093
rect 14791 25037 14847 25093
rect 14885 25037 14941 25093
rect 14979 25037 15035 25093
rect 14509 24955 14565 25011
rect 14603 24955 14659 25011
rect 14697 24955 14753 25011
rect 14791 24955 14847 25011
rect 14885 24955 14941 25011
rect 14979 24955 15035 25011
rect 14509 24873 14565 24929
rect 14603 24873 14659 24929
rect 14697 24873 14753 24929
rect 14791 24873 14847 24929
rect 14885 24873 14941 24929
rect 14979 24873 15035 24929
rect 14509 24791 14565 24847
rect 14603 24791 14659 24847
rect 14697 24791 14753 24847
rect 14791 24791 14847 24847
rect 14885 24791 14941 24847
rect 14979 24791 15035 24847
rect 14509 24709 14565 24765
rect 14603 24709 14659 24765
rect 14697 24709 14753 24765
rect 14791 24709 14847 24765
rect 14885 24709 14941 24765
rect 14979 24709 15035 24765
rect 14509 24627 14565 24683
rect 14603 24627 14659 24683
rect 14697 24627 14753 24683
rect 14791 24627 14847 24683
rect 14885 24627 14941 24683
rect 14979 24627 15035 24683
rect 2170 24548 2226 24604
rect 2252 24548 2308 24604
rect 2334 24548 2390 24604
rect 2416 24548 2472 24604
rect 14509 24545 14565 24601
rect 14603 24545 14659 24601
rect 14697 24545 14753 24601
rect 14791 24545 14847 24601
rect 14885 24545 14941 24601
rect 14979 24545 15035 24601
rect 2170 24466 2226 24522
rect 2252 24466 2308 24522
rect 2334 24466 2390 24522
rect 2416 24466 2472 24522
rect 14509 24463 14565 24519
rect 14603 24463 14659 24519
rect 14697 24463 14753 24519
rect 14791 24463 14847 24519
rect 14885 24463 14941 24519
rect 14979 24463 15035 24519
rect 2170 24384 2226 24440
rect 2252 24384 2308 24440
rect 2334 24384 2390 24440
rect 2416 24384 2472 24440
rect 14509 24381 14565 24437
rect 14603 24381 14659 24437
rect 14697 24381 14753 24437
rect 14791 24381 14847 24437
rect 14885 24381 14941 24437
rect 14979 24381 15035 24437
rect 2170 24302 2226 24358
rect 2252 24302 2308 24358
rect 2334 24302 2390 24358
rect 2416 24302 2472 24358
rect 2170 24220 2226 24276
rect 2252 24220 2308 24276
rect 2334 24220 2390 24276
rect 2416 24220 2472 24276
rect 5425 24267 5481 24323
rect 5506 24267 5562 24323
rect 5587 24267 5643 24323
rect 5668 24267 5724 24323
rect 5749 24267 5805 24323
rect 5830 24267 5886 24323
rect 5911 24267 5967 24323
rect 5992 24267 6048 24323
rect 6073 24267 6129 24323
rect 6154 24267 6210 24323
rect 6235 24267 6291 24323
rect 6316 24267 6372 24323
rect 6397 24267 6453 24323
rect 6478 24267 6534 24323
rect 6559 24267 6615 24323
rect 6640 24267 6696 24323
rect 6721 24267 6777 24323
rect 6802 24267 6858 24323
rect 6883 24267 6939 24323
rect 6964 24267 7020 24323
rect 7045 24267 7101 24323
rect 7126 24267 7182 24323
rect 7207 24267 7263 24323
rect 7288 24267 7344 24323
rect 7369 24267 7425 24323
rect 7450 24267 7506 24323
rect 7531 24267 7587 24323
rect 7612 24267 7668 24323
rect 7693 24267 7749 24323
rect 7774 24267 7830 24323
rect 7855 24267 7911 24323
rect 7936 24267 7992 24323
rect 8017 24267 8073 24323
rect 8098 24267 8154 24323
rect 8179 24267 8235 24323
rect 8260 24267 8316 24323
rect 8341 24267 8397 24323
rect 8422 24267 8478 24323
rect 8503 24267 8559 24323
rect 8584 24267 8640 24323
rect 8665 24267 8721 24323
rect 8746 24267 8802 24323
rect 8827 24267 8883 24323
rect 8908 24267 8964 24323
rect 8989 24267 9045 24323
rect 9070 24267 9126 24323
rect 9151 24267 9207 24323
rect 9232 24267 9288 24323
rect 9313 24267 9369 24323
rect 9394 24267 9450 24323
rect 9475 24267 9531 24323
rect 9556 24267 9612 24323
rect 9637 24267 9693 24323
rect 9718 24267 9774 24323
rect 9799 24267 9855 24323
rect 9880 24267 9936 24323
rect 9961 24267 10017 24323
rect 10042 24267 10098 24323
rect 10123 24267 10179 24323
rect 10204 24267 10260 24323
rect 10285 24267 10341 24323
rect 10366 24267 10422 24323
rect 10447 24267 10503 24323
rect 10528 24267 10584 24323
rect 10609 24267 10665 24323
rect 10690 24267 10746 24323
rect 10771 24267 10827 24323
rect 10852 24267 10908 24323
rect 10933 24267 10989 24323
rect 11014 24267 11070 24323
rect 11095 24267 11151 24323
rect 11176 24267 11232 24323
rect 11257 24267 11313 24323
rect 11338 24267 11394 24323
rect 11419 24267 11475 24323
rect 2170 24138 2226 24194
rect 2252 24138 2308 24194
rect 2334 24138 2390 24194
rect 2416 24138 2472 24194
rect 5425 24187 5481 24243
rect 5506 24187 5562 24243
rect 5587 24187 5643 24243
rect 5668 24187 5724 24243
rect 5749 24187 5805 24243
rect 5830 24187 5886 24243
rect 5911 24187 5967 24243
rect 5992 24187 6048 24243
rect 6073 24187 6129 24243
rect 6154 24187 6210 24243
rect 6235 24187 6291 24243
rect 6316 24187 6372 24243
rect 6397 24187 6453 24243
rect 6478 24187 6534 24243
rect 6559 24187 6615 24243
rect 6640 24187 6696 24243
rect 6721 24187 6777 24243
rect 6802 24187 6858 24243
rect 6883 24187 6939 24243
rect 6964 24187 7020 24243
rect 7045 24187 7101 24243
rect 7126 24187 7182 24243
rect 7207 24187 7263 24243
rect 7288 24187 7344 24243
rect 7369 24187 7425 24243
rect 7450 24187 7506 24243
rect 7531 24187 7587 24243
rect 7612 24187 7668 24243
rect 7693 24187 7749 24243
rect 7774 24187 7830 24243
rect 7855 24187 7911 24243
rect 7936 24187 7992 24243
rect 8017 24187 8073 24243
rect 8098 24187 8154 24243
rect 8179 24187 8235 24243
rect 8260 24187 8316 24243
rect 8341 24187 8397 24243
rect 8422 24187 8478 24243
rect 8503 24187 8559 24243
rect 8584 24187 8640 24243
rect 8665 24187 8721 24243
rect 8746 24187 8802 24243
rect 8827 24187 8883 24243
rect 8908 24187 8964 24243
rect 8989 24187 9045 24243
rect 9070 24187 9126 24243
rect 9151 24187 9207 24243
rect 9232 24187 9288 24243
rect 9313 24187 9369 24243
rect 9394 24187 9450 24243
rect 9475 24187 9531 24243
rect 9556 24187 9612 24243
rect 9637 24187 9693 24243
rect 9718 24187 9774 24243
rect 9799 24187 9855 24243
rect 9880 24187 9936 24243
rect 9961 24187 10017 24243
rect 10042 24187 10098 24243
rect 10123 24187 10179 24243
rect 10204 24187 10260 24243
rect 10285 24187 10341 24243
rect 10366 24187 10422 24243
rect 10447 24187 10503 24243
rect 10528 24187 10584 24243
rect 10609 24187 10665 24243
rect 10690 24187 10746 24243
rect 10771 24187 10827 24243
rect 10852 24187 10908 24243
rect 10933 24187 10989 24243
rect 11014 24187 11070 24243
rect 11095 24187 11151 24243
rect 11176 24187 11232 24243
rect 11257 24187 11313 24243
rect 11338 24187 11394 24243
rect 11419 24187 11475 24243
rect 2170 24056 2226 24112
rect 2252 24056 2308 24112
rect 2334 24056 2390 24112
rect 2416 24056 2472 24112
rect 5425 24107 5481 24163
rect 5506 24107 5562 24163
rect 5587 24107 5643 24163
rect 5668 24107 5724 24163
rect 5749 24107 5805 24163
rect 5830 24107 5886 24163
rect 5911 24107 5967 24163
rect 5992 24107 6048 24163
rect 6073 24107 6129 24163
rect 6154 24107 6210 24163
rect 6235 24107 6291 24163
rect 6316 24107 6372 24163
rect 6397 24107 6453 24163
rect 6478 24107 6534 24163
rect 6559 24107 6615 24163
rect 6640 24107 6696 24163
rect 6721 24107 6777 24163
rect 6802 24107 6858 24163
rect 6883 24107 6939 24163
rect 6964 24107 7020 24163
rect 7045 24107 7101 24163
rect 7126 24107 7182 24163
rect 7207 24107 7263 24163
rect 7288 24107 7344 24163
rect 7369 24107 7425 24163
rect 7450 24107 7506 24163
rect 7531 24107 7587 24163
rect 7612 24107 7668 24163
rect 7693 24107 7749 24163
rect 7774 24107 7830 24163
rect 7855 24107 7911 24163
rect 7936 24107 7992 24163
rect 8017 24107 8073 24163
rect 8098 24107 8154 24163
rect 8179 24107 8235 24163
rect 8260 24107 8316 24163
rect 8341 24107 8397 24163
rect 8422 24107 8478 24163
rect 8503 24107 8559 24163
rect 8584 24107 8640 24163
rect 8665 24107 8721 24163
rect 8746 24107 8802 24163
rect 8827 24107 8883 24163
rect 8908 24107 8964 24163
rect 8989 24107 9045 24163
rect 9070 24107 9126 24163
rect 9151 24107 9207 24163
rect 9232 24107 9288 24163
rect 9313 24107 9369 24163
rect 9394 24107 9450 24163
rect 9475 24107 9531 24163
rect 9556 24107 9612 24163
rect 9637 24107 9693 24163
rect 9718 24107 9774 24163
rect 9799 24107 9855 24163
rect 9880 24107 9936 24163
rect 9961 24107 10017 24163
rect 10042 24107 10098 24163
rect 10123 24107 10179 24163
rect 10204 24107 10260 24163
rect 10285 24107 10341 24163
rect 10366 24107 10422 24163
rect 10447 24107 10503 24163
rect 10528 24107 10584 24163
rect 10609 24107 10665 24163
rect 10690 24107 10746 24163
rect 10771 24107 10827 24163
rect 10852 24107 10908 24163
rect 10933 24107 10989 24163
rect 11014 24107 11070 24163
rect 11095 24107 11151 24163
rect 11176 24107 11232 24163
rect 11257 24107 11313 24163
rect 11338 24107 11394 24163
rect 11419 24107 11475 24163
rect 2170 23974 2226 24030
rect 2252 23974 2308 24030
rect 2334 23974 2390 24030
rect 2416 23974 2472 24030
rect 5425 24027 5481 24083
rect 5506 24027 5562 24083
rect 5587 24027 5643 24083
rect 5668 24027 5724 24083
rect 5749 24027 5805 24083
rect 5830 24027 5886 24083
rect 5911 24027 5967 24083
rect 5992 24027 6048 24083
rect 6073 24027 6129 24083
rect 6154 24027 6210 24083
rect 6235 24027 6291 24083
rect 6316 24027 6372 24083
rect 6397 24027 6453 24083
rect 6478 24027 6534 24083
rect 6559 24027 6615 24083
rect 6640 24027 6696 24083
rect 6721 24027 6777 24083
rect 6802 24027 6858 24083
rect 6883 24027 6939 24083
rect 6964 24027 7020 24083
rect 7045 24027 7101 24083
rect 7126 24027 7182 24083
rect 7207 24027 7263 24083
rect 7288 24027 7344 24083
rect 7369 24027 7425 24083
rect 7450 24027 7506 24083
rect 7531 24027 7587 24083
rect 7612 24027 7668 24083
rect 7693 24027 7749 24083
rect 7774 24027 7830 24083
rect 7855 24027 7911 24083
rect 7936 24027 7992 24083
rect 8017 24027 8073 24083
rect 8098 24027 8154 24083
rect 8179 24027 8235 24083
rect 8260 24027 8316 24083
rect 8341 24027 8397 24083
rect 8422 24027 8478 24083
rect 8503 24027 8559 24083
rect 8584 24027 8640 24083
rect 8665 24027 8721 24083
rect 8746 24027 8802 24083
rect 8827 24027 8883 24083
rect 8908 24027 8964 24083
rect 8989 24027 9045 24083
rect 9070 24027 9126 24083
rect 9151 24027 9207 24083
rect 9232 24027 9288 24083
rect 9313 24027 9369 24083
rect 9394 24027 9450 24083
rect 9475 24027 9531 24083
rect 9556 24027 9612 24083
rect 9637 24027 9693 24083
rect 9718 24027 9774 24083
rect 9799 24027 9855 24083
rect 9880 24027 9936 24083
rect 9961 24027 10017 24083
rect 10042 24027 10098 24083
rect 10123 24027 10179 24083
rect 10204 24027 10260 24083
rect 10285 24027 10341 24083
rect 10366 24027 10422 24083
rect 10447 24027 10503 24083
rect 10528 24027 10584 24083
rect 10609 24027 10665 24083
rect 10690 24027 10746 24083
rect 10771 24027 10827 24083
rect 10852 24027 10908 24083
rect 10933 24027 10989 24083
rect 11014 24027 11070 24083
rect 11095 24027 11151 24083
rect 11176 24027 11232 24083
rect 11257 24027 11313 24083
rect 11338 24027 11394 24083
rect 11419 24027 11475 24083
rect 2170 23892 2226 23948
rect 2252 23892 2308 23948
rect 2334 23892 2390 23948
rect 2416 23892 2472 23948
rect 5425 23947 5481 24003
rect 5506 23947 5562 24003
rect 5587 23947 5643 24003
rect 5668 23947 5724 24003
rect 5749 23947 5805 24003
rect 5830 23947 5886 24003
rect 5911 23947 5967 24003
rect 5992 23947 6048 24003
rect 6073 23947 6129 24003
rect 6154 23947 6210 24003
rect 6235 23947 6291 24003
rect 6316 23947 6372 24003
rect 6397 23947 6453 24003
rect 6478 23947 6534 24003
rect 6559 23947 6615 24003
rect 6640 23947 6696 24003
rect 6721 23947 6777 24003
rect 6802 23947 6858 24003
rect 6883 23947 6939 24003
rect 6964 23947 7020 24003
rect 7045 23947 7101 24003
rect 7126 23947 7182 24003
rect 7207 23947 7263 24003
rect 7288 23947 7344 24003
rect 7369 23947 7425 24003
rect 7450 23947 7506 24003
rect 7531 23947 7587 24003
rect 7612 23947 7668 24003
rect 7693 23947 7749 24003
rect 7774 23947 7830 24003
rect 7855 23947 7911 24003
rect 7936 23947 7992 24003
rect 8017 23947 8073 24003
rect 8098 23947 8154 24003
rect 8179 23947 8235 24003
rect 8260 23947 8316 24003
rect 8341 23947 8397 24003
rect 8422 23947 8478 24003
rect 8503 23947 8559 24003
rect 8584 23947 8640 24003
rect 8665 23947 8721 24003
rect 8746 23947 8802 24003
rect 8827 23947 8883 24003
rect 8908 23947 8964 24003
rect 8989 23947 9045 24003
rect 9070 23947 9126 24003
rect 9151 23947 9207 24003
rect 9232 23947 9288 24003
rect 9313 23947 9369 24003
rect 9394 23947 9450 24003
rect 9475 23947 9531 24003
rect 9556 23947 9612 24003
rect 9637 23947 9693 24003
rect 9718 23947 9774 24003
rect 9799 23947 9855 24003
rect 9880 23947 9936 24003
rect 9961 23947 10017 24003
rect 10042 23947 10098 24003
rect 10123 23947 10179 24003
rect 10204 23947 10260 24003
rect 10285 23947 10341 24003
rect 10366 23947 10422 24003
rect 10447 23947 10503 24003
rect 10528 23947 10584 24003
rect 10609 23947 10665 24003
rect 10690 23947 10746 24003
rect 10771 23947 10827 24003
rect 10852 23947 10908 24003
rect 10933 23947 10989 24003
rect 11014 23947 11070 24003
rect 11095 23947 11151 24003
rect 11176 23947 11232 24003
rect 11257 23947 11313 24003
rect 11338 23947 11394 24003
rect 11419 23947 11475 24003
rect 5425 23867 5481 23923
rect 5506 23867 5562 23923
rect 5587 23867 5643 23923
rect 5668 23867 5724 23923
rect 5749 23867 5805 23923
rect 5830 23867 5886 23923
rect 5911 23867 5967 23923
rect 5992 23867 6048 23923
rect 6073 23867 6129 23923
rect 6154 23867 6210 23923
rect 6235 23867 6291 23923
rect 6316 23867 6372 23923
rect 6397 23867 6453 23923
rect 6478 23867 6534 23923
rect 6559 23867 6615 23923
rect 6640 23867 6696 23923
rect 6721 23867 6777 23923
rect 6802 23867 6858 23923
rect 6883 23867 6939 23923
rect 6964 23867 7020 23923
rect 7045 23867 7101 23923
rect 7126 23867 7182 23923
rect 7207 23867 7263 23923
rect 7288 23867 7344 23923
rect 7369 23867 7425 23923
rect 7450 23867 7506 23923
rect 7531 23867 7587 23923
rect 7612 23867 7668 23923
rect 7693 23867 7749 23923
rect 7774 23867 7830 23923
rect 7855 23867 7911 23923
rect 7936 23867 7992 23923
rect 8017 23867 8073 23923
rect 8098 23867 8154 23923
rect 8179 23867 8235 23923
rect 8260 23867 8316 23923
rect 8341 23867 8397 23923
rect 8422 23867 8478 23923
rect 8503 23867 8559 23923
rect 8584 23867 8640 23923
rect 8665 23867 8721 23923
rect 8746 23867 8802 23923
rect 8827 23867 8883 23923
rect 8908 23867 8964 23923
rect 8989 23867 9045 23923
rect 9070 23867 9126 23923
rect 9151 23867 9207 23923
rect 9232 23867 9288 23923
rect 9313 23867 9369 23923
rect 9394 23867 9450 23923
rect 9475 23867 9531 23923
rect 9556 23867 9612 23923
rect 9637 23867 9693 23923
rect 9718 23867 9774 23923
rect 9799 23867 9855 23923
rect 9880 23867 9936 23923
rect 9961 23867 10017 23923
rect 10042 23867 10098 23923
rect 10123 23867 10179 23923
rect 10204 23867 10260 23923
rect 10285 23867 10341 23923
rect 10366 23867 10422 23923
rect 10447 23867 10503 23923
rect 10528 23867 10584 23923
rect 10609 23867 10665 23923
rect 10690 23867 10746 23923
rect 10771 23867 10827 23923
rect 10852 23867 10908 23923
rect 10933 23867 10989 23923
rect 11014 23867 11070 23923
rect 11095 23867 11151 23923
rect 11176 23867 11232 23923
rect 11257 23867 11313 23923
rect 11338 23867 11394 23923
rect 11419 23867 11475 23923
rect 2170 23810 2226 23866
rect 2252 23810 2308 23866
rect 2334 23810 2390 23866
rect 2416 23810 2472 23866
rect 5425 23787 5481 23843
rect 5506 23787 5562 23843
rect 5587 23787 5643 23843
rect 5668 23787 5724 23843
rect 5749 23787 5805 23843
rect 5830 23787 5886 23843
rect 5911 23787 5967 23843
rect 5992 23787 6048 23843
rect 6073 23787 6129 23843
rect 6154 23787 6210 23843
rect 6235 23787 6291 23843
rect 6316 23787 6372 23843
rect 6397 23787 6453 23843
rect 6478 23787 6534 23843
rect 6559 23787 6615 23843
rect 6640 23787 6696 23843
rect 6721 23787 6777 23843
rect 6802 23787 6858 23843
rect 6883 23787 6939 23843
rect 6964 23787 7020 23843
rect 7045 23787 7101 23843
rect 7126 23787 7182 23843
rect 7207 23787 7263 23843
rect 7288 23787 7344 23843
rect 7369 23787 7425 23843
rect 7450 23787 7506 23843
rect 7531 23787 7587 23843
rect 7612 23787 7668 23843
rect 7693 23787 7749 23843
rect 7774 23787 7830 23843
rect 7855 23787 7911 23843
rect 7936 23787 7992 23843
rect 8017 23787 8073 23843
rect 8098 23787 8154 23843
rect 8179 23787 8235 23843
rect 8260 23787 8316 23843
rect 8341 23787 8397 23843
rect 8422 23787 8478 23843
rect 8503 23787 8559 23843
rect 8584 23787 8640 23843
rect 8665 23787 8721 23843
rect 8746 23787 8802 23843
rect 8827 23787 8883 23843
rect 8908 23787 8964 23843
rect 8989 23787 9045 23843
rect 9070 23787 9126 23843
rect 9151 23787 9207 23843
rect 9232 23787 9288 23843
rect 9313 23787 9369 23843
rect 9394 23787 9450 23843
rect 9475 23787 9531 23843
rect 9556 23787 9612 23843
rect 9637 23787 9693 23843
rect 9718 23787 9774 23843
rect 9799 23787 9855 23843
rect 9880 23787 9936 23843
rect 9961 23787 10017 23843
rect 10042 23787 10098 23843
rect 10123 23787 10179 23843
rect 10204 23787 10260 23843
rect 10285 23787 10341 23843
rect 10366 23787 10422 23843
rect 10447 23787 10503 23843
rect 10528 23787 10584 23843
rect 10609 23787 10665 23843
rect 10690 23787 10746 23843
rect 10771 23787 10827 23843
rect 10852 23787 10908 23843
rect 10933 23787 10989 23843
rect 11014 23787 11070 23843
rect 11095 23787 11151 23843
rect 11176 23787 11232 23843
rect 11257 23787 11313 23843
rect 11338 23787 11394 23843
rect 11419 23787 11475 23843
rect 2170 23728 2226 23784
rect 2252 23728 2308 23784
rect 2334 23728 2390 23784
rect 2416 23728 2472 23784
rect 5425 23707 5481 23763
rect 5506 23707 5562 23763
rect 5587 23707 5643 23763
rect 5668 23707 5724 23763
rect 5749 23707 5805 23763
rect 5830 23707 5886 23763
rect 5911 23707 5967 23763
rect 5992 23707 6048 23763
rect 6073 23707 6129 23763
rect 6154 23707 6210 23763
rect 6235 23707 6291 23763
rect 6316 23707 6372 23763
rect 6397 23707 6453 23763
rect 6478 23707 6534 23763
rect 6559 23707 6615 23763
rect 6640 23707 6696 23763
rect 6721 23707 6777 23763
rect 6802 23707 6858 23763
rect 6883 23707 6939 23763
rect 6964 23707 7020 23763
rect 7045 23707 7101 23763
rect 7126 23707 7182 23763
rect 7207 23707 7263 23763
rect 7288 23707 7344 23763
rect 7369 23707 7425 23763
rect 7450 23707 7506 23763
rect 7531 23707 7587 23763
rect 7612 23707 7668 23763
rect 7693 23707 7749 23763
rect 7774 23707 7830 23763
rect 7855 23707 7911 23763
rect 7936 23707 7992 23763
rect 8017 23707 8073 23763
rect 8098 23707 8154 23763
rect 8179 23707 8235 23763
rect 8260 23707 8316 23763
rect 8341 23707 8397 23763
rect 8422 23707 8478 23763
rect 8503 23707 8559 23763
rect 8584 23707 8640 23763
rect 8665 23707 8721 23763
rect 8746 23707 8802 23763
rect 8827 23707 8883 23763
rect 8908 23707 8964 23763
rect 8989 23707 9045 23763
rect 9070 23707 9126 23763
rect 9151 23707 9207 23763
rect 9232 23707 9288 23763
rect 9313 23707 9369 23763
rect 9394 23707 9450 23763
rect 9475 23707 9531 23763
rect 9556 23707 9612 23763
rect 9637 23707 9693 23763
rect 9718 23707 9774 23763
rect 9799 23707 9855 23763
rect 9880 23707 9936 23763
rect 9961 23707 10017 23763
rect 10042 23707 10098 23763
rect 10123 23707 10179 23763
rect 10204 23707 10260 23763
rect 10285 23707 10341 23763
rect 10366 23707 10422 23763
rect 10447 23707 10503 23763
rect 10528 23707 10584 23763
rect 10609 23707 10665 23763
rect 10690 23707 10746 23763
rect 10771 23707 10827 23763
rect 10852 23707 10908 23763
rect 10933 23707 10989 23763
rect 11014 23707 11070 23763
rect 11095 23707 11151 23763
rect 11176 23707 11232 23763
rect 11257 23707 11313 23763
rect 11338 23707 11394 23763
rect 11419 23707 11475 23763
rect 2170 23646 2226 23702
rect 2252 23646 2308 23702
rect 2334 23646 2390 23702
rect 2416 23646 2472 23702
rect 5425 23627 5481 23683
rect 5506 23627 5562 23683
rect 5587 23627 5643 23683
rect 5668 23627 5724 23683
rect 5749 23627 5805 23683
rect 5830 23627 5886 23683
rect 5911 23627 5967 23683
rect 5992 23627 6048 23683
rect 6073 23627 6129 23683
rect 6154 23627 6210 23683
rect 6235 23627 6291 23683
rect 6316 23627 6372 23683
rect 6397 23627 6453 23683
rect 6478 23627 6534 23683
rect 6559 23627 6615 23683
rect 6640 23627 6696 23683
rect 6721 23627 6777 23683
rect 6802 23627 6858 23683
rect 6883 23627 6939 23683
rect 6964 23627 7020 23683
rect 7045 23627 7101 23683
rect 7126 23627 7182 23683
rect 7207 23627 7263 23683
rect 7288 23627 7344 23683
rect 7369 23627 7425 23683
rect 7450 23627 7506 23683
rect 7531 23627 7587 23683
rect 7612 23627 7668 23683
rect 7693 23627 7749 23683
rect 7774 23627 7830 23683
rect 7855 23627 7911 23683
rect 7936 23627 7992 23683
rect 8017 23627 8073 23683
rect 8098 23627 8154 23683
rect 8179 23627 8235 23683
rect 8260 23627 8316 23683
rect 8341 23627 8397 23683
rect 8422 23627 8478 23683
rect 8503 23627 8559 23683
rect 8584 23627 8640 23683
rect 8665 23627 8721 23683
rect 8746 23627 8802 23683
rect 8827 23627 8883 23683
rect 8908 23627 8964 23683
rect 8989 23627 9045 23683
rect 9070 23627 9126 23683
rect 9151 23627 9207 23683
rect 9232 23627 9288 23683
rect 9313 23627 9369 23683
rect 9394 23627 9450 23683
rect 9475 23627 9531 23683
rect 9556 23627 9612 23683
rect 9637 23627 9693 23683
rect 9718 23627 9774 23683
rect 9799 23627 9855 23683
rect 9880 23627 9936 23683
rect 9961 23627 10017 23683
rect 10042 23627 10098 23683
rect 10123 23627 10179 23683
rect 10204 23627 10260 23683
rect 10285 23627 10341 23683
rect 10366 23627 10422 23683
rect 10447 23627 10503 23683
rect 10528 23627 10584 23683
rect 10609 23627 10665 23683
rect 10690 23627 10746 23683
rect 10771 23627 10827 23683
rect 10852 23627 10908 23683
rect 10933 23627 10989 23683
rect 11014 23627 11070 23683
rect 11095 23627 11151 23683
rect 11176 23627 11232 23683
rect 11257 23627 11313 23683
rect 11338 23627 11394 23683
rect 11419 23627 11475 23683
rect 2170 23564 2226 23620
rect 2252 23564 2308 23620
rect 2334 23564 2390 23620
rect 2416 23564 2472 23620
rect 5425 23547 5481 23603
rect 5506 23547 5562 23603
rect 5587 23547 5643 23603
rect 5668 23547 5724 23603
rect 5749 23547 5805 23603
rect 5830 23547 5886 23603
rect 5911 23547 5967 23603
rect 5992 23547 6048 23603
rect 6073 23547 6129 23603
rect 6154 23547 6210 23603
rect 6235 23547 6291 23603
rect 6316 23547 6372 23603
rect 6397 23547 6453 23603
rect 6478 23547 6534 23603
rect 6559 23547 6615 23603
rect 6640 23547 6696 23603
rect 6721 23547 6777 23603
rect 6802 23547 6858 23603
rect 6883 23547 6939 23603
rect 6964 23547 7020 23603
rect 7045 23547 7101 23603
rect 7126 23547 7182 23603
rect 7207 23547 7263 23603
rect 7288 23547 7344 23603
rect 7369 23547 7425 23603
rect 7450 23547 7506 23603
rect 7531 23547 7587 23603
rect 7612 23547 7668 23603
rect 7693 23547 7749 23603
rect 7774 23547 7830 23603
rect 7855 23547 7911 23603
rect 7936 23547 7992 23603
rect 8017 23547 8073 23603
rect 8098 23547 8154 23603
rect 8179 23547 8235 23603
rect 8260 23547 8316 23603
rect 8341 23547 8397 23603
rect 8422 23547 8478 23603
rect 8503 23547 8559 23603
rect 8584 23547 8640 23603
rect 8665 23547 8721 23603
rect 8746 23547 8802 23603
rect 8827 23547 8883 23603
rect 8908 23547 8964 23603
rect 8989 23547 9045 23603
rect 9070 23547 9126 23603
rect 9151 23547 9207 23603
rect 9232 23547 9288 23603
rect 9313 23547 9369 23603
rect 9394 23547 9450 23603
rect 9475 23547 9531 23603
rect 9556 23547 9612 23603
rect 9637 23547 9693 23603
rect 9718 23547 9774 23603
rect 9799 23547 9855 23603
rect 9880 23547 9936 23603
rect 9961 23547 10017 23603
rect 10042 23547 10098 23603
rect 10123 23547 10179 23603
rect 10204 23547 10260 23603
rect 10285 23547 10341 23603
rect 10366 23547 10422 23603
rect 10447 23547 10503 23603
rect 10528 23547 10584 23603
rect 10609 23547 10665 23603
rect 10690 23547 10746 23603
rect 10771 23547 10827 23603
rect 10852 23547 10908 23603
rect 10933 23547 10989 23603
rect 11014 23547 11070 23603
rect 11095 23547 11151 23603
rect 11176 23547 11232 23603
rect 11257 23547 11313 23603
rect 11338 23547 11394 23603
rect 11419 23547 11475 23603
rect 2170 23482 2226 23538
rect 2252 23482 2308 23538
rect 2334 23482 2390 23538
rect 2416 23482 2472 23538
rect 5425 23467 5481 23523
rect 5506 23467 5562 23523
rect 5587 23467 5643 23523
rect 5668 23467 5724 23523
rect 5749 23467 5805 23523
rect 5830 23467 5886 23523
rect 5911 23467 5967 23523
rect 5992 23467 6048 23523
rect 6073 23467 6129 23523
rect 6154 23467 6210 23523
rect 6235 23467 6291 23523
rect 6316 23467 6372 23523
rect 6397 23467 6453 23523
rect 6478 23467 6534 23523
rect 6559 23467 6615 23523
rect 6640 23467 6696 23523
rect 6721 23467 6777 23523
rect 6802 23467 6858 23523
rect 6883 23467 6939 23523
rect 6964 23467 7020 23523
rect 7045 23467 7101 23523
rect 7126 23467 7182 23523
rect 7207 23467 7263 23523
rect 7288 23467 7344 23523
rect 7369 23467 7425 23523
rect 7450 23467 7506 23523
rect 7531 23467 7587 23523
rect 7612 23467 7668 23523
rect 7693 23467 7749 23523
rect 7774 23467 7830 23523
rect 7855 23467 7911 23523
rect 7936 23467 7992 23523
rect 8017 23467 8073 23523
rect 8098 23467 8154 23523
rect 8179 23467 8235 23523
rect 8260 23467 8316 23523
rect 8341 23467 8397 23523
rect 8422 23467 8478 23523
rect 8503 23467 8559 23523
rect 8584 23467 8640 23523
rect 8665 23467 8721 23523
rect 8746 23467 8802 23523
rect 8827 23467 8883 23523
rect 8908 23467 8964 23523
rect 8989 23467 9045 23523
rect 9070 23467 9126 23523
rect 9151 23467 9207 23523
rect 9232 23467 9288 23523
rect 9313 23467 9369 23523
rect 9394 23467 9450 23523
rect 9475 23467 9531 23523
rect 9556 23467 9612 23523
rect 9637 23467 9693 23523
rect 9718 23467 9774 23523
rect 9799 23467 9855 23523
rect 9880 23467 9936 23523
rect 9961 23467 10017 23523
rect 10042 23467 10098 23523
rect 10123 23467 10179 23523
rect 10204 23467 10260 23523
rect 10285 23467 10341 23523
rect 10366 23467 10422 23523
rect 10447 23467 10503 23523
rect 10528 23467 10584 23523
rect 10609 23467 10665 23523
rect 10690 23467 10746 23523
rect 10771 23467 10827 23523
rect 10852 23467 10908 23523
rect 10933 23467 10989 23523
rect 11014 23467 11070 23523
rect 11095 23467 11151 23523
rect 11176 23467 11232 23523
rect 11257 23467 11313 23523
rect 11338 23467 11394 23523
rect 11419 23467 11475 23523
rect 2170 23400 2226 23456
rect 2252 23400 2308 23456
rect 2334 23400 2390 23456
rect 2416 23400 2472 23456
rect 5425 23387 5481 23443
rect 5506 23387 5562 23443
rect 5587 23387 5643 23443
rect 5668 23387 5724 23443
rect 5749 23387 5805 23443
rect 5830 23387 5886 23443
rect 5911 23387 5967 23443
rect 5992 23387 6048 23443
rect 6073 23387 6129 23443
rect 6154 23387 6210 23443
rect 6235 23387 6291 23443
rect 6316 23387 6372 23443
rect 6397 23387 6453 23443
rect 6478 23387 6534 23443
rect 6559 23387 6615 23443
rect 6640 23387 6696 23443
rect 6721 23387 6777 23443
rect 6802 23387 6858 23443
rect 6883 23387 6939 23443
rect 6964 23387 7020 23443
rect 7045 23387 7101 23443
rect 7126 23387 7182 23443
rect 7207 23387 7263 23443
rect 7288 23387 7344 23443
rect 7369 23387 7425 23443
rect 7450 23387 7506 23443
rect 7531 23387 7587 23443
rect 7612 23387 7668 23443
rect 7693 23387 7749 23443
rect 7774 23387 7830 23443
rect 7855 23387 7911 23443
rect 7936 23387 7992 23443
rect 8017 23387 8073 23443
rect 8098 23387 8154 23443
rect 8179 23387 8235 23443
rect 8260 23387 8316 23443
rect 8341 23387 8397 23443
rect 8422 23387 8478 23443
rect 8503 23387 8559 23443
rect 8584 23387 8640 23443
rect 8665 23387 8721 23443
rect 8746 23387 8802 23443
rect 8827 23387 8883 23443
rect 8908 23387 8964 23443
rect 8989 23387 9045 23443
rect 9070 23387 9126 23443
rect 9151 23387 9207 23443
rect 9232 23387 9288 23443
rect 9313 23387 9369 23443
rect 9394 23387 9450 23443
rect 9475 23387 9531 23443
rect 9556 23387 9612 23443
rect 9637 23387 9693 23443
rect 9718 23387 9774 23443
rect 9799 23387 9855 23443
rect 9880 23387 9936 23443
rect 9961 23387 10017 23443
rect 10042 23387 10098 23443
rect 10123 23387 10179 23443
rect 10204 23387 10260 23443
rect 10285 23387 10341 23443
rect 10366 23387 10422 23443
rect 10447 23387 10503 23443
rect 10528 23387 10584 23443
rect 10609 23387 10665 23443
rect 10690 23387 10746 23443
rect 10771 23387 10827 23443
rect 10852 23387 10908 23443
rect 10933 23387 10989 23443
rect 11014 23387 11070 23443
rect 11095 23387 11151 23443
rect 11176 23387 11232 23443
rect 11257 23387 11313 23443
rect 11338 23387 11394 23443
rect 11419 23387 11475 23443
rect 2170 23318 2226 23374
rect 2252 23318 2308 23374
rect 2334 23318 2390 23374
rect 2416 23318 2472 23374
rect 5425 23307 5481 23363
rect 5506 23307 5562 23363
rect 5587 23307 5643 23363
rect 5668 23307 5724 23363
rect 5749 23307 5805 23363
rect 5830 23307 5886 23363
rect 5911 23307 5967 23363
rect 5992 23307 6048 23363
rect 6073 23307 6129 23363
rect 6154 23307 6210 23363
rect 6235 23307 6291 23363
rect 6316 23307 6372 23363
rect 6397 23307 6453 23363
rect 6478 23307 6534 23363
rect 6559 23307 6615 23363
rect 6640 23307 6696 23363
rect 6721 23307 6777 23363
rect 6802 23307 6858 23363
rect 6883 23307 6939 23363
rect 6964 23307 7020 23363
rect 7045 23307 7101 23363
rect 7126 23307 7182 23363
rect 7207 23307 7263 23363
rect 7288 23307 7344 23363
rect 7369 23307 7425 23363
rect 7450 23307 7506 23363
rect 7531 23307 7587 23363
rect 7612 23307 7668 23363
rect 7693 23307 7749 23363
rect 7774 23307 7830 23363
rect 7855 23307 7911 23363
rect 7936 23307 7992 23363
rect 8017 23307 8073 23363
rect 8098 23307 8154 23363
rect 8179 23307 8235 23363
rect 8260 23307 8316 23363
rect 8341 23307 8397 23363
rect 8422 23307 8478 23363
rect 8503 23307 8559 23363
rect 8584 23307 8640 23363
rect 8665 23307 8721 23363
rect 8746 23307 8802 23363
rect 8827 23307 8883 23363
rect 8908 23307 8964 23363
rect 8989 23307 9045 23363
rect 9070 23307 9126 23363
rect 9151 23307 9207 23363
rect 9232 23307 9288 23363
rect 9313 23307 9369 23363
rect 9394 23307 9450 23363
rect 9475 23307 9531 23363
rect 9556 23307 9612 23363
rect 9637 23307 9693 23363
rect 9718 23307 9774 23363
rect 9799 23307 9855 23363
rect 9880 23307 9936 23363
rect 9961 23307 10017 23363
rect 10042 23307 10098 23363
rect 10123 23307 10179 23363
rect 10204 23307 10260 23363
rect 10285 23307 10341 23363
rect 10366 23307 10422 23363
rect 10447 23307 10503 23363
rect 10528 23307 10584 23363
rect 10609 23307 10665 23363
rect 10690 23307 10746 23363
rect 10771 23307 10827 23363
rect 10852 23307 10908 23363
rect 10933 23307 10989 23363
rect 11014 23307 11070 23363
rect 11095 23307 11151 23363
rect 11176 23307 11232 23363
rect 11257 23307 11313 23363
rect 11338 23307 11394 23363
rect 11419 23307 11475 23363
rect 2170 23236 2226 23292
rect 2252 23236 2308 23292
rect 2334 23236 2390 23292
rect 2416 23236 2472 23292
rect 5425 23227 5481 23283
rect 5506 23227 5562 23283
rect 5587 23227 5643 23283
rect 5668 23227 5724 23283
rect 5749 23227 5805 23283
rect 5830 23227 5886 23283
rect 5911 23227 5967 23283
rect 5992 23227 6048 23283
rect 6073 23227 6129 23283
rect 6154 23227 6210 23283
rect 6235 23227 6291 23283
rect 6316 23227 6372 23283
rect 6397 23227 6453 23283
rect 6478 23227 6534 23283
rect 6559 23227 6615 23283
rect 6640 23227 6696 23283
rect 6721 23227 6777 23283
rect 6802 23227 6858 23283
rect 6883 23227 6939 23283
rect 6964 23227 7020 23283
rect 7045 23227 7101 23283
rect 7126 23227 7182 23283
rect 7207 23227 7263 23283
rect 7288 23227 7344 23283
rect 7369 23227 7425 23283
rect 7450 23227 7506 23283
rect 7531 23227 7587 23283
rect 7612 23227 7668 23283
rect 7693 23227 7749 23283
rect 7774 23227 7830 23283
rect 7855 23227 7911 23283
rect 7936 23227 7992 23283
rect 8017 23227 8073 23283
rect 8098 23227 8154 23283
rect 8179 23227 8235 23283
rect 8260 23227 8316 23283
rect 8341 23227 8397 23283
rect 8422 23227 8478 23283
rect 8503 23227 8559 23283
rect 8584 23227 8640 23283
rect 8665 23227 8721 23283
rect 8746 23227 8802 23283
rect 8827 23227 8883 23283
rect 8908 23227 8964 23283
rect 8989 23227 9045 23283
rect 9070 23227 9126 23283
rect 9151 23227 9207 23283
rect 9232 23227 9288 23283
rect 9313 23227 9369 23283
rect 9394 23227 9450 23283
rect 9475 23227 9531 23283
rect 9556 23227 9612 23283
rect 9637 23227 9693 23283
rect 9718 23227 9774 23283
rect 9799 23227 9855 23283
rect 9880 23227 9936 23283
rect 9961 23227 10017 23283
rect 10042 23227 10098 23283
rect 10123 23227 10179 23283
rect 10204 23227 10260 23283
rect 10285 23227 10341 23283
rect 10366 23227 10422 23283
rect 10447 23227 10503 23283
rect 10528 23227 10584 23283
rect 10609 23227 10665 23283
rect 10690 23227 10746 23283
rect 10771 23227 10827 23283
rect 10852 23227 10908 23283
rect 10933 23227 10989 23283
rect 11014 23227 11070 23283
rect 11095 23227 11151 23283
rect 11176 23227 11232 23283
rect 11257 23227 11313 23283
rect 11338 23227 11394 23283
rect 11419 23227 11475 23283
rect 2170 23154 2226 23210
rect 2252 23154 2308 23210
rect 2334 23154 2390 23210
rect 2416 23154 2472 23210
rect 5425 23147 5481 23203
rect 5506 23147 5562 23203
rect 5587 23147 5643 23203
rect 5668 23147 5724 23203
rect 5749 23147 5805 23203
rect 5830 23147 5886 23203
rect 5911 23147 5967 23203
rect 5992 23147 6048 23203
rect 6073 23147 6129 23203
rect 6154 23147 6210 23203
rect 6235 23147 6291 23203
rect 6316 23147 6372 23203
rect 6397 23147 6453 23203
rect 6478 23147 6534 23203
rect 6559 23147 6615 23203
rect 6640 23147 6696 23203
rect 6721 23147 6777 23203
rect 6802 23147 6858 23203
rect 6883 23147 6939 23203
rect 6964 23147 7020 23203
rect 7045 23147 7101 23203
rect 7126 23147 7182 23203
rect 7207 23147 7263 23203
rect 7288 23147 7344 23203
rect 7369 23147 7425 23203
rect 7450 23147 7506 23203
rect 7531 23147 7587 23203
rect 7612 23147 7668 23203
rect 7693 23147 7749 23203
rect 7774 23147 7830 23203
rect 7855 23147 7911 23203
rect 7936 23147 7992 23203
rect 8017 23147 8073 23203
rect 8098 23147 8154 23203
rect 8179 23147 8235 23203
rect 8260 23147 8316 23203
rect 8341 23147 8397 23203
rect 8422 23147 8478 23203
rect 8503 23147 8559 23203
rect 8584 23147 8640 23203
rect 8665 23147 8721 23203
rect 8746 23147 8802 23203
rect 8827 23147 8883 23203
rect 8908 23147 8964 23203
rect 8989 23147 9045 23203
rect 9070 23147 9126 23203
rect 9151 23147 9207 23203
rect 9232 23147 9288 23203
rect 9313 23147 9369 23203
rect 9394 23147 9450 23203
rect 9475 23147 9531 23203
rect 9556 23147 9612 23203
rect 9637 23147 9693 23203
rect 9718 23147 9774 23203
rect 9799 23147 9855 23203
rect 9880 23147 9936 23203
rect 9961 23147 10017 23203
rect 10042 23147 10098 23203
rect 10123 23147 10179 23203
rect 10204 23147 10260 23203
rect 10285 23147 10341 23203
rect 10366 23147 10422 23203
rect 10447 23147 10503 23203
rect 10528 23147 10584 23203
rect 10609 23147 10665 23203
rect 10690 23147 10746 23203
rect 10771 23147 10827 23203
rect 10852 23147 10908 23203
rect 10933 23147 10989 23203
rect 11014 23147 11070 23203
rect 11095 23147 11151 23203
rect 11176 23147 11232 23203
rect 11257 23147 11313 23203
rect 11338 23147 11394 23203
rect 11419 23147 11475 23203
rect 11500 23147 13076 24323
rect 14509 24299 14565 24355
rect 14603 24299 14659 24355
rect 14697 24299 14753 24355
rect 14791 24299 14847 24355
rect 14885 24299 14941 24355
rect 14979 24299 15035 24355
rect 14509 24217 14565 24273
rect 14603 24217 14659 24273
rect 14697 24217 14753 24273
rect 14791 24217 14847 24273
rect 14885 24217 14941 24273
rect 14979 24217 15035 24273
rect 14509 24135 14565 24191
rect 14603 24135 14659 24191
rect 14697 24135 14753 24191
rect 14791 24135 14847 24191
rect 14885 24135 14941 24191
rect 14979 24135 15035 24191
rect 14509 24053 14565 24109
rect 14603 24053 14659 24109
rect 14697 24053 14753 24109
rect 14791 24053 14847 24109
rect 14885 24053 14941 24109
rect 14979 24053 15035 24109
rect 14509 23971 14565 24027
rect 14603 23971 14659 24027
rect 14697 23971 14753 24027
rect 14791 23971 14847 24027
rect 14885 23971 14941 24027
rect 14979 23971 15035 24027
rect 14509 23889 14565 23945
rect 14603 23889 14659 23945
rect 14697 23889 14753 23945
rect 14791 23889 14847 23945
rect 14885 23889 14941 23945
rect 14979 23889 15035 23945
rect 14509 23807 14565 23863
rect 14603 23807 14659 23863
rect 14697 23807 14753 23863
rect 14791 23807 14847 23863
rect 14885 23807 14941 23863
rect 14979 23807 15035 23863
rect 14509 23725 14565 23781
rect 14603 23725 14659 23781
rect 14697 23725 14753 23781
rect 14791 23725 14847 23781
rect 14885 23725 14941 23781
rect 14979 23725 15035 23781
rect 14509 23643 14565 23699
rect 14603 23643 14659 23699
rect 14697 23643 14753 23699
rect 14791 23643 14847 23699
rect 14885 23643 14941 23699
rect 14979 23643 15035 23699
rect 14509 23561 14565 23617
rect 14603 23561 14659 23617
rect 14697 23561 14753 23617
rect 14791 23561 14847 23617
rect 14885 23561 14941 23617
rect 14979 23561 15035 23617
rect 14509 23479 14565 23535
rect 14603 23479 14659 23535
rect 14697 23479 14753 23535
rect 14791 23479 14847 23535
rect 14885 23479 14941 23535
rect 14979 23479 15035 23535
rect 14509 23397 14565 23453
rect 14603 23397 14659 23453
rect 14697 23397 14753 23453
rect 14791 23397 14847 23453
rect 14885 23397 14941 23453
rect 14979 23397 15035 23453
rect 14509 23315 14565 23371
rect 14603 23315 14659 23371
rect 14697 23315 14753 23371
rect 14791 23315 14847 23371
rect 14885 23315 14941 23371
rect 14979 23315 15035 23371
rect 14509 23233 14565 23289
rect 14603 23233 14659 23289
rect 14697 23233 14753 23289
rect 14791 23233 14847 23289
rect 14885 23233 14941 23289
rect 14979 23233 15035 23289
rect 14509 23151 14565 23207
rect 14603 23151 14659 23207
rect 14697 23151 14753 23207
rect 14791 23151 14847 23207
rect 14885 23151 14941 23207
rect 14979 23151 15035 23207
rect 670 20918 726 20923
rect 794 20918 850 20923
rect 670 20867 712 20918
rect 712 20867 726 20918
rect 794 20867 796 20918
rect 796 20867 848 20918
rect 848 20867 850 20918
rect 670 20802 712 20832
rect 712 20802 726 20832
rect 794 20802 796 20832
rect 796 20802 848 20832
rect 848 20802 850 20832
rect 670 20790 726 20802
rect 794 20790 850 20802
rect 670 20776 712 20790
rect 712 20776 726 20790
rect 670 20738 712 20741
rect 712 20738 726 20741
rect 794 20776 796 20790
rect 796 20776 848 20790
rect 848 20776 850 20790
rect 794 20738 796 20741
rect 796 20738 848 20741
rect 848 20738 850 20741
rect 670 20726 726 20738
rect 794 20726 850 20738
rect 670 20685 712 20726
rect 712 20685 726 20726
rect 794 20685 796 20726
rect 796 20685 848 20726
rect 848 20685 850 20726
rect 670 20610 712 20650
rect 712 20610 726 20650
rect 794 20610 796 20650
rect 796 20610 848 20650
rect 848 20610 850 20650
rect 670 20598 726 20610
rect 794 20598 850 20610
rect 670 20594 712 20598
rect 712 20594 726 20598
rect 670 20546 712 20559
rect 712 20546 726 20559
rect 794 20594 796 20598
rect 796 20594 848 20598
rect 848 20594 850 20598
rect 794 20546 796 20559
rect 796 20546 848 20559
rect 848 20546 850 20559
rect 670 20534 726 20546
rect 794 20534 850 20546
rect 670 20503 712 20534
rect 712 20503 726 20534
rect 794 20503 796 20534
rect 796 20503 848 20534
rect 848 20503 850 20534
rect 670 20418 712 20468
rect 712 20418 726 20468
rect 794 20418 796 20468
rect 796 20418 848 20468
rect 848 20418 850 20468
rect 670 20412 726 20418
rect 794 20412 850 20418
rect 1627 20867 1683 20923
rect 1715 20867 1771 20923
rect 1803 20867 1859 20923
rect 1891 20867 1947 20923
rect 1979 20867 2035 20923
rect 2067 20867 2123 20923
rect 2790 20875 2846 20931
rect 2873 20875 2929 20931
rect 2956 20875 3012 20931
rect 3039 20875 3095 20931
rect 3122 20875 3178 20931
rect 3205 20875 3261 20931
rect 3288 20875 3344 20931
rect 3371 20875 3427 20931
rect 3454 20875 3510 20931
rect 3537 20875 3593 20931
rect 3620 20875 3676 20931
rect 3703 20875 3759 20931
rect 1627 20776 1683 20832
rect 1715 20776 1771 20832
rect 1803 20776 1859 20832
rect 1891 20776 1947 20832
rect 1979 20776 2035 20832
rect 2067 20776 2123 20832
rect 2790 20781 2846 20837
rect 2873 20781 2929 20837
rect 2956 20781 3012 20837
rect 3039 20781 3095 20837
rect 3122 20781 3178 20837
rect 3205 20781 3261 20837
rect 3288 20781 3344 20837
rect 3371 20781 3427 20837
rect 3454 20781 3510 20837
rect 3537 20781 3593 20837
rect 3620 20781 3676 20837
rect 3703 20781 3759 20837
rect 1627 20685 1683 20741
rect 1715 20685 1771 20741
rect 1803 20685 1859 20741
rect 1891 20685 1947 20741
rect 1979 20685 2035 20741
rect 2067 20685 2123 20741
rect 2790 20687 2846 20743
rect 2873 20687 2929 20743
rect 2956 20687 3012 20743
rect 3039 20687 3095 20743
rect 3122 20687 3178 20743
rect 3205 20687 3261 20743
rect 3288 20687 3344 20743
rect 3371 20687 3427 20743
rect 3454 20687 3510 20743
rect 3537 20687 3593 20743
rect 3620 20687 3676 20743
rect 3703 20687 3759 20743
rect 1627 20594 1683 20650
rect 1715 20594 1771 20650
rect 1803 20594 1859 20650
rect 1891 20594 1947 20650
rect 1979 20594 2035 20650
rect 2067 20594 2123 20650
rect 2790 20593 2846 20649
rect 2873 20593 2929 20649
rect 2956 20593 3012 20649
rect 3039 20593 3095 20649
rect 3122 20593 3178 20649
rect 3205 20593 3261 20649
rect 3288 20593 3344 20649
rect 3371 20593 3427 20649
rect 3454 20593 3510 20649
rect 3537 20593 3593 20649
rect 3620 20593 3676 20649
rect 3703 20593 3759 20649
rect 1627 20503 1683 20559
rect 1715 20503 1771 20559
rect 1803 20503 1859 20559
rect 1891 20503 1947 20559
rect 1979 20503 2035 20559
rect 2067 20503 2123 20559
rect 2790 20519 2836 20555
rect 2836 20519 2846 20555
rect 2873 20519 2905 20555
rect 2905 20519 2922 20555
rect 2922 20519 2929 20555
rect 2956 20519 2974 20555
rect 2974 20519 2991 20555
rect 2991 20519 3012 20555
rect 3039 20519 3043 20555
rect 3043 20519 3060 20555
rect 3060 20519 3095 20555
rect 3122 20519 3128 20555
rect 3128 20519 3178 20555
rect 3205 20519 3248 20555
rect 3248 20519 3261 20555
rect 3288 20519 3316 20555
rect 3316 20519 3332 20555
rect 3332 20519 3344 20555
rect 3371 20519 3384 20555
rect 3384 20519 3400 20555
rect 3400 20519 3427 20555
rect 3454 20519 3468 20555
rect 3468 20519 3510 20555
rect 3537 20519 3588 20555
rect 3588 20519 3593 20555
rect 3620 20519 3656 20555
rect 3656 20519 3672 20555
rect 3672 20519 3676 20555
rect 3703 20519 3724 20555
rect 3724 20519 3759 20555
rect 2790 20499 2846 20519
rect 2873 20499 2929 20519
rect 2956 20499 3012 20519
rect 3039 20499 3095 20519
rect 3122 20499 3178 20519
rect 3205 20499 3261 20519
rect 3288 20499 3344 20519
rect 3371 20499 3427 20519
rect 3454 20499 3510 20519
rect 3537 20499 3593 20519
rect 3620 20499 3676 20519
rect 3703 20499 3759 20519
rect 1627 20412 1683 20468
rect 1715 20412 1771 20468
rect 1803 20412 1859 20468
rect 1891 20412 1947 20468
rect 1979 20412 2035 20468
rect 2067 20412 2123 20468
rect 2790 20459 2846 20461
rect 2873 20459 2929 20461
rect 2956 20459 3012 20461
rect 3039 20459 3095 20461
rect 3122 20459 3178 20461
rect 3205 20459 3261 20461
rect 3288 20459 3344 20461
rect 3371 20459 3427 20461
rect 3454 20459 3510 20461
rect 3537 20459 3593 20461
rect 3620 20459 3676 20461
rect 3703 20459 3759 20461
rect 2790 20407 2836 20459
rect 2836 20407 2846 20459
rect 2873 20407 2905 20459
rect 2905 20407 2922 20459
rect 2922 20407 2929 20459
rect 2956 20407 2974 20459
rect 2974 20407 2991 20459
rect 2991 20407 3012 20459
rect 3039 20407 3043 20459
rect 3043 20407 3060 20459
rect 3060 20407 3095 20459
rect 3122 20407 3128 20459
rect 3128 20407 3178 20459
rect 3205 20407 3248 20459
rect 3248 20407 3261 20459
rect 3288 20407 3316 20459
rect 3316 20407 3332 20459
rect 3332 20407 3344 20459
rect 3371 20407 3384 20459
rect 3384 20407 3400 20459
rect 3400 20407 3427 20459
rect 3454 20407 3468 20459
rect 3468 20407 3510 20459
rect 3537 20407 3588 20459
rect 3588 20407 3593 20459
rect 3620 20407 3656 20459
rect 3656 20407 3672 20459
rect 3672 20407 3676 20459
rect 3703 20407 3724 20459
rect 3724 20407 3759 20459
rect 2790 20405 2846 20407
rect 2873 20405 2929 20407
rect 2956 20405 3012 20407
rect 3039 20405 3095 20407
rect 3122 20405 3178 20407
rect 3205 20405 3261 20407
rect 3288 20405 3344 20407
rect 3371 20405 3427 20407
rect 3454 20405 3510 20407
rect 3537 20405 3593 20407
rect 3620 20405 3676 20407
rect 3703 20405 3759 20407
rect 2790 19191 2839 19243
rect 2839 19191 2846 19243
rect 2874 19191 2906 19243
rect 2906 19191 2921 19243
rect 2921 19191 2930 19243
rect 2958 19191 2973 19243
rect 2973 19191 2988 19243
rect 2988 19191 3014 19243
rect 3042 19191 3055 19243
rect 3055 19191 3098 19243
rect 3126 19191 3174 19243
rect 3174 19191 3182 19243
rect 3210 19191 3241 19243
rect 3241 19191 3256 19243
rect 3256 19191 3266 19243
rect 3294 19191 3308 19243
rect 3308 19191 3323 19243
rect 3323 19191 3350 19243
rect 3378 19191 3390 19243
rect 3390 19191 3434 19243
rect 3462 19191 3508 19243
rect 3508 19191 3518 19243
rect 3546 19191 3574 19243
rect 3574 19191 3588 19243
rect 3588 19191 3602 19243
rect 3630 19191 3640 19243
rect 3640 19191 3654 19243
rect 3654 19191 3686 19243
rect 3713 19191 3720 19243
rect 3720 19191 3769 19243
rect 2790 19187 2846 19191
rect 2874 19187 2930 19191
rect 2958 19187 3014 19191
rect 3042 19187 3098 19191
rect 3126 19187 3182 19191
rect 3210 19187 3266 19191
rect 3294 19187 3350 19191
rect 3378 19187 3434 19191
rect 3462 19187 3518 19191
rect 3546 19187 3602 19191
rect 3630 19187 3686 19191
rect 3713 19187 3769 19191
rect 3025 19069 3081 19073
rect 3111 19069 3167 19073
rect 3197 19069 3253 19073
rect 3283 19069 3339 19073
rect 3369 19069 3425 19073
rect 3455 19069 3511 19073
rect 3541 19069 3597 19073
rect 3627 19069 3683 19073
rect 3713 19069 3769 19073
rect 3025 19017 3074 19069
rect 3074 19017 3081 19069
rect 3111 19017 3144 19069
rect 3144 19017 3162 19069
rect 3162 19017 3167 19069
rect 3197 19017 3214 19069
rect 3214 19017 3232 19069
rect 3232 19017 3253 19069
rect 3283 19017 3284 19069
rect 3284 19017 3302 19069
rect 3302 19017 3339 19069
rect 3369 19017 3372 19069
rect 3372 19017 3424 19069
rect 3424 19017 3425 19069
rect 3455 19017 3494 19069
rect 3494 19017 3511 19069
rect 3541 19017 3564 19069
rect 3564 19017 3582 19069
rect 3582 19017 3597 19069
rect 3627 19017 3634 19069
rect 3634 19017 3651 19069
rect 3651 19017 3683 19069
rect 3713 19017 3720 19069
rect 3720 19017 3769 19069
rect 3207 17349 3263 17353
rect 3207 17297 3256 17349
rect 3256 17297 3263 17349
rect 3289 17349 3345 17353
rect 3289 17297 3296 17349
rect 3296 17297 3345 17349
rect 8454 17227 8510 17283
rect 8604 17227 8660 17283
rect 8754 17227 8810 17283
rect 8903 17227 8959 17283
rect 9052 17227 9108 17283
rect 8454 17139 8510 17195
rect 8604 17139 8660 17195
rect 8754 17139 8810 17195
rect 8903 17139 8959 17195
rect 9052 17139 9108 17195
rect 8454 17051 8510 17107
rect 8604 17051 8660 17107
rect 8754 17051 8810 17107
rect 8903 17051 8959 17107
rect 9052 17051 9108 17107
rect 7041 16777 7097 16795
rect 7121 16777 7177 16795
rect 7041 16739 7088 16777
rect 7088 16739 7097 16777
rect 7121 16739 7152 16777
rect 7152 16739 7164 16777
rect 7164 16739 7177 16777
rect 8454 16395 8510 16451
rect 8604 16395 8660 16451
rect 8754 16395 8810 16451
rect 8903 16395 8959 16451
rect 9052 16395 9108 16451
rect 3894 16327 3950 16383
rect 4019 16327 4075 16383
rect 4144 16327 4200 16383
rect 4269 16327 4325 16383
rect 3894 16247 3950 16303
rect 4019 16247 4075 16303
rect 4144 16247 4200 16303
rect 4269 16247 4325 16303
rect 3894 16167 3950 16223
rect 4019 16167 4075 16223
rect 4144 16167 4200 16223
rect 4269 16167 4325 16223
rect 8454 16307 8510 16363
rect 8604 16307 8660 16363
rect 8754 16307 8810 16363
rect 8903 16307 8959 16363
rect 9052 16307 9108 16363
rect 8454 16219 8510 16275
rect 8604 16219 8660 16275
rect 8754 16219 8810 16275
rect 8903 16219 8959 16275
rect 9052 16219 9108 16275
rect 11011 13844 11067 13900
rect 11111 13844 11167 13900
rect 11211 13844 11267 13900
rect 2234 9999 2283 10044
rect 2283 9999 2290 10044
rect 2333 9999 2351 10044
rect 2351 9999 2367 10044
rect 2367 9999 2389 10044
rect 2431 9999 2435 10044
rect 2435 9999 2487 10044
rect 2529 9999 2555 10044
rect 2555 9999 2571 10044
rect 2571 9999 2585 10044
rect 2627 9999 2638 10044
rect 2638 9999 2683 10044
rect 2234 9988 2290 9999
rect 2333 9988 2389 9999
rect 2431 9988 2487 9999
rect 2529 9988 2585 9999
rect 2627 9988 2683 9999
rect 2234 9925 2283 9950
rect 2283 9925 2290 9950
rect 2333 9925 2351 9950
rect 2351 9925 2367 9950
rect 2367 9925 2389 9950
rect 2431 9925 2435 9950
rect 2435 9925 2487 9950
rect 2529 9925 2555 9950
rect 2555 9925 2571 9950
rect 2571 9925 2585 9950
rect 2627 9925 2638 9950
rect 2638 9925 2683 9950
rect 2234 9903 2290 9925
rect 2333 9903 2389 9925
rect 2431 9903 2487 9925
rect 2529 9903 2585 9925
rect 2627 9903 2683 9925
rect 2234 9894 2283 9903
rect 2283 9894 2290 9903
rect 2333 9894 2351 9903
rect 2351 9894 2367 9903
rect 2367 9894 2389 9903
rect 2431 9894 2435 9903
rect 2435 9894 2487 9903
rect 2234 9851 2283 9856
rect 2283 9851 2290 9856
rect 2333 9851 2351 9856
rect 2351 9851 2367 9856
rect 2367 9851 2389 9856
rect 2431 9851 2435 9856
rect 2435 9851 2487 9856
rect 2529 9894 2555 9903
rect 2555 9894 2571 9903
rect 2571 9894 2585 9903
rect 2627 9894 2638 9903
rect 2638 9894 2683 9903
rect 2529 9851 2555 9856
rect 2555 9851 2571 9856
rect 2571 9851 2585 9856
rect 2627 9851 2638 9856
rect 2638 9851 2683 9856
rect 2234 9829 2290 9851
rect 2333 9829 2389 9851
rect 2431 9829 2487 9851
rect 2529 9829 2585 9851
rect 2627 9829 2683 9851
rect 2234 9800 2283 9829
rect 2283 9800 2290 9829
rect 2333 9800 2351 9829
rect 2351 9800 2367 9829
rect 2367 9800 2389 9829
rect 2431 9800 2435 9829
rect 2435 9800 2487 9829
rect 2529 9800 2555 9829
rect 2555 9800 2571 9829
rect 2571 9800 2585 9829
rect 2627 9800 2638 9829
rect 2638 9800 2683 9829
rect 2234 9755 2290 9762
rect 2333 9755 2389 9762
rect 2431 9755 2487 9762
rect 2529 9755 2585 9762
rect 2627 9755 2683 9762
rect 2234 9706 2283 9755
rect 2283 9706 2290 9755
rect 2333 9706 2351 9755
rect 2351 9706 2367 9755
rect 2367 9706 2389 9755
rect 2431 9706 2435 9755
rect 2435 9706 2487 9755
rect 2529 9706 2555 9755
rect 2555 9706 2571 9755
rect 2571 9706 2585 9755
rect 2627 9706 2638 9755
rect 2638 9706 2683 9755
rect 9346 13059 9402 13077
rect 9346 13021 9359 13059
rect 9359 13021 9402 13059
rect 9346 12995 9402 12997
rect 9346 12943 9359 12995
rect 9359 12943 9402 12995
rect 9346 12941 9402 12943
rect 9475 13024 9531 13080
rect 9475 12944 9531 13000
rect 8023 11784 8079 11840
rect 8023 11747 8079 11760
rect 8023 11704 8068 11747
rect 8068 11704 8079 11747
rect 4625 11472 4681 11528
rect 4715 11472 4771 11528
rect 6704 11530 6760 11586
rect 6704 11450 6760 11506
rect 2999 10385 3055 10398
rect 3088 10385 3144 10398
rect 3177 10385 3233 10398
rect 3265 10385 3321 10398
rect 3353 10385 3409 10398
rect 3441 10385 3497 10398
rect 3529 10385 3585 10398
rect 3617 10385 3673 10398
rect 3705 10385 3761 10398
rect 2999 10342 3000 10385
rect 3000 10342 3052 10385
rect 3052 10342 3055 10385
rect 3088 10342 3117 10385
rect 3117 10342 3130 10385
rect 3130 10342 3144 10385
rect 3177 10342 3182 10385
rect 3182 10342 3194 10385
rect 3194 10342 3233 10385
rect 3265 10342 3310 10385
rect 3310 10342 3321 10385
rect 3353 10342 3374 10385
rect 3374 10342 3386 10385
rect 3386 10342 3409 10385
rect 3441 10342 3450 10385
rect 3450 10342 3497 10385
rect 3529 10342 3566 10385
rect 3566 10342 3578 10385
rect 3578 10342 3585 10385
rect 3617 10342 3630 10385
rect 3630 10342 3642 10385
rect 3642 10342 3673 10385
rect 3705 10342 3706 10385
rect 3706 10342 3758 10385
rect 3758 10342 3761 10385
rect 2999 10309 3055 10318
rect 3088 10309 3144 10318
rect 3177 10309 3233 10318
rect 3265 10309 3321 10318
rect 3353 10309 3409 10318
rect 3441 10309 3497 10318
rect 3529 10309 3585 10318
rect 3617 10309 3673 10318
rect 3705 10309 3761 10318
rect 2999 10262 3000 10309
rect 3000 10262 3052 10309
rect 3052 10262 3055 10309
rect 3088 10262 3117 10309
rect 3117 10262 3130 10309
rect 3130 10262 3144 10309
rect 3177 10262 3182 10309
rect 3182 10262 3194 10309
rect 3194 10262 3233 10309
rect 3265 10262 3310 10309
rect 3310 10262 3321 10309
rect 3353 10262 3374 10309
rect 3374 10262 3386 10309
rect 3386 10262 3409 10309
rect 3441 10262 3450 10309
rect 3450 10262 3497 10309
rect 3529 10262 3566 10309
rect 3566 10262 3578 10309
rect 3578 10262 3585 10309
rect 3617 10262 3630 10309
rect 3630 10262 3642 10309
rect 3642 10262 3673 10309
rect 3705 10262 3706 10309
rect 3706 10262 3758 10309
rect 3758 10262 3761 10309
rect 2789 9259 2845 9260
rect 2921 9259 2977 9260
rect 3053 9259 3109 9260
rect 3185 9259 3241 9260
rect 3317 9259 3373 9260
rect 3449 9259 3505 9260
rect 3581 9259 3637 9260
rect 3713 9259 3769 9260
rect 2789 9207 2836 9259
rect 2836 9207 2845 9259
rect 2921 9207 2970 9259
rect 2970 9207 2977 9259
rect 3053 9207 3104 9259
rect 3104 9207 3109 9259
rect 3185 9207 3186 9259
rect 3186 9207 3238 9259
rect 3238 9207 3241 9259
rect 3317 9207 3320 9259
rect 3320 9207 3372 9259
rect 3372 9207 3373 9259
rect 3449 9207 3454 9259
rect 3454 9207 3505 9259
rect 3581 9207 3588 9259
rect 3588 9207 3637 9259
rect 3713 9207 3720 9259
rect 3720 9207 3769 9259
rect 2789 9204 2845 9207
rect 2921 9204 2977 9207
rect 3053 9204 3109 9207
rect 3185 9204 3241 9207
rect 3317 9204 3373 9207
rect 3449 9204 3505 9207
rect 3581 9204 3637 9207
rect 3713 9204 3769 9207
rect 2789 9111 2845 9120
rect 2921 9111 2977 9120
rect 3053 9111 3109 9120
rect 3185 9111 3241 9120
rect 3317 9111 3373 9120
rect 3449 9111 3505 9120
rect 3581 9111 3637 9120
rect 3713 9111 3769 9120
rect 2789 9064 2836 9111
rect 2836 9064 2845 9111
rect 2921 9064 2970 9111
rect 2970 9064 2977 9111
rect 3053 9064 3104 9111
rect 3104 9064 3109 9111
rect 3185 9064 3186 9111
rect 3186 9064 3238 9111
rect 3238 9064 3241 9111
rect 3317 9064 3320 9111
rect 3320 9064 3372 9111
rect 3372 9064 3373 9111
rect 3449 9064 3454 9111
rect 3454 9064 3505 9111
rect 3581 9064 3588 9111
rect 3588 9064 3637 9111
rect 3713 9064 3720 9111
rect 3720 9064 3769 9111
rect 2850 8217 2897 8232
rect 2897 8217 2906 8232
rect 2974 8217 2981 8232
rect 2981 8217 3030 8232
rect 3098 8217 3101 8232
rect 3101 8217 3117 8232
rect 3117 8217 3154 8232
rect 3221 8217 3236 8232
rect 3236 8217 3251 8232
rect 3251 8217 3277 8232
rect 3344 8217 3370 8232
rect 3370 8217 3385 8232
rect 3385 8217 3400 8232
rect 3467 8217 3504 8232
rect 3504 8217 3519 8232
rect 3519 8217 3523 8232
rect 3590 8217 3638 8232
rect 3638 8217 3646 8232
rect 3713 8217 3720 8232
rect 3720 8217 3769 8232
rect 2850 8191 2906 8217
rect 2974 8191 3030 8217
rect 3098 8191 3154 8217
rect 3221 8191 3277 8217
rect 3344 8191 3400 8217
rect 3467 8191 3523 8217
rect 3590 8191 3646 8217
rect 3713 8191 3769 8217
rect 2850 8176 2897 8191
rect 2897 8176 2906 8191
rect 2974 8176 2981 8191
rect 2981 8176 3030 8191
rect 3098 8176 3101 8191
rect 3101 8176 3117 8191
rect 3117 8176 3154 8191
rect 3221 8176 3236 8191
rect 3236 8176 3251 8191
rect 3251 8176 3277 8191
rect 3344 8176 3370 8191
rect 3370 8176 3385 8191
rect 3385 8176 3400 8191
rect 3467 8176 3504 8191
rect 3504 8176 3519 8191
rect 3519 8176 3523 8191
rect 3590 8176 3638 8191
rect 3638 8176 3646 8191
rect 3713 8176 3720 8191
rect 3720 8176 3769 8191
rect 1536 8021 1592 8077
rect 1626 8021 1682 8077
rect 1716 8021 1772 8077
rect 1806 8021 1862 8077
rect 1896 8021 1952 8077
rect 1986 8021 2042 8077
rect 2076 8021 2132 8077
rect 1536 7937 1592 7993
rect 1626 7937 1682 7993
rect 1716 7937 1772 7993
rect 1806 7937 1862 7993
rect 1896 7937 1952 7993
rect 1986 7937 2042 7993
rect 2076 7937 2132 7993
rect 1536 7853 1592 7909
rect 1626 7853 1682 7909
rect 1716 7853 1772 7909
rect 1806 7853 1862 7909
rect 1896 7853 1952 7909
rect 1986 7853 2042 7909
rect 2076 7853 2132 7909
rect 941 2757 997 2813
rect 941 2677 997 2733
rect 1536 7769 1592 7825
rect 1626 7769 1682 7825
rect 1716 7769 1772 7825
rect 1806 7769 1862 7825
rect 1896 7769 1952 7825
rect 1986 7769 2042 7825
rect 2076 7769 2132 7825
rect 1536 7685 1592 7741
rect 1626 7685 1682 7741
rect 1716 7685 1772 7741
rect 1806 7685 1862 7741
rect 1896 7685 1952 7741
rect 1986 7685 2042 7741
rect 2076 7685 2132 7741
rect 1536 7601 1592 7657
rect 1626 7601 1682 7657
rect 1716 7601 1772 7657
rect 1806 7601 1862 7657
rect 1896 7601 1952 7657
rect 1986 7601 2042 7657
rect 2076 7601 2132 7657
rect 1536 7517 1592 7573
rect 1626 7517 1682 7573
rect 1716 7517 1772 7573
rect 1806 7517 1862 7573
rect 1896 7517 1952 7573
rect 1986 7517 2042 7573
rect 2076 7517 2132 7573
rect 1536 7433 1592 7489
rect 1626 7433 1682 7489
rect 1716 7433 1772 7489
rect 1806 7433 1862 7489
rect 1896 7433 1952 7489
rect 1986 7433 2042 7489
rect 2076 7433 2132 7489
rect 1536 7349 1592 7405
rect 1626 7349 1682 7405
rect 1716 7349 1772 7405
rect 1806 7349 1862 7405
rect 1896 7349 1952 7405
rect 1986 7349 2042 7405
rect 2076 7349 2132 7405
rect 1536 7265 1592 7321
rect 1626 7265 1682 7321
rect 1716 7265 1772 7321
rect 1806 7265 1862 7321
rect 1896 7265 1952 7321
rect 1986 7265 2042 7321
rect 2076 7265 2132 7321
rect 1536 7181 1592 7237
rect 1626 7181 1682 7237
rect 1716 7181 1772 7237
rect 1806 7181 1862 7237
rect 1896 7181 1952 7237
rect 1986 7181 2042 7237
rect 2076 7181 2132 7237
rect 1536 7096 1592 7152
rect 1626 7096 1682 7152
rect 1716 7096 1772 7152
rect 1806 7096 1862 7152
rect 1896 7096 1952 7152
rect 1986 7096 2042 7152
rect 2076 7096 2132 7152
rect 1536 7011 1592 7067
rect 1626 7011 1682 7067
rect 1716 7011 1772 7067
rect 1806 7011 1862 7067
rect 1896 7011 1952 7067
rect 1986 7011 2042 7067
rect 2076 7011 2132 7067
rect 1536 6926 1592 6982
rect 1626 6926 1682 6982
rect 1716 6926 1772 6982
rect 1806 6926 1862 6982
rect 1896 6926 1952 6982
rect 1986 6926 2042 6982
rect 2076 6926 2132 6982
rect 1536 6841 1592 6897
rect 1626 6841 1682 6897
rect 1716 6841 1772 6897
rect 1806 6841 1862 6897
rect 1896 6841 1952 6897
rect 1986 6841 2042 6897
rect 2076 6841 2132 6897
rect 1536 6756 1592 6812
rect 1626 6756 1682 6812
rect 1716 6756 1772 6812
rect 1806 6756 1862 6812
rect 1896 6756 1952 6812
rect 1986 6756 2042 6812
rect 2076 6756 2132 6812
rect 1536 6671 1592 6727
rect 1626 6671 1682 6727
rect 1716 6671 1772 6727
rect 1806 6671 1862 6727
rect 1896 6671 1952 6727
rect 1986 6671 2042 6727
rect 2076 6671 2132 6727
rect 1709 6579 1765 6635
rect 1797 6579 1853 6635
rect 1885 6579 1941 6635
rect 1973 6579 2029 6635
rect 2061 6579 2117 6635
rect 1709 6495 1765 6551
rect 1797 6495 1853 6551
rect 1885 6495 1941 6551
rect 1973 6495 2029 6551
rect 2061 6495 2117 6551
rect 1709 6411 1765 6467
rect 1797 6411 1853 6467
rect 1885 6411 1941 6467
rect 1973 6411 2029 6467
rect 2061 6411 2117 6467
rect 1709 6327 1765 6383
rect 1797 6327 1853 6383
rect 1885 6327 1941 6383
rect 1973 6327 2029 6383
rect 2061 6327 2117 6383
rect 1709 6243 1765 6299
rect 1797 6243 1853 6299
rect 1885 6243 1941 6299
rect 1973 6243 2029 6299
rect 2061 6243 2117 6299
rect 1709 6159 1765 6215
rect 1797 6159 1853 6215
rect 1885 6159 1941 6215
rect 1973 6159 2029 6215
rect 2061 6159 2117 6215
rect 1709 6075 1765 6131
rect 1797 6075 1853 6131
rect 1885 6075 1941 6131
rect 1973 6075 2029 6131
rect 2061 6075 2117 6131
rect 1709 5990 1765 6046
rect 1797 5990 1853 6046
rect 1885 5990 1941 6046
rect 1973 5990 2029 6046
rect 2061 5990 2117 6046
rect 1709 5905 1765 5961
rect 1797 5905 1853 5961
rect 1885 5905 1941 5961
rect 1973 5905 2029 5961
rect 2061 5905 2117 5961
rect 1708 5780 1764 5836
rect 1814 5780 1870 5836
rect 1920 5780 1976 5836
rect 1708 5698 1764 5754
rect 1814 5698 1870 5754
rect 1920 5698 1976 5754
rect 1708 5616 1764 5672
rect 1814 5616 1870 5672
rect 1920 5616 1976 5672
rect 1708 5534 1764 5590
rect 1814 5534 1870 5590
rect 1920 5534 1976 5590
rect 1708 5452 1764 5508
rect 1814 5452 1870 5508
rect 1920 5452 1976 5508
rect 1708 5370 1764 5426
rect 1814 5370 1870 5426
rect 1920 5370 1976 5426
rect 1708 5287 1764 5343
rect 1814 5287 1870 5343
rect 1920 5287 1976 5343
rect 1709 5172 1765 5228
rect 1797 5172 1853 5228
rect 1885 5172 1941 5228
rect 1973 5172 2029 5228
rect 2061 5172 2117 5228
rect 1709 5092 1765 5148
rect 1797 5092 1853 5148
rect 1885 5092 1941 5148
rect 1973 5092 2029 5148
rect 2061 5092 2117 5148
rect 1709 5012 1765 5068
rect 1797 5012 1853 5068
rect 1885 5012 1941 5068
rect 1973 5012 2029 5068
rect 2061 5012 2117 5068
rect 1709 4932 1765 4988
rect 1797 4932 1853 4988
rect 1885 4932 1941 4988
rect 1973 4932 2029 4988
rect 2061 4932 2117 4988
rect 1709 4852 1765 4908
rect 1797 4852 1853 4908
rect 1885 4852 1941 4908
rect 1973 4852 2029 4908
rect 2061 4852 2117 4908
rect 1709 4772 1765 4828
rect 1797 4772 1853 4828
rect 1885 4772 1941 4828
rect 1973 4772 2029 4828
rect 2061 4772 2117 4828
rect 1709 4691 1765 4747
rect 1797 4691 1853 4747
rect 1885 4691 1941 4747
rect 1973 4691 2029 4747
rect 2061 4691 2117 4747
rect 1709 4610 1765 4666
rect 1797 4610 1853 4666
rect 1885 4610 1941 4666
rect 1973 4610 2029 4666
rect 2061 4610 2117 4666
rect 1709 4529 1765 4585
rect 1797 4529 1853 4585
rect 1885 4529 1941 4585
rect 1973 4529 2029 4585
rect 2061 4529 2117 4585
rect 1709 4448 1765 4504
rect 1797 4448 1853 4504
rect 1885 4448 1941 4504
rect 1973 4448 2029 4504
rect 2061 4448 2117 4504
rect 1709 4367 1765 4423
rect 1797 4367 1853 4423
rect 1885 4367 1941 4423
rect 1973 4367 2029 4423
rect 2061 4367 2117 4423
rect 1709 4286 1765 4342
rect 1797 4286 1853 4342
rect 1885 4286 1941 4342
rect 1973 4286 2029 4342
rect 2061 4286 2117 4342
rect 1709 4205 1765 4261
rect 1797 4205 1853 4261
rect 1885 4205 1941 4261
rect 1973 4205 2029 4261
rect 2061 4205 2117 4261
rect 1709 4124 1765 4180
rect 1797 4124 1853 4180
rect 1885 4124 1941 4180
rect 1973 4124 2029 4180
rect 2061 4124 2117 4180
rect 1709 4043 1765 4099
rect 1797 4043 1853 4099
rect 1885 4043 1941 4099
rect 1973 4043 2029 4099
rect 2061 4043 2117 4099
rect 1709 3962 1765 4018
rect 1797 3962 1853 4018
rect 1885 3962 1941 4018
rect 1973 3962 2029 4018
rect 2061 3962 2117 4018
rect 1709 3881 1765 3937
rect 1797 3881 1853 3937
rect 1885 3881 1941 3937
rect 1973 3881 2029 3937
rect 2061 3881 2117 3937
rect 1507 1646 1563 1652
rect 1507 1596 1551 1646
rect 1551 1596 1563 1646
rect 1590 1646 1646 1652
rect 1590 1596 1603 1646
rect 1603 1596 1646 1646
rect 1507 1456 1551 1506
rect 1551 1456 1563 1506
rect 1507 1450 1563 1456
rect 1590 1456 1603 1506
rect 1603 1456 1646 1506
rect 1590 1450 1646 1456
rect 1789 1651 1845 1653
rect 1789 1599 1838 1651
rect 1838 1599 1845 1651
rect 1789 1597 1845 1599
rect 1789 1503 1845 1507
rect 1789 1451 1838 1503
rect 1838 1451 1845 1503
rect 288 274 344 330
rect 288 194 344 250
rect 11015 10281 11059 10326
rect 11059 10281 11071 10326
rect 11116 10281 11133 10326
rect 11133 10281 11155 10326
rect 11155 10281 11172 10326
rect 11216 10281 11229 10326
rect 11229 10281 11272 10326
rect 11015 10270 11071 10281
rect 11116 10270 11172 10281
rect 11216 10270 11272 10281
rect 11015 10205 11071 10216
rect 11116 10205 11172 10216
rect 11216 10205 11272 10216
rect 11015 10160 11059 10205
rect 11059 10160 11071 10205
rect 11116 10160 11133 10205
rect 11133 10160 11155 10205
rect 11155 10160 11172 10205
rect 11216 10160 11229 10205
rect 11229 10160 11272 10205
rect 7872 10028 7928 10030
rect 7872 9976 7874 10028
rect 7874 9976 7886 10028
rect 7886 9976 7928 10028
rect 7872 9974 7928 9976
rect 7872 9894 7928 9950
rect 9682 9932 9738 9988
rect 9682 9907 9738 9908
rect 9682 9855 9706 9907
rect 9706 9855 9718 9907
rect 9718 9855 9738 9907
rect 9682 9852 9738 9855
rect 10956 9448 10968 9471
rect 10968 9448 11012 9471
rect 11039 9448 11086 9471
rect 11086 9448 11095 9471
rect 11122 9448 11151 9471
rect 11151 9448 11164 9471
rect 11164 9448 11178 9471
rect 10956 9426 11012 9448
rect 11039 9426 11095 9448
rect 11122 9426 11178 9448
rect 10956 9415 10968 9426
rect 10968 9415 11012 9426
rect 10956 9374 10968 9387
rect 10968 9374 11012 9387
rect 11039 9415 11086 9426
rect 11086 9415 11095 9426
rect 11122 9415 11151 9426
rect 11151 9415 11164 9426
rect 11164 9415 11178 9426
rect 11039 9374 11086 9387
rect 11086 9374 11095 9387
rect 11122 9374 11151 9387
rect 11151 9374 11164 9387
rect 11164 9374 11178 9387
rect 10956 9352 11012 9374
rect 11039 9352 11095 9374
rect 11122 9352 11178 9374
rect 10956 9331 10968 9352
rect 10968 9331 11012 9352
rect 11039 9331 11086 9352
rect 11086 9331 11095 9352
rect 11122 9331 11151 9352
rect 11151 9331 11164 9352
rect 11164 9331 11178 9352
rect 9121 9209 9177 9265
rect 9217 9209 9273 9265
rect 9313 9209 9369 9265
rect 9409 9209 9465 9265
rect 9505 9209 9561 9265
rect 9121 9122 9177 9178
rect 9217 9122 9273 9178
rect 9313 9122 9369 9178
rect 9409 9122 9465 9178
rect 9505 9122 9561 9178
rect 9121 9035 9177 9091
rect 9217 9035 9273 9091
rect 9313 9035 9369 9091
rect 9409 9035 9465 9091
rect 9505 9035 9561 9091
rect 9121 8948 9177 9004
rect 9217 8948 9273 9004
rect 9313 8948 9369 9004
rect 9409 8948 9465 9004
rect 9505 8948 9561 9004
rect 9121 8861 9177 8917
rect 9217 8861 9273 8917
rect 9313 8861 9369 8917
rect 9409 8861 9465 8917
rect 9505 8861 9561 8917
rect 9121 8774 9177 8830
rect 9217 8774 9273 8830
rect 9313 8774 9369 8830
rect 9409 8774 9465 8830
rect 9505 8774 9561 8830
rect 9121 8686 9177 8742
rect 9217 8686 9273 8742
rect 9313 8686 9369 8742
rect 9409 8686 9465 8742
rect 9505 8686 9561 8742
rect 9121 8598 9177 8654
rect 9217 8598 9273 8654
rect 9313 8598 9369 8654
rect 9409 8598 9465 8654
rect 9505 8598 9561 8654
rect 9121 8510 9177 8566
rect 9217 8510 9273 8566
rect 9313 8510 9369 8566
rect 9409 8510 9465 8566
rect 9505 8510 9561 8566
rect 9121 8422 9177 8478
rect 9217 8422 9273 8478
rect 9313 8422 9369 8478
rect 9409 8422 9465 8478
rect 9505 8422 9561 8478
rect 9121 8334 9177 8390
rect 9217 8334 9273 8390
rect 9313 8334 9369 8390
rect 9409 8334 9465 8390
rect 9505 8334 9561 8390
rect 10506 8217 10554 8235
rect 10554 8217 10562 8235
rect 10506 8191 10562 8217
rect 10506 8179 10554 8191
rect 10554 8179 10562 8191
rect 10587 8217 10591 8235
rect 10591 8217 10643 8235
rect 10587 8191 10643 8217
rect 10587 8179 10591 8191
rect 10591 8179 10643 8191
rect 10668 8217 10680 8235
rect 10680 8217 10724 8235
rect 10668 8191 10724 8217
rect 10668 8179 10680 8191
rect 10680 8179 10724 8191
rect 13577 8257 13633 8313
rect 13661 8257 13717 8313
rect 13745 8257 13801 8313
rect 13829 8298 13872 8313
rect 13872 8298 13885 8313
rect 13912 8298 13944 8313
rect 13944 8298 13964 8313
rect 13964 8298 13968 8313
rect 13995 8298 14016 8313
rect 14016 8298 14036 8313
rect 14036 8298 14051 8313
rect 13829 8272 13885 8298
rect 13912 8272 13968 8298
rect 13995 8272 14051 8298
rect 13829 8257 13872 8272
rect 13872 8257 13885 8272
rect 13912 8257 13944 8272
rect 13944 8257 13964 8272
rect 13964 8257 13968 8272
rect 13995 8257 14016 8272
rect 14016 8257 14036 8272
rect 14036 8257 14051 8272
rect 14141 8127 14197 8183
rect 14285 8127 14341 8183
rect 14141 8046 14197 8102
rect 14285 8046 14341 8102
rect 14141 7965 14197 8021
rect 14285 7965 14341 8021
rect 14141 7884 14197 7940
rect 14285 7884 14341 7940
rect 14141 7803 14197 7859
rect 14285 7803 14341 7859
rect 14141 7722 14197 7778
rect 14285 7722 14341 7778
rect 14141 7641 14197 7697
rect 14285 7641 14341 7697
rect 14141 7560 14197 7616
rect 14285 7560 14341 7616
rect 14141 7479 14197 7535
rect 14285 7479 14341 7535
rect 14141 7398 14197 7454
rect 14285 7398 14341 7454
rect 14141 7317 14197 7373
rect 14285 7317 14341 7373
rect 14141 7235 14197 7291
rect 14285 7235 14341 7291
rect 14141 7153 14197 7209
rect 14285 7153 14341 7209
rect 14141 7071 14197 7127
rect 14285 7071 14341 7127
rect 14141 6989 14197 7045
rect 14285 6989 14341 7045
rect 14141 6907 14197 6963
rect 14285 6907 14341 6963
rect 14141 6825 14197 6881
rect 14285 6825 14341 6881
rect 14141 6743 14197 6799
rect 14285 6743 14341 6799
rect 14141 6661 14197 6717
rect 14285 6661 14341 6717
rect 14141 6579 14197 6635
rect 14285 6579 14341 6635
rect 14141 6497 14197 6553
rect 14285 6497 14341 6553
rect 14141 6415 14197 6471
rect 14285 6415 14341 6471
rect 14141 6333 14197 6389
rect 14285 6333 14341 6389
rect 3674 2594 3685 2639
rect 3685 2594 3702 2639
rect 3702 2594 3730 2639
rect 3756 2594 3771 2639
rect 3771 2594 3812 2639
rect 3837 2594 3840 2639
rect 3840 2594 3892 2639
rect 3892 2594 3893 2639
rect 3918 2594 3961 2639
rect 3961 2594 3974 2639
rect 3999 2594 4030 2639
rect 4030 2594 4047 2639
rect 4047 2594 4055 2639
rect 4080 2594 4099 2639
rect 4099 2594 4116 2639
rect 4116 2594 4136 2639
rect 4161 2594 4168 2639
rect 4168 2594 4185 2639
rect 4185 2594 4217 2639
rect 4242 2594 4254 2639
rect 4254 2594 4298 2639
rect 3674 2583 3730 2594
rect 3756 2583 3812 2594
rect 3837 2583 3893 2594
rect 3918 2583 3974 2594
rect 3999 2583 4055 2594
rect 4080 2583 4136 2594
rect 4161 2583 4217 2594
rect 4242 2583 4298 2594
rect 3674 2502 3730 2509
rect 3756 2502 3812 2509
rect 3837 2502 3893 2509
rect 3918 2502 3974 2509
rect 3999 2502 4055 2509
rect 4080 2502 4136 2509
rect 4161 2502 4217 2509
rect 4242 2502 4298 2509
rect 3674 2453 3685 2502
rect 3685 2453 3702 2502
rect 3702 2453 3730 2502
rect 3756 2453 3771 2502
rect 3771 2453 3812 2502
rect 3837 2453 3840 2502
rect 3840 2453 3892 2502
rect 3892 2453 3893 2502
rect 3918 2453 3961 2502
rect 3961 2453 3974 2502
rect 3999 2453 4030 2502
rect 4030 2453 4047 2502
rect 4047 2453 4055 2502
rect 4080 2453 4099 2502
rect 4099 2453 4116 2502
rect 4116 2453 4136 2502
rect 4161 2453 4168 2502
rect 4168 2453 4185 2502
rect 4185 2453 4217 2502
rect 4242 2453 4254 2502
rect 4254 2453 4298 2502
rect 2788 1086 2844 1087
rect 2889 1086 2945 1087
rect 2990 1086 3046 1087
rect 3091 1086 3147 1087
rect 3192 1086 3248 1087
rect 3293 1086 3349 1087
rect 1388 255 1444 256
rect 1475 255 1531 256
rect 1562 255 1618 256
rect 1388 203 1440 255
rect 1440 203 1444 255
rect 1475 203 1492 255
rect 1492 203 1531 255
rect 1562 203 1600 255
rect 1600 203 1618 255
rect 1388 200 1444 203
rect 1475 200 1531 203
rect 1562 200 1618 203
rect 1648 255 1704 256
rect 1734 255 1790 256
rect 1820 255 1876 256
rect 1906 255 1962 256
rect 1992 255 2048 256
rect 1648 203 1656 255
rect 1656 203 1704 255
rect 1734 203 1764 255
rect 1764 203 1790 255
rect 1820 203 1871 255
rect 1871 203 1876 255
rect 1906 203 1923 255
rect 1923 203 1962 255
rect 1992 203 2030 255
rect 2030 203 2048 255
rect 1648 200 1704 203
rect 1734 200 1790 203
rect 1820 200 1876 203
rect 1906 200 1962 203
rect 1992 200 2048 203
rect 2078 255 2134 256
rect 2078 203 2085 255
rect 2085 203 2134 255
rect 2078 200 2134 203
rect 1388 107 1444 110
rect 1475 107 1531 110
rect 1562 107 1618 110
rect 1388 55 1440 107
rect 1440 55 1444 107
rect 1475 55 1492 107
rect 1492 55 1531 107
rect 1562 55 1600 107
rect 1600 55 1618 107
rect 1388 54 1444 55
rect 1475 54 1531 55
rect 1562 54 1618 55
rect 1648 107 1704 110
rect 1734 107 1790 110
rect 1820 107 1876 110
rect 1906 107 1962 110
rect 1992 107 2048 110
rect 1648 55 1656 107
rect 1656 55 1704 107
rect 1734 55 1764 107
rect 1764 55 1790 107
rect 1820 55 1871 107
rect 1871 55 1876 107
rect 1906 55 1923 107
rect 1923 55 1962 107
rect 1992 55 2030 107
rect 2030 55 2048 107
rect 1648 54 1704 55
rect 1734 54 1790 55
rect 1820 54 1876 55
rect 1906 54 1962 55
rect 1992 54 2048 55
rect 2078 107 2134 110
rect 2078 55 2085 107
rect 2085 55 2134 107
rect 2078 54 2134 55
rect 2788 1034 2837 1086
rect 2837 1034 2844 1086
rect 2889 1034 2909 1086
rect 2909 1034 2928 1086
rect 2928 1034 2945 1086
rect 2990 1034 2999 1086
rect 2999 1034 3046 1086
rect 3091 1034 3122 1086
rect 3122 1034 3141 1086
rect 3141 1034 3147 1086
rect 3192 1034 3193 1086
rect 3193 1034 3212 1086
rect 3212 1034 3248 1086
rect 3293 1034 3335 1086
rect 3335 1034 3349 1086
rect 2788 1031 2844 1034
rect 2889 1031 2945 1034
rect 2990 1031 3046 1034
rect 3091 1031 3147 1034
rect 3192 1031 3248 1034
rect 3293 1031 3349 1034
rect 2788 934 2844 937
rect 2889 934 2945 937
rect 2990 934 3046 937
rect 3091 934 3147 937
rect 3192 934 3248 937
rect 3293 934 3349 937
rect 2788 882 2837 934
rect 2837 882 2844 934
rect 2889 882 2909 934
rect 2909 882 2928 934
rect 2928 882 2945 934
rect 2990 882 2999 934
rect 2999 882 3046 934
rect 3091 882 3122 934
rect 3122 882 3141 934
rect 3141 882 3147 934
rect 3192 882 3193 934
rect 3193 882 3212 934
rect 3212 882 3248 934
rect 3293 882 3335 934
rect 3335 882 3349 934
rect 2788 881 2844 882
rect 2889 881 2945 882
rect 2990 881 3046 882
rect 3091 881 3147 882
rect 3192 881 3248 882
rect 3293 881 3349 882
rect 4857 1651 4913 1653
rect 4940 1651 4996 1653
rect 5023 1651 5079 1653
rect 5106 1651 5162 1653
rect 5188 1651 5244 1653
rect 4857 1599 4906 1651
rect 4906 1599 4913 1651
rect 4940 1599 4975 1651
rect 4975 1599 4991 1651
rect 4991 1599 4996 1651
rect 5023 1599 5043 1651
rect 5043 1599 5059 1651
rect 5059 1599 5079 1651
rect 5106 1599 5111 1651
rect 5111 1599 5127 1651
rect 5127 1599 5162 1651
rect 5188 1599 5195 1651
rect 5195 1599 5244 1651
rect 4857 1597 4913 1599
rect 4940 1597 4996 1599
rect 5023 1597 5079 1599
rect 5106 1597 5162 1599
rect 5188 1597 5244 1599
rect 4857 1503 4913 1507
rect 4940 1503 4996 1507
rect 5023 1503 5079 1507
rect 5106 1503 5162 1507
rect 5188 1503 5244 1507
rect 4857 1451 4906 1503
rect 4906 1451 4913 1503
rect 4940 1451 4975 1503
rect 4975 1451 4991 1503
rect 4991 1451 4996 1503
rect 5023 1451 5043 1503
rect 5043 1451 5059 1503
rect 5059 1451 5079 1503
rect 5106 1451 5111 1503
rect 5111 1451 5127 1503
rect 5127 1451 5162 1503
rect 5188 1451 5195 1503
rect 5195 1451 5244 1503
rect 4862 713 5238 1409
rect 6847 3089 6903 3145
rect 6931 3089 6987 3145
rect 7015 3089 7071 3145
rect 6847 2966 6903 3022
rect 6931 2966 6987 3022
rect 7015 2966 7071 3022
rect 6847 2843 6903 2899
rect 6931 2843 6987 2899
rect 7015 2843 7071 2899
rect 6847 2720 6903 2776
rect 6931 2720 6987 2776
rect 7015 2720 7071 2776
rect 6847 2597 6903 2653
rect 6931 2597 6987 2653
rect 7015 2597 7071 2653
rect 6847 2474 6903 2530
rect 6931 2474 6987 2530
rect 7015 2474 7071 2530
rect 6847 2351 6903 2407
rect 6931 2351 6987 2407
rect 7015 2351 7071 2407
rect 6847 2228 6903 2284
rect 6931 2228 6987 2284
rect 7015 2228 7071 2284
rect 8615 3089 8671 3145
rect 8719 3089 8775 3145
rect 8615 2967 8671 3023
rect 8719 2967 8775 3023
rect 8615 2845 8671 2901
rect 8719 2845 8775 2901
rect 8615 2723 8671 2779
rect 8719 2723 8775 2779
rect 8615 2601 8671 2657
rect 8719 2601 8775 2657
rect 8615 2479 8671 2535
rect 8719 2479 8775 2535
rect 10522 2595 10564 2637
rect 10564 2595 10578 2637
rect 10614 2595 10631 2637
rect 10631 2595 10670 2637
rect 10522 2581 10578 2595
rect 10614 2581 10670 2595
rect 10706 2595 10707 2637
rect 10707 2595 10759 2637
rect 10759 2595 10762 2637
rect 10798 2595 10832 2637
rect 10832 2595 10853 2637
rect 10853 2595 10854 2637
rect 10890 2595 10905 2637
rect 10905 2595 10926 2637
rect 10926 2595 10946 2637
rect 10982 2595 10999 2637
rect 10999 2595 11038 2637
rect 10706 2581 10762 2595
rect 10798 2581 10854 2595
rect 10890 2581 10946 2595
rect 10982 2581 11038 2595
rect 10522 2503 10578 2515
rect 10614 2503 10670 2515
rect 10522 2459 10564 2503
rect 10564 2459 10578 2503
rect 10614 2459 10631 2503
rect 10631 2459 10670 2503
rect 10706 2503 10762 2515
rect 10798 2503 10854 2515
rect 10890 2503 10946 2515
rect 10982 2503 11038 2515
rect 10706 2459 10707 2503
rect 10707 2459 10759 2503
rect 10759 2459 10762 2503
rect 10798 2459 10832 2503
rect 10832 2459 10853 2503
rect 10853 2459 10854 2503
rect 10890 2459 10905 2503
rect 10905 2459 10926 2503
rect 10926 2459 10946 2503
rect 10982 2459 10999 2503
rect 10999 2459 11038 2503
rect 8615 2356 8671 2412
rect 8719 2356 8775 2412
rect 6847 2105 6903 2161
rect 6931 2105 6987 2161
rect 7015 2105 7071 2161
rect 6847 1982 6903 2038
rect 6931 1982 6987 2038
rect 7015 1982 7071 2038
rect 6847 1859 6903 1915
rect 6931 1859 6987 1915
rect 7015 1859 7071 1915
rect 8615 2233 8671 2289
rect 8719 2233 8775 2289
rect 8615 2110 8671 2166
rect 8719 2110 8775 2166
rect 8615 1987 8671 2043
rect 8719 1987 8775 2043
rect 4862 632 4918 688
rect 4942 632 4998 688
rect 5022 632 5078 688
rect 5102 632 5158 688
rect 5182 632 5238 688
rect 4862 551 4918 607
rect 4942 551 4998 607
rect 5022 551 5078 607
rect 5102 551 5158 607
rect 5182 551 5238 607
rect 4862 470 4918 526
rect 4942 470 4998 526
rect 5022 470 5078 526
rect 5102 470 5158 526
rect 5182 470 5238 526
rect 4862 389 4918 445
rect 4942 389 4998 445
rect 5022 389 5078 445
rect 5102 389 5158 445
rect 5182 389 5238 445
rect 4862 308 4918 364
rect 4942 308 4998 364
rect 5022 308 5078 364
rect 5102 308 5158 364
rect 5182 308 5238 364
rect 4608 256 4664 257
rect 4691 256 4747 257
rect 4774 256 4830 257
rect 4608 204 4660 256
rect 4660 204 4664 256
rect 4691 204 4712 256
rect 4712 204 4747 256
rect 4774 204 4819 256
rect 4819 204 4830 256
rect 4608 201 4664 204
rect 4691 201 4747 204
rect 4774 201 4830 204
rect 4857 256 4913 257
rect 4940 256 4996 257
rect 5023 256 5079 257
rect 5106 256 5162 257
rect 4857 204 4874 256
rect 4874 204 4913 256
rect 4940 204 4981 256
rect 4981 204 4996 256
rect 5023 204 5033 256
rect 5033 204 5079 256
rect 5106 204 5140 256
rect 5140 204 5162 256
rect 4857 201 4913 204
rect 4940 201 4996 204
rect 5023 201 5079 204
rect 5106 201 5162 204
rect 5188 256 5244 257
rect 5188 204 5195 256
rect 5195 204 5244 256
rect 5188 201 5244 204
rect 4608 108 4664 111
rect 4691 108 4747 111
rect 4774 108 4830 111
rect 4608 56 4660 108
rect 4660 56 4664 108
rect 4691 56 4712 108
rect 4712 56 4747 108
rect 4774 56 4819 108
rect 4819 56 4830 108
rect 4608 55 4664 56
rect 4691 55 4747 56
rect 4774 55 4830 56
rect 4857 108 4913 111
rect 4940 108 4996 111
rect 5023 108 5079 111
rect 5106 108 5162 111
rect 4857 56 4874 108
rect 4874 56 4913 108
rect 4940 56 4981 108
rect 4981 56 4996 108
rect 5023 56 5033 108
rect 5033 56 5079 108
rect 5106 56 5140 108
rect 5140 56 5162 108
rect 4857 55 4913 56
rect 4940 55 4996 56
rect 5023 55 5079 56
rect 5106 55 5162 56
rect 5188 108 5244 111
rect 5188 56 5195 108
rect 5195 56 5244 108
rect 5188 55 5244 56
rect 9776 709 9828 758
rect 9828 709 9832 758
rect 9776 702 9832 709
rect 9776 645 9828 678
rect 9828 645 9832 678
rect 9776 622 9832 645
rect 10519 1038 10563 1076
rect 10563 1038 10575 1076
rect 10600 1038 10629 1076
rect 10629 1038 10643 1076
rect 10643 1038 10656 1076
rect 10681 1038 10695 1076
rect 10695 1038 10708 1076
rect 10708 1038 10737 1076
rect 10763 1038 10773 1076
rect 10773 1038 10819 1076
rect 15594 1430 15650 1486
rect 15594 1348 15650 1404
rect 15594 1266 15650 1322
rect 10519 1020 10575 1038
rect 10600 1020 10656 1038
rect 10681 1020 10737 1038
rect 10763 1020 10819 1038
rect 10519 958 10563 994
rect 10563 958 10575 994
rect 10600 958 10629 994
rect 10629 958 10643 994
rect 10643 958 10656 994
rect 10681 958 10695 994
rect 10695 958 10708 994
rect 10708 958 10737 994
rect 10763 958 10773 994
rect 10773 958 10819 994
rect 10519 938 10575 958
rect 10600 938 10656 958
rect 10681 938 10737 958
rect 10763 938 10819 958
rect 10519 878 10563 912
rect 10563 878 10575 912
rect 10600 878 10629 912
rect 10629 878 10643 912
rect 10643 878 10656 912
rect 10681 878 10695 912
rect 10695 878 10708 912
rect 10708 878 10737 912
rect 10763 878 10773 912
rect 10773 878 10819 912
rect 10519 856 10575 878
rect 10600 856 10656 878
rect 10681 856 10737 878
rect 10763 856 10819 878
rect 10519 774 10575 830
rect 10600 774 10656 830
rect 10681 774 10737 830
rect 10763 774 10819 830
rect 10519 692 10575 748
rect 10600 692 10656 748
rect 10681 692 10737 748
rect 10763 692 10819 748
rect 10519 610 10575 666
rect 10600 610 10656 666
rect 10681 610 10737 666
rect 10763 610 10819 666
rect 9888 374 9944 430
rect 9968 374 10024 430
rect 10519 528 10575 584
rect 10600 528 10656 584
rect 10681 528 10737 584
rect 10763 528 10819 584
rect 13012 483 13068 539
rect 13102 483 13158 539
rect 10347 237 10403 293
rect 10427 237 10483 293
rect 13317 239 13373 295
rect 13407 239 13463 295
rect 9927 109 9983 165
rect 10007 109 10063 165
rect 15487 237 15543 293
rect 15577 237 15633 293
<< metal3 >>
rect 1054 39995 11350 40000
rect 1054 39950 1903 39995
rect 1054 39894 1361 39950
rect 1417 39894 1443 39950
rect 1499 39894 1525 39950
rect 1581 39894 1607 39950
rect 1663 39894 1689 39950
rect 1745 39939 1903 39950
rect 1959 39939 1984 39995
rect 2040 39939 2065 39995
rect 2121 39939 2146 39995
rect 2202 39939 2227 39995
rect 2283 39939 2308 39995
rect 2364 39939 2389 39995
rect 2445 39939 2470 39995
rect 2526 39939 2551 39995
rect 2607 39939 2632 39995
rect 2688 39939 2713 39995
rect 2769 39939 2794 39995
rect 2850 39939 2875 39995
rect 2931 39939 2956 39995
rect 3012 39939 3037 39995
rect 3093 39939 3118 39995
rect 1745 39915 3118 39939
rect 1745 39894 1903 39915
rect 1054 39868 1903 39894
rect 1054 39812 1361 39868
rect 1417 39812 1443 39868
rect 1499 39812 1525 39868
rect 1581 39812 1607 39868
rect 1663 39812 1689 39868
rect 1745 39859 1903 39868
rect 1959 39859 1984 39915
rect 2040 39859 2065 39915
rect 2121 39859 2146 39915
rect 2202 39859 2227 39915
rect 2283 39859 2308 39915
rect 2364 39859 2389 39915
rect 2445 39859 2470 39915
rect 2526 39859 2551 39915
rect 2607 39859 2632 39915
rect 2688 39859 2713 39915
rect 2769 39859 2794 39915
rect 2850 39859 2875 39915
rect 2931 39859 2956 39915
rect 3012 39859 3037 39915
rect 3093 39859 3118 39915
rect 1745 39835 3118 39859
rect 1745 39812 1903 39835
rect 1054 39786 1903 39812
rect 1054 39730 1361 39786
rect 1417 39730 1443 39786
rect 1499 39730 1525 39786
rect 1581 39730 1607 39786
rect 1663 39730 1689 39786
rect 1745 39779 1903 39786
rect 1959 39779 1984 39835
rect 2040 39779 2065 39835
rect 2121 39779 2146 39835
rect 2202 39779 2227 39835
rect 2283 39779 2308 39835
rect 2364 39779 2389 39835
rect 2445 39779 2470 39835
rect 2526 39779 2551 39835
rect 2607 39779 2632 39835
rect 2688 39779 2713 39835
rect 2769 39779 2794 39835
rect 2850 39779 2875 39835
rect 2931 39779 2956 39835
rect 3012 39779 3037 39835
rect 3093 39779 3118 39835
rect 1745 39755 3118 39779
rect 1745 39730 1903 39755
rect 1054 39704 1903 39730
rect 1054 39648 1361 39704
rect 1417 39648 1443 39704
rect 1499 39648 1525 39704
rect 1581 39648 1607 39704
rect 1663 39648 1689 39704
rect 1745 39699 1903 39704
rect 1959 39699 1984 39755
rect 2040 39699 2065 39755
rect 2121 39699 2146 39755
rect 2202 39699 2227 39755
rect 2283 39699 2308 39755
rect 2364 39699 2389 39755
rect 2445 39699 2470 39755
rect 2526 39699 2551 39755
rect 2607 39699 2632 39755
rect 2688 39699 2713 39755
rect 2769 39699 2794 39755
rect 2850 39699 2875 39755
rect 2931 39699 2956 39755
rect 3012 39699 3037 39755
rect 3093 39699 3118 39755
rect 1745 39675 3118 39699
rect 1745 39648 1903 39675
rect 1054 39622 1903 39648
rect 1054 39566 1361 39622
rect 1417 39566 1443 39622
rect 1499 39566 1525 39622
rect 1581 39566 1607 39622
rect 1663 39566 1689 39622
rect 1745 39619 1903 39622
rect 1959 39619 1984 39675
rect 2040 39619 2065 39675
rect 2121 39619 2146 39675
rect 2202 39619 2227 39675
rect 2283 39619 2308 39675
rect 2364 39619 2389 39675
rect 2445 39619 2470 39675
rect 2526 39619 2551 39675
rect 2607 39619 2632 39675
rect 2688 39619 2713 39675
rect 2769 39619 2794 39675
rect 2850 39619 2875 39675
rect 2931 39619 2956 39675
rect 3012 39619 3037 39675
rect 3093 39619 3118 39675
rect 1745 39595 3118 39619
rect 1745 39566 1903 39595
rect 1054 39540 1903 39566
rect 1054 39484 1361 39540
rect 1417 39484 1443 39540
rect 1499 39484 1525 39540
rect 1581 39484 1607 39540
rect 1663 39484 1689 39540
rect 1745 39539 1903 39540
rect 1959 39539 1984 39595
rect 2040 39539 2065 39595
rect 2121 39539 2146 39595
rect 2202 39539 2227 39595
rect 2283 39539 2308 39595
rect 2364 39539 2389 39595
rect 2445 39539 2470 39595
rect 2526 39539 2551 39595
rect 2607 39539 2632 39595
rect 2688 39539 2713 39595
rect 2769 39539 2794 39595
rect 2850 39539 2875 39595
rect 2931 39539 2956 39595
rect 3012 39539 3037 39595
rect 3093 39539 3118 39595
rect 11334 39539 11350 39995
rect 1745 39519 11350 39539
rect 14399 39995 15371 40000
rect 14399 39939 14411 39995
rect 14467 39939 14492 39995
rect 14548 39939 14573 39995
rect 14629 39939 14654 39995
rect 14710 39939 14735 39995
rect 14791 39939 14816 39995
rect 14872 39939 14897 39995
rect 14953 39939 14977 39995
rect 15033 39939 15057 39995
rect 15113 39939 15137 39995
rect 15193 39939 15217 39995
rect 15273 39939 15297 39995
rect 15353 39939 15371 39995
rect 14399 39899 15371 39939
rect 14399 39843 14411 39899
rect 14467 39843 14492 39899
rect 14548 39843 14573 39899
rect 14629 39843 14654 39899
rect 14710 39843 14735 39899
rect 14791 39843 14816 39899
rect 14872 39843 14897 39899
rect 14953 39843 14977 39899
rect 15033 39843 15057 39899
rect 15113 39843 15137 39899
rect 15193 39843 15217 39899
rect 15273 39843 15297 39899
rect 15353 39843 15371 39899
rect 14399 39803 15371 39843
rect 14399 39747 14411 39803
rect 14467 39747 14492 39803
rect 14548 39747 14573 39803
rect 14629 39747 14654 39803
rect 14710 39747 14735 39803
rect 14791 39747 14816 39803
rect 14872 39747 14897 39803
rect 14953 39747 14977 39803
rect 15033 39747 15057 39803
rect 15113 39747 15137 39803
rect 15193 39747 15217 39803
rect 15273 39747 15297 39803
rect 15353 39747 15371 39803
rect 1745 39484 2415 39519
rect 1054 39458 2415 39484
rect 1054 39402 1361 39458
rect 1417 39402 1443 39458
rect 1499 39402 1525 39458
rect 1581 39402 1607 39458
rect 1663 39402 1689 39458
rect 1745 39402 2415 39458
rect 1054 39389 2415 39402
tri 2415 39389 2545 39519 nw
rect 1054 39376 2397 39389
rect 1054 39320 1361 39376
rect 1417 39320 1443 39376
rect 1499 39320 1525 39376
rect 1581 39320 1607 39376
rect 1663 39320 1689 39376
rect 1745 39371 2397 39376
tri 2397 39371 2415 39389 nw
rect 12587 39372 13005 39389
rect 1745 39320 2054 39371
rect 1054 39294 2054 39320
rect 1054 39238 1361 39294
rect 1417 39238 1443 39294
rect 1499 39238 1525 39294
rect 1581 39238 1607 39294
rect 1663 39238 1689 39294
rect 1745 39238 2054 39294
rect 1054 39212 2054 39238
rect 1054 39156 1361 39212
rect 1417 39156 1443 39212
rect 1499 39156 1525 39212
rect 1581 39156 1607 39212
rect 1663 39156 1689 39212
rect 1745 39156 2054 39212
rect 1054 39130 2054 39156
rect 1054 39074 1361 39130
rect 1417 39074 1443 39130
rect 1499 39074 1525 39130
rect 1581 39074 1607 39130
rect 1663 39074 1689 39130
rect 1745 39074 2054 39130
rect 1054 39048 2054 39074
rect 1054 38992 1361 39048
rect 1417 38992 1443 39048
rect 1499 38992 1525 39048
rect 1581 38992 1607 39048
rect 1663 38992 1689 39048
rect 1745 38992 2054 39048
tri 2054 39028 2397 39371 nw
rect 5106 39365 6298 39371
rect 5106 39301 5110 39365
rect 5174 39301 5190 39365
rect 5254 39301 5270 39365
rect 5334 39301 5350 39365
rect 5414 39301 5430 39365
rect 5494 39301 5510 39365
rect 5574 39301 5590 39365
rect 5654 39301 5670 39365
rect 5734 39301 5750 39365
rect 5814 39301 5830 39365
rect 5894 39301 5910 39365
rect 5974 39301 5990 39365
rect 6054 39301 6070 39365
rect 6134 39301 6150 39365
rect 6214 39301 6230 39365
rect 6294 39301 6298 39365
rect 5106 39284 6298 39301
rect 5106 39220 5110 39284
rect 5174 39220 5190 39284
rect 5254 39220 5270 39284
rect 5334 39220 5350 39284
rect 5414 39220 5430 39284
rect 5494 39220 5510 39284
rect 5574 39220 5590 39284
rect 5654 39220 5670 39284
rect 5734 39220 5750 39284
rect 5814 39220 5830 39284
rect 5894 39220 5910 39284
rect 5974 39220 5990 39284
rect 6054 39220 6070 39284
rect 6134 39220 6150 39284
rect 6214 39220 6230 39284
rect 6294 39220 6298 39284
rect 5106 39203 6298 39220
rect 5106 39139 5110 39203
rect 5174 39139 5190 39203
rect 5254 39139 5270 39203
rect 5334 39139 5350 39203
rect 5414 39139 5430 39203
rect 5494 39139 5510 39203
rect 5574 39139 5590 39203
rect 5654 39139 5670 39203
rect 5734 39139 5750 39203
rect 5814 39139 5830 39203
rect 5894 39139 5910 39203
rect 5974 39139 5990 39203
rect 6054 39139 6070 39203
rect 6134 39139 6150 39203
rect 6214 39139 6230 39203
rect 6294 39139 6298 39203
rect 5106 39122 6298 39139
rect 5106 39058 5110 39122
rect 5174 39058 5190 39122
rect 5254 39058 5270 39122
rect 5334 39058 5350 39122
rect 5414 39058 5430 39122
rect 5494 39058 5510 39122
rect 5574 39058 5590 39122
rect 5654 39058 5670 39122
rect 5734 39058 5750 39122
rect 5814 39058 5830 39122
rect 5894 39058 5910 39122
rect 5974 39058 5990 39122
rect 6054 39058 6070 39122
rect 6134 39058 6150 39122
rect 6214 39058 6230 39122
rect 6294 39058 6298 39122
rect 5106 39041 6298 39058
rect 1054 38966 2054 38992
rect 1054 38910 1361 38966
rect 1417 38910 1443 38966
rect 1499 38910 1525 38966
rect 1581 38910 1607 38966
rect 1663 38910 1689 38966
rect 1745 38910 2054 38966
rect 1054 38884 2054 38910
rect 1054 38828 1361 38884
rect 1417 38828 1443 38884
rect 1499 38828 1525 38884
rect 1581 38828 1607 38884
rect 1663 38828 1689 38884
rect 1745 38828 2054 38884
rect 1054 38802 2054 38828
rect 1054 38746 1361 38802
rect 1417 38746 1443 38802
rect 1499 38746 1525 38802
rect 1581 38746 1607 38802
rect 1663 38746 1689 38802
rect 1745 38746 2054 38802
rect 1054 38720 2054 38746
rect 1054 38664 1361 38720
rect 1417 38664 1443 38720
rect 1499 38664 1525 38720
rect 1581 38664 1607 38720
rect 1663 38664 1689 38720
rect 1745 38664 2054 38720
rect 1054 38638 2054 38664
rect 1054 38582 1361 38638
rect 1417 38582 1443 38638
rect 1499 38582 1525 38638
rect 1581 38582 1607 38638
rect 1663 38582 1689 38638
rect 1745 38582 2054 38638
rect 1054 38556 2054 38582
rect 1054 38500 1361 38556
rect 1417 38500 1443 38556
rect 1499 38500 1525 38556
rect 1581 38500 1607 38556
rect 1663 38500 1689 38556
rect 1745 38500 2054 38556
rect 1054 38474 2054 38500
rect 1054 38418 1361 38474
rect 1417 38418 1443 38474
rect 1499 38418 1525 38474
rect 1581 38418 1607 38474
rect 1663 38418 1689 38474
rect 1745 38418 2054 38474
rect 1054 38392 2054 38418
rect 1054 38336 1361 38392
rect 1417 38336 1443 38392
rect 1499 38336 1525 38392
rect 1581 38336 1607 38392
rect 1663 38336 1689 38392
rect 1745 38336 2054 38392
rect 1054 38310 2054 38336
rect 1054 38254 1361 38310
rect 1417 38254 1443 38310
rect 1499 38254 1525 38310
rect 1581 38254 1607 38310
rect 1663 38254 1689 38310
rect 1745 38254 2054 38310
rect 1054 38228 2054 38254
rect 1054 38172 1361 38228
rect 1417 38172 1443 38228
rect 1499 38172 1525 38228
rect 1581 38172 1607 38228
rect 1663 38172 1689 38228
rect 1745 38172 2054 38228
rect 1054 38146 2054 38172
rect 1054 38090 1361 38146
rect 1417 38090 1443 38146
rect 1499 38090 1525 38146
rect 1581 38090 1607 38146
rect 1663 38090 1689 38146
rect 1745 38090 2054 38146
rect 1054 38064 2054 38090
rect 1054 38008 1361 38064
rect 1417 38008 1443 38064
rect 1499 38008 1525 38064
rect 1581 38008 1607 38064
rect 1663 38008 1689 38064
rect 1745 38008 2054 38064
rect 1054 37981 2054 38008
rect 1054 37925 1361 37981
rect 1417 37925 1443 37981
rect 1499 37925 1525 37981
rect 1581 37925 1607 37981
rect 1663 37925 1689 37981
rect 1745 37925 2054 37981
rect 1054 37898 2054 37925
rect 1054 37842 1361 37898
rect 1417 37842 1443 37898
rect 1499 37842 1525 37898
rect 1581 37842 1607 37898
rect 1663 37842 1689 37898
rect 1745 37842 2054 37898
rect 1054 37815 2054 37842
rect 1054 37759 1361 37815
rect 1417 37759 1443 37815
rect 1499 37759 1525 37815
rect 1581 37759 1607 37815
rect 1663 37759 1689 37815
rect 1745 37759 2054 37815
rect 1054 37732 2054 37759
rect 1054 37676 1361 37732
rect 1417 37676 1443 37732
rect 1499 37676 1525 37732
rect 1581 37676 1607 37732
rect 1663 37676 1689 37732
rect 1745 37676 2054 37732
rect 1054 37649 2054 37676
rect 1054 37593 1361 37649
rect 1417 37593 1443 37649
rect 1499 37593 1525 37649
rect 1581 37593 1607 37649
rect 1663 37593 1689 37649
rect 1745 37593 2054 37649
rect 1054 37566 2054 37593
rect 1054 37510 1361 37566
rect 1417 37510 1443 37566
rect 1499 37510 1525 37566
rect 1581 37510 1607 37566
rect 1663 37510 1689 37566
rect 1745 37510 2054 37566
rect 1054 37483 2054 37510
rect 1054 37427 1361 37483
rect 1417 37427 1443 37483
rect 1499 37427 1525 37483
rect 1581 37427 1607 37483
rect 1663 37427 1689 37483
rect 1745 37427 2054 37483
rect 1054 37400 2054 37427
rect 1054 37344 1361 37400
rect 1417 37344 1443 37400
rect 1499 37344 1525 37400
rect 1581 37344 1607 37400
rect 1663 37344 1689 37400
rect 1745 37344 2054 37400
rect 1054 37317 2054 37344
rect 1054 37261 1361 37317
rect 1417 37261 1443 37317
rect 1499 37261 1525 37317
rect 1581 37261 1607 37317
rect 1663 37261 1689 37317
rect 1745 37261 2054 37317
rect 1054 37234 2054 37261
rect 1054 37178 1361 37234
rect 1417 37178 1443 37234
rect 1499 37178 1525 37234
rect 1581 37178 1607 37234
rect 1663 37178 1689 37234
rect 1745 37178 2054 37234
tri 612 36229 617 36234 se
rect 617 36229 913 36234
tri 556 36173 612 36229 se
rect 612 36173 837 36229
rect 893 36173 913 36229
tri 532 36149 556 36173 se
rect 556 36149 913 36173
tri 476 36093 532 36149 se
rect 532 36093 837 36149
rect 893 36093 913 36149
tri 464 36081 476 36093 se
rect 476 36088 913 36093
rect 476 36081 638 36088
tri 638 36081 645 36088 nw
tri 443 36060 464 36081 se
rect 464 36060 617 36081
tri 617 36060 638 36081 nw
tri 408 36025 443 36060 se
rect 443 36025 582 36060
tri 582 36025 617 36060 nw
tri 346 35963 408 36025 se
rect 408 35963 520 36025
tri 520 35963 582 36025 nw
tri 290 35907 346 35963 se
rect 346 35907 464 35963
tri 464 35907 520 35963 nw
tri 269 35886 290 35907 se
rect 290 35886 443 35907
tri 443 35886 464 35907 nw
tri 228 35845 269 35886 se
rect 269 35845 402 35886
tri 402 35845 443 35886 nw
tri 172 35789 228 35845 se
rect 228 35789 346 35845
tri 346 35789 402 35845 nw
tri 95 35712 172 35789 se
rect 172 35712 269 35789
tri 269 35712 346 35789 nw
tri 80 35697 95 35712 se
rect 95 35697 254 35712
tri 254 35697 269 35712 nw
rect 80 0 204 35697
tri 204 35647 254 35697 nw
rect 292 35618 656 35629
rect 292 35562 298 35618
rect 354 35562 396 35618
rect 452 35562 494 35618
rect 550 35562 592 35618
rect 648 35562 656 35618
rect 292 35538 656 35562
rect 292 35482 298 35538
rect 354 35482 396 35538
rect 452 35482 494 35538
rect 550 35482 592 35538
rect 648 35482 656 35538
rect 292 35458 656 35482
rect 292 35402 298 35458
rect 354 35402 396 35458
rect 452 35402 494 35458
rect 550 35402 592 35458
rect 648 35402 656 35458
rect 292 35378 656 35402
rect 292 35322 298 35378
rect 354 35322 396 35378
rect 452 35322 494 35378
rect 550 35322 592 35378
rect 648 35322 656 35378
rect 292 35298 656 35322
rect 292 35242 298 35298
rect 354 35242 396 35298
rect 452 35242 494 35298
rect 550 35242 592 35298
rect 648 35242 656 35298
rect 292 35218 656 35242
rect 292 35162 298 35218
rect 354 35162 396 35218
rect 452 35162 494 35218
rect 550 35162 592 35218
rect 648 35162 656 35218
rect 292 35138 656 35162
rect 292 35082 298 35138
rect 354 35082 396 35138
rect 452 35082 494 35138
rect 550 35082 592 35138
rect 648 35082 656 35138
rect 292 35058 656 35082
rect 292 35002 298 35058
rect 354 35002 396 35058
rect 452 35002 494 35058
rect 550 35002 592 35058
rect 648 35002 656 35058
rect 292 34978 656 35002
rect 292 34922 298 34978
rect 354 34922 396 34978
rect 452 34922 494 34978
rect 550 34922 592 34978
rect 648 34922 656 34978
rect 292 34898 656 34922
rect 292 34842 298 34898
rect 354 34842 396 34898
rect 452 34842 494 34898
rect 550 34842 592 34898
rect 648 34842 656 34898
rect 292 34818 656 34842
rect 292 34762 298 34818
rect 354 34762 396 34818
rect 452 34762 494 34818
rect 550 34762 592 34818
rect 648 34762 656 34818
rect 292 34738 656 34762
rect 292 34682 298 34738
rect 354 34682 396 34738
rect 452 34682 494 34738
rect 550 34682 592 34738
rect 648 34682 656 34738
rect 292 34658 656 34682
rect 292 34602 298 34658
rect 354 34602 396 34658
rect 452 34602 494 34658
rect 550 34602 592 34658
rect 648 34602 656 34658
rect 292 34578 656 34602
rect 292 34522 298 34578
rect 354 34522 396 34578
rect 452 34522 494 34578
rect 550 34522 592 34578
rect 648 34522 656 34578
rect 292 34498 656 34522
rect 292 34442 298 34498
rect 354 34442 396 34498
rect 452 34442 494 34498
rect 550 34442 592 34498
rect 648 34442 656 34498
rect 292 34418 656 34442
rect 292 34362 298 34418
rect 354 34362 396 34418
rect 452 34362 494 34418
rect 550 34362 592 34418
rect 648 34362 656 34418
rect 292 34338 656 34362
rect 292 34282 298 34338
rect 354 34282 396 34338
rect 452 34282 494 34338
rect 550 34282 592 34338
rect 648 34282 656 34338
rect 292 34258 656 34282
rect 292 34202 298 34258
rect 354 34202 396 34258
rect 452 34202 494 34258
rect 550 34202 592 34258
rect 648 34202 656 34258
rect 292 34178 656 34202
rect 292 34122 298 34178
rect 354 34122 396 34178
rect 452 34122 494 34178
rect 550 34122 592 34178
rect 648 34122 656 34178
rect 292 34098 656 34122
rect 292 34042 298 34098
rect 354 34042 396 34098
rect 452 34042 494 34098
rect 550 34042 592 34098
rect 648 34042 656 34098
rect 292 34018 656 34042
rect 292 33962 298 34018
rect 354 33962 396 34018
rect 452 33962 494 34018
rect 550 33962 592 34018
rect 648 33962 656 34018
rect 292 33938 656 33962
rect 292 33882 298 33938
rect 354 33882 396 33938
rect 452 33882 494 33938
rect 550 33882 592 33938
rect 648 33882 656 33938
rect 292 33858 656 33882
rect 292 33802 298 33858
rect 354 33802 396 33858
rect 452 33802 494 33858
rect 550 33802 592 33858
rect 648 33802 656 33858
rect 292 33778 656 33802
rect 292 33722 298 33778
rect 354 33722 396 33778
rect 452 33722 494 33778
rect 550 33722 592 33778
rect 648 33722 656 33778
rect 292 33698 656 33722
rect 292 33642 298 33698
rect 354 33642 396 33698
rect 452 33642 494 33698
rect 550 33642 592 33698
rect 648 33642 656 33698
rect 292 33618 656 33642
rect 292 33562 298 33618
rect 354 33562 396 33618
rect 452 33562 494 33618
rect 550 33562 592 33618
rect 648 33562 656 33618
rect 292 33538 656 33562
rect 292 33482 298 33538
rect 354 33482 396 33538
rect 452 33482 494 33538
rect 550 33482 592 33538
rect 648 33482 656 33538
rect 292 33458 656 33482
rect 292 33402 298 33458
rect 354 33402 396 33458
rect 452 33402 494 33458
rect 550 33402 592 33458
rect 648 33402 656 33458
rect 292 33378 656 33402
rect 292 33322 298 33378
rect 354 33322 396 33378
rect 452 33322 494 33378
rect 550 33322 592 33378
rect 648 33322 656 33378
rect 292 33298 656 33322
rect 292 33242 298 33298
rect 354 33242 396 33298
rect 452 33242 494 33298
rect 550 33242 592 33298
rect 648 33242 656 33298
rect 292 33218 656 33242
rect 292 33162 298 33218
rect 354 33162 396 33218
rect 452 33162 494 33218
rect 550 33162 592 33218
rect 648 33162 656 33218
rect 292 33138 656 33162
rect 292 33082 298 33138
rect 354 33082 396 33138
rect 452 33082 494 33138
rect 550 33082 592 33138
rect 648 33082 656 33138
rect 292 33058 656 33082
rect 292 33002 298 33058
rect 354 33002 396 33058
rect 452 33002 494 33058
rect 550 33002 592 33058
rect 648 33002 656 33058
rect 292 32978 656 33002
rect 292 32922 298 32978
rect 354 32922 396 32978
rect 452 32922 494 32978
rect 550 32922 592 32978
rect 648 32922 656 32978
rect 292 32898 656 32922
rect 292 32842 298 32898
rect 354 32842 396 32898
rect 452 32842 494 32898
rect 550 32842 592 32898
rect 648 32842 656 32898
rect 292 32818 656 32842
rect 292 32762 298 32818
rect 354 32762 396 32818
rect 452 32762 494 32818
rect 550 32762 592 32818
rect 648 32762 656 32818
rect 292 32738 656 32762
rect 292 32682 298 32738
rect 354 32682 396 32738
rect 452 32682 494 32738
rect 550 32682 592 32738
rect 648 32682 656 32738
rect 292 32658 656 32682
rect 292 32602 298 32658
rect 354 32602 396 32658
rect 452 32602 494 32658
rect 550 32602 592 32658
rect 648 32602 656 32658
rect 292 32578 656 32602
rect 292 32522 298 32578
rect 354 32522 396 32578
rect 452 32522 494 32578
rect 550 32522 592 32578
rect 648 32522 656 32578
rect 292 32498 656 32522
rect 292 32442 298 32498
rect 354 32442 396 32498
rect 452 32442 494 32498
rect 550 32442 592 32498
rect 648 32442 656 32498
rect 292 32418 656 32442
rect 292 32362 298 32418
rect 354 32362 396 32418
rect 452 32362 494 32418
rect 550 32362 592 32418
rect 648 32362 656 32418
rect 292 32338 656 32362
rect 292 32282 298 32338
rect 354 32282 396 32338
rect 452 32282 494 32338
rect 550 32282 592 32338
rect 648 32282 656 32338
rect 292 32258 656 32282
rect 292 32202 298 32258
rect 354 32202 396 32258
rect 452 32202 494 32258
rect 550 32202 592 32258
rect 648 32202 656 32258
rect 292 32177 656 32202
rect 292 32121 298 32177
rect 354 32121 396 32177
rect 452 32121 494 32177
rect 550 32121 592 32177
rect 648 32121 656 32177
rect 292 32096 656 32121
rect 292 32040 298 32096
rect 354 32040 396 32096
rect 452 32040 494 32096
rect 550 32040 592 32096
rect 648 32040 656 32096
rect 292 32015 656 32040
rect 292 31959 298 32015
rect 354 31959 396 32015
rect 452 31959 494 32015
rect 550 31959 592 32015
rect 648 31959 656 32015
rect 292 31934 656 31959
rect 292 31878 298 31934
rect 354 31878 396 31934
rect 452 31878 494 31934
rect 550 31878 592 31934
rect 648 31878 656 31934
rect 292 31853 656 31878
rect 292 31797 298 31853
rect 354 31797 396 31853
rect 452 31797 494 31853
rect 550 31797 592 31853
rect 648 31797 656 31853
rect 292 31772 656 31797
rect 292 31716 298 31772
rect 354 31716 396 31772
rect 452 31716 494 31772
rect 550 31716 592 31772
rect 648 31716 656 31772
rect 292 31691 656 31716
rect 292 31635 298 31691
rect 354 31635 396 31691
rect 452 31635 494 31691
rect 550 31635 592 31691
rect 648 31635 656 31691
rect 292 31610 656 31635
rect 292 31554 298 31610
rect 354 31554 396 31610
rect 452 31554 494 31610
rect 550 31554 592 31610
rect 648 31554 656 31610
rect 292 31529 656 31554
rect 292 31473 298 31529
rect 354 31473 396 31529
rect 452 31473 494 31529
rect 550 31473 592 31529
rect 648 31473 656 31529
rect 292 31448 656 31473
rect 292 31392 298 31448
rect 354 31392 396 31448
rect 452 31392 494 31448
rect 550 31392 592 31448
rect 648 31392 656 31448
rect 292 31367 656 31392
rect 292 31311 298 31367
rect 354 31311 396 31367
rect 452 31311 494 31367
rect 550 31311 592 31367
rect 648 31311 656 31367
rect 292 31286 656 31311
rect 292 31230 298 31286
rect 354 31230 396 31286
rect 452 31230 494 31286
rect 550 31230 592 31286
rect 648 31230 656 31286
rect 292 31205 656 31230
rect 292 31149 298 31205
rect 354 31149 396 31205
rect 452 31149 494 31205
rect 550 31149 592 31205
rect 648 31149 656 31205
rect 292 31124 656 31149
rect 292 31068 298 31124
rect 354 31068 396 31124
rect 452 31068 494 31124
rect 550 31068 592 31124
rect 648 31068 656 31124
rect 292 31043 656 31068
rect 292 30987 298 31043
rect 354 30987 396 31043
rect 452 30987 494 31043
rect 550 30987 592 31043
rect 648 30987 656 31043
rect 292 30962 656 30987
rect 292 30906 298 30962
rect 354 30906 396 30962
rect 452 30906 494 30962
rect 550 30906 592 30962
rect 648 30906 656 30962
rect 292 30881 656 30906
rect 292 30825 298 30881
rect 354 30825 396 30881
rect 452 30825 494 30881
rect 550 30825 592 30881
rect 648 30825 656 30881
rect 292 30800 656 30825
rect 292 30744 298 30800
rect 354 30744 396 30800
rect 452 30744 494 30800
rect 550 30744 592 30800
rect 648 30744 656 30800
rect 292 30719 656 30744
rect 292 30663 298 30719
rect 354 30663 396 30719
rect 452 30663 494 30719
rect 550 30663 592 30719
rect 648 30663 656 30719
rect 292 30638 656 30663
rect 292 30582 298 30638
rect 354 30582 396 30638
rect 452 30582 494 30638
rect 550 30582 592 30638
rect 648 30582 656 30638
rect 292 30557 656 30582
rect 292 30501 298 30557
rect 354 30501 396 30557
rect 452 30501 494 30557
rect 550 30501 592 30557
rect 648 30501 656 30557
rect 292 30476 656 30501
rect 292 30420 298 30476
rect 354 30420 396 30476
rect 452 30420 494 30476
rect 550 30420 592 30476
rect 648 30420 656 30476
rect 292 30395 656 30420
rect 292 30339 298 30395
rect 354 30339 396 30395
rect 452 30339 494 30395
rect 550 30339 592 30395
rect 648 30339 656 30395
rect 292 30314 656 30339
rect 292 30258 298 30314
rect 354 30258 396 30314
rect 452 30258 494 30314
rect 550 30258 592 30314
rect 648 30258 656 30314
rect 292 30233 656 30258
rect 292 30177 298 30233
rect 354 30177 396 30233
rect 452 30177 494 30233
rect 550 30177 592 30233
rect 648 30177 656 30233
rect 292 30152 656 30177
rect 292 30096 298 30152
rect 354 30096 396 30152
rect 452 30096 494 30152
rect 550 30096 592 30152
rect 648 30096 656 30152
rect 292 30071 656 30096
rect 292 30015 298 30071
rect 354 30015 396 30071
rect 452 30015 494 30071
rect 550 30015 592 30071
rect 648 30015 656 30071
rect 292 29990 656 30015
rect 292 29934 298 29990
rect 354 29934 396 29990
rect 452 29934 494 29990
rect 550 29934 592 29990
rect 648 29934 656 29990
rect 292 29909 656 29934
rect 292 29853 298 29909
rect 354 29853 396 29909
rect 452 29853 494 29909
rect 550 29853 592 29909
rect 648 29853 656 29909
rect 292 29828 656 29853
rect 292 29772 298 29828
rect 354 29772 396 29828
rect 452 29772 494 29828
rect 550 29772 592 29828
rect 648 29772 656 29828
rect 292 29747 656 29772
rect 292 29691 298 29747
rect 354 29691 396 29747
rect 452 29691 494 29747
rect 550 29691 592 29747
rect 648 29691 656 29747
rect 292 29666 656 29691
rect 292 29610 298 29666
rect 354 29610 396 29666
rect 452 29610 494 29666
rect 550 29610 592 29666
rect 648 29610 656 29666
rect 292 29585 656 29610
rect 292 29529 298 29585
rect 354 29529 396 29585
rect 452 29529 494 29585
rect 550 29529 592 29585
rect 648 29529 656 29585
rect 292 29504 656 29529
rect 292 29448 298 29504
rect 354 29448 396 29504
rect 452 29448 494 29504
rect 550 29448 592 29504
rect 648 29448 656 29504
rect 292 29423 656 29448
rect 292 29367 298 29423
rect 354 29367 396 29423
rect 452 29367 494 29423
rect 550 29367 592 29423
rect 648 29367 656 29423
rect 292 29342 656 29367
rect 292 29286 298 29342
rect 354 29286 396 29342
rect 452 29286 494 29342
rect 550 29286 592 29342
rect 648 29286 656 29342
rect 292 29261 656 29286
rect 292 29205 298 29261
rect 354 29205 396 29261
rect 452 29205 494 29261
rect 550 29205 592 29261
rect 648 29205 656 29261
rect 292 29180 656 29205
rect 292 29124 298 29180
rect 354 29124 396 29180
rect 452 29124 494 29180
rect 550 29124 592 29180
rect 648 29124 656 29180
rect 292 29099 656 29124
rect 292 29043 298 29099
rect 354 29043 396 29099
rect 452 29043 494 29099
rect 550 29043 592 29099
rect 648 29043 656 29099
rect 292 28015 656 29043
rect 292 27959 299 28015
rect 355 27959 393 28015
rect 449 27959 487 28015
rect 543 27959 581 28015
rect 637 27959 656 28015
rect 292 27933 656 27959
rect 292 27877 299 27933
rect 355 27877 393 27933
rect 449 27877 487 27933
rect 543 27877 581 27933
rect 637 27877 656 27933
rect 292 27851 656 27877
rect 292 27795 299 27851
rect 355 27795 393 27851
rect 449 27795 487 27851
rect 543 27795 581 27851
rect 637 27795 656 27851
rect 292 27769 656 27795
rect 292 27713 299 27769
rect 355 27713 393 27769
rect 449 27713 487 27769
rect 543 27713 581 27769
rect 637 27713 656 27769
rect 292 27687 656 27713
rect 292 27631 299 27687
rect 355 27631 393 27687
rect 449 27631 487 27687
rect 543 27631 581 27687
rect 637 27631 656 27687
rect 292 27605 656 27631
rect 292 27549 299 27605
rect 355 27549 393 27605
rect 449 27549 487 27605
rect 543 27549 581 27605
rect 637 27549 656 27605
rect 292 27523 656 27549
rect 292 27467 299 27523
rect 355 27467 393 27523
rect 449 27467 487 27523
rect 543 27467 581 27523
rect 637 27467 656 27523
rect 292 27441 656 27467
rect 292 27385 299 27441
rect 355 27385 393 27441
rect 449 27385 487 27441
rect 543 27385 581 27441
rect 637 27385 656 27441
rect 292 27359 656 27385
rect 292 27303 299 27359
rect 355 27303 393 27359
rect 449 27303 487 27359
rect 543 27303 581 27359
rect 637 27303 656 27359
rect 292 27277 656 27303
rect 292 27221 299 27277
rect 355 27221 393 27277
rect 449 27221 487 27277
rect 543 27221 581 27277
rect 637 27221 656 27277
rect 292 27195 656 27221
rect 292 27139 299 27195
rect 355 27139 393 27195
rect 449 27139 487 27195
rect 543 27139 581 27195
rect 637 27139 656 27195
rect 292 27112 656 27139
rect 292 27056 299 27112
rect 355 27056 393 27112
rect 449 27056 487 27112
rect 543 27056 581 27112
rect 637 27056 656 27112
rect 292 27029 656 27056
rect 292 26973 299 27029
rect 355 26973 393 27029
rect 449 26973 487 27029
rect 543 26973 581 27029
rect 637 26973 656 27029
rect 292 26946 656 26973
rect 292 26890 299 26946
rect 355 26890 393 26946
rect 449 26890 487 26946
rect 543 26890 581 26946
rect 637 26890 656 26946
rect 292 26863 656 26890
rect 292 26807 299 26863
rect 355 26807 393 26863
rect 449 26807 487 26863
rect 543 26807 581 26863
rect 637 26807 656 26863
rect 292 26780 656 26807
rect 292 26724 299 26780
rect 355 26724 393 26780
rect 449 26724 487 26780
rect 543 26724 581 26780
rect 637 26724 656 26780
rect 292 26697 656 26724
rect 292 26641 299 26697
rect 355 26641 393 26697
rect 449 26641 487 26697
rect 543 26641 581 26697
rect 637 26641 656 26697
rect 292 26614 656 26641
rect 292 26558 299 26614
rect 355 26558 393 26614
rect 449 26558 487 26614
rect 543 26558 581 26614
rect 637 26558 656 26614
rect 292 26531 656 26558
rect 292 26475 299 26531
rect 355 26475 393 26531
rect 449 26475 487 26531
rect 543 26475 581 26531
rect 637 26475 656 26531
rect 292 26448 656 26475
rect 292 26392 299 26448
rect 355 26392 393 26448
rect 449 26392 487 26448
rect 543 26392 581 26448
rect 637 26392 656 26448
rect 292 26365 656 26392
rect 1054 33517 2054 37178
rect 5106 38977 5110 39041
rect 5174 38977 5190 39041
rect 5254 38977 5270 39041
rect 5334 38977 5350 39041
rect 5414 38977 5430 39041
rect 5494 38977 5510 39041
rect 5574 38977 5590 39041
rect 5654 38977 5670 39041
rect 5734 38977 5750 39041
rect 5814 38977 5830 39041
rect 5894 38977 5910 39041
rect 5974 38977 5990 39041
rect 6054 38977 6070 39041
rect 6134 38977 6150 39041
rect 6214 38977 6230 39041
rect 6294 38977 6298 39041
rect 5106 38960 6298 38977
rect 5106 38896 5110 38960
rect 5174 38896 5190 38960
rect 5254 38896 5270 38960
rect 5334 38896 5350 38960
rect 5414 38896 5430 38960
rect 5494 38896 5510 38960
rect 5574 38896 5590 38960
rect 5654 38896 5670 38960
rect 5734 38896 5750 38960
rect 5814 38896 5830 38960
rect 5894 38896 5910 38960
rect 5974 38896 5990 38960
rect 6054 38896 6070 38960
rect 6134 38896 6150 38960
rect 6214 38896 6230 38960
rect 6294 38896 6298 38960
rect 5106 38879 6298 38896
rect 5106 38815 5110 38879
rect 5174 38815 5190 38879
rect 5254 38815 5270 38879
rect 5334 38815 5350 38879
rect 5414 38815 5430 38879
rect 5494 38815 5510 38879
rect 5574 38815 5590 38879
rect 5654 38815 5670 38879
rect 5734 38815 5750 38879
rect 5814 38815 5830 38879
rect 5894 38815 5910 38879
rect 5974 38815 5990 38879
rect 6054 38815 6070 38879
rect 6134 38815 6150 38879
rect 6214 38815 6230 38879
rect 6294 38815 6298 38879
rect 5106 38798 6298 38815
rect 5106 38734 5110 38798
rect 5174 38734 5190 38798
rect 5254 38734 5270 38798
rect 5334 38734 5350 38798
rect 5414 38734 5430 38798
rect 5494 38734 5510 38798
rect 5574 38734 5590 38798
rect 5654 38734 5670 38798
rect 5734 38734 5750 38798
rect 5814 38734 5830 38798
rect 5894 38734 5910 38798
rect 5974 38734 5990 38798
rect 6054 38734 6070 38798
rect 6134 38734 6150 38798
rect 6214 38734 6230 38798
rect 6294 38734 6298 38798
rect 5106 38717 6298 38734
rect 5106 38653 5110 38717
rect 5174 38653 5190 38717
rect 5254 38653 5270 38717
rect 5334 38653 5350 38717
rect 5414 38653 5430 38717
rect 5494 38653 5510 38717
rect 5574 38653 5590 38717
rect 5654 38653 5670 38717
rect 5734 38653 5750 38717
rect 5814 38653 5830 38717
rect 5894 38653 5910 38717
rect 5974 38653 5990 38717
rect 6054 38653 6070 38717
rect 6134 38653 6150 38717
rect 6214 38653 6230 38717
rect 6294 38653 6298 38717
rect 5106 38636 6298 38653
rect 5106 38572 5110 38636
rect 5174 38572 5190 38636
rect 5254 38572 5270 38636
rect 5334 38572 5350 38636
rect 5414 38572 5430 38636
rect 5494 38572 5510 38636
rect 5574 38572 5590 38636
rect 5654 38572 5670 38636
rect 5734 38572 5750 38636
rect 5814 38572 5830 38636
rect 5894 38572 5910 38636
rect 5974 38572 5990 38636
rect 6054 38572 6070 38636
rect 6134 38572 6150 38636
rect 6214 38572 6230 38636
rect 6294 38572 6298 38636
rect 5106 38555 6298 38572
rect 5106 38491 5110 38555
rect 5174 38491 5190 38555
rect 5254 38491 5270 38555
rect 5334 38491 5350 38555
rect 5414 38491 5430 38555
rect 5494 38491 5510 38555
rect 5574 38491 5590 38555
rect 5654 38491 5670 38555
rect 5734 38491 5750 38555
rect 5814 38491 5830 38555
rect 5894 38491 5910 38555
rect 5974 38491 5990 38555
rect 6054 38491 6070 38555
rect 6134 38491 6150 38555
rect 6214 38491 6230 38555
rect 6294 38491 6298 38555
rect 5106 38474 6298 38491
rect 5106 38410 5110 38474
rect 5174 38410 5190 38474
rect 5254 38410 5270 38474
rect 5334 38410 5350 38474
rect 5414 38410 5430 38474
rect 5494 38410 5510 38474
rect 5574 38410 5590 38474
rect 5654 38410 5670 38474
rect 5734 38410 5750 38474
rect 5814 38410 5830 38474
rect 5894 38410 5910 38474
rect 5974 38410 5990 38474
rect 6054 38410 6070 38474
rect 6134 38410 6150 38474
rect 6214 38410 6230 38474
rect 6294 38410 6298 38474
rect 5106 38393 6298 38410
rect 5106 38329 5110 38393
rect 5174 38329 5190 38393
rect 5254 38329 5270 38393
rect 5334 38329 5350 38393
rect 5414 38329 5430 38393
rect 5494 38329 5510 38393
rect 5574 38329 5590 38393
rect 5654 38329 5670 38393
rect 5734 38329 5750 38393
rect 5814 38329 5830 38393
rect 5894 38329 5910 38393
rect 5974 38329 5990 38393
rect 6054 38329 6070 38393
rect 6134 38329 6150 38393
rect 6214 38329 6230 38393
rect 6294 38329 6298 38393
rect 5106 38312 6298 38329
rect 5106 38248 5110 38312
rect 5174 38248 5190 38312
rect 5254 38248 5270 38312
rect 5334 38248 5350 38312
rect 5414 38248 5430 38312
rect 5494 38248 5510 38312
rect 5574 38248 5590 38312
rect 5654 38248 5670 38312
rect 5734 38248 5750 38312
rect 5814 38248 5830 38312
rect 5894 38248 5910 38312
rect 5974 38248 5990 38312
rect 6054 38248 6070 38312
rect 6134 38248 6150 38312
rect 6214 38248 6230 38312
rect 6294 38248 6298 38312
rect 5106 38231 6298 38248
rect 5106 38167 5110 38231
rect 5174 38167 5190 38231
rect 5254 38167 5270 38231
rect 5334 38167 5350 38231
rect 5414 38167 5430 38231
rect 5494 38167 5510 38231
rect 5574 38167 5590 38231
rect 5654 38167 5670 38231
rect 5734 38167 5750 38231
rect 5814 38167 5830 38231
rect 5894 38167 5910 38231
rect 5974 38167 5990 38231
rect 6054 38167 6070 38231
rect 6134 38167 6150 38231
rect 6214 38167 6230 38231
rect 6294 38167 6298 38231
rect 5106 38150 6298 38167
rect 5106 38086 5110 38150
rect 5174 38086 5190 38150
rect 5254 38086 5270 38150
rect 5334 38086 5350 38150
rect 5414 38086 5430 38150
rect 5494 38086 5510 38150
rect 5574 38086 5590 38150
rect 5654 38086 5670 38150
rect 5734 38086 5750 38150
rect 5814 38086 5830 38150
rect 5894 38086 5910 38150
rect 5974 38086 5990 38150
rect 6054 38086 6070 38150
rect 6134 38086 6150 38150
rect 6214 38086 6230 38150
rect 6294 38086 6298 38150
rect 5106 38069 6298 38086
rect 5106 38005 5110 38069
rect 5174 38005 5190 38069
rect 5254 38005 5270 38069
rect 5334 38005 5350 38069
rect 5414 38005 5430 38069
rect 5494 38005 5510 38069
rect 5574 38005 5590 38069
rect 5654 38005 5670 38069
rect 5734 38005 5750 38069
rect 5814 38005 5830 38069
rect 5894 38005 5910 38069
rect 5974 38005 5990 38069
rect 6054 38005 6070 38069
rect 6134 38005 6150 38069
rect 6214 38005 6230 38069
rect 6294 38005 6298 38069
rect 5106 37988 6298 38005
rect 5106 37924 5110 37988
rect 5174 37924 5190 37988
rect 5254 37924 5270 37988
rect 5334 37924 5350 37988
rect 5414 37924 5430 37988
rect 5494 37924 5510 37988
rect 5574 37924 5590 37988
rect 5654 37924 5670 37988
rect 5734 37924 5750 37988
rect 5814 37924 5830 37988
rect 5894 37924 5910 37988
rect 5974 37924 5990 37988
rect 6054 37924 6070 37988
rect 6134 37924 6150 37988
rect 6214 37924 6230 37988
rect 6294 37924 6298 37988
rect 5106 37907 6298 37924
rect 5106 37843 5110 37907
rect 5174 37843 5190 37907
rect 5254 37843 5270 37907
rect 5334 37843 5350 37907
rect 5414 37843 5430 37907
rect 5494 37843 5510 37907
rect 5574 37843 5590 37907
rect 5654 37843 5670 37907
rect 5734 37843 5750 37907
rect 5814 37843 5830 37907
rect 5894 37843 5910 37907
rect 5974 37843 5990 37907
rect 6054 37843 6070 37907
rect 6134 37843 6150 37907
rect 6214 37843 6230 37907
rect 6294 37843 6298 37907
rect 5106 37826 6298 37843
rect 5106 37762 5110 37826
rect 5174 37762 5190 37826
rect 5254 37762 5270 37826
rect 5334 37762 5350 37826
rect 5414 37762 5430 37826
rect 5494 37762 5510 37826
rect 5574 37762 5590 37826
rect 5654 37762 5670 37826
rect 5734 37762 5750 37826
rect 5814 37762 5830 37826
rect 5894 37762 5910 37826
rect 5974 37762 5990 37826
rect 6054 37762 6070 37826
rect 6134 37762 6150 37826
rect 6214 37762 6230 37826
rect 6294 37762 6298 37826
rect 5106 37745 6298 37762
rect 5106 37681 5110 37745
rect 5174 37681 5190 37745
rect 5254 37681 5270 37745
rect 5334 37681 5350 37745
rect 5414 37681 5430 37745
rect 5494 37681 5510 37745
rect 5574 37681 5590 37745
rect 5654 37681 5670 37745
rect 5734 37681 5750 37745
rect 5814 37681 5830 37745
rect 5894 37681 5910 37745
rect 5974 37681 5990 37745
rect 6054 37681 6070 37745
rect 6134 37681 6150 37745
rect 6214 37681 6230 37745
rect 6294 37681 6298 37745
rect 5106 37664 6298 37681
rect 5106 37600 5110 37664
rect 5174 37600 5190 37664
rect 5254 37600 5270 37664
rect 5334 37600 5350 37664
rect 5414 37600 5430 37664
rect 5494 37600 5510 37664
rect 5574 37600 5590 37664
rect 5654 37600 5670 37664
rect 5734 37600 5750 37664
rect 5814 37600 5830 37664
rect 5894 37600 5910 37664
rect 5974 37600 5990 37664
rect 6054 37600 6070 37664
rect 6134 37600 6150 37664
rect 6214 37600 6230 37664
rect 6294 37600 6298 37664
rect 5106 37583 6298 37600
rect 5106 37519 5110 37583
rect 5174 37519 5190 37583
rect 5254 37519 5270 37583
rect 5334 37519 5350 37583
rect 5414 37519 5430 37583
rect 5494 37519 5510 37583
rect 5574 37519 5590 37583
rect 5654 37519 5670 37583
rect 5734 37519 5750 37583
rect 5814 37519 5830 37583
rect 5894 37519 5910 37583
rect 5974 37519 5990 37583
rect 6054 37519 6070 37583
rect 6134 37519 6150 37583
rect 6214 37519 6230 37583
rect 6294 37519 6298 37583
rect 5106 37502 6298 37519
rect 5106 37438 5110 37502
rect 5174 37438 5190 37502
rect 5254 37438 5270 37502
rect 5334 37438 5350 37502
rect 5414 37438 5430 37502
rect 5494 37438 5510 37502
rect 5574 37438 5590 37502
rect 5654 37438 5670 37502
rect 5734 37438 5750 37502
rect 5814 37438 5830 37502
rect 5894 37438 5910 37502
rect 5974 37438 5990 37502
rect 6054 37438 6070 37502
rect 6134 37438 6150 37502
rect 6214 37438 6230 37502
rect 6294 37438 6298 37502
rect 5106 37421 6298 37438
rect 5106 37357 5110 37421
rect 5174 37357 5190 37421
rect 5254 37357 5270 37421
rect 5334 37357 5350 37421
rect 5414 37357 5430 37421
rect 5494 37357 5510 37421
rect 5574 37357 5590 37421
rect 5654 37357 5670 37421
rect 5734 37357 5750 37421
rect 5814 37357 5830 37421
rect 5894 37357 5910 37421
rect 5974 37357 5990 37421
rect 6054 37357 6070 37421
rect 6134 37357 6150 37421
rect 6214 37357 6230 37421
rect 6294 37357 6298 37421
rect 5106 37340 6298 37357
rect 5106 37276 5110 37340
rect 5174 37276 5190 37340
rect 5254 37276 5270 37340
rect 5334 37276 5350 37340
rect 5414 37276 5430 37340
rect 5494 37276 5510 37340
rect 5574 37276 5590 37340
rect 5654 37276 5670 37340
rect 5734 37276 5750 37340
rect 5814 37276 5830 37340
rect 5894 37276 5910 37340
rect 5974 37276 5990 37340
rect 6054 37276 6070 37340
rect 6134 37276 6150 37340
rect 6214 37276 6230 37340
rect 6294 37276 6298 37340
rect 5106 37259 6298 37276
rect 5106 37195 5110 37259
rect 5174 37195 5190 37259
rect 5254 37195 5270 37259
rect 5334 37195 5350 37259
rect 5414 37195 5430 37259
rect 5494 37195 5510 37259
rect 5574 37195 5590 37259
rect 5654 37195 5670 37259
rect 5734 37195 5750 37259
rect 5814 37195 5830 37259
rect 5894 37195 5910 37259
rect 5974 37195 5990 37259
rect 6054 37195 6070 37259
rect 6134 37195 6150 37259
rect 6214 37195 6230 37259
rect 6294 37195 6298 37259
rect 5106 37178 6298 37195
rect 5106 37114 5110 37178
rect 5174 37114 5190 37178
rect 5254 37114 5270 37178
rect 5334 37114 5350 37178
rect 5414 37114 5430 37178
rect 5494 37114 5510 37178
rect 5574 37114 5590 37178
rect 5654 37114 5670 37178
rect 5734 37114 5750 37178
rect 5814 37114 5830 37178
rect 5894 37114 5910 37178
rect 5974 37114 5990 37178
rect 6054 37114 6070 37178
rect 6134 37114 6150 37178
rect 6214 37114 6230 37178
rect 6294 37114 6298 37178
rect 5106 37097 6298 37114
rect 5106 37033 5110 37097
rect 5174 37033 5190 37097
rect 5254 37033 5270 37097
rect 5334 37033 5350 37097
rect 5414 37033 5430 37097
rect 5494 37033 5510 37097
rect 5574 37033 5590 37097
rect 5654 37033 5670 37097
rect 5734 37033 5750 37097
rect 5814 37033 5830 37097
rect 5894 37033 5910 37097
rect 5974 37033 5990 37097
rect 6054 37033 6070 37097
rect 6134 37033 6150 37097
rect 6214 37033 6230 37097
rect 6294 37033 6298 37097
rect 5106 37016 6298 37033
rect 5106 36952 5110 37016
rect 5174 36952 5190 37016
rect 5254 36952 5270 37016
rect 5334 36952 5350 37016
rect 5414 36952 5430 37016
rect 5494 36952 5510 37016
rect 5574 36952 5590 37016
rect 5654 36952 5670 37016
rect 5734 36952 5750 37016
rect 5814 36952 5830 37016
rect 5894 36952 5910 37016
rect 5974 36952 5990 37016
rect 6054 36952 6070 37016
rect 6134 36952 6150 37016
rect 6214 36952 6230 37016
rect 6294 36952 6298 37016
rect 5106 36935 6298 36952
rect 5106 36871 5110 36935
rect 5174 36871 5190 36935
rect 5254 36871 5270 36935
rect 5334 36871 5350 36935
rect 5414 36871 5430 36935
rect 5494 36871 5510 36935
rect 5574 36871 5590 36935
rect 5654 36871 5670 36935
rect 5734 36871 5750 36935
rect 5814 36871 5830 36935
rect 5894 36871 5910 36935
rect 5974 36871 5990 36935
rect 6054 36871 6070 36935
rect 6134 36871 6150 36935
rect 6214 36871 6230 36935
rect 6294 36871 6298 36935
rect 5106 36854 6298 36871
rect 5106 36790 5110 36854
rect 5174 36790 5190 36854
rect 5254 36790 5270 36854
rect 5334 36790 5350 36854
rect 5414 36790 5430 36854
rect 5494 36790 5510 36854
rect 5574 36790 5590 36854
rect 5654 36790 5670 36854
rect 5734 36790 5750 36854
rect 5814 36790 5830 36854
rect 5894 36790 5910 36854
rect 5974 36790 5990 36854
rect 6054 36790 6070 36854
rect 6134 36790 6150 36854
rect 6214 36790 6230 36854
rect 6294 36790 6298 36854
rect 5106 36773 6298 36790
rect 5106 36709 5110 36773
rect 5174 36709 5190 36773
rect 5254 36709 5270 36773
rect 5334 36709 5350 36773
rect 5414 36709 5430 36773
rect 5494 36709 5510 36773
rect 5574 36709 5590 36773
rect 5654 36709 5670 36773
rect 5734 36709 5750 36773
rect 5814 36709 5830 36773
rect 5894 36709 5910 36773
rect 5974 36709 5990 36773
rect 6054 36709 6070 36773
rect 6134 36709 6150 36773
rect 6214 36709 6230 36773
rect 6294 36709 6298 36773
rect 5106 36692 6298 36709
rect 5106 36628 5110 36692
rect 5174 36628 5190 36692
rect 5254 36628 5270 36692
rect 5334 36628 5350 36692
rect 5414 36628 5430 36692
rect 5494 36628 5510 36692
rect 5574 36628 5590 36692
rect 5654 36628 5670 36692
rect 5734 36628 5750 36692
rect 5814 36628 5830 36692
rect 5894 36628 5910 36692
rect 5974 36628 5990 36692
rect 6054 36628 6070 36692
rect 6134 36628 6150 36692
rect 6214 36628 6230 36692
rect 6294 36628 6298 36692
rect 5106 36611 6298 36628
rect 5106 36547 5110 36611
rect 5174 36547 5190 36611
rect 5254 36547 5270 36611
rect 5334 36547 5350 36611
rect 5414 36547 5430 36611
rect 5494 36547 5510 36611
rect 5574 36547 5590 36611
rect 5654 36547 5670 36611
rect 5734 36547 5750 36611
rect 5814 36547 5830 36611
rect 5894 36547 5910 36611
rect 5974 36547 5990 36611
rect 6054 36547 6070 36611
rect 6134 36547 6150 36611
rect 6214 36547 6230 36611
rect 6294 36547 6298 36611
rect 5106 36530 6298 36547
rect 5106 36466 5110 36530
rect 5174 36466 5190 36530
rect 5254 36466 5270 36530
rect 5334 36466 5350 36530
rect 5414 36466 5430 36530
rect 5494 36466 5510 36530
rect 5574 36466 5590 36530
rect 5654 36466 5670 36530
rect 5734 36466 5750 36530
rect 5814 36466 5830 36530
rect 5894 36466 5910 36530
rect 5974 36466 5990 36530
rect 6054 36466 6070 36530
rect 6134 36466 6150 36530
rect 6214 36466 6230 36530
rect 6294 36466 6298 36530
rect 5106 36449 6298 36466
rect 4077 36366 4723 36386
rect 4077 36310 4089 36366
rect 4145 36310 4231 36366
rect 4287 36310 4372 36366
rect 4428 36310 4513 36366
rect 4569 36310 4654 36366
rect 4710 36310 4723 36366
rect 4077 36266 4723 36310
rect 4077 36210 4089 36266
rect 4145 36210 4231 36266
rect 4287 36210 4372 36266
rect 4428 36210 4513 36266
rect 4569 36210 4654 36266
rect 4710 36210 4723 36266
rect 1054 28506 2024 33517
tri 2024 33487 2054 33517 nw
rect 2781 36081 3778 36133
rect 2781 36025 2792 36081
rect 2848 36025 2924 36081
rect 2980 36025 3056 36081
rect 3112 36025 3187 36081
rect 3243 36025 3318 36081
rect 3374 36025 3449 36081
rect 3505 36025 3580 36081
rect 3636 36025 3711 36081
rect 3767 36025 3778 36081
rect 2781 35963 3778 36025
rect 2781 35907 2792 35963
rect 2848 35907 2924 35963
rect 2980 35907 3056 35963
rect 3112 35907 3187 35963
rect 3243 35907 3318 35963
rect 3374 35907 3449 35963
rect 3505 35907 3580 35963
rect 3636 35907 3711 35963
rect 3767 35907 3778 35963
rect 2781 35845 3778 35907
rect 2781 35789 2792 35845
rect 2848 35789 2924 35845
rect 2980 35789 3056 35845
rect 3112 35789 3187 35845
rect 3243 35789 3318 35845
rect 3374 35789 3449 35845
rect 3505 35789 3580 35845
rect 3636 35789 3711 35845
rect 3767 35789 3778 35845
rect 2132 31167 2496 31173
rect 2196 31103 2232 31167
rect 2296 31103 2332 31167
rect 2396 31103 2432 31167
rect 2132 31085 2496 31103
rect 2196 31021 2232 31085
rect 2296 31021 2332 31085
rect 2396 31021 2432 31085
rect 2132 31003 2496 31021
rect 2196 30939 2232 31003
rect 2296 30939 2332 31003
rect 2396 30939 2432 31003
rect 2132 30921 2496 30939
rect 2196 30857 2232 30921
rect 2296 30857 2332 30921
rect 2396 30857 2432 30921
rect 2132 30839 2496 30857
rect 2196 30775 2232 30839
rect 2296 30775 2332 30839
rect 2396 30775 2432 30839
rect 2132 30757 2496 30775
rect 2196 30693 2232 30757
rect 2296 30693 2332 30757
rect 2396 30693 2432 30757
rect 2132 30675 2496 30693
rect 2196 30611 2232 30675
rect 2296 30611 2332 30675
rect 2396 30611 2432 30675
rect 2132 30593 2496 30611
rect 2196 30529 2232 30593
rect 2296 30529 2332 30593
rect 2396 30529 2432 30593
rect 2132 30511 2496 30529
rect 2196 30447 2232 30511
rect 2296 30447 2332 30511
rect 2396 30447 2432 30511
rect 2132 30429 2496 30447
rect 2196 30365 2232 30429
rect 2296 30365 2332 30429
rect 2396 30365 2432 30429
rect 2132 30347 2496 30365
rect 2196 30283 2232 30347
rect 2296 30283 2332 30347
rect 2396 30283 2432 30347
rect 2132 30282 2139 30283
rect 2195 30282 2237 30283
rect 2293 30282 2335 30283
rect 2391 30282 2433 30283
rect 2489 30282 2496 30283
rect 2132 30264 2496 30282
rect 2196 30200 2232 30264
rect 2296 30200 2332 30264
rect 2396 30200 2432 30264
rect 2132 30199 2139 30200
rect 2195 30199 2237 30200
rect 2293 30199 2335 30200
rect 2391 30199 2433 30200
rect 2489 30199 2496 30200
rect 2132 30181 2496 30199
rect 2196 30117 2232 30181
rect 2296 30117 2332 30181
rect 2396 30117 2432 30181
rect 2132 30116 2139 30117
rect 2195 30116 2237 30117
rect 2293 30116 2335 30117
rect 2391 30116 2433 30117
rect 2489 30116 2496 30117
rect 2132 30098 2496 30116
rect 2196 30034 2232 30098
rect 2296 30034 2332 30098
rect 2396 30034 2432 30098
rect 2132 30033 2139 30034
rect 2195 30033 2237 30034
rect 2293 30033 2335 30034
rect 2391 30033 2433 30034
rect 2489 30033 2496 30034
rect 2132 30015 2496 30033
rect 2196 29951 2232 30015
rect 2296 29951 2332 30015
rect 2396 29951 2432 30015
rect 2132 29950 2139 29951
rect 2195 29950 2237 29951
rect 2293 29950 2335 29951
rect 2391 29950 2433 29951
rect 2489 29950 2496 29951
rect 2132 29932 2496 29950
rect 2196 29868 2232 29932
rect 2296 29868 2332 29932
rect 2396 29868 2432 29932
rect 2132 29867 2139 29868
rect 2195 29867 2237 29868
rect 2293 29867 2335 29868
rect 2391 29867 2433 29868
rect 2489 29867 2496 29868
rect 2132 29849 2496 29867
rect 2196 29785 2232 29849
rect 2296 29785 2332 29849
rect 2396 29785 2432 29849
rect 2132 29784 2139 29785
rect 2195 29784 2237 29785
rect 2293 29784 2335 29785
rect 2391 29784 2433 29785
rect 2489 29784 2496 29785
rect 2132 29766 2496 29784
rect 2196 29702 2232 29766
rect 2296 29702 2332 29766
rect 2396 29702 2432 29766
rect 2132 29701 2139 29702
rect 2195 29701 2237 29702
rect 2293 29701 2335 29702
rect 2391 29701 2433 29702
rect 2489 29701 2496 29702
rect 2132 29683 2496 29701
rect 2196 29619 2232 29683
rect 2296 29619 2332 29683
rect 2396 29619 2432 29683
rect 2132 29618 2139 29619
rect 2195 29618 2237 29619
rect 2293 29618 2335 29619
rect 2391 29618 2433 29619
rect 2489 29618 2496 29619
rect 2132 29600 2496 29618
rect 2196 29536 2232 29600
rect 2296 29536 2332 29600
rect 2396 29536 2432 29600
rect 2132 29535 2139 29536
rect 2195 29535 2237 29536
rect 2293 29535 2335 29536
rect 2391 29535 2433 29536
rect 2489 29535 2496 29536
rect 2132 29517 2496 29535
rect 2196 29453 2232 29517
rect 2296 29453 2332 29517
rect 2396 29453 2432 29517
rect 2132 29452 2139 29453
rect 2195 29452 2237 29453
rect 2293 29452 2335 29453
rect 2391 29452 2433 29453
rect 2489 29452 2496 29453
rect 2132 29434 2496 29452
rect 2196 29370 2232 29434
rect 2296 29370 2332 29434
rect 2396 29370 2432 29434
rect 2132 29369 2139 29370
rect 2195 29369 2237 29370
rect 2293 29369 2335 29370
rect 2391 29369 2433 29370
rect 2489 29369 2496 29370
rect 2132 29351 2496 29369
rect 2196 29287 2232 29351
rect 2296 29287 2332 29351
rect 2396 29287 2432 29351
rect 2132 29286 2139 29287
rect 2195 29286 2237 29287
rect 2293 29286 2335 29287
rect 2391 29286 2433 29287
rect 2489 29286 2496 29287
rect 2132 29268 2496 29286
rect 2196 29204 2232 29268
rect 2296 29204 2332 29268
rect 2396 29204 2432 29268
rect 2132 29203 2139 29204
rect 2195 29203 2237 29204
rect 2293 29203 2335 29204
rect 2391 29203 2433 29204
rect 2489 29203 2496 29204
rect 2132 29185 2496 29203
rect 2196 29121 2232 29185
rect 2296 29121 2332 29185
rect 2396 29121 2432 29185
rect 2132 29120 2139 29121
rect 2195 29120 2237 29121
rect 2293 29120 2335 29121
rect 2391 29120 2433 29121
rect 2489 29120 2496 29121
rect 2132 29102 2496 29120
rect 2196 29038 2232 29102
rect 2296 29038 2332 29102
rect 2396 29038 2432 29102
rect 2132 29037 2139 29038
rect 2195 29037 2237 29038
rect 2293 29037 2335 29038
rect 2391 29037 2433 29038
rect 2489 29037 2496 29038
rect 2132 29019 2496 29037
rect 2196 28955 2232 29019
rect 2296 28955 2332 29019
rect 2396 28955 2432 29019
rect 2132 28954 2139 28955
rect 2195 28954 2237 28955
rect 2293 28954 2335 28955
rect 2391 28954 2433 28955
rect 2489 28954 2496 28955
rect 2132 28936 2496 28954
rect 2196 28872 2232 28936
rect 2296 28872 2332 28936
rect 2396 28872 2432 28936
rect 2132 28871 2139 28872
rect 2195 28871 2237 28872
rect 2293 28871 2335 28872
rect 2391 28871 2433 28872
rect 2489 28871 2496 28872
rect 2132 28866 2496 28871
rect 2781 28562 3778 35789
rect 4077 34681 4723 36210
rect 4077 34617 4083 34681
rect 4147 34617 4165 34681
rect 4229 34617 4247 34681
rect 4311 34617 4329 34681
rect 4393 34617 4410 34681
rect 4474 34617 4491 34681
rect 4555 34617 4572 34681
rect 4636 34617 4653 34681
rect 4717 34617 4723 34681
rect 4077 34593 4723 34617
rect 4077 34529 4083 34593
rect 4147 34529 4165 34593
rect 4229 34529 4247 34593
rect 4311 34529 4329 34593
rect 4393 34529 4410 34593
rect 4474 34529 4491 34593
rect 4555 34529 4572 34593
rect 4636 34529 4653 34593
rect 4717 34529 4723 34593
rect 4077 34505 4723 34529
rect 4077 34441 4083 34505
rect 4147 34441 4165 34505
rect 4229 34441 4247 34505
rect 4311 34441 4329 34505
rect 4393 34441 4410 34505
rect 4474 34441 4491 34505
rect 4555 34441 4572 34505
rect 4636 34441 4653 34505
rect 4717 34441 4723 34505
rect 4077 34417 4723 34441
rect 4077 34353 4083 34417
rect 4147 34353 4165 34417
rect 4229 34353 4247 34417
rect 4311 34353 4329 34417
rect 4393 34353 4410 34417
rect 4474 34353 4491 34417
rect 4555 34353 4572 34417
rect 4636 34353 4653 34417
rect 4717 34353 4723 34417
rect 4077 34329 4723 34353
rect 4077 34265 4083 34329
rect 4147 34265 4165 34329
rect 4229 34265 4247 34329
rect 4311 34265 4329 34329
rect 4393 34265 4410 34329
rect 4474 34265 4491 34329
rect 4555 34265 4572 34329
rect 4636 34265 4653 34329
rect 4717 34265 4723 34329
rect 4077 34241 4723 34265
rect 4077 34177 4083 34241
rect 4147 34177 4165 34241
rect 4229 34177 4247 34241
rect 4311 34177 4329 34241
rect 4393 34177 4410 34241
rect 4474 34177 4491 34241
rect 4555 34177 4572 34241
rect 4636 34177 4653 34241
rect 4717 34177 4723 34241
rect 4077 34172 4723 34177
rect 5106 36385 5110 36449
rect 5174 36385 5190 36449
rect 5254 36385 5270 36449
rect 5334 36385 5350 36449
rect 5414 36385 5430 36449
rect 5494 36385 5510 36449
rect 5574 36385 5590 36449
rect 5654 36385 5670 36449
rect 5734 36385 5750 36449
rect 5814 36385 5830 36449
rect 5894 36385 5910 36449
rect 5974 36385 5990 36449
rect 6054 36385 6070 36449
rect 6134 36385 6150 36449
rect 6214 36385 6230 36449
rect 6294 36385 6298 36449
rect 5106 36368 6298 36385
rect 5106 36304 5110 36368
rect 5174 36304 5190 36368
rect 5254 36304 5270 36368
rect 5334 36304 5350 36368
rect 5414 36304 5430 36368
rect 5494 36304 5510 36368
rect 5574 36304 5590 36368
rect 5654 36304 5670 36368
rect 5734 36304 5750 36368
rect 5814 36304 5830 36368
rect 5894 36304 5910 36368
rect 5974 36304 5990 36368
rect 6054 36304 6070 36368
rect 6134 36304 6150 36368
rect 6214 36304 6230 36368
rect 6294 36304 6298 36368
rect 5106 36287 6298 36304
rect 5106 36223 5110 36287
rect 5174 36223 5190 36287
rect 5254 36223 5270 36287
rect 5334 36223 5350 36287
rect 5414 36223 5430 36287
rect 5494 36223 5510 36287
rect 5574 36223 5590 36287
rect 5654 36223 5670 36287
rect 5734 36223 5750 36287
rect 5814 36223 5830 36287
rect 5894 36223 5910 36287
rect 5974 36223 5990 36287
rect 6054 36223 6070 36287
rect 6134 36223 6150 36287
rect 6214 36223 6230 36287
rect 6294 36223 6298 36287
rect 5106 36206 6298 36223
rect 5106 36142 5110 36206
rect 5174 36142 5190 36206
rect 5254 36142 5270 36206
rect 5334 36142 5350 36206
rect 5414 36142 5430 36206
rect 5494 36142 5510 36206
rect 5574 36142 5590 36206
rect 5654 36142 5670 36206
rect 5734 36142 5750 36206
rect 5814 36142 5830 36206
rect 5894 36142 5910 36206
rect 5974 36142 5990 36206
rect 6054 36142 6070 36206
rect 6134 36142 6150 36206
rect 6214 36142 6230 36206
rect 6294 36142 6298 36206
rect 5106 36124 6298 36142
rect 5106 36060 5110 36124
rect 5174 36060 5190 36124
rect 5254 36060 5270 36124
rect 5334 36060 5350 36124
rect 5414 36060 5430 36124
rect 5494 36060 5510 36124
rect 5574 36060 5590 36124
rect 5654 36060 5670 36124
rect 5734 36060 5750 36124
rect 5814 36060 5830 36124
rect 5894 36060 5910 36124
rect 5974 36060 5990 36124
rect 6054 36060 6070 36124
rect 6134 36060 6150 36124
rect 6214 36060 6230 36124
rect 6294 36060 6298 36124
rect 5106 36042 6298 36060
rect 5106 35978 5110 36042
rect 5174 35978 5190 36042
rect 5254 35978 5270 36042
rect 5334 35978 5350 36042
rect 5414 35978 5430 36042
rect 5494 35978 5510 36042
rect 5574 35978 5590 36042
rect 5654 35978 5670 36042
rect 5734 35978 5750 36042
rect 5814 35978 5830 36042
rect 5894 35978 5910 36042
rect 5974 35978 5990 36042
rect 6054 35978 6070 36042
rect 6134 35978 6150 36042
rect 6214 35978 6230 36042
rect 6294 35978 6298 36042
rect 5106 35960 6298 35978
rect 5106 35896 5110 35960
rect 5174 35896 5190 35960
rect 5254 35896 5270 35960
rect 5334 35896 5350 35960
rect 5414 35896 5430 35960
rect 5494 35896 5510 35960
rect 5574 35896 5590 35960
rect 5654 35896 5670 35960
rect 5734 35896 5750 35960
rect 5814 35896 5830 35960
rect 5894 35896 5910 35960
rect 5974 35896 5990 35960
rect 6054 35896 6070 35960
rect 6134 35896 6150 35960
rect 6214 35896 6230 35960
rect 6294 35896 6298 35960
rect 5106 35878 6298 35896
rect 5106 35814 5110 35878
rect 5174 35814 5190 35878
rect 5254 35814 5270 35878
rect 5334 35814 5350 35878
rect 5414 35814 5430 35878
rect 5494 35814 5510 35878
rect 5574 35814 5590 35878
rect 5654 35814 5670 35878
rect 5734 35814 5750 35878
rect 5814 35814 5830 35878
rect 5894 35814 5910 35878
rect 5974 35814 5990 35878
rect 6054 35814 6070 35878
rect 6134 35814 6150 35878
rect 6214 35814 6230 35878
rect 6294 35814 6298 35878
rect 5106 35796 6298 35814
rect 5106 35732 5110 35796
rect 5174 35732 5190 35796
rect 5254 35732 5270 35796
rect 5334 35732 5350 35796
rect 5414 35732 5430 35796
rect 5494 35732 5510 35796
rect 5574 35732 5590 35796
rect 5654 35732 5670 35796
rect 5734 35732 5750 35796
rect 5814 35732 5830 35796
rect 5894 35732 5910 35796
rect 5974 35732 5990 35796
rect 6054 35732 6070 35796
rect 6134 35732 6150 35796
rect 6214 35732 6230 35796
rect 6294 35732 6298 35796
rect 5106 35714 6298 35732
rect 5106 35650 5110 35714
rect 5174 35650 5190 35714
rect 5254 35650 5270 35714
rect 5334 35650 5350 35714
rect 5414 35650 5430 35714
rect 5494 35650 5510 35714
rect 5574 35650 5590 35714
rect 5654 35650 5670 35714
rect 5734 35650 5750 35714
rect 5814 35650 5830 35714
rect 5894 35650 5910 35714
rect 5974 35650 5990 35714
rect 6054 35650 6070 35714
rect 6134 35650 6150 35714
rect 6214 35650 6230 35714
rect 6294 35650 6298 35714
rect 5106 35632 6298 35650
rect 5106 35568 5110 35632
rect 5174 35568 5190 35632
rect 5254 35568 5270 35632
rect 5334 35568 5350 35632
rect 5414 35568 5430 35632
rect 5494 35568 5510 35632
rect 5574 35568 5590 35632
rect 5654 35568 5670 35632
rect 5734 35568 5750 35632
rect 5814 35568 5830 35632
rect 5894 35568 5910 35632
rect 5974 35568 5990 35632
rect 6054 35568 6070 35632
rect 6134 35568 6150 35632
rect 6214 35568 6230 35632
rect 6294 35568 6298 35632
rect 5106 35550 6298 35568
rect 5106 35486 5110 35550
rect 5174 35486 5190 35550
rect 5254 35486 5270 35550
rect 5334 35486 5350 35550
rect 5414 35486 5430 35550
rect 5494 35486 5510 35550
rect 5574 35486 5590 35550
rect 5654 35486 5670 35550
rect 5734 35486 5750 35550
rect 5814 35486 5830 35550
rect 5894 35486 5910 35550
rect 5974 35486 5990 35550
rect 6054 35486 6070 35550
rect 6134 35486 6150 35550
rect 6214 35486 6230 35550
rect 6294 35486 6298 35550
rect 5106 35468 6298 35486
rect 5106 35404 5110 35468
rect 5174 35404 5190 35468
rect 5254 35404 5270 35468
rect 5334 35404 5350 35468
rect 5414 35404 5430 35468
rect 5494 35404 5510 35468
rect 5574 35404 5590 35468
rect 5654 35404 5670 35468
rect 5734 35404 5750 35468
rect 5814 35404 5830 35468
rect 5894 35404 5910 35468
rect 5974 35404 5990 35468
rect 6054 35404 6070 35468
rect 6134 35404 6150 35468
rect 6214 35404 6230 35468
rect 6294 35404 6298 35468
rect 5106 35386 6298 35404
rect 5106 35322 5110 35386
rect 5174 35322 5190 35386
rect 5254 35322 5270 35386
rect 5334 35322 5350 35386
rect 5414 35322 5430 35386
rect 5494 35322 5510 35386
rect 5574 35322 5590 35386
rect 5654 35322 5670 35386
rect 5734 35322 5750 35386
rect 5814 35322 5830 35386
rect 5894 35322 5910 35386
rect 5974 35322 5990 35386
rect 6054 35322 6070 35386
rect 6134 35322 6150 35386
rect 6214 35322 6230 35386
rect 6294 35322 6298 35386
rect 5106 35304 6298 35322
rect 5106 35240 5110 35304
rect 5174 35240 5190 35304
rect 5254 35240 5270 35304
rect 5334 35240 5350 35304
rect 5414 35240 5430 35304
rect 5494 35240 5510 35304
rect 5574 35240 5590 35304
rect 5654 35240 5670 35304
rect 5734 35240 5750 35304
rect 5814 35240 5830 35304
rect 5894 35240 5910 35304
rect 5974 35240 5990 35304
rect 6054 35240 6070 35304
rect 6134 35240 6150 35304
rect 6214 35240 6230 35304
rect 6294 35240 6298 35304
rect 5106 35222 6298 35240
rect 5106 35158 5110 35222
rect 5174 35158 5190 35222
rect 5254 35158 5270 35222
rect 5334 35158 5350 35222
rect 5414 35158 5430 35222
rect 5494 35158 5510 35222
rect 5574 35158 5590 35222
rect 5654 35158 5670 35222
rect 5734 35158 5750 35222
rect 5814 35158 5830 35222
rect 5894 35158 5910 35222
rect 5974 35158 5990 35222
rect 6054 35158 6070 35222
rect 6134 35158 6150 35222
rect 6214 35158 6230 35222
rect 6294 35158 6298 35222
rect 5106 32613 6298 35158
rect 5106 32557 5112 32613
rect 5168 32557 5193 32613
rect 5249 32557 5273 32613
rect 5329 32557 5353 32613
rect 5409 32557 5433 32613
rect 5489 32557 5513 32613
rect 5569 32557 5593 32613
rect 5649 32557 5673 32613
rect 5729 32557 5753 32613
rect 5809 32557 5833 32613
rect 5889 32557 5913 32613
rect 5969 32557 5993 32613
rect 6049 32557 6073 32613
rect 6129 32557 6153 32613
rect 6209 32557 6233 32613
rect 6289 32557 6298 32613
rect 5106 32531 6298 32557
rect 5106 32475 5112 32531
rect 5168 32475 5193 32531
rect 5249 32475 5273 32531
rect 5329 32475 5353 32531
rect 5409 32475 5433 32531
rect 5489 32475 5513 32531
rect 5569 32475 5593 32531
rect 5649 32475 5673 32531
rect 5729 32475 5753 32531
rect 5809 32475 5833 32531
rect 5889 32475 5913 32531
rect 5969 32475 5993 32531
rect 6049 32475 6073 32531
rect 6129 32475 6153 32531
rect 6209 32475 6233 32531
rect 6289 32475 6298 32531
rect 5106 32449 6298 32475
rect 5106 32393 5112 32449
rect 5168 32393 5193 32449
rect 5249 32393 5273 32449
rect 5329 32393 5353 32449
rect 5409 32393 5433 32449
rect 5489 32393 5513 32449
rect 5569 32393 5593 32449
rect 5649 32393 5673 32449
rect 5729 32393 5753 32449
rect 5809 32393 5833 32449
rect 5889 32393 5913 32449
rect 5969 32393 5993 32449
rect 6049 32393 6073 32449
rect 6129 32393 6153 32449
rect 6209 32393 6233 32449
rect 6289 32393 6298 32449
rect 5106 32367 6298 32393
rect 5106 32311 5112 32367
rect 5168 32311 5193 32367
rect 5249 32311 5273 32367
rect 5329 32311 5353 32367
rect 5409 32311 5433 32367
rect 5489 32311 5513 32367
rect 5569 32311 5593 32367
rect 5649 32311 5673 32367
rect 5729 32311 5753 32367
rect 5809 32311 5833 32367
rect 5889 32311 5913 32367
rect 5969 32311 5993 32367
rect 6049 32311 6073 32367
rect 6129 32311 6153 32367
rect 6209 32311 6233 32367
rect 6289 32311 6298 32367
rect 5106 32285 6298 32311
rect 5106 32229 5112 32285
rect 5168 32229 5193 32285
rect 5249 32229 5273 32285
rect 5329 32229 5353 32285
rect 5409 32229 5433 32285
rect 5489 32229 5513 32285
rect 5569 32229 5593 32285
rect 5649 32229 5673 32285
rect 5729 32229 5753 32285
rect 5809 32229 5833 32285
rect 5889 32229 5913 32285
rect 5969 32229 5993 32285
rect 6049 32229 6073 32285
rect 6129 32229 6153 32285
rect 6209 32229 6233 32285
rect 6289 32229 6298 32285
rect 5106 32203 6298 32229
rect 5106 32147 5112 32203
rect 5168 32147 5193 32203
rect 5249 32147 5273 32203
rect 5329 32147 5353 32203
rect 5409 32147 5433 32203
rect 5489 32147 5513 32203
rect 5569 32147 5593 32203
rect 5649 32147 5673 32203
rect 5729 32147 5753 32203
rect 5809 32147 5833 32203
rect 5889 32147 5913 32203
rect 5969 32147 5993 32203
rect 6049 32147 6073 32203
rect 6129 32147 6153 32203
rect 6209 32147 6233 32203
rect 6289 32147 6298 32203
rect 5106 32121 6298 32147
rect 5106 32065 5112 32121
rect 5168 32065 5193 32121
rect 5249 32065 5273 32121
rect 5329 32065 5353 32121
rect 5409 32065 5433 32121
rect 5489 32065 5513 32121
rect 5569 32065 5593 32121
rect 5649 32065 5673 32121
rect 5729 32065 5753 32121
rect 5809 32065 5833 32121
rect 5889 32065 5913 32121
rect 5969 32065 5993 32121
rect 6049 32065 6073 32121
rect 6129 32065 6153 32121
rect 6209 32065 6233 32121
rect 6289 32065 6298 32121
rect 5106 32039 6298 32065
rect 5106 31983 5112 32039
rect 5168 31983 5193 32039
rect 5249 31983 5273 32039
rect 5329 31983 5353 32039
rect 5409 31983 5433 32039
rect 5489 31983 5513 32039
rect 5569 31983 5593 32039
rect 5649 31983 5673 32039
rect 5729 31983 5753 32039
rect 5809 31983 5833 32039
rect 5889 31983 5913 32039
rect 5969 31983 5993 32039
rect 6049 31983 6073 32039
rect 6129 31983 6153 32039
rect 6209 31983 6233 32039
rect 6289 31983 6298 32039
rect 5106 31957 6298 31983
rect 5106 31901 5112 31957
rect 5168 31901 5193 31957
rect 5249 31901 5273 31957
rect 5329 31901 5353 31957
rect 5409 31901 5433 31957
rect 5489 31901 5513 31957
rect 5569 31901 5593 31957
rect 5649 31901 5673 31957
rect 5729 31901 5753 31957
rect 5809 31901 5833 31957
rect 5889 31901 5913 31957
rect 5969 31901 5993 31957
rect 6049 31901 6073 31957
rect 6129 31901 6153 31957
rect 6209 31901 6233 31957
rect 6289 31901 6298 31957
rect 5106 31875 6298 31901
rect 5106 31819 5112 31875
rect 5168 31819 5193 31875
rect 5249 31819 5273 31875
rect 5329 31819 5353 31875
rect 5409 31819 5433 31875
rect 5489 31819 5513 31875
rect 5569 31819 5593 31875
rect 5649 31819 5673 31875
rect 5729 31819 5753 31875
rect 5809 31819 5833 31875
rect 5889 31819 5913 31875
rect 5969 31819 5993 31875
rect 6049 31819 6073 31875
rect 6129 31819 6153 31875
rect 6209 31819 6233 31875
rect 6289 31819 6298 31875
rect 5106 31793 6298 31819
rect 5106 31737 5112 31793
rect 5168 31737 5193 31793
rect 5249 31737 5273 31793
rect 5329 31737 5353 31793
rect 5409 31737 5433 31793
rect 5489 31737 5513 31793
rect 5569 31737 5593 31793
rect 5649 31737 5673 31793
rect 5729 31737 5753 31793
rect 5809 31737 5833 31793
rect 5889 31737 5913 31793
rect 5969 31737 5993 31793
rect 6049 31737 6073 31793
rect 6129 31737 6153 31793
rect 6209 31737 6233 31793
rect 6289 31737 6298 31793
rect 5106 31711 6298 31737
rect 5106 31655 5112 31711
rect 5168 31655 5193 31711
rect 5249 31655 5273 31711
rect 5329 31655 5353 31711
rect 5409 31655 5433 31711
rect 5489 31655 5513 31711
rect 5569 31655 5593 31711
rect 5649 31655 5673 31711
rect 5729 31655 5753 31711
rect 5809 31655 5833 31711
rect 5889 31655 5913 31711
rect 5969 31655 5993 31711
rect 6049 31655 6073 31711
rect 6129 31655 6153 31711
rect 6209 31655 6233 31711
rect 6289 31655 6298 31711
rect 5106 31629 6298 31655
rect 5106 31573 5112 31629
rect 5168 31573 5193 31629
rect 5249 31573 5273 31629
rect 5329 31573 5353 31629
rect 5409 31573 5433 31629
rect 5489 31573 5513 31629
rect 5569 31573 5593 31629
rect 5649 31573 5673 31629
rect 5729 31573 5753 31629
rect 5809 31573 5833 31629
rect 5889 31573 5913 31629
rect 5969 31573 5993 31629
rect 6049 31573 6073 31629
rect 6129 31573 6153 31629
rect 6209 31573 6233 31629
rect 6289 31573 6298 31629
rect 5106 31547 6298 31573
rect 5106 31491 5112 31547
rect 5168 31491 5193 31547
rect 5249 31491 5273 31547
rect 5329 31491 5353 31547
rect 5409 31491 5433 31547
rect 5489 31491 5513 31547
rect 5569 31491 5593 31547
rect 5649 31491 5673 31547
rect 5729 31491 5753 31547
rect 5809 31491 5833 31547
rect 5889 31491 5913 31547
rect 5969 31491 5993 31547
rect 6049 31491 6073 31547
rect 6129 31491 6153 31547
rect 6209 31491 6233 31547
rect 6289 31491 6298 31547
rect 5106 31478 6298 31491
rect 6599 39365 7795 39371
rect 6599 39301 6607 39365
rect 6671 39301 6687 39365
rect 6751 39301 6767 39365
rect 6831 39301 6847 39365
rect 6911 39301 6927 39365
rect 6991 39301 7007 39365
rect 7071 39301 7087 39365
rect 7151 39301 7167 39365
rect 7231 39301 7247 39365
rect 7311 39301 7327 39365
rect 7391 39301 7407 39365
rect 7471 39301 7487 39365
rect 7551 39301 7567 39365
rect 7631 39301 7647 39365
rect 7711 39301 7727 39365
rect 7791 39301 7795 39365
rect 6599 39284 7795 39301
rect 6599 39220 6607 39284
rect 6671 39220 6687 39284
rect 6751 39220 6767 39284
rect 6831 39220 6847 39284
rect 6911 39220 6927 39284
rect 6991 39220 7007 39284
rect 7071 39220 7087 39284
rect 7151 39220 7167 39284
rect 7231 39220 7247 39284
rect 7311 39220 7327 39284
rect 7391 39220 7407 39284
rect 7471 39220 7487 39284
rect 7551 39220 7567 39284
rect 7631 39220 7647 39284
rect 7711 39220 7727 39284
rect 7791 39220 7795 39284
rect 6599 39203 7795 39220
rect 6599 39139 6607 39203
rect 6671 39139 6687 39203
rect 6751 39139 6767 39203
rect 6831 39139 6847 39203
rect 6911 39139 6927 39203
rect 6991 39139 7007 39203
rect 7071 39139 7087 39203
rect 7151 39139 7167 39203
rect 7231 39139 7247 39203
rect 7311 39139 7327 39203
rect 7391 39139 7407 39203
rect 7471 39139 7487 39203
rect 7551 39139 7567 39203
rect 7631 39139 7647 39203
rect 7711 39139 7727 39203
rect 7791 39139 7795 39203
rect 6599 39122 7795 39139
rect 6599 39058 6607 39122
rect 6671 39058 6687 39122
rect 6751 39058 6767 39122
rect 6831 39058 6847 39122
rect 6911 39058 6927 39122
rect 6991 39058 7007 39122
rect 7071 39058 7087 39122
rect 7151 39058 7167 39122
rect 7231 39058 7247 39122
rect 7311 39058 7327 39122
rect 7391 39058 7407 39122
rect 7471 39058 7487 39122
rect 7551 39058 7567 39122
rect 7631 39058 7647 39122
rect 7711 39058 7727 39122
rect 7791 39058 7795 39122
rect 6599 39041 7795 39058
rect 6599 38977 6607 39041
rect 6671 38977 6687 39041
rect 6751 38977 6767 39041
rect 6831 38977 6847 39041
rect 6911 38977 6927 39041
rect 6991 38977 7007 39041
rect 7071 38977 7087 39041
rect 7151 38977 7167 39041
rect 7231 38977 7247 39041
rect 7311 38977 7327 39041
rect 7391 38977 7407 39041
rect 7471 38977 7487 39041
rect 7551 38977 7567 39041
rect 7631 38977 7647 39041
rect 7711 38977 7727 39041
rect 7791 38977 7795 39041
rect 6599 38960 7795 38977
rect 6599 38896 6607 38960
rect 6671 38896 6687 38960
rect 6751 38896 6767 38960
rect 6831 38896 6847 38960
rect 6911 38896 6927 38960
rect 6991 38896 7007 38960
rect 7071 38896 7087 38960
rect 7151 38896 7167 38960
rect 7231 38896 7247 38960
rect 7311 38896 7327 38960
rect 7391 38896 7407 38960
rect 7471 38896 7487 38960
rect 7551 38896 7567 38960
rect 7631 38896 7647 38960
rect 7711 38896 7727 38960
rect 7791 38896 7795 38960
rect 6599 38879 7795 38896
rect 6599 38815 6607 38879
rect 6671 38815 6687 38879
rect 6751 38815 6767 38879
rect 6831 38815 6847 38879
rect 6911 38815 6927 38879
rect 6991 38815 7007 38879
rect 7071 38815 7087 38879
rect 7151 38815 7167 38879
rect 7231 38815 7247 38879
rect 7311 38815 7327 38879
rect 7391 38815 7407 38879
rect 7471 38815 7487 38879
rect 7551 38815 7567 38879
rect 7631 38815 7647 38879
rect 7711 38815 7727 38879
rect 7791 38815 7795 38879
rect 6599 38798 7795 38815
rect 6599 38734 6607 38798
rect 6671 38734 6687 38798
rect 6751 38734 6767 38798
rect 6831 38734 6847 38798
rect 6911 38734 6927 38798
rect 6991 38734 7007 38798
rect 7071 38734 7087 38798
rect 7151 38734 7167 38798
rect 7231 38734 7247 38798
rect 7311 38734 7327 38798
rect 7391 38734 7407 38798
rect 7471 38734 7487 38798
rect 7551 38734 7567 38798
rect 7631 38734 7647 38798
rect 7711 38734 7727 38798
rect 7791 38734 7795 38798
rect 6599 38717 7795 38734
rect 6599 38653 6607 38717
rect 6671 38653 6687 38717
rect 6751 38653 6767 38717
rect 6831 38653 6847 38717
rect 6911 38653 6927 38717
rect 6991 38653 7007 38717
rect 7071 38653 7087 38717
rect 7151 38653 7167 38717
rect 7231 38653 7247 38717
rect 7311 38653 7327 38717
rect 7391 38653 7407 38717
rect 7471 38653 7487 38717
rect 7551 38653 7567 38717
rect 7631 38653 7647 38717
rect 7711 38653 7727 38717
rect 7791 38653 7795 38717
rect 6599 38636 7795 38653
rect 6599 38572 6607 38636
rect 6671 38572 6687 38636
rect 6751 38572 6767 38636
rect 6831 38572 6847 38636
rect 6911 38572 6927 38636
rect 6991 38572 7007 38636
rect 7071 38572 7087 38636
rect 7151 38572 7167 38636
rect 7231 38572 7247 38636
rect 7311 38572 7327 38636
rect 7391 38572 7407 38636
rect 7471 38572 7487 38636
rect 7551 38572 7567 38636
rect 7631 38572 7647 38636
rect 7711 38572 7727 38636
rect 7791 38572 7795 38636
rect 6599 38555 7795 38572
rect 6599 38491 6607 38555
rect 6671 38491 6687 38555
rect 6751 38491 6767 38555
rect 6831 38491 6847 38555
rect 6911 38491 6927 38555
rect 6991 38491 7007 38555
rect 7071 38491 7087 38555
rect 7151 38491 7167 38555
rect 7231 38491 7247 38555
rect 7311 38491 7327 38555
rect 7391 38491 7407 38555
rect 7471 38491 7487 38555
rect 7551 38491 7567 38555
rect 7631 38491 7647 38555
rect 7711 38491 7727 38555
rect 7791 38491 7795 38555
rect 6599 38474 7795 38491
rect 6599 38410 6607 38474
rect 6671 38410 6687 38474
rect 6751 38410 6767 38474
rect 6831 38410 6847 38474
rect 6911 38410 6927 38474
rect 6991 38410 7007 38474
rect 7071 38410 7087 38474
rect 7151 38410 7167 38474
rect 7231 38410 7247 38474
rect 7311 38410 7327 38474
rect 7391 38410 7407 38474
rect 7471 38410 7487 38474
rect 7551 38410 7567 38474
rect 7631 38410 7647 38474
rect 7711 38410 7727 38474
rect 7791 38410 7795 38474
rect 6599 38393 7795 38410
rect 6599 38329 6607 38393
rect 6671 38329 6687 38393
rect 6751 38329 6767 38393
rect 6831 38329 6847 38393
rect 6911 38329 6927 38393
rect 6991 38329 7007 38393
rect 7071 38329 7087 38393
rect 7151 38329 7167 38393
rect 7231 38329 7247 38393
rect 7311 38329 7327 38393
rect 7391 38329 7407 38393
rect 7471 38329 7487 38393
rect 7551 38329 7567 38393
rect 7631 38329 7647 38393
rect 7711 38329 7727 38393
rect 7791 38329 7795 38393
rect 6599 38312 7795 38329
rect 6599 38248 6607 38312
rect 6671 38248 6687 38312
rect 6751 38248 6767 38312
rect 6831 38248 6847 38312
rect 6911 38248 6927 38312
rect 6991 38248 7007 38312
rect 7071 38248 7087 38312
rect 7151 38248 7167 38312
rect 7231 38248 7247 38312
rect 7311 38248 7327 38312
rect 7391 38248 7407 38312
rect 7471 38248 7487 38312
rect 7551 38248 7567 38312
rect 7631 38248 7647 38312
rect 7711 38248 7727 38312
rect 7791 38248 7795 38312
rect 6599 38231 7795 38248
rect 6599 38167 6607 38231
rect 6671 38167 6687 38231
rect 6751 38167 6767 38231
rect 6831 38167 6847 38231
rect 6911 38167 6927 38231
rect 6991 38167 7007 38231
rect 7071 38167 7087 38231
rect 7151 38167 7167 38231
rect 7231 38167 7247 38231
rect 7311 38167 7327 38231
rect 7391 38167 7407 38231
rect 7471 38167 7487 38231
rect 7551 38167 7567 38231
rect 7631 38167 7647 38231
rect 7711 38167 7727 38231
rect 7791 38167 7795 38231
rect 6599 38150 7795 38167
rect 6599 38086 6607 38150
rect 6671 38086 6687 38150
rect 6751 38086 6767 38150
rect 6831 38086 6847 38150
rect 6911 38086 6927 38150
rect 6991 38086 7007 38150
rect 7071 38086 7087 38150
rect 7151 38086 7167 38150
rect 7231 38086 7247 38150
rect 7311 38086 7327 38150
rect 7391 38086 7407 38150
rect 7471 38086 7487 38150
rect 7551 38086 7567 38150
rect 7631 38086 7647 38150
rect 7711 38086 7727 38150
rect 7791 38086 7795 38150
rect 6599 38069 7795 38086
rect 6599 38005 6607 38069
rect 6671 38005 6687 38069
rect 6751 38005 6767 38069
rect 6831 38005 6847 38069
rect 6911 38005 6927 38069
rect 6991 38005 7007 38069
rect 7071 38005 7087 38069
rect 7151 38005 7167 38069
rect 7231 38005 7247 38069
rect 7311 38005 7327 38069
rect 7391 38005 7407 38069
rect 7471 38005 7487 38069
rect 7551 38005 7567 38069
rect 7631 38005 7647 38069
rect 7711 38005 7727 38069
rect 7791 38005 7795 38069
rect 6599 37988 7795 38005
rect 6599 37924 6607 37988
rect 6671 37924 6687 37988
rect 6751 37924 6767 37988
rect 6831 37924 6847 37988
rect 6911 37924 6927 37988
rect 6991 37924 7007 37988
rect 7071 37924 7087 37988
rect 7151 37924 7167 37988
rect 7231 37924 7247 37988
rect 7311 37924 7327 37988
rect 7391 37924 7407 37988
rect 7471 37924 7487 37988
rect 7551 37924 7567 37988
rect 7631 37924 7647 37988
rect 7711 37924 7727 37988
rect 7791 37924 7795 37988
rect 6599 37907 7795 37924
rect 6599 37843 6607 37907
rect 6671 37843 6687 37907
rect 6751 37843 6767 37907
rect 6831 37843 6847 37907
rect 6911 37843 6927 37907
rect 6991 37843 7007 37907
rect 7071 37843 7087 37907
rect 7151 37843 7167 37907
rect 7231 37843 7247 37907
rect 7311 37843 7327 37907
rect 7391 37843 7407 37907
rect 7471 37843 7487 37907
rect 7551 37843 7567 37907
rect 7631 37843 7647 37907
rect 7711 37843 7727 37907
rect 7791 37843 7795 37907
rect 6599 37826 7795 37843
rect 6599 37762 6607 37826
rect 6671 37762 6687 37826
rect 6751 37762 6767 37826
rect 6831 37762 6847 37826
rect 6911 37762 6927 37826
rect 6991 37762 7007 37826
rect 7071 37762 7087 37826
rect 7151 37762 7167 37826
rect 7231 37762 7247 37826
rect 7311 37762 7327 37826
rect 7391 37762 7407 37826
rect 7471 37762 7487 37826
rect 7551 37762 7567 37826
rect 7631 37762 7647 37826
rect 7711 37762 7727 37826
rect 7791 37762 7795 37826
rect 6599 37745 7795 37762
rect 6599 37681 6607 37745
rect 6671 37681 6687 37745
rect 6751 37681 6767 37745
rect 6831 37681 6847 37745
rect 6911 37681 6927 37745
rect 6991 37681 7007 37745
rect 7071 37681 7087 37745
rect 7151 37681 7167 37745
rect 7231 37681 7247 37745
rect 7311 37681 7327 37745
rect 7391 37681 7407 37745
rect 7471 37681 7487 37745
rect 7551 37681 7567 37745
rect 7631 37681 7647 37745
rect 7711 37681 7727 37745
rect 7791 37681 7795 37745
rect 6599 37664 7795 37681
rect 6599 37600 6607 37664
rect 6671 37600 6687 37664
rect 6751 37600 6767 37664
rect 6831 37600 6847 37664
rect 6911 37600 6927 37664
rect 6991 37600 7007 37664
rect 7071 37600 7087 37664
rect 7151 37600 7167 37664
rect 7231 37600 7247 37664
rect 7311 37600 7327 37664
rect 7391 37600 7407 37664
rect 7471 37600 7487 37664
rect 7551 37600 7567 37664
rect 7631 37600 7647 37664
rect 7711 37600 7727 37664
rect 7791 37600 7795 37664
rect 6599 37583 7795 37600
rect 6599 37519 6607 37583
rect 6671 37519 6687 37583
rect 6751 37519 6767 37583
rect 6831 37519 6847 37583
rect 6911 37519 6927 37583
rect 6991 37519 7007 37583
rect 7071 37519 7087 37583
rect 7151 37519 7167 37583
rect 7231 37519 7247 37583
rect 7311 37519 7327 37583
rect 7391 37519 7407 37583
rect 7471 37519 7487 37583
rect 7551 37519 7567 37583
rect 7631 37519 7647 37583
rect 7711 37519 7727 37583
rect 7791 37519 7795 37583
rect 6599 37502 7795 37519
rect 6599 37438 6607 37502
rect 6671 37438 6687 37502
rect 6751 37438 6767 37502
rect 6831 37438 6847 37502
rect 6911 37438 6927 37502
rect 6991 37438 7007 37502
rect 7071 37438 7087 37502
rect 7151 37438 7167 37502
rect 7231 37438 7247 37502
rect 7311 37438 7327 37502
rect 7391 37438 7407 37502
rect 7471 37438 7487 37502
rect 7551 37438 7567 37502
rect 7631 37438 7647 37502
rect 7711 37438 7727 37502
rect 7791 37438 7795 37502
rect 6599 37421 7795 37438
rect 6599 37357 6607 37421
rect 6671 37357 6687 37421
rect 6751 37357 6767 37421
rect 6831 37357 6847 37421
rect 6911 37357 6927 37421
rect 6991 37357 7007 37421
rect 7071 37357 7087 37421
rect 7151 37357 7167 37421
rect 7231 37357 7247 37421
rect 7311 37357 7327 37421
rect 7391 37357 7407 37421
rect 7471 37357 7487 37421
rect 7551 37357 7567 37421
rect 7631 37357 7647 37421
rect 7711 37357 7727 37421
rect 7791 37357 7795 37421
rect 6599 37340 7795 37357
rect 6599 37276 6607 37340
rect 6671 37276 6687 37340
rect 6751 37276 6767 37340
rect 6831 37276 6847 37340
rect 6911 37276 6927 37340
rect 6991 37276 7007 37340
rect 7071 37276 7087 37340
rect 7151 37276 7167 37340
rect 7231 37276 7247 37340
rect 7311 37276 7327 37340
rect 7391 37276 7407 37340
rect 7471 37276 7487 37340
rect 7551 37276 7567 37340
rect 7631 37276 7647 37340
rect 7711 37276 7727 37340
rect 7791 37276 7795 37340
rect 6599 37259 7795 37276
rect 6599 37195 6607 37259
rect 6671 37195 6687 37259
rect 6751 37195 6767 37259
rect 6831 37195 6847 37259
rect 6911 37195 6927 37259
rect 6991 37195 7007 37259
rect 7071 37195 7087 37259
rect 7151 37195 7167 37259
rect 7231 37195 7247 37259
rect 7311 37195 7327 37259
rect 7391 37195 7407 37259
rect 7471 37195 7487 37259
rect 7551 37195 7567 37259
rect 7631 37195 7647 37259
rect 7711 37195 7727 37259
rect 7791 37195 7795 37259
rect 6599 37178 7795 37195
rect 6599 37114 6607 37178
rect 6671 37114 6687 37178
rect 6751 37114 6767 37178
rect 6831 37114 6847 37178
rect 6911 37114 6927 37178
rect 6991 37114 7007 37178
rect 7071 37114 7087 37178
rect 7151 37114 7167 37178
rect 7231 37114 7247 37178
rect 7311 37114 7327 37178
rect 7391 37114 7407 37178
rect 7471 37114 7487 37178
rect 7551 37114 7567 37178
rect 7631 37114 7647 37178
rect 7711 37114 7727 37178
rect 7791 37114 7795 37178
rect 6599 37097 7795 37114
rect 6599 37033 6607 37097
rect 6671 37033 6687 37097
rect 6751 37033 6767 37097
rect 6831 37033 6847 37097
rect 6911 37033 6927 37097
rect 6991 37033 7007 37097
rect 7071 37033 7087 37097
rect 7151 37033 7167 37097
rect 7231 37033 7247 37097
rect 7311 37033 7327 37097
rect 7391 37033 7407 37097
rect 7471 37033 7487 37097
rect 7551 37033 7567 37097
rect 7631 37033 7647 37097
rect 7711 37033 7727 37097
rect 7791 37033 7795 37097
rect 6599 37016 7795 37033
rect 6599 36952 6607 37016
rect 6671 36952 6687 37016
rect 6751 36952 6767 37016
rect 6831 36952 6847 37016
rect 6911 36952 6927 37016
rect 6991 36952 7007 37016
rect 7071 36952 7087 37016
rect 7151 36952 7167 37016
rect 7231 36952 7247 37016
rect 7311 36952 7327 37016
rect 7391 36952 7407 37016
rect 7471 36952 7487 37016
rect 7551 36952 7567 37016
rect 7631 36952 7647 37016
rect 7711 36952 7727 37016
rect 7791 36952 7795 37016
rect 6599 36935 7795 36952
rect 6599 36871 6607 36935
rect 6671 36871 6687 36935
rect 6751 36871 6767 36935
rect 6831 36871 6847 36935
rect 6911 36871 6927 36935
rect 6991 36871 7007 36935
rect 7071 36871 7087 36935
rect 7151 36871 7167 36935
rect 7231 36871 7247 36935
rect 7311 36871 7327 36935
rect 7391 36871 7407 36935
rect 7471 36871 7487 36935
rect 7551 36871 7567 36935
rect 7631 36871 7647 36935
rect 7711 36871 7727 36935
rect 7791 36871 7795 36935
rect 6599 36854 7795 36871
rect 6599 36790 6607 36854
rect 6671 36790 6687 36854
rect 6751 36790 6767 36854
rect 6831 36790 6847 36854
rect 6911 36790 6927 36854
rect 6991 36790 7007 36854
rect 7071 36790 7087 36854
rect 7151 36790 7167 36854
rect 7231 36790 7247 36854
rect 7311 36790 7327 36854
rect 7391 36790 7407 36854
rect 7471 36790 7487 36854
rect 7551 36790 7567 36854
rect 7631 36790 7647 36854
rect 7711 36790 7727 36854
rect 7791 36790 7795 36854
rect 6599 36773 7795 36790
rect 6599 36709 6607 36773
rect 6671 36709 6687 36773
rect 6751 36709 6767 36773
rect 6831 36709 6847 36773
rect 6911 36709 6927 36773
rect 6991 36709 7007 36773
rect 7071 36709 7087 36773
rect 7151 36709 7167 36773
rect 7231 36709 7247 36773
rect 7311 36709 7327 36773
rect 7391 36709 7407 36773
rect 7471 36709 7487 36773
rect 7551 36709 7567 36773
rect 7631 36709 7647 36773
rect 7711 36709 7727 36773
rect 7791 36709 7795 36773
rect 6599 36692 7795 36709
rect 6599 36628 6607 36692
rect 6671 36628 6687 36692
rect 6751 36628 6767 36692
rect 6831 36628 6847 36692
rect 6911 36628 6927 36692
rect 6991 36628 7007 36692
rect 7071 36628 7087 36692
rect 7151 36628 7167 36692
rect 7231 36628 7247 36692
rect 7311 36628 7327 36692
rect 7391 36628 7407 36692
rect 7471 36628 7487 36692
rect 7551 36628 7567 36692
rect 7631 36628 7647 36692
rect 7711 36628 7727 36692
rect 7791 36628 7795 36692
rect 6599 36611 7795 36628
rect 6599 36547 6607 36611
rect 6671 36547 6687 36611
rect 6751 36547 6767 36611
rect 6831 36547 6847 36611
rect 6911 36547 6927 36611
rect 6991 36547 7007 36611
rect 7071 36547 7087 36611
rect 7151 36547 7167 36611
rect 7231 36547 7247 36611
rect 7311 36547 7327 36611
rect 7391 36547 7407 36611
rect 7471 36547 7487 36611
rect 7551 36547 7567 36611
rect 7631 36547 7647 36611
rect 7711 36547 7727 36611
rect 7791 36547 7795 36611
rect 6599 36530 7795 36547
rect 6599 36466 6607 36530
rect 6671 36466 6687 36530
rect 6751 36466 6767 36530
rect 6831 36466 6847 36530
rect 6911 36466 6927 36530
rect 6991 36466 7007 36530
rect 7071 36466 7087 36530
rect 7151 36466 7167 36530
rect 7231 36466 7247 36530
rect 7311 36466 7327 36530
rect 7391 36466 7407 36530
rect 7471 36466 7487 36530
rect 7551 36466 7567 36530
rect 7631 36466 7647 36530
rect 7711 36466 7727 36530
rect 7791 36466 7795 36530
rect 6599 36449 7795 36466
rect 6599 36385 6607 36449
rect 6671 36385 6687 36449
rect 6751 36385 6767 36449
rect 6831 36385 6847 36449
rect 6911 36385 6927 36449
rect 6991 36385 7007 36449
rect 7071 36385 7087 36449
rect 7151 36385 7167 36449
rect 7231 36385 7247 36449
rect 7311 36385 7327 36449
rect 7391 36385 7407 36449
rect 7471 36385 7487 36449
rect 7551 36385 7567 36449
rect 7631 36385 7647 36449
rect 7711 36385 7727 36449
rect 7791 36385 7795 36449
rect 6599 36368 7795 36385
rect 6599 36304 6607 36368
rect 6671 36304 6687 36368
rect 6751 36304 6767 36368
rect 6831 36304 6847 36368
rect 6911 36304 6927 36368
rect 6991 36304 7007 36368
rect 7071 36304 7087 36368
rect 7151 36304 7167 36368
rect 7231 36304 7247 36368
rect 7311 36304 7327 36368
rect 7391 36304 7407 36368
rect 7471 36304 7487 36368
rect 7551 36304 7567 36368
rect 7631 36304 7647 36368
rect 7711 36304 7727 36368
rect 7791 36304 7795 36368
rect 6599 36287 7795 36304
rect 6599 36223 6607 36287
rect 6671 36223 6687 36287
rect 6751 36223 6767 36287
rect 6831 36223 6847 36287
rect 6911 36223 6927 36287
rect 6991 36223 7007 36287
rect 7071 36223 7087 36287
rect 7151 36223 7167 36287
rect 7231 36223 7247 36287
rect 7311 36223 7327 36287
rect 7391 36223 7407 36287
rect 7471 36223 7487 36287
rect 7551 36223 7567 36287
rect 7631 36223 7647 36287
rect 7711 36223 7727 36287
rect 7791 36223 7795 36287
rect 6599 36206 7795 36223
rect 6599 36142 6607 36206
rect 6671 36142 6687 36206
rect 6751 36142 6767 36206
rect 6831 36142 6847 36206
rect 6911 36142 6927 36206
rect 6991 36142 7007 36206
rect 7071 36142 7087 36206
rect 7151 36142 7167 36206
rect 7231 36142 7247 36206
rect 7311 36142 7327 36206
rect 7391 36142 7407 36206
rect 7471 36142 7487 36206
rect 7551 36142 7567 36206
rect 7631 36142 7647 36206
rect 7711 36142 7727 36206
rect 7791 36142 7795 36206
rect 6599 36124 7795 36142
rect 6599 36060 6607 36124
rect 6671 36060 6687 36124
rect 6751 36060 6767 36124
rect 6831 36060 6847 36124
rect 6911 36060 6927 36124
rect 6991 36060 7007 36124
rect 7071 36060 7087 36124
rect 7151 36060 7167 36124
rect 7231 36060 7247 36124
rect 7311 36060 7327 36124
rect 7391 36060 7407 36124
rect 7471 36060 7487 36124
rect 7551 36060 7567 36124
rect 7631 36060 7647 36124
rect 7711 36060 7727 36124
rect 7791 36060 7795 36124
rect 6599 36042 7795 36060
rect 6599 35978 6607 36042
rect 6671 35978 6687 36042
rect 6751 35978 6767 36042
rect 6831 35978 6847 36042
rect 6911 35978 6927 36042
rect 6991 35978 7007 36042
rect 7071 35978 7087 36042
rect 7151 35978 7167 36042
rect 7231 35978 7247 36042
rect 7311 35978 7327 36042
rect 7391 35978 7407 36042
rect 7471 35978 7487 36042
rect 7551 35978 7567 36042
rect 7631 35978 7647 36042
rect 7711 35978 7727 36042
rect 7791 35978 7795 36042
rect 6599 35960 7795 35978
rect 6599 35896 6607 35960
rect 6671 35896 6687 35960
rect 6751 35896 6767 35960
rect 6831 35896 6847 35960
rect 6911 35896 6927 35960
rect 6991 35896 7007 35960
rect 7071 35896 7087 35960
rect 7151 35896 7167 35960
rect 7231 35896 7247 35960
rect 7311 35896 7327 35960
rect 7391 35896 7407 35960
rect 7471 35896 7487 35960
rect 7551 35896 7567 35960
rect 7631 35896 7647 35960
rect 7711 35896 7727 35960
rect 7791 35896 7795 35960
rect 6599 35878 7795 35896
rect 6599 35814 6607 35878
rect 6671 35814 6687 35878
rect 6751 35814 6767 35878
rect 6831 35814 6847 35878
rect 6911 35814 6927 35878
rect 6991 35814 7007 35878
rect 7071 35814 7087 35878
rect 7151 35814 7167 35878
rect 7231 35814 7247 35878
rect 7311 35814 7327 35878
rect 7391 35814 7407 35878
rect 7471 35814 7487 35878
rect 7551 35814 7567 35878
rect 7631 35814 7647 35878
rect 7711 35814 7727 35878
rect 7791 35814 7795 35878
rect 6599 35796 7795 35814
rect 6599 35732 6607 35796
rect 6671 35732 6687 35796
rect 6751 35732 6767 35796
rect 6831 35732 6847 35796
rect 6911 35732 6927 35796
rect 6991 35732 7007 35796
rect 7071 35732 7087 35796
rect 7151 35732 7167 35796
rect 7231 35732 7247 35796
rect 7311 35732 7327 35796
rect 7391 35732 7407 35796
rect 7471 35732 7487 35796
rect 7551 35732 7567 35796
rect 7631 35732 7647 35796
rect 7711 35732 7727 35796
rect 7791 35732 7795 35796
rect 6599 35714 7795 35732
rect 6599 35650 6607 35714
rect 6671 35650 6687 35714
rect 6751 35650 6767 35714
rect 6831 35650 6847 35714
rect 6911 35650 6927 35714
rect 6991 35650 7007 35714
rect 7071 35650 7087 35714
rect 7151 35650 7167 35714
rect 7231 35650 7247 35714
rect 7311 35650 7327 35714
rect 7391 35650 7407 35714
rect 7471 35650 7487 35714
rect 7551 35650 7567 35714
rect 7631 35650 7647 35714
rect 7711 35650 7727 35714
rect 7791 35650 7795 35714
rect 6599 35632 7795 35650
rect 6599 35568 6607 35632
rect 6671 35568 6687 35632
rect 6751 35568 6767 35632
rect 6831 35568 6847 35632
rect 6911 35568 6927 35632
rect 6991 35568 7007 35632
rect 7071 35568 7087 35632
rect 7151 35568 7167 35632
rect 7231 35568 7247 35632
rect 7311 35568 7327 35632
rect 7391 35568 7407 35632
rect 7471 35568 7487 35632
rect 7551 35568 7567 35632
rect 7631 35568 7647 35632
rect 7711 35568 7727 35632
rect 7791 35568 7795 35632
rect 6599 35550 7795 35568
rect 6599 35486 6607 35550
rect 6671 35486 6687 35550
rect 6751 35486 6767 35550
rect 6831 35486 6847 35550
rect 6911 35486 6927 35550
rect 6991 35486 7007 35550
rect 7071 35486 7087 35550
rect 7151 35486 7167 35550
rect 7231 35486 7247 35550
rect 7311 35486 7327 35550
rect 7391 35486 7407 35550
rect 7471 35486 7487 35550
rect 7551 35486 7567 35550
rect 7631 35486 7647 35550
rect 7711 35486 7727 35550
rect 7791 35486 7795 35550
rect 6599 35468 7795 35486
rect 6599 35404 6607 35468
rect 6671 35404 6687 35468
rect 6751 35404 6767 35468
rect 6831 35404 6847 35468
rect 6911 35404 6927 35468
rect 6991 35404 7007 35468
rect 7071 35404 7087 35468
rect 7151 35404 7167 35468
rect 7231 35404 7247 35468
rect 7311 35404 7327 35468
rect 7391 35404 7407 35468
rect 7471 35404 7487 35468
rect 7551 35404 7567 35468
rect 7631 35404 7647 35468
rect 7711 35404 7727 35468
rect 7791 35404 7795 35468
rect 6599 35386 7795 35404
rect 6599 35322 6607 35386
rect 6671 35322 6687 35386
rect 6751 35322 6767 35386
rect 6831 35322 6847 35386
rect 6911 35322 6927 35386
rect 6991 35322 7007 35386
rect 7071 35322 7087 35386
rect 7151 35322 7167 35386
rect 7231 35322 7247 35386
rect 7311 35322 7327 35386
rect 7391 35322 7407 35386
rect 7471 35322 7487 35386
rect 7551 35322 7567 35386
rect 7631 35322 7647 35386
rect 7711 35322 7727 35386
rect 7791 35322 7795 35386
rect 6599 35304 7795 35322
rect 6599 35240 6607 35304
rect 6671 35240 6687 35304
rect 6751 35240 6767 35304
rect 6831 35240 6847 35304
rect 6911 35240 6927 35304
rect 6991 35240 7007 35304
rect 7071 35240 7087 35304
rect 7151 35240 7167 35304
rect 7231 35240 7247 35304
rect 7311 35240 7327 35304
rect 7391 35240 7407 35304
rect 7471 35240 7487 35304
rect 7551 35240 7567 35304
rect 7631 35240 7647 35304
rect 7711 35240 7727 35304
rect 7791 35240 7795 35304
rect 6599 35222 7795 35240
rect 6599 35158 6607 35222
rect 6671 35158 6687 35222
rect 6751 35158 6767 35222
rect 6831 35158 6847 35222
rect 6911 35158 6927 35222
rect 6991 35158 7007 35222
rect 7071 35158 7087 35222
rect 7151 35158 7167 35222
rect 7231 35158 7247 35222
rect 7311 35158 7327 35222
rect 7391 35158 7407 35222
rect 7471 35158 7487 35222
rect 7551 35158 7567 35222
rect 7631 35158 7647 35222
rect 7711 35158 7727 35222
rect 7791 35158 7795 35222
rect 6599 32613 7795 35158
rect 6599 32557 6610 32613
rect 6666 32557 6691 32613
rect 6747 32557 6772 32613
rect 6828 32557 6853 32613
rect 6909 32557 6934 32613
rect 6990 32557 7014 32613
rect 7070 32557 7094 32613
rect 7150 32557 7174 32613
rect 7230 32557 7254 32613
rect 7310 32557 7334 32613
rect 7390 32557 7414 32613
rect 7470 32557 7494 32613
rect 7550 32557 7574 32613
rect 7630 32557 7654 32613
rect 7710 32557 7734 32613
rect 7790 32557 7795 32613
rect 6599 32531 7795 32557
rect 6599 32475 6610 32531
rect 6666 32475 6691 32531
rect 6747 32475 6772 32531
rect 6828 32475 6853 32531
rect 6909 32475 6934 32531
rect 6990 32475 7014 32531
rect 7070 32475 7094 32531
rect 7150 32475 7174 32531
rect 7230 32475 7254 32531
rect 7310 32475 7334 32531
rect 7390 32475 7414 32531
rect 7470 32475 7494 32531
rect 7550 32475 7574 32531
rect 7630 32475 7654 32531
rect 7710 32475 7734 32531
rect 7790 32475 7795 32531
rect 6599 32449 7795 32475
rect 6599 32393 6610 32449
rect 6666 32393 6691 32449
rect 6747 32393 6772 32449
rect 6828 32393 6853 32449
rect 6909 32393 6934 32449
rect 6990 32393 7014 32449
rect 7070 32393 7094 32449
rect 7150 32393 7174 32449
rect 7230 32393 7254 32449
rect 7310 32393 7334 32449
rect 7390 32393 7414 32449
rect 7470 32393 7494 32449
rect 7550 32393 7574 32449
rect 7630 32393 7654 32449
rect 7710 32393 7734 32449
rect 7790 32393 7795 32449
rect 6599 32367 7795 32393
rect 6599 32311 6610 32367
rect 6666 32311 6691 32367
rect 6747 32311 6772 32367
rect 6828 32311 6853 32367
rect 6909 32311 6934 32367
rect 6990 32311 7014 32367
rect 7070 32311 7094 32367
rect 7150 32311 7174 32367
rect 7230 32311 7254 32367
rect 7310 32311 7334 32367
rect 7390 32311 7414 32367
rect 7470 32311 7494 32367
rect 7550 32311 7574 32367
rect 7630 32311 7654 32367
rect 7710 32311 7734 32367
rect 7790 32311 7795 32367
rect 6599 32285 7795 32311
rect 6599 32229 6610 32285
rect 6666 32229 6691 32285
rect 6747 32229 6772 32285
rect 6828 32229 6853 32285
rect 6909 32229 6934 32285
rect 6990 32229 7014 32285
rect 7070 32229 7094 32285
rect 7150 32229 7174 32285
rect 7230 32229 7254 32285
rect 7310 32229 7334 32285
rect 7390 32229 7414 32285
rect 7470 32229 7494 32285
rect 7550 32229 7574 32285
rect 7630 32229 7654 32285
rect 7710 32229 7734 32285
rect 7790 32229 7795 32285
rect 6599 32203 7795 32229
rect 6599 32147 6610 32203
rect 6666 32147 6691 32203
rect 6747 32147 6772 32203
rect 6828 32147 6853 32203
rect 6909 32147 6934 32203
rect 6990 32147 7014 32203
rect 7070 32147 7094 32203
rect 7150 32147 7174 32203
rect 7230 32147 7254 32203
rect 7310 32147 7334 32203
rect 7390 32147 7414 32203
rect 7470 32147 7494 32203
rect 7550 32147 7574 32203
rect 7630 32147 7654 32203
rect 7710 32147 7734 32203
rect 7790 32147 7795 32203
rect 6599 32121 7795 32147
rect 6599 32065 6610 32121
rect 6666 32065 6691 32121
rect 6747 32065 6772 32121
rect 6828 32065 6853 32121
rect 6909 32065 6934 32121
rect 6990 32065 7014 32121
rect 7070 32065 7094 32121
rect 7150 32065 7174 32121
rect 7230 32065 7254 32121
rect 7310 32065 7334 32121
rect 7390 32065 7414 32121
rect 7470 32065 7494 32121
rect 7550 32065 7574 32121
rect 7630 32065 7654 32121
rect 7710 32065 7734 32121
rect 7790 32065 7795 32121
rect 6599 32039 7795 32065
rect 6599 31983 6610 32039
rect 6666 31983 6691 32039
rect 6747 31983 6772 32039
rect 6828 31983 6853 32039
rect 6909 31983 6934 32039
rect 6990 31983 7014 32039
rect 7070 31983 7094 32039
rect 7150 31983 7174 32039
rect 7230 31983 7254 32039
rect 7310 31983 7334 32039
rect 7390 31983 7414 32039
rect 7470 31983 7494 32039
rect 7550 31983 7574 32039
rect 7630 31983 7654 32039
rect 7710 31983 7734 32039
rect 7790 31983 7795 32039
rect 6599 31957 7795 31983
rect 6599 31901 6610 31957
rect 6666 31901 6691 31957
rect 6747 31901 6772 31957
rect 6828 31901 6853 31957
rect 6909 31901 6934 31957
rect 6990 31901 7014 31957
rect 7070 31901 7094 31957
rect 7150 31901 7174 31957
rect 7230 31901 7254 31957
rect 7310 31901 7334 31957
rect 7390 31901 7414 31957
rect 7470 31901 7494 31957
rect 7550 31901 7574 31957
rect 7630 31901 7654 31957
rect 7710 31901 7734 31957
rect 7790 31901 7795 31957
rect 6599 31875 7795 31901
rect 6599 31819 6610 31875
rect 6666 31819 6691 31875
rect 6747 31819 6772 31875
rect 6828 31819 6853 31875
rect 6909 31819 6934 31875
rect 6990 31819 7014 31875
rect 7070 31819 7094 31875
rect 7150 31819 7174 31875
rect 7230 31819 7254 31875
rect 7310 31819 7334 31875
rect 7390 31819 7414 31875
rect 7470 31819 7494 31875
rect 7550 31819 7574 31875
rect 7630 31819 7654 31875
rect 7710 31819 7734 31875
rect 7790 31819 7795 31875
rect 6599 31793 7795 31819
rect 6599 31737 6610 31793
rect 6666 31737 6691 31793
rect 6747 31737 6772 31793
rect 6828 31737 6853 31793
rect 6909 31737 6934 31793
rect 6990 31737 7014 31793
rect 7070 31737 7094 31793
rect 7150 31737 7174 31793
rect 7230 31737 7254 31793
rect 7310 31737 7334 31793
rect 7390 31737 7414 31793
rect 7470 31737 7494 31793
rect 7550 31737 7574 31793
rect 7630 31737 7654 31793
rect 7710 31737 7734 31793
rect 7790 31737 7795 31793
rect 6599 31711 7795 31737
rect 6599 31655 6610 31711
rect 6666 31655 6691 31711
rect 6747 31655 6772 31711
rect 6828 31655 6853 31711
rect 6909 31655 6934 31711
rect 6990 31655 7014 31711
rect 7070 31655 7094 31711
rect 7150 31655 7174 31711
rect 7230 31655 7254 31711
rect 7310 31655 7334 31711
rect 7390 31655 7414 31711
rect 7470 31655 7494 31711
rect 7550 31655 7574 31711
rect 7630 31655 7654 31711
rect 7710 31655 7734 31711
rect 7790 31655 7795 31711
rect 6599 31629 7795 31655
rect 6599 31573 6610 31629
rect 6666 31573 6691 31629
rect 6747 31573 6772 31629
rect 6828 31573 6853 31629
rect 6909 31573 6934 31629
rect 6990 31573 7014 31629
rect 7070 31573 7094 31629
rect 7150 31573 7174 31629
rect 7230 31573 7254 31629
rect 7310 31573 7334 31629
rect 7390 31573 7414 31629
rect 7470 31573 7494 31629
rect 7550 31573 7574 31629
rect 7630 31573 7654 31629
rect 7710 31573 7734 31629
rect 7790 31573 7795 31629
rect 6599 31547 7795 31573
rect 6599 31491 6610 31547
rect 6666 31491 6691 31547
rect 6747 31491 6772 31547
rect 6828 31491 6853 31547
rect 6909 31491 6934 31547
rect 6990 31491 7014 31547
rect 7070 31491 7094 31547
rect 7150 31491 7174 31547
rect 7230 31491 7254 31547
rect 7310 31491 7334 31547
rect 7390 31491 7414 31547
rect 7470 31491 7494 31547
rect 7550 31491 7574 31547
rect 7630 31491 7654 31547
rect 7710 31491 7734 31547
rect 7790 31491 7795 31547
rect 6599 31478 7795 31491
rect 8096 39365 9292 39371
rect 8096 39301 8100 39365
rect 8164 39301 8180 39365
rect 8244 39301 8260 39365
rect 8324 39301 8340 39365
rect 8404 39301 8420 39365
rect 8484 39301 8500 39365
rect 8564 39301 8580 39365
rect 8644 39301 8660 39365
rect 8724 39301 8740 39365
rect 8804 39301 8820 39365
rect 8884 39301 8900 39365
rect 8964 39301 8980 39365
rect 9044 39301 9060 39365
rect 9124 39301 9140 39365
rect 9204 39301 9220 39365
rect 9284 39301 9292 39365
rect 8096 39284 9292 39301
rect 8096 39220 8100 39284
rect 8164 39220 8180 39284
rect 8244 39220 8260 39284
rect 8324 39220 8340 39284
rect 8404 39220 8420 39284
rect 8484 39220 8500 39284
rect 8564 39220 8580 39284
rect 8644 39220 8660 39284
rect 8724 39220 8740 39284
rect 8804 39220 8820 39284
rect 8884 39220 8900 39284
rect 8964 39220 8980 39284
rect 9044 39220 9060 39284
rect 9124 39220 9140 39284
rect 9204 39220 9220 39284
rect 9284 39220 9292 39284
rect 8096 39203 9292 39220
rect 8096 39139 8100 39203
rect 8164 39139 8180 39203
rect 8244 39139 8260 39203
rect 8324 39139 8340 39203
rect 8404 39139 8420 39203
rect 8484 39139 8500 39203
rect 8564 39139 8580 39203
rect 8644 39139 8660 39203
rect 8724 39139 8740 39203
rect 8804 39139 8820 39203
rect 8884 39139 8900 39203
rect 8964 39139 8980 39203
rect 9044 39139 9060 39203
rect 9124 39139 9140 39203
rect 9204 39139 9220 39203
rect 9284 39139 9292 39203
rect 8096 39122 9292 39139
rect 8096 39058 8100 39122
rect 8164 39058 8180 39122
rect 8244 39058 8260 39122
rect 8324 39058 8340 39122
rect 8404 39058 8420 39122
rect 8484 39058 8500 39122
rect 8564 39058 8580 39122
rect 8644 39058 8660 39122
rect 8724 39058 8740 39122
rect 8804 39058 8820 39122
rect 8884 39058 8900 39122
rect 8964 39058 8980 39122
rect 9044 39058 9060 39122
rect 9124 39058 9140 39122
rect 9204 39058 9220 39122
rect 9284 39058 9292 39122
rect 8096 39041 9292 39058
rect 8096 38977 8100 39041
rect 8164 38977 8180 39041
rect 8244 38977 8260 39041
rect 8324 38977 8340 39041
rect 8404 38977 8420 39041
rect 8484 38977 8500 39041
rect 8564 38977 8580 39041
rect 8644 38977 8660 39041
rect 8724 38977 8740 39041
rect 8804 38977 8820 39041
rect 8884 38977 8900 39041
rect 8964 38977 8980 39041
rect 9044 38977 9060 39041
rect 9124 38977 9140 39041
rect 9204 38977 9220 39041
rect 9284 38977 9292 39041
rect 8096 38960 9292 38977
rect 8096 38896 8100 38960
rect 8164 38896 8180 38960
rect 8244 38896 8260 38960
rect 8324 38896 8340 38960
rect 8404 38896 8420 38960
rect 8484 38896 8500 38960
rect 8564 38896 8580 38960
rect 8644 38896 8660 38960
rect 8724 38896 8740 38960
rect 8804 38896 8820 38960
rect 8884 38896 8900 38960
rect 8964 38896 8980 38960
rect 9044 38896 9060 38960
rect 9124 38896 9140 38960
rect 9204 38896 9220 38960
rect 9284 38896 9292 38960
rect 8096 38879 9292 38896
rect 8096 38815 8100 38879
rect 8164 38815 8180 38879
rect 8244 38815 8260 38879
rect 8324 38815 8340 38879
rect 8404 38815 8420 38879
rect 8484 38815 8500 38879
rect 8564 38815 8580 38879
rect 8644 38815 8660 38879
rect 8724 38815 8740 38879
rect 8804 38815 8820 38879
rect 8884 38815 8900 38879
rect 8964 38815 8980 38879
rect 9044 38815 9060 38879
rect 9124 38815 9140 38879
rect 9204 38815 9220 38879
rect 9284 38815 9292 38879
rect 8096 38798 9292 38815
rect 8096 38734 8100 38798
rect 8164 38734 8180 38798
rect 8244 38734 8260 38798
rect 8324 38734 8340 38798
rect 8404 38734 8420 38798
rect 8484 38734 8500 38798
rect 8564 38734 8580 38798
rect 8644 38734 8660 38798
rect 8724 38734 8740 38798
rect 8804 38734 8820 38798
rect 8884 38734 8900 38798
rect 8964 38734 8980 38798
rect 9044 38734 9060 38798
rect 9124 38734 9140 38798
rect 9204 38734 9220 38798
rect 9284 38734 9292 38798
rect 8096 38717 9292 38734
rect 8096 38653 8100 38717
rect 8164 38653 8180 38717
rect 8244 38653 8260 38717
rect 8324 38653 8340 38717
rect 8404 38653 8420 38717
rect 8484 38653 8500 38717
rect 8564 38653 8580 38717
rect 8644 38653 8660 38717
rect 8724 38653 8740 38717
rect 8804 38653 8820 38717
rect 8884 38653 8900 38717
rect 8964 38653 8980 38717
rect 9044 38653 9060 38717
rect 9124 38653 9140 38717
rect 9204 38653 9220 38717
rect 9284 38653 9292 38717
rect 8096 38636 9292 38653
rect 8096 38572 8100 38636
rect 8164 38572 8180 38636
rect 8244 38572 8260 38636
rect 8324 38572 8340 38636
rect 8404 38572 8420 38636
rect 8484 38572 8500 38636
rect 8564 38572 8580 38636
rect 8644 38572 8660 38636
rect 8724 38572 8740 38636
rect 8804 38572 8820 38636
rect 8884 38572 8900 38636
rect 8964 38572 8980 38636
rect 9044 38572 9060 38636
rect 9124 38572 9140 38636
rect 9204 38572 9220 38636
rect 9284 38572 9292 38636
rect 8096 38555 9292 38572
rect 8096 38491 8100 38555
rect 8164 38491 8180 38555
rect 8244 38491 8260 38555
rect 8324 38491 8340 38555
rect 8404 38491 8420 38555
rect 8484 38491 8500 38555
rect 8564 38491 8580 38555
rect 8644 38491 8660 38555
rect 8724 38491 8740 38555
rect 8804 38491 8820 38555
rect 8884 38491 8900 38555
rect 8964 38491 8980 38555
rect 9044 38491 9060 38555
rect 9124 38491 9140 38555
rect 9204 38491 9220 38555
rect 9284 38491 9292 38555
rect 8096 38474 9292 38491
rect 8096 38410 8100 38474
rect 8164 38410 8180 38474
rect 8244 38410 8260 38474
rect 8324 38410 8340 38474
rect 8404 38410 8420 38474
rect 8484 38410 8500 38474
rect 8564 38410 8580 38474
rect 8644 38410 8660 38474
rect 8724 38410 8740 38474
rect 8804 38410 8820 38474
rect 8884 38410 8900 38474
rect 8964 38410 8980 38474
rect 9044 38410 9060 38474
rect 9124 38410 9140 38474
rect 9204 38410 9220 38474
rect 9284 38410 9292 38474
rect 8096 38393 9292 38410
rect 8096 38329 8100 38393
rect 8164 38329 8180 38393
rect 8244 38329 8260 38393
rect 8324 38329 8340 38393
rect 8404 38329 8420 38393
rect 8484 38329 8500 38393
rect 8564 38329 8580 38393
rect 8644 38329 8660 38393
rect 8724 38329 8740 38393
rect 8804 38329 8820 38393
rect 8884 38329 8900 38393
rect 8964 38329 8980 38393
rect 9044 38329 9060 38393
rect 9124 38329 9140 38393
rect 9204 38329 9220 38393
rect 9284 38329 9292 38393
rect 8096 38312 9292 38329
rect 8096 38248 8100 38312
rect 8164 38248 8180 38312
rect 8244 38248 8260 38312
rect 8324 38248 8340 38312
rect 8404 38248 8420 38312
rect 8484 38248 8500 38312
rect 8564 38248 8580 38312
rect 8644 38248 8660 38312
rect 8724 38248 8740 38312
rect 8804 38248 8820 38312
rect 8884 38248 8900 38312
rect 8964 38248 8980 38312
rect 9044 38248 9060 38312
rect 9124 38248 9140 38312
rect 9204 38248 9220 38312
rect 9284 38248 9292 38312
rect 8096 38231 9292 38248
rect 8096 38167 8100 38231
rect 8164 38167 8180 38231
rect 8244 38167 8260 38231
rect 8324 38167 8340 38231
rect 8404 38167 8420 38231
rect 8484 38167 8500 38231
rect 8564 38167 8580 38231
rect 8644 38167 8660 38231
rect 8724 38167 8740 38231
rect 8804 38167 8820 38231
rect 8884 38167 8900 38231
rect 8964 38167 8980 38231
rect 9044 38167 9060 38231
rect 9124 38167 9140 38231
rect 9204 38167 9220 38231
rect 9284 38167 9292 38231
rect 8096 38150 9292 38167
rect 8096 38086 8100 38150
rect 8164 38086 8180 38150
rect 8244 38086 8260 38150
rect 8324 38086 8340 38150
rect 8404 38086 8420 38150
rect 8484 38086 8500 38150
rect 8564 38086 8580 38150
rect 8644 38086 8660 38150
rect 8724 38086 8740 38150
rect 8804 38086 8820 38150
rect 8884 38086 8900 38150
rect 8964 38086 8980 38150
rect 9044 38086 9060 38150
rect 9124 38086 9140 38150
rect 9204 38086 9220 38150
rect 9284 38086 9292 38150
rect 8096 38069 9292 38086
rect 8096 38005 8100 38069
rect 8164 38005 8180 38069
rect 8244 38005 8260 38069
rect 8324 38005 8340 38069
rect 8404 38005 8420 38069
rect 8484 38005 8500 38069
rect 8564 38005 8580 38069
rect 8644 38005 8660 38069
rect 8724 38005 8740 38069
rect 8804 38005 8820 38069
rect 8884 38005 8900 38069
rect 8964 38005 8980 38069
rect 9044 38005 9060 38069
rect 9124 38005 9140 38069
rect 9204 38005 9220 38069
rect 9284 38005 9292 38069
rect 8096 37988 9292 38005
rect 8096 37924 8100 37988
rect 8164 37924 8180 37988
rect 8244 37924 8260 37988
rect 8324 37924 8340 37988
rect 8404 37924 8420 37988
rect 8484 37924 8500 37988
rect 8564 37924 8580 37988
rect 8644 37924 8660 37988
rect 8724 37924 8740 37988
rect 8804 37924 8820 37988
rect 8884 37924 8900 37988
rect 8964 37924 8980 37988
rect 9044 37924 9060 37988
rect 9124 37924 9140 37988
rect 9204 37924 9220 37988
rect 9284 37924 9292 37988
rect 8096 37907 9292 37924
rect 8096 37843 8100 37907
rect 8164 37843 8180 37907
rect 8244 37843 8260 37907
rect 8324 37843 8340 37907
rect 8404 37843 8420 37907
rect 8484 37843 8500 37907
rect 8564 37843 8580 37907
rect 8644 37843 8660 37907
rect 8724 37843 8740 37907
rect 8804 37843 8820 37907
rect 8884 37843 8900 37907
rect 8964 37843 8980 37907
rect 9044 37843 9060 37907
rect 9124 37843 9140 37907
rect 9204 37843 9220 37907
rect 9284 37843 9292 37907
rect 8096 37826 9292 37843
rect 8096 37762 8100 37826
rect 8164 37762 8180 37826
rect 8244 37762 8260 37826
rect 8324 37762 8340 37826
rect 8404 37762 8420 37826
rect 8484 37762 8500 37826
rect 8564 37762 8580 37826
rect 8644 37762 8660 37826
rect 8724 37762 8740 37826
rect 8804 37762 8820 37826
rect 8884 37762 8900 37826
rect 8964 37762 8980 37826
rect 9044 37762 9060 37826
rect 9124 37762 9140 37826
rect 9204 37762 9220 37826
rect 9284 37762 9292 37826
rect 8096 37745 9292 37762
rect 8096 37681 8100 37745
rect 8164 37681 8180 37745
rect 8244 37681 8260 37745
rect 8324 37681 8340 37745
rect 8404 37681 8420 37745
rect 8484 37681 8500 37745
rect 8564 37681 8580 37745
rect 8644 37681 8660 37745
rect 8724 37681 8740 37745
rect 8804 37681 8820 37745
rect 8884 37681 8900 37745
rect 8964 37681 8980 37745
rect 9044 37681 9060 37745
rect 9124 37681 9140 37745
rect 9204 37681 9220 37745
rect 9284 37681 9292 37745
rect 8096 37664 9292 37681
rect 8096 37600 8100 37664
rect 8164 37600 8180 37664
rect 8244 37600 8260 37664
rect 8324 37600 8340 37664
rect 8404 37600 8420 37664
rect 8484 37600 8500 37664
rect 8564 37600 8580 37664
rect 8644 37600 8660 37664
rect 8724 37600 8740 37664
rect 8804 37600 8820 37664
rect 8884 37600 8900 37664
rect 8964 37600 8980 37664
rect 9044 37600 9060 37664
rect 9124 37600 9140 37664
rect 9204 37600 9220 37664
rect 9284 37600 9292 37664
rect 8096 37583 9292 37600
rect 8096 37519 8100 37583
rect 8164 37519 8180 37583
rect 8244 37519 8260 37583
rect 8324 37519 8340 37583
rect 8404 37519 8420 37583
rect 8484 37519 8500 37583
rect 8564 37519 8580 37583
rect 8644 37519 8660 37583
rect 8724 37519 8740 37583
rect 8804 37519 8820 37583
rect 8884 37519 8900 37583
rect 8964 37519 8980 37583
rect 9044 37519 9060 37583
rect 9124 37519 9140 37583
rect 9204 37519 9220 37583
rect 9284 37519 9292 37583
rect 8096 37502 9292 37519
rect 8096 37438 8100 37502
rect 8164 37438 8180 37502
rect 8244 37438 8260 37502
rect 8324 37438 8340 37502
rect 8404 37438 8420 37502
rect 8484 37438 8500 37502
rect 8564 37438 8580 37502
rect 8644 37438 8660 37502
rect 8724 37438 8740 37502
rect 8804 37438 8820 37502
rect 8884 37438 8900 37502
rect 8964 37438 8980 37502
rect 9044 37438 9060 37502
rect 9124 37438 9140 37502
rect 9204 37438 9220 37502
rect 9284 37438 9292 37502
rect 8096 37421 9292 37438
rect 8096 37357 8100 37421
rect 8164 37357 8180 37421
rect 8244 37357 8260 37421
rect 8324 37357 8340 37421
rect 8404 37357 8420 37421
rect 8484 37357 8500 37421
rect 8564 37357 8580 37421
rect 8644 37357 8660 37421
rect 8724 37357 8740 37421
rect 8804 37357 8820 37421
rect 8884 37357 8900 37421
rect 8964 37357 8980 37421
rect 9044 37357 9060 37421
rect 9124 37357 9140 37421
rect 9204 37357 9220 37421
rect 9284 37357 9292 37421
rect 8096 37340 9292 37357
rect 8096 37276 8100 37340
rect 8164 37276 8180 37340
rect 8244 37276 8260 37340
rect 8324 37276 8340 37340
rect 8404 37276 8420 37340
rect 8484 37276 8500 37340
rect 8564 37276 8580 37340
rect 8644 37276 8660 37340
rect 8724 37276 8740 37340
rect 8804 37276 8820 37340
rect 8884 37276 8900 37340
rect 8964 37276 8980 37340
rect 9044 37276 9060 37340
rect 9124 37276 9140 37340
rect 9204 37276 9220 37340
rect 9284 37276 9292 37340
rect 8096 37259 9292 37276
rect 8096 37195 8100 37259
rect 8164 37195 8180 37259
rect 8244 37195 8260 37259
rect 8324 37195 8340 37259
rect 8404 37195 8420 37259
rect 8484 37195 8500 37259
rect 8564 37195 8580 37259
rect 8644 37195 8660 37259
rect 8724 37195 8740 37259
rect 8804 37195 8820 37259
rect 8884 37195 8900 37259
rect 8964 37195 8980 37259
rect 9044 37195 9060 37259
rect 9124 37195 9140 37259
rect 9204 37195 9220 37259
rect 9284 37195 9292 37259
rect 8096 37178 9292 37195
rect 8096 37114 8100 37178
rect 8164 37114 8180 37178
rect 8244 37114 8260 37178
rect 8324 37114 8340 37178
rect 8404 37114 8420 37178
rect 8484 37114 8500 37178
rect 8564 37114 8580 37178
rect 8644 37114 8660 37178
rect 8724 37114 8740 37178
rect 8804 37114 8820 37178
rect 8884 37114 8900 37178
rect 8964 37114 8980 37178
rect 9044 37114 9060 37178
rect 9124 37114 9140 37178
rect 9204 37114 9220 37178
rect 9284 37114 9292 37178
rect 8096 37097 9292 37114
rect 8096 37033 8100 37097
rect 8164 37033 8180 37097
rect 8244 37033 8260 37097
rect 8324 37033 8340 37097
rect 8404 37033 8420 37097
rect 8484 37033 8500 37097
rect 8564 37033 8580 37097
rect 8644 37033 8660 37097
rect 8724 37033 8740 37097
rect 8804 37033 8820 37097
rect 8884 37033 8900 37097
rect 8964 37033 8980 37097
rect 9044 37033 9060 37097
rect 9124 37033 9140 37097
rect 9204 37033 9220 37097
rect 9284 37033 9292 37097
rect 8096 37016 9292 37033
rect 8096 36952 8100 37016
rect 8164 36952 8180 37016
rect 8244 36952 8260 37016
rect 8324 36952 8340 37016
rect 8404 36952 8420 37016
rect 8484 36952 8500 37016
rect 8564 36952 8580 37016
rect 8644 36952 8660 37016
rect 8724 36952 8740 37016
rect 8804 36952 8820 37016
rect 8884 36952 8900 37016
rect 8964 36952 8980 37016
rect 9044 36952 9060 37016
rect 9124 36952 9140 37016
rect 9204 36952 9220 37016
rect 9284 36952 9292 37016
rect 8096 36935 9292 36952
rect 8096 36871 8100 36935
rect 8164 36871 8180 36935
rect 8244 36871 8260 36935
rect 8324 36871 8340 36935
rect 8404 36871 8420 36935
rect 8484 36871 8500 36935
rect 8564 36871 8580 36935
rect 8644 36871 8660 36935
rect 8724 36871 8740 36935
rect 8804 36871 8820 36935
rect 8884 36871 8900 36935
rect 8964 36871 8980 36935
rect 9044 36871 9060 36935
rect 9124 36871 9140 36935
rect 9204 36871 9220 36935
rect 9284 36871 9292 36935
rect 8096 36854 9292 36871
rect 8096 36790 8100 36854
rect 8164 36790 8180 36854
rect 8244 36790 8260 36854
rect 8324 36790 8340 36854
rect 8404 36790 8420 36854
rect 8484 36790 8500 36854
rect 8564 36790 8580 36854
rect 8644 36790 8660 36854
rect 8724 36790 8740 36854
rect 8804 36790 8820 36854
rect 8884 36790 8900 36854
rect 8964 36790 8980 36854
rect 9044 36790 9060 36854
rect 9124 36790 9140 36854
rect 9204 36790 9220 36854
rect 9284 36790 9292 36854
rect 8096 36773 9292 36790
rect 8096 36709 8100 36773
rect 8164 36709 8180 36773
rect 8244 36709 8260 36773
rect 8324 36709 8340 36773
rect 8404 36709 8420 36773
rect 8484 36709 8500 36773
rect 8564 36709 8580 36773
rect 8644 36709 8660 36773
rect 8724 36709 8740 36773
rect 8804 36709 8820 36773
rect 8884 36709 8900 36773
rect 8964 36709 8980 36773
rect 9044 36709 9060 36773
rect 9124 36709 9140 36773
rect 9204 36709 9220 36773
rect 9284 36709 9292 36773
rect 8096 36692 9292 36709
rect 8096 36628 8100 36692
rect 8164 36628 8180 36692
rect 8244 36628 8260 36692
rect 8324 36628 8340 36692
rect 8404 36628 8420 36692
rect 8484 36628 8500 36692
rect 8564 36628 8580 36692
rect 8644 36628 8660 36692
rect 8724 36628 8740 36692
rect 8804 36628 8820 36692
rect 8884 36628 8900 36692
rect 8964 36628 8980 36692
rect 9044 36628 9060 36692
rect 9124 36628 9140 36692
rect 9204 36628 9220 36692
rect 9284 36628 9292 36692
rect 8096 36611 9292 36628
rect 8096 36547 8100 36611
rect 8164 36547 8180 36611
rect 8244 36547 8260 36611
rect 8324 36547 8340 36611
rect 8404 36547 8420 36611
rect 8484 36547 8500 36611
rect 8564 36547 8580 36611
rect 8644 36547 8660 36611
rect 8724 36547 8740 36611
rect 8804 36547 8820 36611
rect 8884 36547 8900 36611
rect 8964 36547 8980 36611
rect 9044 36547 9060 36611
rect 9124 36547 9140 36611
rect 9204 36547 9220 36611
rect 9284 36547 9292 36611
rect 8096 36530 9292 36547
rect 8096 36466 8100 36530
rect 8164 36466 8180 36530
rect 8244 36466 8260 36530
rect 8324 36466 8340 36530
rect 8404 36466 8420 36530
rect 8484 36466 8500 36530
rect 8564 36466 8580 36530
rect 8644 36466 8660 36530
rect 8724 36466 8740 36530
rect 8804 36466 8820 36530
rect 8884 36466 8900 36530
rect 8964 36466 8980 36530
rect 9044 36466 9060 36530
rect 9124 36466 9140 36530
rect 9204 36466 9220 36530
rect 9284 36466 9292 36530
rect 8096 36449 9292 36466
rect 8096 36385 8100 36449
rect 8164 36385 8180 36449
rect 8244 36385 8260 36449
rect 8324 36385 8340 36449
rect 8404 36385 8420 36449
rect 8484 36385 8500 36449
rect 8564 36385 8580 36449
rect 8644 36385 8660 36449
rect 8724 36385 8740 36449
rect 8804 36385 8820 36449
rect 8884 36385 8900 36449
rect 8964 36385 8980 36449
rect 9044 36385 9060 36449
rect 9124 36385 9140 36449
rect 9204 36385 9220 36449
rect 9284 36385 9292 36449
rect 8096 36368 9292 36385
rect 8096 36304 8100 36368
rect 8164 36304 8180 36368
rect 8244 36304 8260 36368
rect 8324 36304 8340 36368
rect 8404 36304 8420 36368
rect 8484 36304 8500 36368
rect 8564 36304 8580 36368
rect 8644 36304 8660 36368
rect 8724 36304 8740 36368
rect 8804 36304 8820 36368
rect 8884 36304 8900 36368
rect 8964 36304 8980 36368
rect 9044 36304 9060 36368
rect 9124 36304 9140 36368
rect 9204 36304 9220 36368
rect 9284 36304 9292 36368
rect 8096 36287 9292 36304
rect 8096 36223 8100 36287
rect 8164 36223 8180 36287
rect 8244 36223 8260 36287
rect 8324 36223 8340 36287
rect 8404 36223 8420 36287
rect 8484 36223 8500 36287
rect 8564 36223 8580 36287
rect 8644 36223 8660 36287
rect 8724 36223 8740 36287
rect 8804 36223 8820 36287
rect 8884 36223 8900 36287
rect 8964 36223 8980 36287
rect 9044 36223 9060 36287
rect 9124 36223 9140 36287
rect 9204 36223 9220 36287
rect 9284 36223 9292 36287
rect 8096 36206 9292 36223
rect 8096 36142 8100 36206
rect 8164 36142 8180 36206
rect 8244 36142 8260 36206
rect 8324 36142 8340 36206
rect 8404 36142 8420 36206
rect 8484 36142 8500 36206
rect 8564 36142 8580 36206
rect 8644 36142 8660 36206
rect 8724 36142 8740 36206
rect 8804 36142 8820 36206
rect 8884 36142 8900 36206
rect 8964 36142 8980 36206
rect 9044 36142 9060 36206
rect 9124 36142 9140 36206
rect 9204 36142 9220 36206
rect 9284 36142 9292 36206
rect 8096 36124 9292 36142
rect 8096 36060 8100 36124
rect 8164 36060 8180 36124
rect 8244 36060 8260 36124
rect 8324 36060 8340 36124
rect 8404 36060 8420 36124
rect 8484 36060 8500 36124
rect 8564 36060 8580 36124
rect 8644 36060 8660 36124
rect 8724 36060 8740 36124
rect 8804 36060 8820 36124
rect 8884 36060 8900 36124
rect 8964 36060 8980 36124
rect 9044 36060 9060 36124
rect 9124 36060 9140 36124
rect 9204 36060 9220 36124
rect 9284 36060 9292 36124
rect 8096 36042 9292 36060
rect 8096 35978 8100 36042
rect 8164 35978 8180 36042
rect 8244 35978 8260 36042
rect 8324 35978 8340 36042
rect 8404 35978 8420 36042
rect 8484 35978 8500 36042
rect 8564 35978 8580 36042
rect 8644 35978 8660 36042
rect 8724 35978 8740 36042
rect 8804 35978 8820 36042
rect 8884 35978 8900 36042
rect 8964 35978 8980 36042
rect 9044 35978 9060 36042
rect 9124 35978 9140 36042
rect 9204 35978 9220 36042
rect 9284 35978 9292 36042
rect 8096 35960 9292 35978
rect 8096 35896 8100 35960
rect 8164 35896 8180 35960
rect 8244 35896 8260 35960
rect 8324 35896 8340 35960
rect 8404 35896 8420 35960
rect 8484 35896 8500 35960
rect 8564 35896 8580 35960
rect 8644 35896 8660 35960
rect 8724 35896 8740 35960
rect 8804 35896 8820 35960
rect 8884 35896 8900 35960
rect 8964 35896 8980 35960
rect 9044 35896 9060 35960
rect 9124 35896 9140 35960
rect 9204 35896 9220 35960
rect 9284 35896 9292 35960
rect 8096 35878 9292 35896
rect 8096 35814 8100 35878
rect 8164 35814 8180 35878
rect 8244 35814 8260 35878
rect 8324 35814 8340 35878
rect 8404 35814 8420 35878
rect 8484 35814 8500 35878
rect 8564 35814 8580 35878
rect 8644 35814 8660 35878
rect 8724 35814 8740 35878
rect 8804 35814 8820 35878
rect 8884 35814 8900 35878
rect 8964 35814 8980 35878
rect 9044 35814 9060 35878
rect 9124 35814 9140 35878
rect 9204 35814 9220 35878
rect 9284 35814 9292 35878
rect 8096 35796 9292 35814
rect 8096 35732 8100 35796
rect 8164 35732 8180 35796
rect 8244 35732 8260 35796
rect 8324 35732 8340 35796
rect 8404 35732 8420 35796
rect 8484 35732 8500 35796
rect 8564 35732 8580 35796
rect 8644 35732 8660 35796
rect 8724 35732 8740 35796
rect 8804 35732 8820 35796
rect 8884 35732 8900 35796
rect 8964 35732 8980 35796
rect 9044 35732 9060 35796
rect 9124 35732 9140 35796
rect 9204 35732 9220 35796
rect 9284 35732 9292 35796
rect 8096 35714 9292 35732
rect 8096 35650 8100 35714
rect 8164 35650 8180 35714
rect 8244 35650 8260 35714
rect 8324 35650 8340 35714
rect 8404 35650 8420 35714
rect 8484 35650 8500 35714
rect 8564 35650 8580 35714
rect 8644 35650 8660 35714
rect 8724 35650 8740 35714
rect 8804 35650 8820 35714
rect 8884 35650 8900 35714
rect 8964 35650 8980 35714
rect 9044 35650 9060 35714
rect 9124 35650 9140 35714
rect 9204 35650 9220 35714
rect 9284 35650 9292 35714
rect 8096 35632 9292 35650
rect 8096 35568 8100 35632
rect 8164 35568 8180 35632
rect 8244 35568 8260 35632
rect 8324 35568 8340 35632
rect 8404 35568 8420 35632
rect 8484 35568 8500 35632
rect 8564 35568 8580 35632
rect 8644 35568 8660 35632
rect 8724 35568 8740 35632
rect 8804 35568 8820 35632
rect 8884 35568 8900 35632
rect 8964 35568 8980 35632
rect 9044 35568 9060 35632
rect 9124 35568 9140 35632
rect 9204 35568 9220 35632
rect 9284 35568 9292 35632
rect 8096 35550 9292 35568
rect 8096 35486 8100 35550
rect 8164 35486 8180 35550
rect 8244 35486 8260 35550
rect 8324 35486 8340 35550
rect 8404 35486 8420 35550
rect 8484 35486 8500 35550
rect 8564 35486 8580 35550
rect 8644 35486 8660 35550
rect 8724 35486 8740 35550
rect 8804 35486 8820 35550
rect 8884 35486 8900 35550
rect 8964 35486 8980 35550
rect 9044 35486 9060 35550
rect 9124 35486 9140 35550
rect 9204 35486 9220 35550
rect 9284 35486 9292 35550
rect 8096 35468 9292 35486
rect 8096 35404 8100 35468
rect 8164 35404 8180 35468
rect 8244 35404 8260 35468
rect 8324 35404 8340 35468
rect 8404 35404 8420 35468
rect 8484 35404 8500 35468
rect 8564 35404 8580 35468
rect 8644 35404 8660 35468
rect 8724 35404 8740 35468
rect 8804 35404 8820 35468
rect 8884 35404 8900 35468
rect 8964 35404 8980 35468
rect 9044 35404 9060 35468
rect 9124 35404 9140 35468
rect 9204 35404 9220 35468
rect 9284 35404 9292 35468
rect 8096 35386 9292 35404
rect 8096 35322 8100 35386
rect 8164 35322 8180 35386
rect 8244 35322 8260 35386
rect 8324 35322 8340 35386
rect 8404 35322 8420 35386
rect 8484 35322 8500 35386
rect 8564 35322 8580 35386
rect 8644 35322 8660 35386
rect 8724 35322 8740 35386
rect 8804 35322 8820 35386
rect 8884 35322 8900 35386
rect 8964 35322 8980 35386
rect 9044 35322 9060 35386
rect 9124 35322 9140 35386
rect 9204 35322 9220 35386
rect 9284 35322 9292 35386
rect 8096 35304 9292 35322
rect 8096 35240 8100 35304
rect 8164 35240 8180 35304
rect 8244 35240 8260 35304
rect 8324 35240 8340 35304
rect 8404 35240 8420 35304
rect 8484 35240 8500 35304
rect 8564 35240 8580 35304
rect 8644 35240 8660 35304
rect 8724 35240 8740 35304
rect 8804 35240 8820 35304
rect 8884 35240 8900 35304
rect 8964 35240 8980 35304
rect 9044 35240 9060 35304
rect 9124 35240 9140 35304
rect 9204 35240 9220 35304
rect 9284 35240 9292 35304
rect 8096 35222 9292 35240
rect 8096 35158 8100 35222
rect 8164 35158 8180 35222
rect 8244 35158 8260 35222
rect 8324 35158 8340 35222
rect 8404 35158 8420 35222
rect 8484 35158 8500 35222
rect 8564 35158 8580 35222
rect 8644 35158 8660 35222
rect 8724 35158 8740 35222
rect 8804 35158 8820 35222
rect 8884 35158 8900 35222
rect 8964 35158 8980 35222
rect 9044 35158 9060 35222
rect 9124 35158 9140 35222
rect 9204 35158 9220 35222
rect 9284 35158 9292 35222
rect 8096 32613 9292 35158
rect 8096 32557 8107 32613
rect 8163 32557 8188 32613
rect 8244 32557 8269 32613
rect 8325 32557 8350 32613
rect 8406 32557 8431 32613
rect 8487 32557 8511 32613
rect 8567 32557 8591 32613
rect 8647 32557 8671 32613
rect 8727 32557 8751 32613
rect 8807 32557 8831 32613
rect 8887 32557 8911 32613
rect 8967 32557 8991 32613
rect 9047 32557 9071 32613
rect 9127 32557 9151 32613
rect 9207 32557 9231 32613
rect 9287 32557 9292 32613
rect 8096 32531 9292 32557
rect 8096 32475 8107 32531
rect 8163 32475 8188 32531
rect 8244 32475 8269 32531
rect 8325 32475 8350 32531
rect 8406 32475 8431 32531
rect 8487 32475 8511 32531
rect 8567 32475 8591 32531
rect 8647 32475 8671 32531
rect 8727 32475 8751 32531
rect 8807 32475 8831 32531
rect 8887 32475 8911 32531
rect 8967 32475 8991 32531
rect 9047 32475 9071 32531
rect 9127 32475 9151 32531
rect 9207 32475 9231 32531
rect 9287 32475 9292 32531
rect 8096 32449 9292 32475
rect 8096 32393 8107 32449
rect 8163 32393 8188 32449
rect 8244 32393 8269 32449
rect 8325 32393 8350 32449
rect 8406 32393 8431 32449
rect 8487 32393 8511 32449
rect 8567 32393 8591 32449
rect 8647 32393 8671 32449
rect 8727 32393 8751 32449
rect 8807 32393 8831 32449
rect 8887 32393 8911 32449
rect 8967 32393 8991 32449
rect 9047 32393 9071 32449
rect 9127 32393 9151 32449
rect 9207 32393 9231 32449
rect 9287 32393 9292 32449
rect 8096 32367 9292 32393
rect 8096 32311 8107 32367
rect 8163 32311 8188 32367
rect 8244 32311 8269 32367
rect 8325 32311 8350 32367
rect 8406 32311 8431 32367
rect 8487 32311 8511 32367
rect 8567 32311 8591 32367
rect 8647 32311 8671 32367
rect 8727 32311 8751 32367
rect 8807 32311 8831 32367
rect 8887 32311 8911 32367
rect 8967 32311 8991 32367
rect 9047 32311 9071 32367
rect 9127 32311 9151 32367
rect 9207 32311 9231 32367
rect 9287 32311 9292 32367
rect 8096 32285 9292 32311
rect 8096 32229 8107 32285
rect 8163 32229 8188 32285
rect 8244 32229 8269 32285
rect 8325 32229 8350 32285
rect 8406 32229 8431 32285
rect 8487 32229 8511 32285
rect 8567 32229 8591 32285
rect 8647 32229 8671 32285
rect 8727 32229 8751 32285
rect 8807 32229 8831 32285
rect 8887 32229 8911 32285
rect 8967 32229 8991 32285
rect 9047 32229 9071 32285
rect 9127 32229 9151 32285
rect 9207 32229 9231 32285
rect 9287 32229 9292 32285
rect 8096 32203 9292 32229
rect 8096 32147 8107 32203
rect 8163 32147 8188 32203
rect 8244 32147 8269 32203
rect 8325 32147 8350 32203
rect 8406 32147 8431 32203
rect 8487 32147 8511 32203
rect 8567 32147 8591 32203
rect 8647 32147 8671 32203
rect 8727 32147 8751 32203
rect 8807 32147 8831 32203
rect 8887 32147 8911 32203
rect 8967 32147 8991 32203
rect 9047 32147 9071 32203
rect 9127 32147 9151 32203
rect 9207 32147 9231 32203
rect 9287 32147 9292 32203
rect 8096 32121 9292 32147
rect 8096 32065 8107 32121
rect 8163 32065 8188 32121
rect 8244 32065 8269 32121
rect 8325 32065 8350 32121
rect 8406 32065 8431 32121
rect 8487 32065 8511 32121
rect 8567 32065 8591 32121
rect 8647 32065 8671 32121
rect 8727 32065 8751 32121
rect 8807 32065 8831 32121
rect 8887 32065 8911 32121
rect 8967 32065 8991 32121
rect 9047 32065 9071 32121
rect 9127 32065 9151 32121
rect 9207 32065 9231 32121
rect 9287 32065 9292 32121
rect 8096 32039 9292 32065
rect 8096 31983 8107 32039
rect 8163 31983 8188 32039
rect 8244 31983 8269 32039
rect 8325 31983 8350 32039
rect 8406 31983 8431 32039
rect 8487 31983 8511 32039
rect 8567 31983 8591 32039
rect 8647 31983 8671 32039
rect 8727 31983 8751 32039
rect 8807 31983 8831 32039
rect 8887 31983 8911 32039
rect 8967 31983 8991 32039
rect 9047 31983 9071 32039
rect 9127 31983 9151 32039
rect 9207 31983 9231 32039
rect 9287 31983 9292 32039
rect 8096 31957 9292 31983
rect 8096 31901 8107 31957
rect 8163 31901 8188 31957
rect 8244 31901 8269 31957
rect 8325 31901 8350 31957
rect 8406 31901 8431 31957
rect 8487 31901 8511 31957
rect 8567 31901 8591 31957
rect 8647 31901 8671 31957
rect 8727 31901 8751 31957
rect 8807 31901 8831 31957
rect 8887 31901 8911 31957
rect 8967 31901 8991 31957
rect 9047 31901 9071 31957
rect 9127 31901 9151 31957
rect 9207 31901 9231 31957
rect 9287 31901 9292 31957
rect 8096 31875 9292 31901
rect 8096 31819 8107 31875
rect 8163 31819 8188 31875
rect 8244 31819 8269 31875
rect 8325 31819 8350 31875
rect 8406 31819 8431 31875
rect 8487 31819 8511 31875
rect 8567 31819 8591 31875
rect 8647 31819 8671 31875
rect 8727 31819 8751 31875
rect 8807 31819 8831 31875
rect 8887 31819 8911 31875
rect 8967 31819 8991 31875
rect 9047 31819 9071 31875
rect 9127 31819 9151 31875
rect 9207 31819 9231 31875
rect 9287 31819 9292 31875
rect 8096 31793 9292 31819
rect 8096 31737 8107 31793
rect 8163 31737 8188 31793
rect 8244 31737 8269 31793
rect 8325 31737 8350 31793
rect 8406 31737 8431 31793
rect 8487 31737 8511 31793
rect 8567 31737 8591 31793
rect 8647 31737 8671 31793
rect 8727 31737 8751 31793
rect 8807 31737 8831 31793
rect 8887 31737 8911 31793
rect 8967 31737 8991 31793
rect 9047 31737 9071 31793
rect 9127 31737 9151 31793
rect 9207 31737 9231 31793
rect 9287 31737 9292 31793
rect 8096 31711 9292 31737
rect 8096 31655 8107 31711
rect 8163 31655 8188 31711
rect 8244 31655 8269 31711
rect 8325 31655 8350 31711
rect 8406 31655 8431 31711
rect 8487 31655 8511 31711
rect 8567 31655 8591 31711
rect 8647 31655 8671 31711
rect 8727 31655 8751 31711
rect 8807 31655 8831 31711
rect 8887 31655 8911 31711
rect 8967 31655 8991 31711
rect 9047 31655 9071 31711
rect 9127 31655 9151 31711
rect 9207 31655 9231 31711
rect 9287 31655 9292 31711
rect 8096 31629 9292 31655
rect 8096 31573 8107 31629
rect 8163 31573 8188 31629
rect 8244 31573 8269 31629
rect 8325 31573 8350 31629
rect 8406 31573 8431 31629
rect 8487 31573 8511 31629
rect 8567 31573 8591 31629
rect 8647 31573 8671 31629
rect 8727 31573 8751 31629
rect 8807 31573 8831 31629
rect 8887 31573 8911 31629
rect 8967 31573 8991 31629
rect 9047 31573 9071 31629
rect 9127 31573 9151 31629
rect 9207 31573 9231 31629
rect 9287 31573 9292 31629
rect 8096 31547 9292 31573
rect 8096 31491 8107 31547
rect 8163 31491 8188 31547
rect 8244 31491 8269 31547
rect 8325 31491 8350 31547
rect 8406 31491 8431 31547
rect 8487 31491 8511 31547
rect 8567 31491 8591 31547
rect 8647 31491 8671 31547
rect 8727 31491 8751 31547
rect 8807 31491 8831 31547
rect 8887 31491 8911 31547
rect 8967 31491 8991 31547
rect 9047 31491 9071 31547
rect 9127 31491 9151 31547
rect 9207 31491 9231 31547
rect 9287 31491 9292 31547
rect 8096 31478 9292 31491
rect 9593 39365 10789 39371
rect 9593 39301 9597 39365
rect 9661 39301 9677 39365
rect 9741 39301 9757 39365
rect 9821 39301 9837 39365
rect 9901 39301 9917 39365
rect 9981 39301 9997 39365
rect 10061 39301 10077 39365
rect 10141 39301 10157 39365
rect 10221 39301 10237 39365
rect 10301 39301 10317 39365
rect 10381 39301 10397 39365
rect 10461 39301 10477 39365
rect 10541 39301 10557 39365
rect 10621 39301 10637 39365
rect 10701 39301 10717 39365
rect 10781 39301 10789 39365
rect 9593 39284 10789 39301
rect 9593 39220 9597 39284
rect 9661 39220 9677 39284
rect 9741 39220 9757 39284
rect 9821 39220 9837 39284
rect 9901 39220 9917 39284
rect 9981 39220 9997 39284
rect 10061 39220 10077 39284
rect 10141 39220 10157 39284
rect 10221 39220 10237 39284
rect 10301 39220 10317 39284
rect 10381 39220 10397 39284
rect 10461 39220 10477 39284
rect 10541 39220 10557 39284
rect 10621 39220 10637 39284
rect 10701 39220 10717 39284
rect 10781 39220 10789 39284
rect 9593 39203 10789 39220
rect 9593 39139 9597 39203
rect 9661 39139 9677 39203
rect 9741 39139 9757 39203
rect 9821 39139 9837 39203
rect 9901 39139 9917 39203
rect 9981 39139 9997 39203
rect 10061 39139 10077 39203
rect 10141 39139 10157 39203
rect 10221 39139 10237 39203
rect 10301 39139 10317 39203
rect 10381 39139 10397 39203
rect 10461 39139 10477 39203
rect 10541 39139 10557 39203
rect 10621 39139 10637 39203
rect 10701 39139 10717 39203
rect 10781 39139 10789 39203
rect 9593 39122 10789 39139
rect 9593 39058 9597 39122
rect 9661 39058 9677 39122
rect 9741 39058 9757 39122
rect 9821 39058 9837 39122
rect 9901 39058 9917 39122
rect 9981 39058 9997 39122
rect 10061 39058 10077 39122
rect 10141 39058 10157 39122
rect 10221 39058 10237 39122
rect 10301 39058 10317 39122
rect 10381 39058 10397 39122
rect 10461 39058 10477 39122
rect 10541 39058 10557 39122
rect 10621 39058 10637 39122
rect 10701 39058 10717 39122
rect 10781 39058 10789 39122
rect 9593 39041 10789 39058
rect 9593 38977 9597 39041
rect 9661 38977 9677 39041
rect 9741 38977 9757 39041
rect 9821 38977 9837 39041
rect 9901 38977 9917 39041
rect 9981 38977 9997 39041
rect 10061 38977 10077 39041
rect 10141 38977 10157 39041
rect 10221 38977 10237 39041
rect 10301 38977 10317 39041
rect 10381 38977 10397 39041
rect 10461 38977 10477 39041
rect 10541 38977 10557 39041
rect 10621 38977 10637 39041
rect 10701 38977 10717 39041
rect 10781 38977 10789 39041
rect 9593 38960 10789 38977
rect 9593 38896 9597 38960
rect 9661 38896 9677 38960
rect 9741 38896 9757 38960
rect 9821 38896 9837 38960
rect 9901 38896 9917 38960
rect 9981 38896 9997 38960
rect 10061 38896 10077 38960
rect 10141 38896 10157 38960
rect 10221 38896 10237 38960
rect 10301 38896 10317 38960
rect 10381 38896 10397 38960
rect 10461 38896 10477 38960
rect 10541 38896 10557 38960
rect 10621 38896 10637 38960
rect 10701 38896 10717 38960
rect 10781 38896 10789 38960
rect 9593 38879 10789 38896
rect 9593 38815 9597 38879
rect 9661 38815 9677 38879
rect 9741 38815 9757 38879
rect 9821 38815 9837 38879
rect 9901 38815 9917 38879
rect 9981 38815 9997 38879
rect 10061 38815 10077 38879
rect 10141 38815 10157 38879
rect 10221 38815 10237 38879
rect 10301 38815 10317 38879
rect 10381 38815 10397 38879
rect 10461 38815 10477 38879
rect 10541 38815 10557 38879
rect 10621 38815 10637 38879
rect 10701 38815 10717 38879
rect 10781 38815 10789 38879
rect 9593 38798 10789 38815
rect 9593 38734 9597 38798
rect 9661 38734 9677 38798
rect 9741 38734 9757 38798
rect 9821 38734 9837 38798
rect 9901 38734 9917 38798
rect 9981 38734 9997 38798
rect 10061 38734 10077 38798
rect 10141 38734 10157 38798
rect 10221 38734 10237 38798
rect 10301 38734 10317 38798
rect 10381 38734 10397 38798
rect 10461 38734 10477 38798
rect 10541 38734 10557 38798
rect 10621 38734 10637 38798
rect 10701 38734 10717 38798
rect 10781 38734 10789 38798
rect 9593 38717 10789 38734
rect 9593 38653 9597 38717
rect 9661 38653 9677 38717
rect 9741 38653 9757 38717
rect 9821 38653 9837 38717
rect 9901 38653 9917 38717
rect 9981 38653 9997 38717
rect 10061 38653 10077 38717
rect 10141 38653 10157 38717
rect 10221 38653 10237 38717
rect 10301 38653 10317 38717
rect 10381 38653 10397 38717
rect 10461 38653 10477 38717
rect 10541 38653 10557 38717
rect 10621 38653 10637 38717
rect 10701 38653 10717 38717
rect 10781 38653 10789 38717
rect 9593 38636 10789 38653
rect 9593 38572 9597 38636
rect 9661 38572 9677 38636
rect 9741 38572 9757 38636
rect 9821 38572 9837 38636
rect 9901 38572 9917 38636
rect 9981 38572 9997 38636
rect 10061 38572 10077 38636
rect 10141 38572 10157 38636
rect 10221 38572 10237 38636
rect 10301 38572 10317 38636
rect 10381 38572 10397 38636
rect 10461 38572 10477 38636
rect 10541 38572 10557 38636
rect 10621 38572 10637 38636
rect 10701 38572 10717 38636
rect 10781 38572 10789 38636
rect 9593 38555 10789 38572
rect 9593 38491 9597 38555
rect 9661 38491 9677 38555
rect 9741 38491 9757 38555
rect 9821 38491 9837 38555
rect 9901 38491 9917 38555
rect 9981 38491 9997 38555
rect 10061 38491 10077 38555
rect 10141 38491 10157 38555
rect 10221 38491 10237 38555
rect 10301 38491 10317 38555
rect 10381 38491 10397 38555
rect 10461 38491 10477 38555
rect 10541 38491 10557 38555
rect 10621 38491 10637 38555
rect 10701 38491 10717 38555
rect 10781 38491 10789 38555
rect 9593 38474 10789 38491
rect 9593 38410 9597 38474
rect 9661 38410 9677 38474
rect 9741 38410 9757 38474
rect 9821 38410 9837 38474
rect 9901 38410 9917 38474
rect 9981 38410 9997 38474
rect 10061 38410 10077 38474
rect 10141 38410 10157 38474
rect 10221 38410 10237 38474
rect 10301 38410 10317 38474
rect 10381 38410 10397 38474
rect 10461 38410 10477 38474
rect 10541 38410 10557 38474
rect 10621 38410 10637 38474
rect 10701 38410 10717 38474
rect 10781 38410 10789 38474
rect 9593 38393 10789 38410
rect 9593 38329 9597 38393
rect 9661 38329 9677 38393
rect 9741 38329 9757 38393
rect 9821 38329 9837 38393
rect 9901 38329 9917 38393
rect 9981 38329 9997 38393
rect 10061 38329 10077 38393
rect 10141 38329 10157 38393
rect 10221 38329 10237 38393
rect 10301 38329 10317 38393
rect 10381 38329 10397 38393
rect 10461 38329 10477 38393
rect 10541 38329 10557 38393
rect 10621 38329 10637 38393
rect 10701 38329 10717 38393
rect 10781 38329 10789 38393
rect 9593 38312 10789 38329
rect 9593 38248 9597 38312
rect 9661 38248 9677 38312
rect 9741 38248 9757 38312
rect 9821 38248 9837 38312
rect 9901 38248 9917 38312
rect 9981 38248 9997 38312
rect 10061 38248 10077 38312
rect 10141 38248 10157 38312
rect 10221 38248 10237 38312
rect 10301 38248 10317 38312
rect 10381 38248 10397 38312
rect 10461 38248 10477 38312
rect 10541 38248 10557 38312
rect 10621 38248 10637 38312
rect 10701 38248 10717 38312
rect 10781 38248 10789 38312
rect 9593 38231 10789 38248
rect 9593 38167 9597 38231
rect 9661 38167 9677 38231
rect 9741 38167 9757 38231
rect 9821 38167 9837 38231
rect 9901 38167 9917 38231
rect 9981 38167 9997 38231
rect 10061 38167 10077 38231
rect 10141 38167 10157 38231
rect 10221 38167 10237 38231
rect 10301 38167 10317 38231
rect 10381 38167 10397 38231
rect 10461 38167 10477 38231
rect 10541 38167 10557 38231
rect 10621 38167 10637 38231
rect 10701 38167 10717 38231
rect 10781 38167 10789 38231
rect 9593 38150 10789 38167
rect 9593 38086 9597 38150
rect 9661 38086 9677 38150
rect 9741 38086 9757 38150
rect 9821 38086 9837 38150
rect 9901 38086 9917 38150
rect 9981 38086 9997 38150
rect 10061 38086 10077 38150
rect 10141 38086 10157 38150
rect 10221 38086 10237 38150
rect 10301 38086 10317 38150
rect 10381 38086 10397 38150
rect 10461 38086 10477 38150
rect 10541 38086 10557 38150
rect 10621 38086 10637 38150
rect 10701 38086 10717 38150
rect 10781 38086 10789 38150
rect 9593 38069 10789 38086
rect 9593 38005 9597 38069
rect 9661 38005 9677 38069
rect 9741 38005 9757 38069
rect 9821 38005 9837 38069
rect 9901 38005 9917 38069
rect 9981 38005 9997 38069
rect 10061 38005 10077 38069
rect 10141 38005 10157 38069
rect 10221 38005 10237 38069
rect 10301 38005 10317 38069
rect 10381 38005 10397 38069
rect 10461 38005 10477 38069
rect 10541 38005 10557 38069
rect 10621 38005 10637 38069
rect 10701 38005 10717 38069
rect 10781 38005 10789 38069
rect 9593 37988 10789 38005
rect 9593 37924 9597 37988
rect 9661 37924 9677 37988
rect 9741 37924 9757 37988
rect 9821 37924 9837 37988
rect 9901 37924 9917 37988
rect 9981 37924 9997 37988
rect 10061 37924 10077 37988
rect 10141 37924 10157 37988
rect 10221 37924 10237 37988
rect 10301 37924 10317 37988
rect 10381 37924 10397 37988
rect 10461 37924 10477 37988
rect 10541 37924 10557 37988
rect 10621 37924 10637 37988
rect 10701 37924 10717 37988
rect 10781 37924 10789 37988
rect 9593 37907 10789 37924
rect 9593 37843 9597 37907
rect 9661 37843 9677 37907
rect 9741 37843 9757 37907
rect 9821 37843 9837 37907
rect 9901 37843 9917 37907
rect 9981 37843 9997 37907
rect 10061 37843 10077 37907
rect 10141 37843 10157 37907
rect 10221 37843 10237 37907
rect 10301 37843 10317 37907
rect 10381 37843 10397 37907
rect 10461 37843 10477 37907
rect 10541 37843 10557 37907
rect 10621 37843 10637 37907
rect 10701 37843 10717 37907
rect 10781 37843 10789 37907
rect 9593 37826 10789 37843
rect 9593 37762 9597 37826
rect 9661 37762 9677 37826
rect 9741 37762 9757 37826
rect 9821 37762 9837 37826
rect 9901 37762 9917 37826
rect 9981 37762 9997 37826
rect 10061 37762 10077 37826
rect 10141 37762 10157 37826
rect 10221 37762 10237 37826
rect 10301 37762 10317 37826
rect 10381 37762 10397 37826
rect 10461 37762 10477 37826
rect 10541 37762 10557 37826
rect 10621 37762 10637 37826
rect 10701 37762 10717 37826
rect 10781 37762 10789 37826
rect 9593 37745 10789 37762
rect 9593 37681 9597 37745
rect 9661 37681 9677 37745
rect 9741 37681 9757 37745
rect 9821 37681 9837 37745
rect 9901 37681 9917 37745
rect 9981 37681 9997 37745
rect 10061 37681 10077 37745
rect 10141 37681 10157 37745
rect 10221 37681 10237 37745
rect 10301 37681 10317 37745
rect 10381 37681 10397 37745
rect 10461 37681 10477 37745
rect 10541 37681 10557 37745
rect 10621 37681 10637 37745
rect 10701 37681 10717 37745
rect 10781 37681 10789 37745
rect 9593 37664 10789 37681
rect 9593 37600 9597 37664
rect 9661 37600 9677 37664
rect 9741 37600 9757 37664
rect 9821 37600 9837 37664
rect 9901 37600 9917 37664
rect 9981 37600 9997 37664
rect 10061 37600 10077 37664
rect 10141 37600 10157 37664
rect 10221 37600 10237 37664
rect 10301 37600 10317 37664
rect 10381 37600 10397 37664
rect 10461 37600 10477 37664
rect 10541 37600 10557 37664
rect 10621 37600 10637 37664
rect 10701 37600 10717 37664
rect 10781 37600 10789 37664
rect 9593 37583 10789 37600
rect 9593 37519 9597 37583
rect 9661 37519 9677 37583
rect 9741 37519 9757 37583
rect 9821 37519 9837 37583
rect 9901 37519 9917 37583
rect 9981 37519 9997 37583
rect 10061 37519 10077 37583
rect 10141 37519 10157 37583
rect 10221 37519 10237 37583
rect 10301 37519 10317 37583
rect 10381 37519 10397 37583
rect 10461 37519 10477 37583
rect 10541 37519 10557 37583
rect 10621 37519 10637 37583
rect 10701 37519 10717 37583
rect 10781 37519 10789 37583
rect 9593 37502 10789 37519
rect 9593 37438 9597 37502
rect 9661 37438 9677 37502
rect 9741 37438 9757 37502
rect 9821 37438 9837 37502
rect 9901 37438 9917 37502
rect 9981 37438 9997 37502
rect 10061 37438 10077 37502
rect 10141 37438 10157 37502
rect 10221 37438 10237 37502
rect 10301 37438 10317 37502
rect 10381 37438 10397 37502
rect 10461 37438 10477 37502
rect 10541 37438 10557 37502
rect 10621 37438 10637 37502
rect 10701 37438 10717 37502
rect 10781 37438 10789 37502
rect 9593 37421 10789 37438
rect 9593 37357 9597 37421
rect 9661 37357 9677 37421
rect 9741 37357 9757 37421
rect 9821 37357 9837 37421
rect 9901 37357 9917 37421
rect 9981 37357 9997 37421
rect 10061 37357 10077 37421
rect 10141 37357 10157 37421
rect 10221 37357 10237 37421
rect 10301 37357 10317 37421
rect 10381 37357 10397 37421
rect 10461 37357 10477 37421
rect 10541 37357 10557 37421
rect 10621 37357 10637 37421
rect 10701 37357 10717 37421
rect 10781 37357 10789 37421
rect 9593 37340 10789 37357
rect 9593 37276 9597 37340
rect 9661 37276 9677 37340
rect 9741 37276 9757 37340
rect 9821 37276 9837 37340
rect 9901 37276 9917 37340
rect 9981 37276 9997 37340
rect 10061 37276 10077 37340
rect 10141 37276 10157 37340
rect 10221 37276 10237 37340
rect 10301 37276 10317 37340
rect 10381 37276 10397 37340
rect 10461 37276 10477 37340
rect 10541 37276 10557 37340
rect 10621 37276 10637 37340
rect 10701 37276 10717 37340
rect 10781 37276 10789 37340
rect 9593 37259 10789 37276
rect 9593 37195 9597 37259
rect 9661 37195 9677 37259
rect 9741 37195 9757 37259
rect 9821 37195 9837 37259
rect 9901 37195 9917 37259
rect 9981 37195 9997 37259
rect 10061 37195 10077 37259
rect 10141 37195 10157 37259
rect 10221 37195 10237 37259
rect 10301 37195 10317 37259
rect 10381 37195 10397 37259
rect 10461 37195 10477 37259
rect 10541 37195 10557 37259
rect 10621 37195 10637 37259
rect 10701 37195 10717 37259
rect 10781 37195 10789 37259
rect 9593 37178 10789 37195
rect 9593 37114 9597 37178
rect 9661 37114 9677 37178
rect 9741 37114 9757 37178
rect 9821 37114 9837 37178
rect 9901 37114 9917 37178
rect 9981 37114 9997 37178
rect 10061 37114 10077 37178
rect 10141 37114 10157 37178
rect 10221 37114 10237 37178
rect 10301 37114 10317 37178
rect 10381 37114 10397 37178
rect 10461 37114 10477 37178
rect 10541 37114 10557 37178
rect 10621 37114 10637 37178
rect 10701 37114 10717 37178
rect 10781 37114 10789 37178
rect 9593 37097 10789 37114
rect 9593 37033 9597 37097
rect 9661 37033 9677 37097
rect 9741 37033 9757 37097
rect 9821 37033 9837 37097
rect 9901 37033 9917 37097
rect 9981 37033 9997 37097
rect 10061 37033 10077 37097
rect 10141 37033 10157 37097
rect 10221 37033 10237 37097
rect 10301 37033 10317 37097
rect 10381 37033 10397 37097
rect 10461 37033 10477 37097
rect 10541 37033 10557 37097
rect 10621 37033 10637 37097
rect 10701 37033 10717 37097
rect 10781 37033 10789 37097
rect 9593 37016 10789 37033
rect 9593 36952 9597 37016
rect 9661 36952 9677 37016
rect 9741 36952 9757 37016
rect 9821 36952 9837 37016
rect 9901 36952 9917 37016
rect 9981 36952 9997 37016
rect 10061 36952 10077 37016
rect 10141 36952 10157 37016
rect 10221 36952 10237 37016
rect 10301 36952 10317 37016
rect 10381 36952 10397 37016
rect 10461 36952 10477 37016
rect 10541 36952 10557 37016
rect 10621 36952 10637 37016
rect 10701 36952 10717 37016
rect 10781 36952 10789 37016
rect 9593 36935 10789 36952
rect 9593 36871 9597 36935
rect 9661 36871 9677 36935
rect 9741 36871 9757 36935
rect 9821 36871 9837 36935
rect 9901 36871 9917 36935
rect 9981 36871 9997 36935
rect 10061 36871 10077 36935
rect 10141 36871 10157 36935
rect 10221 36871 10237 36935
rect 10301 36871 10317 36935
rect 10381 36871 10397 36935
rect 10461 36871 10477 36935
rect 10541 36871 10557 36935
rect 10621 36871 10637 36935
rect 10701 36871 10717 36935
rect 10781 36871 10789 36935
rect 9593 36854 10789 36871
rect 9593 36790 9597 36854
rect 9661 36790 9677 36854
rect 9741 36790 9757 36854
rect 9821 36790 9837 36854
rect 9901 36790 9917 36854
rect 9981 36790 9997 36854
rect 10061 36790 10077 36854
rect 10141 36790 10157 36854
rect 10221 36790 10237 36854
rect 10301 36790 10317 36854
rect 10381 36790 10397 36854
rect 10461 36790 10477 36854
rect 10541 36790 10557 36854
rect 10621 36790 10637 36854
rect 10701 36790 10717 36854
rect 10781 36790 10789 36854
rect 9593 36773 10789 36790
rect 9593 36709 9597 36773
rect 9661 36709 9677 36773
rect 9741 36709 9757 36773
rect 9821 36709 9837 36773
rect 9901 36709 9917 36773
rect 9981 36709 9997 36773
rect 10061 36709 10077 36773
rect 10141 36709 10157 36773
rect 10221 36709 10237 36773
rect 10301 36709 10317 36773
rect 10381 36709 10397 36773
rect 10461 36709 10477 36773
rect 10541 36709 10557 36773
rect 10621 36709 10637 36773
rect 10701 36709 10717 36773
rect 10781 36709 10789 36773
rect 9593 36692 10789 36709
rect 9593 36628 9597 36692
rect 9661 36628 9677 36692
rect 9741 36628 9757 36692
rect 9821 36628 9837 36692
rect 9901 36628 9917 36692
rect 9981 36628 9997 36692
rect 10061 36628 10077 36692
rect 10141 36628 10157 36692
rect 10221 36628 10237 36692
rect 10301 36628 10317 36692
rect 10381 36628 10397 36692
rect 10461 36628 10477 36692
rect 10541 36628 10557 36692
rect 10621 36628 10637 36692
rect 10701 36628 10717 36692
rect 10781 36628 10789 36692
rect 9593 36611 10789 36628
rect 9593 36547 9597 36611
rect 9661 36547 9677 36611
rect 9741 36547 9757 36611
rect 9821 36547 9837 36611
rect 9901 36547 9917 36611
rect 9981 36547 9997 36611
rect 10061 36547 10077 36611
rect 10141 36547 10157 36611
rect 10221 36547 10237 36611
rect 10301 36547 10317 36611
rect 10381 36547 10397 36611
rect 10461 36547 10477 36611
rect 10541 36547 10557 36611
rect 10621 36547 10637 36611
rect 10701 36547 10717 36611
rect 10781 36547 10789 36611
rect 9593 36530 10789 36547
rect 9593 36466 9597 36530
rect 9661 36466 9677 36530
rect 9741 36466 9757 36530
rect 9821 36466 9837 36530
rect 9901 36466 9917 36530
rect 9981 36466 9997 36530
rect 10061 36466 10077 36530
rect 10141 36466 10157 36530
rect 10221 36466 10237 36530
rect 10301 36466 10317 36530
rect 10381 36466 10397 36530
rect 10461 36466 10477 36530
rect 10541 36466 10557 36530
rect 10621 36466 10637 36530
rect 10701 36466 10717 36530
rect 10781 36466 10789 36530
rect 9593 36449 10789 36466
rect 9593 36385 9597 36449
rect 9661 36385 9677 36449
rect 9741 36385 9757 36449
rect 9821 36385 9837 36449
rect 9901 36385 9917 36449
rect 9981 36385 9997 36449
rect 10061 36385 10077 36449
rect 10141 36385 10157 36449
rect 10221 36385 10237 36449
rect 10301 36385 10317 36449
rect 10381 36385 10397 36449
rect 10461 36385 10477 36449
rect 10541 36385 10557 36449
rect 10621 36385 10637 36449
rect 10701 36385 10717 36449
rect 10781 36385 10789 36449
rect 9593 36368 10789 36385
rect 9593 36304 9597 36368
rect 9661 36304 9677 36368
rect 9741 36304 9757 36368
rect 9821 36304 9837 36368
rect 9901 36304 9917 36368
rect 9981 36304 9997 36368
rect 10061 36304 10077 36368
rect 10141 36304 10157 36368
rect 10221 36304 10237 36368
rect 10301 36304 10317 36368
rect 10381 36304 10397 36368
rect 10461 36304 10477 36368
rect 10541 36304 10557 36368
rect 10621 36304 10637 36368
rect 10701 36304 10717 36368
rect 10781 36304 10789 36368
rect 9593 36287 10789 36304
rect 9593 36223 9597 36287
rect 9661 36223 9677 36287
rect 9741 36223 9757 36287
rect 9821 36223 9837 36287
rect 9901 36223 9917 36287
rect 9981 36223 9997 36287
rect 10061 36223 10077 36287
rect 10141 36223 10157 36287
rect 10221 36223 10237 36287
rect 10301 36223 10317 36287
rect 10381 36223 10397 36287
rect 10461 36223 10477 36287
rect 10541 36223 10557 36287
rect 10621 36223 10637 36287
rect 10701 36223 10717 36287
rect 10781 36223 10789 36287
rect 9593 36206 10789 36223
rect 9593 36142 9597 36206
rect 9661 36142 9677 36206
rect 9741 36142 9757 36206
rect 9821 36142 9837 36206
rect 9901 36142 9917 36206
rect 9981 36142 9997 36206
rect 10061 36142 10077 36206
rect 10141 36142 10157 36206
rect 10221 36142 10237 36206
rect 10301 36142 10317 36206
rect 10381 36142 10397 36206
rect 10461 36142 10477 36206
rect 10541 36142 10557 36206
rect 10621 36142 10637 36206
rect 10701 36142 10717 36206
rect 10781 36142 10789 36206
rect 9593 36124 10789 36142
rect 9593 36060 9597 36124
rect 9661 36060 9677 36124
rect 9741 36060 9757 36124
rect 9821 36060 9837 36124
rect 9901 36060 9917 36124
rect 9981 36060 9997 36124
rect 10061 36060 10077 36124
rect 10141 36060 10157 36124
rect 10221 36060 10237 36124
rect 10301 36060 10317 36124
rect 10381 36060 10397 36124
rect 10461 36060 10477 36124
rect 10541 36060 10557 36124
rect 10621 36060 10637 36124
rect 10701 36060 10717 36124
rect 10781 36060 10789 36124
rect 9593 36042 10789 36060
rect 9593 35978 9597 36042
rect 9661 35978 9677 36042
rect 9741 35978 9757 36042
rect 9821 35978 9837 36042
rect 9901 35978 9917 36042
rect 9981 35978 9997 36042
rect 10061 35978 10077 36042
rect 10141 35978 10157 36042
rect 10221 35978 10237 36042
rect 10301 35978 10317 36042
rect 10381 35978 10397 36042
rect 10461 35978 10477 36042
rect 10541 35978 10557 36042
rect 10621 35978 10637 36042
rect 10701 35978 10717 36042
rect 10781 35978 10789 36042
rect 9593 35960 10789 35978
rect 9593 35896 9597 35960
rect 9661 35896 9677 35960
rect 9741 35896 9757 35960
rect 9821 35896 9837 35960
rect 9901 35896 9917 35960
rect 9981 35896 9997 35960
rect 10061 35896 10077 35960
rect 10141 35896 10157 35960
rect 10221 35896 10237 35960
rect 10301 35896 10317 35960
rect 10381 35896 10397 35960
rect 10461 35896 10477 35960
rect 10541 35896 10557 35960
rect 10621 35896 10637 35960
rect 10701 35896 10717 35960
rect 10781 35896 10789 35960
rect 9593 35878 10789 35896
rect 9593 35814 9597 35878
rect 9661 35814 9677 35878
rect 9741 35814 9757 35878
rect 9821 35814 9837 35878
rect 9901 35814 9917 35878
rect 9981 35814 9997 35878
rect 10061 35814 10077 35878
rect 10141 35814 10157 35878
rect 10221 35814 10237 35878
rect 10301 35814 10317 35878
rect 10381 35814 10397 35878
rect 10461 35814 10477 35878
rect 10541 35814 10557 35878
rect 10621 35814 10637 35878
rect 10701 35814 10717 35878
rect 10781 35814 10789 35878
rect 9593 35796 10789 35814
rect 9593 35732 9597 35796
rect 9661 35732 9677 35796
rect 9741 35732 9757 35796
rect 9821 35732 9837 35796
rect 9901 35732 9917 35796
rect 9981 35732 9997 35796
rect 10061 35732 10077 35796
rect 10141 35732 10157 35796
rect 10221 35732 10237 35796
rect 10301 35732 10317 35796
rect 10381 35732 10397 35796
rect 10461 35732 10477 35796
rect 10541 35732 10557 35796
rect 10621 35732 10637 35796
rect 10701 35732 10717 35796
rect 10781 35732 10789 35796
rect 9593 35714 10789 35732
rect 9593 35650 9597 35714
rect 9661 35650 9677 35714
rect 9741 35650 9757 35714
rect 9821 35650 9837 35714
rect 9901 35650 9917 35714
rect 9981 35650 9997 35714
rect 10061 35650 10077 35714
rect 10141 35650 10157 35714
rect 10221 35650 10237 35714
rect 10301 35650 10317 35714
rect 10381 35650 10397 35714
rect 10461 35650 10477 35714
rect 10541 35650 10557 35714
rect 10621 35650 10637 35714
rect 10701 35650 10717 35714
rect 10781 35650 10789 35714
rect 9593 35632 10789 35650
rect 9593 35568 9597 35632
rect 9661 35568 9677 35632
rect 9741 35568 9757 35632
rect 9821 35568 9837 35632
rect 9901 35568 9917 35632
rect 9981 35568 9997 35632
rect 10061 35568 10077 35632
rect 10141 35568 10157 35632
rect 10221 35568 10237 35632
rect 10301 35568 10317 35632
rect 10381 35568 10397 35632
rect 10461 35568 10477 35632
rect 10541 35568 10557 35632
rect 10621 35568 10637 35632
rect 10701 35568 10717 35632
rect 10781 35568 10789 35632
rect 9593 35550 10789 35568
rect 9593 35486 9597 35550
rect 9661 35486 9677 35550
rect 9741 35486 9757 35550
rect 9821 35486 9837 35550
rect 9901 35486 9917 35550
rect 9981 35486 9997 35550
rect 10061 35486 10077 35550
rect 10141 35486 10157 35550
rect 10221 35486 10237 35550
rect 10301 35486 10317 35550
rect 10381 35486 10397 35550
rect 10461 35486 10477 35550
rect 10541 35486 10557 35550
rect 10621 35486 10637 35550
rect 10701 35486 10717 35550
rect 10781 35486 10789 35550
rect 9593 35468 10789 35486
rect 9593 35404 9597 35468
rect 9661 35404 9677 35468
rect 9741 35404 9757 35468
rect 9821 35404 9837 35468
rect 9901 35404 9917 35468
rect 9981 35404 9997 35468
rect 10061 35404 10077 35468
rect 10141 35404 10157 35468
rect 10221 35404 10237 35468
rect 10301 35404 10317 35468
rect 10381 35404 10397 35468
rect 10461 35404 10477 35468
rect 10541 35404 10557 35468
rect 10621 35404 10637 35468
rect 10701 35404 10717 35468
rect 10781 35404 10789 35468
rect 9593 35386 10789 35404
rect 9593 35322 9597 35386
rect 9661 35322 9677 35386
rect 9741 35322 9757 35386
rect 9821 35322 9837 35386
rect 9901 35322 9917 35386
rect 9981 35322 9997 35386
rect 10061 35322 10077 35386
rect 10141 35322 10157 35386
rect 10221 35322 10237 35386
rect 10301 35322 10317 35386
rect 10381 35322 10397 35386
rect 10461 35322 10477 35386
rect 10541 35322 10557 35386
rect 10621 35322 10637 35386
rect 10701 35322 10717 35386
rect 10781 35322 10789 35386
rect 9593 35304 10789 35322
rect 9593 35240 9597 35304
rect 9661 35240 9677 35304
rect 9741 35240 9757 35304
rect 9821 35240 9837 35304
rect 9901 35240 9917 35304
rect 9981 35240 9997 35304
rect 10061 35240 10077 35304
rect 10141 35240 10157 35304
rect 10221 35240 10237 35304
rect 10301 35240 10317 35304
rect 10381 35240 10397 35304
rect 10461 35240 10477 35304
rect 10541 35240 10557 35304
rect 10621 35240 10637 35304
rect 10701 35240 10717 35304
rect 10781 35240 10789 35304
rect 9593 35222 10789 35240
rect 9593 35158 9597 35222
rect 9661 35158 9677 35222
rect 9741 35158 9757 35222
rect 9821 35158 9837 35222
rect 9901 35158 9917 35222
rect 9981 35158 9997 35222
rect 10061 35158 10077 35222
rect 10141 35158 10157 35222
rect 10221 35158 10237 35222
rect 10301 35158 10317 35222
rect 10381 35158 10397 35222
rect 10461 35158 10477 35222
rect 10541 35158 10557 35222
rect 10621 35158 10637 35222
rect 10701 35158 10717 35222
rect 10781 35158 10789 35222
rect 9593 32613 10789 35158
rect 9593 32557 9604 32613
rect 9660 32557 9685 32613
rect 9741 32557 9766 32613
rect 9822 32557 9847 32613
rect 9903 32557 9928 32613
rect 9984 32557 10008 32613
rect 10064 32557 10088 32613
rect 10144 32557 10168 32613
rect 10224 32557 10248 32613
rect 10304 32557 10328 32613
rect 10384 32557 10408 32613
rect 10464 32557 10488 32613
rect 10544 32557 10568 32613
rect 10624 32557 10648 32613
rect 10704 32557 10728 32613
rect 10784 32557 10789 32613
rect 9593 32531 10789 32557
rect 9593 32475 9604 32531
rect 9660 32475 9685 32531
rect 9741 32475 9766 32531
rect 9822 32475 9847 32531
rect 9903 32475 9928 32531
rect 9984 32475 10008 32531
rect 10064 32475 10088 32531
rect 10144 32475 10168 32531
rect 10224 32475 10248 32531
rect 10304 32475 10328 32531
rect 10384 32475 10408 32531
rect 10464 32475 10488 32531
rect 10544 32475 10568 32531
rect 10624 32475 10648 32531
rect 10704 32475 10728 32531
rect 10784 32475 10789 32531
rect 9593 32449 10789 32475
rect 9593 32393 9604 32449
rect 9660 32393 9685 32449
rect 9741 32393 9766 32449
rect 9822 32393 9847 32449
rect 9903 32393 9928 32449
rect 9984 32393 10008 32449
rect 10064 32393 10088 32449
rect 10144 32393 10168 32449
rect 10224 32393 10248 32449
rect 10304 32393 10328 32449
rect 10384 32393 10408 32449
rect 10464 32393 10488 32449
rect 10544 32393 10568 32449
rect 10624 32393 10648 32449
rect 10704 32393 10728 32449
rect 10784 32393 10789 32449
rect 9593 32367 10789 32393
rect 9593 32311 9604 32367
rect 9660 32311 9685 32367
rect 9741 32311 9766 32367
rect 9822 32311 9847 32367
rect 9903 32311 9928 32367
rect 9984 32311 10008 32367
rect 10064 32311 10088 32367
rect 10144 32311 10168 32367
rect 10224 32311 10248 32367
rect 10304 32311 10328 32367
rect 10384 32311 10408 32367
rect 10464 32311 10488 32367
rect 10544 32311 10568 32367
rect 10624 32311 10648 32367
rect 10704 32311 10728 32367
rect 10784 32311 10789 32367
rect 9593 32285 10789 32311
rect 9593 32229 9604 32285
rect 9660 32229 9685 32285
rect 9741 32229 9766 32285
rect 9822 32229 9847 32285
rect 9903 32229 9928 32285
rect 9984 32229 10008 32285
rect 10064 32229 10088 32285
rect 10144 32229 10168 32285
rect 10224 32229 10248 32285
rect 10304 32229 10328 32285
rect 10384 32229 10408 32285
rect 10464 32229 10488 32285
rect 10544 32229 10568 32285
rect 10624 32229 10648 32285
rect 10704 32229 10728 32285
rect 10784 32229 10789 32285
rect 9593 32203 10789 32229
rect 9593 32147 9604 32203
rect 9660 32147 9685 32203
rect 9741 32147 9766 32203
rect 9822 32147 9847 32203
rect 9903 32147 9928 32203
rect 9984 32147 10008 32203
rect 10064 32147 10088 32203
rect 10144 32147 10168 32203
rect 10224 32147 10248 32203
rect 10304 32147 10328 32203
rect 10384 32147 10408 32203
rect 10464 32147 10488 32203
rect 10544 32147 10568 32203
rect 10624 32147 10648 32203
rect 10704 32147 10728 32203
rect 10784 32147 10789 32203
rect 9593 32121 10789 32147
rect 9593 32065 9604 32121
rect 9660 32065 9685 32121
rect 9741 32065 9766 32121
rect 9822 32065 9847 32121
rect 9903 32065 9928 32121
rect 9984 32065 10008 32121
rect 10064 32065 10088 32121
rect 10144 32065 10168 32121
rect 10224 32065 10248 32121
rect 10304 32065 10328 32121
rect 10384 32065 10408 32121
rect 10464 32065 10488 32121
rect 10544 32065 10568 32121
rect 10624 32065 10648 32121
rect 10704 32065 10728 32121
rect 10784 32065 10789 32121
rect 9593 32039 10789 32065
rect 9593 31983 9604 32039
rect 9660 31983 9685 32039
rect 9741 31983 9766 32039
rect 9822 31983 9847 32039
rect 9903 31983 9928 32039
rect 9984 31983 10008 32039
rect 10064 31983 10088 32039
rect 10144 31983 10168 32039
rect 10224 31983 10248 32039
rect 10304 31983 10328 32039
rect 10384 31983 10408 32039
rect 10464 31983 10488 32039
rect 10544 31983 10568 32039
rect 10624 31983 10648 32039
rect 10704 31983 10728 32039
rect 10784 31983 10789 32039
rect 9593 31957 10789 31983
rect 9593 31901 9604 31957
rect 9660 31901 9685 31957
rect 9741 31901 9766 31957
rect 9822 31901 9847 31957
rect 9903 31901 9928 31957
rect 9984 31901 10008 31957
rect 10064 31901 10088 31957
rect 10144 31901 10168 31957
rect 10224 31901 10248 31957
rect 10304 31901 10328 31957
rect 10384 31901 10408 31957
rect 10464 31901 10488 31957
rect 10544 31901 10568 31957
rect 10624 31901 10648 31957
rect 10704 31901 10728 31957
rect 10784 31901 10789 31957
rect 9593 31875 10789 31901
rect 9593 31819 9604 31875
rect 9660 31819 9685 31875
rect 9741 31819 9766 31875
rect 9822 31819 9847 31875
rect 9903 31819 9928 31875
rect 9984 31819 10008 31875
rect 10064 31819 10088 31875
rect 10144 31819 10168 31875
rect 10224 31819 10248 31875
rect 10304 31819 10328 31875
rect 10384 31819 10408 31875
rect 10464 31819 10488 31875
rect 10544 31819 10568 31875
rect 10624 31819 10648 31875
rect 10704 31819 10728 31875
rect 10784 31819 10789 31875
rect 9593 31793 10789 31819
rect 9593 31737 9604 31793
rect 9660 31737 9685 31793
rect 9741 31737 9766 31793
rect 9822 31737 9847 31793
rect 9903 31737 9928 31793
rect 9984 31737 10008 31793
rect 10064 31737 10088 31793
rect 10144 31737 10168 31793
rect 10224 31737 10248 31793
rect 10304 31737 10328 31793
rect 10384 31737 10408 31793
rect 10464 31737 10488 31793
rect 10544 31737 10568 31793
rect 10624 31737 10648 31793
rect 10704 31737 10728 31793
rect 10784 31737 10789 31793
rect 9593 31711 10789 31737
rect 9593 31655 9604 31711
rect 9660 31655 9685 31711
rect 9741 31655 9766 31711
rect 9822 31655 9847 31711
rect 9903 31655 9928 31711
rect 9984 31655 10008 31711
rect 10064 31655 10088 31711
rect 10144 31655 10168 31711
rect 10224 31655 10248 31711
rect 10304 31655 10328 31711
rect 10384 31655 10408 31711
rect 10464 31655 10488 31711
rect 10544 31655 10568 31711
rect 10624 31655 10648 31711
rect 10704 31655 10728 31711
rect 10784 31655 10789 31711
rect 9593 31629 10789 31655
rect 9593 31573 9604 31629
rect 9660 31573 9685 31629
rect 9741 31573 9766 31629
rect 9822 31573 9847 31629
rect 9903 31573 9928 31629
rect 9984 31573 10008 31629
rect 10064 31573 10088 31629
rect 10144 31573 10168 31629
rect 10224 31573 10248 31629
rect 10304 31573 10328 31629
rect 10384 31573 10408 31629
rect 10464 31573 10488 31629
rect 10544 31573 10568 31629
rect 10624 31573 10648 31629
rect 10704 31573 10728 31629
rect 10784 31573 10789 31629
rect 9593 31547 10789 31573
rect 9593 31491 9604 31547
rect 9660 31491 9685 31547
rect 9741 31491 9766 31547
rect 9822 31491 9847 31547
rect 9903 31491 9928 31547
rect 9984 31491 10008 31547
rect 10064 31491 10088 31547
rect 10144 31491 10168 31547
rect 10224 31491 10248 31547
rect 10304 31491 10328 31547
rect 10384 31491 10408 31547
rect 10464 31491 10488 31547
rect 10544 31491 10568 31547
rect 10624 31491 10648 31547
rect 10704 31491 10728 31547
rect 10784 31491 10789 31547
rect 9593 31478 10789 31491
rect 11090 39365 12286 39371
rect 11090 39301 11098 39365
rect 11162 39301 11178 39365
rect 11242 39301 11258 39365
rect 11322 39301 11338 39365
rect 11402 39301 11418 39365
rect 11482 39301 11498 39365
rect 11562 39301 11578 39365
rect 11642 39301 11658 39365
rect 11722 39301 11738 39365
rect 11802 39301 11818 39365
rect 11882 39301 11898 39365
rect 11962 39301 11978 39365
rect 12042 39301 12058 39365
rect 12122 39301 12138 39365
rect 12202 39301 12218 39365
rect 12282 39301 12286 39365
rect 11090 39284 12286 39301
rect 11090 39220 11098 39284
rect 11162 39220 11178 39284
rect 11242 39220 11258 39284
rect 11322 39220 11338 39284
rect 11402 39220 11418 39284
rect 11482 39220 11498 39284
rect 11562 39220 11578 39284
rect 11642 39220 11658 39284
rect 11722 39220 11738 39284
rect 11802 39220 11818 39284
rect 11882 39220 11898 39284
rect 11962 39220 11978 39284
rect 12042 39220 12058 39284
rect 12122 39220 12138 39284
rect 12202 39220 12218 39284
rect 12282 39220 12286 39284
rect 11090 39203 12286 39220
rect 11090 39139 11098 39203
rect 11162 39139 11178 39203
rect 11242 39139 11258 39203
rect 11322 39139 11338 39203
rect 11402 39139 11418 39203
rect 11482 39139 11498 39203
rect 11562 39139 11578 39203
rect 11642 39139 11658 39203
rect 11722 39139 11738 39203
rect 11802 39139 11818 39203
rect 11882 39139 11898 39203
rect 11962 39139 11978 39203
rect 12042 39139 12058 39203
rect 12122 39139 12138 39203
rect 12202 39139 12218 39203
rect 12282 39139 12286 39203
rect 11090 39122 12286 39139
rect 11090 39058 11098 39122
rect 11162 39058 11178 39122
rect 11242 39058 11258 39122
rect 11322 39058 11338 39122
rect 11402 39058 11418 39122
rect 11482 39058 11498 39122
rect 11562 39058 11578 39122
rect 11642 39058 11658 39122
rect 11722 39058 11738 39122
rect 11802 39058 11818 39122
rect 11882 39058 11898 39122
rect 11962 39058 11978 39122
rect 12042 39058 12058 39122
rect 12122 39058 12138 39122
rect 12202 39058 12218 39122
rect 12282 39058 12286 39122
rect 11090 39041 12286 39058
rect 11090 38977 11098 39041
rect 11162 38977 11178 39041
rect 11242 38977 11258 39041
rect 11322 38977 11338 39041
rect 11402 38977 11418 39041
rect 11482 38977 11498 39041
rect 11562 38977 11578 39041
rect 11642 38977 11658 39041
rect 11722 38977 11738 39041
rect 11802 38977 11818 39041
rect 11882 38977 11898 39041
rect 11962 38977 11978 39041
rect 12042 38977 12058 39041
rect 12122 38977 12138 39041
rect 12202 38977 12218 39041
rect 12282 38977 12286 39041
rect 11090 38960 12286 38977
rect 11090 38896 11098 38960
rect 11162 38896 11178 38960
rect 11242 38896 11258 38960
rect 11322 38896 11338 38960
rect 11402 38896 11418 38960
rect 11482 38896 11498 38960
rect 11562 38896 11578 38960
rect 11642 38896 11658 38960
rect 11722 38896 11738 38960
rect 11802 38896 11818 38960
rect 11882 38896 11898 38960
rect 11962 38896 11978 38960
rect 12042 38896 12058 38960
rect 12122 38896 12138 38960
rect 12202 38896 12218 38960
rect 12282 38896 12286 38960
rect 11090 38879 12286 38896
rect 11090 38815 11098 38879
rect 11162 38815 11178 38879
rect 11242 38815 11258 38879
rect 11322 38815 11338 38879
rect 11402 38815 11418 38879
rect 11482 38815 11498 38879
rect 11562 38815 11578 38879
rect 11642 38815 11658 38879
rect 11722 38815 11738 38879
rect 11802 38815 11818 38879
rect 11882 38815 11898 38879
rect 11962 38815 11978 38879
rect 12042 38815 12058 38879
rect 12122 38815 12138 38879
rect 12202 38815 12218 38879
rect 12282 38815 12286 38879
rect 11090 38798 12286 38815
rect 11090 38734 11098 38798
rect 11162 38734 11178 38798
rect 11242 38734 11258 38798
rect 11322 38734 11338 38798
rect 11402 38734 11418 38798
rect 11482 38734 11498 38798
rect 11562 38734 11578 38798
rect 11642 38734 11658 38798
rect 11722 38734 11738 38798
rect 11802 38734 11818 38798
rect 11882 38734 11898 38798
rect 11962 38734 11978 38798
rect 12042 38734 12058 38798
rect 12122 38734 12138 38798
rect 12202 38734 12218 38798
rect 12282 38734 12286 38798
rect 11090 38717 12286 38734
rect 11090 38653 11098 38717
rect 11162 38653 11178 38717
rect 11242 38653 11258 38717
rect 11322 38653 11338 38717
rect 11402 38653 11418 38717
rect 11482 38653 11498 38717
rect 11562 38653 11578 38717
rect 11642 38653 11658 38717
rect 11722 38653 11738 38717
rect 11802 38653 11818 38717
rect 11882 38653 11898 38717
rect 11962 38653 11978 38717
rect 12042 38653 12058 38717
rect 12122 38653 12138 38717
rect 12202 38653 12218 38717
rect 12282 38653 12286 38717
rect 11090 38636 12286 38653
rect 11090 38572 11098 38636
rect 11162 38572 11178 38636
rect 11242 38572 11258 38636
rect 11322 38572 11338 38636
rect 11402 38572 11418 38636
rect 11482 38572 11498 38636
rect 11562 38572 11578 38636
rect 11642 38572 11658 38636
rect 11722 38572 11738 38636
rect 11802 38572 11818 38636
rect 11882 38572 11898 38636
rect 11962 38572 11978 38636
rect 12042 38572 12058 38636
rect 12122 38572 12138 38636
rect 12202 38572 12218 38636
rect 12282 38572 12286 38636
rect 11090 38555 12286 38572
rect 11090 38491 11098 38555
rect 11162 38491 11178 38555
rect 11242 38491 11258 38555
rect 11322 38491 11338 38555
rect 11402 38491 11418 38555
rect 11482 38491 11498 38555
rect 11562 38491 11578 38555
rect 11642 38491 11658 38555
rect 11722 38491 11738 38555
rect 11802 38491 11818 38555
rect 11882 38491 11898 38555
rect 11962 38491 11978 38555
rect 12042 38491 12058 38555
rect 12122 38491 12138 38555
rect 12202 38491 12218 38555
rect 12282 38491 12286 38555
rect 11090 38474 12286 38491
rect 11090 38410 11098 38474
rect 11162 38410 11178 38474
rect 11242 38410 11258 38474
rect 11322 38410 11338 38474
rect 11402 38410 11418 38474
rect 11482 38410 11498 38474
rect 11562 38410 11578 38474
rect 11642 38410 11658 38474
rect 11722 38410 11738 38474
rect 11802 38410 11818 38474
rect 11882 38410 11898 38474
rect 11962 38410 11978 38474
rect 12042 38410 12058 38474
rect 12122 38410 12138 38474
rect 12202 38410 12218 38474
rect 12282 38410 12286 38474
rect 11090 38393 12286 38410
rect 11090 38329 11098 38393
rect 11162 38329 11178 38393
rect 11242 38329 11258 38393
rect 11322 38329 11338 38393
rect 11402 38329 11418 38393
rect 11482 38329 11498 38393
rect 11562 38329 11578 38393
rect 11642 38329 11658 38393
rect 11722 38329 11738 38393
rect 11802 38329 11818 38393
rect 11882 38329 11898 38393
rect 11962 38329 11978 38393
rect 12042 38329 12058 38393
rect 12122 38329 12138 38393
rect 12202 38329 12218 38393
rect 12282 38329 12286 38393
rect 11090 38312 12286 38329
rect 11090 38248 11098 38312
rect 11162 38248 11178 38312
rect 11242 38248 11258 38312
rect 11322 38248 11338 38312
rect 11402 38248 11418 38312
rect 11482 38248 11498 38312
rect 11562 38248 11578 38312
rect 11642 38248 11658 38312
rect 11722 38248 11738 38312
rect 11802 38248 11818 38312
rect 11882 38248 11898 38312
rect 11962 38248 11978 38312
rect 12042 38248 12058 38312
rect 12122 38248 12138 38312
rect 12202 38248 12218 38312
rect 12282 38248 12286 38312
rect 11090 38231 12286 38248
rect 11090 38167 11098 38231
rect 11162 38167 11178 38231
rect 11242 38167 11258 38231
rect 11322 38167 11338 38231
rect 11402 38167 11418 38231
rect 11482 38167 11498 38231
rect 11562 38167 11578 38231
rect 11642 38167 11658 38231
rect 11722 38167 11738 38231
rect 11802 38167 11818 38231
rect 11882 38167 11898 38231
rect 11962 38167 11978 38231
rect 12042 38167 12058 38231
rect 12122 38167 12138 38231
rect 12202 38167 12218 38231
rect 12282 38167 12286 38231
rect 11090 38150 12286 38167
rect 11090 38086 11098 38150
rect 11162 38086 11178 38150
rect 11242 38086 11258 38150
rect 11322 38086 11338 38150
rect 11402 38086 11418 38150
rect 11482 38086 11498 38150
rect 11562 38086 11578 38150
rect 11642 38086 11658 38150
rect 11722 38086 11738 38150
rect 11802 38086 11818 38150
rect 11882 38086 11898 38150
rect 11962 38086 11978 38150
rect 12042 38086 12058 38150
rect 12122 38086 12138 38150
rect 12202 38086 12218 38150
rect 12282 38086 12286 38150
rect 11090 38069 12286 38086
rect 11090 38005 11098 38069
rect 11162 38005 11178 38069
rect 11242 38005 11258 38069
rect 11322 38005 11338 38069
rect 11402 38005 11418 38069
rect 11482 38005 11498 38069
rect 11562 38005 11578 38069
rect 11642 38005 11658 38069
rect 11722 38005 11738 38069
rect 11802 38005 11818 38069
rect 11882 38005 11898 38069
rect 11962 38005 11978 38069
rect 12042 38005 12058 38069
rect 12122 38005 12138 38069
rect 12202 38005 12218 38069
rect 12282 38005 12286 38069
rect 11090 37988 12286 38005
rect 11090 37924 11098 37988
rect 11162 37924 11178 37988
rect 11242 37924 11258 37988
rect 11322 37924 11338 37988
rect 11402 37924 11418 37988
rect 11482 37924 11498 37988
rect 11562 37924 11578 37988
rect 11642 37924 11658 37988
rect 11722 37924 11738 37988
rect 11802 37924 11818 37988
rect 11882 37924 11898 37988
rect 11962 37924 11978 37988
rect 12042 37924 12058 37988
rect 12122 37924 12138 37988
rect 12202 37924 12218 37988
rect 12282 37924 12286 37988
rect 11090 37907 12286 37924
rect 11090 37843 11098 37907
rect 11162 37843 11178 37907
rect 11242 37843 11258 37907
rect 11322 37843 11338 37907
rect 11402 37843 11418 37907
rect 11482 37843 11498 37907
rect 11562 37843 11578 37907
rect 11642 37843 11658 37907
rect 11722 37843 11738 37907
rect 11802 37843 11818 37907
rect 11882 37843 11898 37907
rect 11962 37843 11978 37907
rect 12042 37843 12058 37907
rect 12122 37843 12138 37907
rect 12202 37843 12218 37907
rect 12282 37843 12286 37907
rect 11090 37826 12286 37843
rect 11090 37762 11098 37826
rect 11162 37762 11178 37826
rect 11242 37762 11258 37826
rect 11322 37762 11338 37826
rect 11402 37762 11418 37826
rect 11482 37762 11498 37826
rect 11562 37762 11578 37826
rect 11642 37762 11658 37826
rect 11722 37762 11738 37826
rect 11802 37762 11818 37826
rect 11882 37762 11898 37826
rect 11962 37762 11978 37826
rect 12042 37762 12058 37826
rect 12122 37762 12138 37826
rect 12202 37762 12218 37826
rect 12282 37762 12286 37826
rect 11090 37745 12286 37762
rect 11090 37681 11098 37745
rect 11162 37681 11178 37745
rect 11242 37681 11258 37745
rect 11322 37681 11338 37745
rect 11402 37681 11418 37745
rect 11482 37681 11498 37745
rect 11562 37681 11578 37745
rect 11642 37681 11658 37745
rect 11722 37681 11738 37745
rect 11802 37681 11818 37745
rect 11882 37681 11898 37745
rect 11962 37681 11978 37745
rect 12042 37681 12058 37745
rect 12122 37681 12138 37745
rect 12202 37681 12218 37745
rect 12282 37681 12286 37745
rect 11090 37664 12286 37681
rect 11090 37600 11098 37664
rect 11162 37600 11178 37664
rect 11242 37600 11258 37664
rect 11322 37600 11338 37664
rect 11402 37600 11418 37664
rect 11482 37600 11498 37664
rect 11562 37600 11578 37664
rect 11642 37600 11658 37664
rect 11722 37600 11738 37664
rect 11802 37600 11818 37664
rect 11882 37600 11898 37664
rect 11962 37600 11978 37664
rect 12042 37600 12058 37664
rect 12122 37600 12138 37664
rect 12202 37600 12218 37664
rect 12282 37600 12286 37664
rect 11090 37583 12286 37600
rect 11090 37519 11098 37583
rect 11162 37519 11178 37583
rect 11242 37519 11258 37583
rect 11322 37519 11338 37583
rect 11402 37519 11418 37583
rect 11482 37519 11498 37583
rect 11562 37519 11578 37583
rect 11642 37519 11658 37583
rect 11722 37519 11738 37583
rect 11802 37519 11818 37583
rect 11882 37519 11898 37583
rect 11962 37519 11978 37583
rect 12042 37519 12058 37583
rect 12122 37519 12138 37583
rect 12202 37519 12218 37583
rect 12282 37519 12286 37583
rect 11090 37502 12286 37519
rect 11090 37438 11098 37502
rect 11162 37438 11178 37502
rect 11242 37438 11258 37502
rect 11322 37438 11338 37502
rect 11402 37438 11418 37502
rect 11482 37438 11498 37502
rect 11562 37438 11578 37502
rect 11642 37438 11658 37502
rect 11722 37438 11738 37502
rect 11802 37438 11818 37502
rect 11882 37438 11898 37502
rect 11962 37438 11978 37502
rect 12042 37438 12058 37502
rect 12122 37438 12138 37502
rect 12202 37438 12218 37502
rect 12282 37438 12286 37502
rect 11090 37421 12286 37438
rect 11090 37357 11098 37421
rect 11162 37357 11178 37421
rect 11242 37357 11258 37421
rect 11322 37357 11338 37421
rect 11402 37357 11418 37421
rect 11482 37357 11498 37421
rect 11562 37357 11578 37421
rect 11642 37357 11658 37421
rect 11722 37357 11738 37421
rect 11802 37357 11818 37421
rect 11882 37357 11898 37421
rect 11962 37357 11978 37421
rect 12042 37357 12058 37421
rect 12122 37357 12138 37421
rect 12202 37357 12218 37421
rect 12282 37357 12286 37421
rect 11090 37340 12286 37357
rect 11090 37276 11098 37340
rect 11162 37276 11178 37340
rect 11242 37276 11258 37340
rect 11322 37276 11338 37340
rect 11402 37276 11418 37340
rect 11482 37276 11498 37340
rect 11562 37276 11578 37340
rect 11642 37276 11658 37340
rect 11722 37276 11738 37340
rect 11802 37276 11818 37340
rect 11882 37276 11898 37340
rect 11962 37276 11978 37340
rect 12042 37276 12058 37340
rect 12122 37276 12138 37340
rect 12202 37276 12218 37340
rect 12282 37276 12286 37340
rect 11090 37259 12286 37276
rect 11090 37195 11098 37259
rect 11162 37195 11178 37259
rect 11242 37195 11258 37259
rect 11322 37195 11338 37259
rect 11402 37195 11418 37259
rect 11482 37195 11498 37259
rect 11562 37195 11578 37259
rect 11642 37195 11658 37259
rect 11722 37195 11738 37259
rect 11802 37195 11818 37259
rect 11882 37195 11898 37259
rect 11962 37195 11978 37259
rect 12042 37195 12058 37259
rect 12122 37195 12138 37259
rect 12202 37195 12218 37259
rect 12282 37195 12286 37259
rect 11090 37178 12286 37195
rect 11090 37114 11098 37178
rect 11162 37114 11178 37178
rect 11242 37114 11258 37178
rect 11322 37114 11338 37178
rect 11402 37114 11418 37178
rect 11482 37114 11498 37178
rect 11562 37114 11578 37178
rect 11642 37114 11658 37178
rect 11722 37114 11738 37178
rect 11802 37114 11818 37178
rect 11882 37114 11898 37178
rect 11962 37114 11978 37178
rect 12042 37114 12058 37178
rect 12122 37114 12138 37178
rect 12202 37114 12218 37178
rect 12282 37114 12286 37178
rect 11090 37097 12286 37114
rect 11090 37033 11098 37097
rect 11162 37033 11178 37097
rect 11242 37033 11258 37097
rect 11322 37033 11338 37097
rect 11402 37033 11418 37097
rect 11482 37033 11498 37097
rect 11562 37033 11578 37097
rect 11642 37033 11658 37097
rect 11722 37033 11738 37097
rect 11802 37033 11818 37097
rect 11882 37033 11898 37097
rect 11962 37033 11978 37097
rect 12042 37033 12058 37097
rect 12122 37033 12138 37097
rect 12202 37033 12218 37097
rect 12282 37033 12286 37097
rect 11090 37016 12286 37033
rect 11090 36952 11098 37016
rect 11162 36952 11178 37016
rect 11242 36952 11258 37016
rect 11322 36952 11338 37016
rect 11402 36952 11418 37016
rect 11482 36952 11498 37016
rect 11562 36952 11578 37016
rect 11642 36952 11658 37016
rect 11722 36952 11738 37016
rect 11802 36952 11818 37016
rect 11882 36952 11898 37016
rect 11962 36952 11978 37016
rect 12042 36952 12058 37016
rect 12122 36952 12138 37016
rect 12202 36952 12218 37016
rect 12282 36952 12286 37016
rect 11090 36935 12286 36952
rect 11090 36871 11098 36935
rect 11162 36871 11178 36935
rect 11242 36871 11258 36935
rect 11322 36871 11338 36935
rect 11402 36871 11418 36935
rect 11482 36871 11498 36935
rect 11562 36871 11578 36935
rect 11642 36871 11658 36935
rect 11722 36871 11738 36935
rect 11802 36871 11818 36935
rect 11882 36871 11898 36935
rect 11962 36871 11978 36935
rect 12042 36871 12058 36935
rect 12122 36871 12138 36935
rect 12202 36871 12218 36935
rect 12282 36871 12286 36935
rect 11090 36854 12286 36871
rect 11090 36790 11098 36854
rect 11162 36790 11178 36854
rect 11242 36790 11258 36854
rect 11322 36790 11338 36854
rect 11402 36790 11418 36854
rect 11482 36790 11498 36854
rect 11562 36790 11578 36854
rect 11642 36790 11658 36854
rect 11722 36790 11738 36854
rect 11802 36790 11818 36854
rect 11882 36790 11898 36854
rect 11962 36790 11978 36854
rect 12042 36790 12058 36854
rect 12122 36790 12138 36854
rect 12202 36790 12218 36854
rect 12282 36790 12286 36854
rect 11090 36773 12286 36790
rect 11090 36709 11098 36773
rect 11162 36709 11178 36773
rect 11242 36709 11258 36773
rect 11322 36709 11338 36773
rect 11402 36709 11418 36773
rect 11482 36709 11498 36773
rect 11562 36709 11578 36773
rect 11642 36709 11658 36773
rect 11722 36709 11738 36773
rect 11802 36709 11818 36773
rect 11882 36709 11898 36773
rect 11962 36709 11978 36773
rect 12042 36709 12058 36773
rect 12122 36709 12138 36773
rect 12202 36709 12218 36773
rect 12282 36709 12286 36773
rect 11090 36692 12286 36709
rect 11090 36628 11098 36692
rect 11162 36628 11178 36692
rect 11242 36628 11258 36692
rect 11322 36628 11338 36692
rect 11402 36628 11418 36692
rect 11482 36628 11498 36692
rect 11562 36628 11578 36692
rect 11642 36628 11658 36692
rect 11722 36628 11738 36692
rect 11802 36628 11818 36692
rect 11882 36628 11898 36692
rect 11962 36628 11978 36692
rect 12042 36628 12058 36692
rect 12122 36628 12138 36692
rect 12202 36628 12218 36692
rect 12282 36628 12286 36692
rect 11090 36611 12286 36628
rect 11090 36547 11098 36611
rect 11162 36547 11178 36611
rect 11242 36547 11258 36611
rect 11322 36547 11338 36611
rect 11402 36547 11418 36611
rect 11482 36547 11498 36611
rect 11562 36547 11578 36611
rect 11642 36547 11658 36611
rect 11722 36547 11738 36611
rect 11802 36547 11818 36611
rect 11882 36547 11898 36611
rect 11962 36547 11978 36611
rect 12042 36547 12058 36611
rect 12122 36547 12138 36611
rect 12202 36547 12218 36611
rect 12282 36547 12286 36611
rect 11090 36530 12286 36547
rect 11090 36466 11098 36530
rect 11162 36466 11178 36530
rect 11242 36466 11258 36530
rect 11322 36466 11338 36530
rect 11402 36466 11418 36530
rect 11482 36466 11498 36530
rect 11562 36466 11578 36530
rect 11642 36466 11658 36530
rect 11722 36466 11738 36530
rect 11802 36466 11818 36530
rect 11882 36466 11898 36530
rect 11962 36466 11978 36530
rect 12042 36466 12058 36530
rect 12122 36466 12138 36530
rect 12202 36466 12218 36530
rect 12282 36466 12286 36530
rect 11090 36449 12286 36466
rect 11090 36385 11098 36449
rect 11162 36385 11178 36449
rect 11242 36385 11258 36449
rect 11322 36385 11338 36449
rect 11402 36385 11418 36449
rect 11482 36385 11498 36449
rect 11562 36385 11578 36449
rect 11642 36385 11658 36449
rect 11722 36385 11738 36449
rect 11802 36385 11818 36449
rect 11882 36385 11898 36449
rect 11962 36385 11978 36449
rect 12042 36385 12058 36449
rect 12122 36385 12138 36449
rect 12202 36385 12218 36449
rect 12282 36385 12286 36449
rect 11090 36368 12286 36385
rect 11090 36304 11098 36368
rect 11162 36304 11178 36368
rect 11242 36304 11258 36368
rect 11322 36304 11338 36368
rect 11402 36304 11418 36368
rect 11482 36304 11498 36368
rect 11562 36304 11578 36368
rect 11642 36304 11658 36368
rect 11722 36304 11738 36368
rect 11802 36304 11818 36368
rect 11882 36304 11898 36368
rect 11962 36304 11978 36368
rect 12042 36304 12058 36368
rect 12122 36304 12138 36368
rect 12202 36304 12218 36368
rect 12282 36304 12286 36368
rect 11090 36287 12286 36304
rect 11090 36223 11098 36287
rect 11162 36223 11178 36287
rect 11242 36223 11258 36287
rect 11322 36223 11338 36287
rect 11402 36223 11418 36287
rect 11482 36223 11498 36287
rect 11562 36223 11578 36287
rect 11642 36223 11658 36287
rect 11722 36223 11738 36287
rect 11802 36223 11818 36287
rect 11882 36223 11898 36287
rect 11962 36223 11978 36287
rect 12042 36223 12058 36287
rect 12122 36223 12138 36287
rect 12202 36223 12218 36287
rect 12282 36223 12286 36287
rect 11090 36206 12286 36223
rect 11090 36142 11098 36206
rect 11162 36142 11178 36206
rect 11242 36142 11258 36206
rect 11322 36142 11338 36206
rect 11402 36142 11418 36206
rect 11482 36142 11498 36206
rect 11562 36142 11578 36206
rect 11642 36142 11658 36206
rect 11722 36142 11738 36206
rect 11802 36142 11818 36206
rect 11882 36142 11898 36206
rect 11962 36142 11978 36206
rect 12042 36142 12058 36206
rect 12122 36142 12138 36206
rect 12202 36142 12218 36206
rect 12282 36142 12286 36206
rect 11090 36124 12286 36142
rect 11090 36060 11098 36124
rect 11162 36060 11178 36124
rect 11242 36060 11258 36124
rect 11322 36060 11338 36124
rect 11402 36060 11418 36124
rect 11482 36060 11498 36124
rect 11562 36060 11578 36124
rect 11642 36060 11658 36124
rect 11722 36060 11738 36124
rect 11802 36060 11818 36124
rect 11882 36060 11898 36124
rect 11962 36060 11978 36124
rect 12042 36060 12058 36124
rect 12122 36060 12138 36124
rect 12202 36060 12218 36124
rect 12282 36060 12286 36124
rect 11090 36042 12286 36060
rect 11090 35978 11098 36042
rect 11162 35978 11178 36042
rect 11242 35978 11258 36042
rect 11322 35978 11338 36042
rect 11402 35978 11418 36042
rect 11482 35978 11498 36042
rect 11562 35978 11578 36042
rect 11642 35978 11658 36042
rect 11722 35978 11738 36042
rect 11802 35978 11818 36042
rect 11882 35978 11898 36042
rect 11962 35978 11978 36042
rect 12042 35978 12058 36042
rect 12122 35978 12138 36042
rect 12202 35978 12218 36042
rect 12282 35978 12286 36042
rect 11090 35960 12286 35978
rect 11090 35896 11098 35960
rect 11162 35896 11178 35960
rect 11242 35896 11258 35960
rect 11322 35896 11338 35960
rect 11402 35896 11418 35960
rect 11482 35896 11498 35960
rect 11562 35896 11578 35960
rect 11642 35896 11658 35960
rect 11722 35896 11738 35960
rect 11802 35896 11818 35960
rect 11882 35896 11898 35960
rect 11962 35896 11978 35960
rect 12042 35896 12058 35960
rect 12122 35896 12138 35960
rect 12202 35896 12218 35960
rect 12282 35896 12286 35960
rect 11090 35878 12286 35896
rect 11090 35814 11098 35878
rect 11162 35814 11178 35878
rect 11242 35814 11258 35878
rect 11322 35814 11338 35878
rect 11402 35814 11418 35878
rect 11482 35814 11498 35878
rect 11562 35814 11578 35878
rect 11642 35814 11658 35878
rect 11722 35814 11738 35878
rect 11802 35814 11818 35878
rect 11882 35814 11898 35878
rect 11962 35814 11978 35878
rect 12042 35814 12058 35878
rect 12122 35814 12138 35878
rect 12202 35814 12218 35878
rect 12282 35814 12286 35878
rect 11090 35796 12286 35814
rect 11090 35732 11098 35796
rect 11162 35732 11178 35796
rect 11242 35732 11258 35796
rect 11322 35732 11338 35796
rect 11402 35732 11418 35796
rect 11482 35732 11498 35796
rect 11562 35732 11578 35796
rect 11642 35732 11658 35796
rect 11722 35732 11738 35796
rect 11802 35732 11818 35796
rect 11882 35732 11898 35796
rect 11962 35732 11978 35796
rect 12042 35732 12058 35796
rect 12122 35732 12138 35796
rect 12202 35732 12218 35796
rect 12282 35732 12286 35796
rect 11090 35714 12286 35732
rect 11090 35650 11098 35714
rect 11162 35650 11178 35714
rect 11242 35650 11258 35714
rect 11322 35650 11338 35714
rect 11402 35650 11418 35714
rect 11482 35650 11498 35714
rect 11562 35650 11578 35714
rect 11642 35650 11658 35714
rect 11722 35650 11738 35714
rect 11802 35650 11818 35714
rect 11882 35650 11898 35714
rect 11962 35650 11978 35714
rect 12042 35650 12058 35714
rect 12122 35650 12138 35714
rect 12202 35650 12218 35714
rect 12282 35650 12286 35714
rect 11090 35632 12286 35650
rect 11090 35568 11098 35632
rect 11162 35568 11178 35632
rect 11242 35568 11258 35632
rect 11322 35568 11338 35632
rect 11402 35568 11418 35632
rect 11482 35568 11498 35632
rect 11562 35568 11578 35632
rect 11642 35568 11658 35632
rect 11722 35568 11738 35632
rect 11802 35568 11818 35632
rect 11882 35568 11898 35632
rect 11962 35568 11978 35632
rect 12042 35568 12058 35632
rect 12122 35568 12138 35632
rect 12202 35568 12218 35632
rect 12282 35568 12286 35632
rect 11090 35550 12286 35568
rect 11090 35486 11098 35550
rect 11162 35486 11178 35550
rect 11242 35486 11258 35550
rect 11322 35486 11338 35550
rect 11402 35486 11418 35550
rect 11482 35486 11498 35550
rect 11562 35486 11578 35550
rect 11642 35486 11658 35550
rect 11722 35486 11738 35550
rect 11802 35486 11818 35550
rect 11882 35486 11898 35550
rect 11962 35486 11978 35550
rect 12042 35486 12058 35550
rect 12122 35486 12138 35550
rect 12202 35486 12218 35550
rect 12282 35486 12286 35550
rect 11090 35468 12286 35486
rect 11090 35404 11098 35468
rect 11162 35404 11178 35468
rect 11242 35404 11258 35468
rect 11322 35404 11338 35468
rect 11402 35404 11418 35468
rect 11482 35404 11498 35468
rect 11562 35404 11578 35468
rect 11642 35404 11658 35468
rect 11722 35404 11738 35468
rect 11802 35404 11818 35468
rect 11882 35404 11898 35468
rect 11962 35404 11978 35468
rect 12042 35404 12058 35468
rect 12122 35404 12138 35468
rect 12202 35404 12218 35468
rect 12282 35404 12286 35468
rect 11090 35386 12286 35404
rect 11090 35322 11098 35386
rect 11162 35322 11178 35386
rect 11242 35322 11258 35386
rect 11322 35322 11338 35386
rect 11402 35322 11418 35386
rect 11482 35322 11498 35386
rect 11562 35322 11578 35386
rect 11642 35322 11658 35386
rect 11722 35322 11738 35386
rect 11802 35322 11818 35386
rect 11882 35322 11898 35386
rect 11962 35322 11978 35386
rect 12042 35322 12058 35386
rect 12122 35322 12138 35386
rect 12202 35322 12218 35386
rect 12282 35322 12286 35386
rect 11090 35304 12286 35322
rect 11090 35240 11098 35304
rect 11162 35240 11178 35304
rect 11242 35240 11258 35304
rect 11322 35240 11338 35304
rect 11402 35240 11418 35304
rect 11482 35240 11498 35304
rect 11562 35240 11578 35304
rect 11642 35240 11658 35304
rect 11722 35240 11738 35304
rect 11802 35240 11818 35304
rect 11882 35240 11898 35304
rect 11962 35240 11978 35304
rect 12042 35240 12058 35304
rect 12122 35240 12138 35304
rect 12202 35240 12218 35304
rect 12282 35240 12286 35304
rect 11090 35222 12286 35240
rect 11090 35158 11098 35222
rect 11162 35158 11178 35222
rect 11242 35158 11258 35222
rect 11322 35158 11338 35222
rect 11402 35158 11418 35222
rect 11482 35158 11498 35222
rect 11562 35158 11578 35222
rect 11642 35158 11658 35222
rect 11722 35158 11738 35222
rect 11802 35158 11818 35222
rect 11882 35158 11898 35222
rect 11962 35158 11978 35222
rect 12042 35158 12058 35222
rect 12122 35158 12138 35222
rect 12202 35158 12218 35222
rect 12282 35158 12286 35222
rect 11090 32613 12286 35158
rect 11090 32557 11101 32613
rect 11157 32557 11182 32613
rect 11238 32557 11263 32613
rect 11319 32557 11344 32613
rect 11400 32557 11425 32613
rect 11481 32557 11505 32613
rect 11561 32557 11585 32613
rect 11641 32557 11665 32613
rect 11721 32557 11745 32613
rect 11801 32557 11825 32613
rect 11881 32557 11905 32613
rect 11961 32557 11985 32613
rect 12041 32557 12065 32613
rect 12121 32557 12145 32613
rect 12201 32557 12225 32613
rect 12281 32557 12286 32613
rect 11090 32531 12286 32557
rect 11090 32475 11101 32531
rect 11157 32475 11182 32531
rect 11238 32475 11263 32531
rect 11319 32475 11344 32531
rect 11400 32475 11425 32531
rect 11481 32475 11505 32531
rect 11561 32475 11585 32531
rect 11641 32475 11665 32531
rect 11721 32475 11745 32531
rect 11801 32475 11825 32531
rect 11881 32475 11905 32531
rect 11961 32475 11985 32531
rect 12041 32475 12065 32531
rect 12121 32475 12145 32531
rect 12201 32475 12225 32531
rect 12281 32475 12286 32531
rect 11090 32449 12286 32475
rect 11090 32393 11101 32449
rect 11157 32393 11182 32449
rect 11238 32393 11263 32449
rect 11319 32393 11344 32449
rect 11400 32393 11425 32449
rect 11481 32393 11505 32449
rect 11561 32393 11585 32449
rect 11641 32393 11665 32449
rect 11721 32393 11745 32449
rect 11801 32393 11825 32449
rect 11881 32393 11905 32449
rect 11961 32393 11985 32449
rect 12041 32393 12065 32449
rect 12121 32393 12145 32449
rect 12201 32393 12225 32449
rect 12281 32393 12286 32449
rect 11090 32367 12286 32393
rect 11090 32311 11101 32367
rect 11157 32311 11182 32367
rect 11238 32311 11263 32367
rect 11319 32311 11344 32367
rect 11400 32311 11425 32367
rect 11481 32311 11505 32367
rect 11561 32311 11585 32367
rect 11641 32311 11665 32367
rect 11721 32311 11745 32367
rect 11801 32311 11825 32367
rect 11881 32311 11905 32367
rect 11961 32311 11985 32367
rect 12041 32311 12065 32367
rect 12121 32311 12145 32367
rect 12201 32311 12225 32367
rect 12281 32311 12286 32367
rect 11090 32285 12286 32311
rect 11090 32229 11101 32285
rect 11157 32229 11182 32285
rect 11238 32229 11263 32285
rect 11319 32229 11344 32285
rect 11400 32229 11425 32285
rect 11481 32229 11505 32285
rect 11561 32229 11585 32285
rect 11641 32229 11665 32285
rect 11721 32229 11745 32285
rect 11801 32229 11825 32285
rect 11881 32229 11905 32285
rect 11961 32229 11985 32285
rect 12041 32229 12065 32285
rect 12121 32229 12145 32285
rect 12201 32229 12225 32285
rect 12281 32229 12286 32285
rect 11090 32203 12286 32229
rect 11090 32147 11101 32203
rect 11157 32147 11182 32203
rect 11238 32147 11263 32203
rect 11319 32147 11344 32203
rect 11400 32147 11425 32203
rect 11481 32147 11505 32203
rect 11561 32147 11585 32203
rect 11641 32147 11665 32203
rect 11721 32147 11745 32203
rect 11801 32147 11825 32203
rect 11881 32147 11905 32203
rect 11961 32147 11985 32203
rect 12041 32147 12065 32203
rect 12121 32147 12145 32203
rect 12201 32147 12225 32203
rect 12281 32147 12286 32203
rect 11090 32121 12286 32147
rect 11090 32065 11101 32121
rect 11157 32065 11182 32121
rect 11238 32065 11263 32121
rect 11319 32065 11344 32121
rect 11400 32065 11425 32121
rect 11481 32065 11505 32121
rect 11561 32065 11585 32121
rect 11641 32065 11665 32121
rect 11721 32065 11745 32121
rect 11801 32065 11825 32121
rect 11881 32065 11905 32121
rect 11961 32065 11985 32121
rect 12041 32065 12065 32121
rect 12121 32065 12145 32121
rect 12201 32065 12225 32121
rect 12281 32065 12286 32121
rect 11090 32039 12286 32065
rect 11090 31983 11101 32039
rect 11157 31983 11182 32039
rect 11238 31983 11263 32039
rect 11319 31983 11344 32039
rect 11400 31983 11425 32039
rect 11481 31983 11505 32039
rect 11561 31983 11585 32039
rect 11641 31983 11665 32039
rect 11721 31983 11745 32039
rect 11801 31983 11825 32039
rect 11881 31983 11905 32039
rect 11961 31983 11985 32039
rect 12041 31983 12065 32039
rect 12121 31983 12145 32039
rect 12201 31983 12225 32039
rect 12281 31983 12286 32039
rect 11090 31957 12286 31983
rect 11090 31901 11101 31957
rect 11157 31901 11182 31957
rect 11238 31901 11263 31957
rect 11319 31901 11344 31957
rect 11400 31901 11425 31957
rect 11481 31901 11505 31957
rect 11561 31901 11585 31957
rect 11641 31901 11665 31957
rect 11721 31901 11745 31957
rect 11801 31901 11825 31957
rect 11881 31901 11905 31957
rect 11961 31901 11985 31957
rect 12041 31901 12065 31957
rect 12121 31901 12145 31957
rect 12201 31901 12225 31957
rect 12281 31901 12286 31957
rect 11090 31875 12286 31901
rect 11090 31819 11101 31875
rect 11157 31819 11182 31875
rect 11238 31819 11263 31875
rect 11319 31819 11344 31875
rect 11400 31819 11425 31875
rect 11481 31819 11505 31875
rect 11561 31819 11585 31875
rect 11641 31819 11665 31875
rect 11721 31819 11745 31875
rect 11801 31819 11825 31875
rect 11881 31819 11905 31875
rect 11961 31819 11985 31875
rect 12041 31819 12065 31875
rect 12121 31819 12145 31875
rect 12201 31819 12225 31875
rect 12281 31819 12286 31875
rect 11090 31793 12286 31819
rect 11090 31737 11101 31793
rect 11157 31737 11182 31793
rect 11238 31737 11263 31793
rect 11319 31737 11344 31793
rect 11400 31737 11425 31793
rect 11481 31737 11505 31793
rect 11561 31737 11585 31793
rect 11641 31737 11665 31793
rect 11721 31737 11745 31793
rect 11801 31737 11825 31793
rect 11881 31737 11905 31793
rect 11961 31737 11985 31793
rect 12041 31737 12065 31793
rect 12121 31737 12145 31793
rect 12201 31737 12225 31793
rect 12281 31737 12286 31793
rect 11090 31711 12286 31737
rect 11090 31655 11101 31711
rect 11157 31655 11182 31711
rect 11238 31655 11263 31711
rect 11319 31655 11344 31711
rect 11400 31655 11425 31711
rect 11481 31655 11505 31711
rect 11561 31655 11585 31711
rect 11641 31655 11665 31711
rect 11721 31655 11745 31711
rect 11801 31655 11825 31711
rect 11881 31655 11905 31711
rect 11961 31655 11985 31711
rect 12041 31655 12065 31711
rect 12121 31655 12145 31711
rect 12201 31655 12225 31711
rect 12281 31655 12286 31711
rect 11090 31629 12286 31655
rect 11090 31573 11101 31629
rect 11157 31573 11182 31629
rect 11238 31573 11263 31629
rect 11319 31573 11344 31629
rect 11400 31573 11425 31629
rect 11481 31573 11505 31629
rect 11561 31573 11585 31629
rect 11641 31573 11665 31629
rect 11721 31573 11745 31629
rect 11801 31573 11825 31629
rect 11881 31573 11905 31629
rect 11961 31573 11985 31629
rect 12041 31573 12065 31629
rect 12121 31573 12145 31629
rect 12201 31573 12225 31629
rect 12281 31573 12286 31629
rect 11090 31547 12286 31573
rect 11090 31491 11101 31547
rect 11157 31491 11182 31547
rect 11238 31491 11263 31547
rect 11319 31491 11344 31547
rect 11400 31491 11425 31547
rect 11481 31491 11505 31547
rect 11561 31491 11585 31547
rect 11641 31491 11665 31547
rect 11721 31491 11745 31547
rect 11801 31491 11825 31547
rect 11881 31491 11905 31547
rect 11961 31491 11985 31547
rect 12041 31491 12065 31547
rect 12121 31491 12145 31547
rect 12201 31491 12225 31547
rect 12281 31491 12286 31547
rect 11090 31478 12286 31491
rect 12587 39308 12588 39372
rect 12652 39308 12676 39372
rect 12740 39308 12764 39372
rect 12828 39308 12852 39372
rect 12916 39308 12940 39372
rect 13004 39308 13005 39372
rect 12587 39292 13005 39308
rect 12587 39228 12588 39292
rect 12652 39228 12676 39292
rect 12740 39228 12764 39292
rect 12828 39228 12852 39292
rect 12916 39228 12940 39292
rect 13004 39228 13005 39292
rect 12587 39212 13005 39228
rect 12587 39148 12588 39212
rect 12652 39148 12676 39212
rect 12740 39148 12764 39212
rect 12828 39148 12852 39212
rect 12916 39148 12940 39212
rect 13004 39148 13005 39212
rect 12587 39132 13005 39148
rect 12587 39068 12588 39132
rect 12652 39068 12676 39132
rect 12740 39068 12764 39132
rect 12828 39068 12852 39132
rect 12916 39068 12940 39132
rect 13004 39068 13005 39132
rect 12587 39052 13005 39068
rect 12587 38988 12588 39052
rect 12652 38988 12676 39052
rect 12740 38988 12764 39052
rect 12828 38988 12852 39052
rect 12916 38988 12940 39052
rect 13004 38988 13005 39052
rect 12587 38972 13005 38988
rect 12587 38908 12588 38972
rect 12652 38908 12676 38972
rect 12740 38908 12764 38972
rect 12828 38908 12852 38972
rect 12916 38908 12940 38972
rect 13004 38908 13005 38972
rect 12587 38892 13005 38908
rect 12587 38828 12588 38892
rect 12652 38828 12676 38892
rect 12740 38828 12764 38892
rect 12828 38828 12852 38892
rect 12916 38828 12940 38892
rect 13004 38828 13005 38892
rect 12587 38812 13005 38828
rect 12587 38748 12588 38812
rect 12652 38748 12676 38812
rect 12740 38748 12764 38812
rect 12828 38748 12852 38812
rect 12916 38748 12940 38812
rect 13004 38748 13005 38812
rect 12587 38731 13005 38748
rect 12587 38667 12588 38731
rect 12652 38667 12676 38731
rect 12740 38667 12764 38731
rect 12828 38667 12852 38731
rect 12916 38667 12940 38731
rect 13004 38667 13005 38731
rect 12587 38650 13005 38667
rect 12587 38586 12588 38650
rect 12652 38586 12676 38650
rect 12740 38586 12764 38650
rect 12828 38586 12852 38650
rect 12916 38586 12940 38650
rect 13004 38586 13005 38650
rect 12587 38569 13005 38586
rect 12587 38505 12588 38569
rect 12652 38505 12676 38569
rect 12740 38505 12764 38569
rect 12828 38505 12852 38569
rect 12916 38505 12940 38569
rect 13004 38505 13005 38569
rect 12587 38488 13005 38505
rect 12587 38424 12588 38488
rect 12652 38424 12676 38488
rect 12740 38424 12764 38488
rect 12828 38424 12852 38488
rect 12916 38424 12940 38488
rect 13004 38424 13005 38488
rect 12587 38407 13005 38424
rect 12587 38343 12588 38407
rect 12652 38343 12676 38407
rect 12740 38343 12764 38407
rect 12828 38343 12852 38407
rect 12916 38343 12940 38407
rect 13004 38343 13005 38407
rect 12587 38326 13005 38343
rect 12587 38262 12588 38326
rect 12652 38262 12676 38326
rect 12740 38262 12764 38326
rect 12828 38262 12852 38326
rect 12916 38262 12940 38326
rect 13004 38262 13005 38326
rect 12587 38245 13005 38262
rect 12587 38181 12588 38245
rect 12652 38181 12676 38245
rect 12740 38181 12764 38245
rect 12828 38181 12852 38245
rect 12916 38181 12940 38245
rect 13004 38181 13005 38245
rect 12587 38164 13005 38181
rect 12587 38100 12588 38164
rect 12652 38100 12676 38164
rect 12740 38100 12764 38164
rect 12828 38100 12852 38164
rect 12916 38100 12940 38164
rect 13004 38100 13005 38164
rect 12587 38083 13005 38100
rect 12587 38019 12588 38083
rect 12652 38019 12676 38083
rect 12740 38019 12764 38083
rect 12828 38019 12852 38083
rect 12916 38019 12940 38083
rect 13004 38019 13005 38083
rect 12587 38002 13005 38019
rect 12587 37938 12588 38002
rect 12652 37938 12676 38002
rect 12740 37938 12764 38002
rect 12828 37938 12852 38002
rect 12916 37938 12940 38002
rect 13004 37938 13005 38002
rect 12587 37921 13005 37938
rect 12587 37857 12588 37921
rect 12652 37857 12676 37921
rect 12740 37857 12764 37921
rect 12828 37857 12852 37921
rect 12916 37857 12940 37921
rect 13004 37857 13005 37921
rect 12587 37840 13005 37857
rect 12587 37776 12588 37840
rect 12652 37776 12676 37840
rect 12740 37776 12764 37840
rect 12828 37776 12852 37840
rect 12916 37776 12940 37840
rect 13004 37776 13005 37840
rect 12587 37759 13005 37776
rect 12587 37695 12588 37759
rect 12652 37695 12676 37759
rect 12740 37695 12764 37759
rect 12828 37695 12852 37759
rect 12916 37695 12940 37759
rect 13004 37695 13005 37759
rect 12587 37678 13005 37695
rect 12587 37614 12588 37678
rect 12652 37614 12676 37678
rect 12740 37614 12764 37678
rect 12828 37614 12852 37678
rect 12916 37614 12940 37678
rect 13004 37614 13005 37678
rect 12587 37597 13005 37614
rect 12587 37533 12588 37597
rect 12652 37533 12676 37597
rect 12740 37533 12764 37597
rect 12828 37533 12852 37597
rect 12916 37533 12940 37597
rect 13004 37533 13005 37597
rect 12587 37516 13005 37533
rect 12587 37452 12588 37516
rect 12652 37452 12676 37516
rect 12740 37452 12764 37516
rect 12828 37452 12852 37516
rect 12916 37452 12940 37516
rect 13004 37452 13005 37516
rect 12587 37435 13005 37452
rect 12587 37371 12588 37435
rect 12652 37371 12676 37435
rect 12740 37371 12764 37435
rect 12828 37371 12852 37435
rect 12916 37371 12940 37435
rect 13004 37371 13005 37435
rect 12587 37354 13005 37371
rect 12587 37290 12588 37354
rect 12652 37290 12676 37354
rect 12740 37290 12764 37354
rect 12828 37290 12852 37354
rect 12916 37290 12940 37354
rect 13004 37290 13005 37354
rect 12587 37273 13005 37290
rect 12587 37209 12588 37273
rect 12652 37209 12676 37273
rect 12740 37209 12764 37273
rect 12828 37209 12852 37273
rect 12916 37209 12940 37273
rect 13004 37209 13005 37273
rect 12587 37192 13005 37209
rect 12587 37128 12588 37192
rect 12652 37128 12676 37192
rect 12740 37128 12764 37192
rect 12828 37128 12852 37192
rect 12916 37128 12940 37192
rect 13004 37128 13005 37192
rect 12587 37111 13005 37128
rect 12587 37047 12588 37111
rect 12652 37047 12676 37111
rect 12740 37047 12764 37111
rect 12828 37047 12852 37111
rect 12916 37047 12940 37111
rect 13004 37047 13005 37111
rect 12587 37030 13005 37047
rect 12587 36966 12588 37030
rect 12652 36966 12676 37030
rect 12740 36966 12764 37030
rect 12828 36966 12852 37030
rect 12916 36966 12940 37030
rect 13004 36966 13005 37030
rect 12587 36949 13005 36966
rect 12587 36885 12588 36949
rect 12652 36885 12676 36949
rect 12740 36885 12764 36949
rect 12828 36885 12852 36949
rect 12916 36885 12940 36949
rect 13004 36885 13005 36949
rect 12587 36868 13005 36885
rect 12587 36804 12588 36868
rect 12652 36804 12676 36868
rect 12740 36804 12764 36868
rect 12828 36804 12852 36868
rect 12916 36804 12940 36868
rect 13004 36804 13005 36868
rect 12587 36787 13005 36804
rect 12587 36723 12588 36787
rect 12652 36723 12676 36787
rect 12740 36723 12764 36787
rect 12828 36723 12852 36787
rect 12916 36723 12940 36787
rect 13004 36723 13005 36787
rect 12587 36706 13005 36723
rect 12587 36642 12588 36706
rect 12652 36642 12676 36706
rect 12740 36642 12764 36706
rect 12828 36642 12852 36706
rect 12916 36642 12940 36706
rect 13004 36642 13005 36706
rect 12587 36625 13005 36642
rect 12587 36561 12588 36625
rect 12652 36561 12676 36625
rect 12740 36561 12764 36625
rect 12828 36561 12852 36625
rect 12916 36561 12940 36625
rect 13004 36561 13005 36625
rect 12587 36544 13005 36561
rect 12587 36480 12588 36544
rect 12652 36480 12676 36544
rect 12740 36480 12764 36544
rect 12828 36480 12852 36544
rect 12916 36480 12940 36544
rect 13004 36480 13005 36544
rect 12587 36463 13005 36480
rect 12587 36399 12588 36463
rect 12652 36399 12676 36463
rect 12740 36399 12764 36463
rect 12828 36399 12852 36463
rect 12916 36399 12940 36463
rect 13004 36399 13005 36463
rect 12587 36382 13005 36399
rect 12587 36318 12588 36382
rect 12652 36318 12676 36382
rect 12740 36318 12764 36382
rect 12828 36318 12852 36382
rect 12916 36318 12940 36382
rect 13004 36318 13005 36382
rect 12587 36301 13005 36318
rect 12587 36237 12588 36301
rect 12652 36237 12676 36301
rect 12740 36237 12764 36301
rect 12828 36237 12852 36301
rect 12916 36237 12940 36301
rect 13004 36237 13005 36301
rect 12587 36220 13005 36237
rect 12587 36156 12588 36220
rect 12652 36156 12676 36220
rect 12740 36156 12764 36220
rect 12828 36156 12852 36220
rect 12916 36156 12940 36220
rect 13004 36156 13005 36220
rect 12587 36139 13005 36156
rect 12587 36075 12588 36139
rect 12652 36075 12676 36139
rect 12740 36075 12764 36139
rect 12828 36075 12852 36139
rect 12916 36075 12940 36139
rect 13004 36075 13005 36139
rect 12587 36058 13005 36075
rect 12587 35994 12588 36058
rect 12652 35994 12676 36058
rect 12740 35994 12764 36058
rect 12828 35994 12852 36058
rect 12916 35994 12940 36058
rect 13004 35994 13005 36058
rect 12587 35977 13005 35994
rect 12587 35913 12588 35977
rect 12652 35913 12676 35977
rect 12740 35913 12764 35977
rect 12828 35913 12852 35977
rect 12916 35913 12940 35977
rect 13004 35913 13005 35977
rect 12587 35851 13005 35913
tri 13005 35851 13156 36002 sw
rect 12587 35787 12598 35851
rect 12662 35787 12682 35851
rect 12746 35787 12766 35851
rect 12830 35787 12850 35851
rect 12914 35787 12933 35851
rect 12997 35787 13016 35851
rect 13080 35787 13099 35851
rect 13163 35787 13182 35851
rect 13246 35787 13264 35851
rect 12587 35767 13264 35787
rect 12587 35703 12598 35767
rect 12662 35703 12682 35767
rect 12746 35703 12766 35767
rect 12830 35703 12850 35767
rect 12914 35703 12933 35767
rect 12997 35703 13016 35767
rect 13080 35703 13099 35767
rect 13163 35703 13182 35767
rect 13246 35703 13264 35767
rect 12587 35683 13264 35703
rect 12587 35619 12598 35683
rect 12662 35619 12682 35683
rect 12746 35619 12766 35683
rect 12830 35619 12850 35683
rect 12914 35619 12933 35683
rect 12997 35619 13016 35683
rect 13080 35619 13099 35683
rect 13163 35619 13182 35683
rect 13246 35619 13264 35683
rect 12587 35599 13264 35619
rect 12587 35535 12598 35599
rect 12662 35535 12682 35599
rect 12746 35535 12766 35599
rect 12830 35535 12850 35599
rect 12914 35535 12933 35599
rect 12997 35535 13016 35599
rect 13080 35535 13099 35599
rect 13163 35535 13182 35599
rect 13246 35535 13264 35599
rect 12587 35515 13264 35535
rect 12587 35451 12598 35515
rect 12662 35451 12682 35515
rect 12746 35451 12766 35515
rect 12830 35451 12850 35515
rect 12914 35451 12933 35515
rect 12997 35451 13016 35515
rect 13080 35451 13099 35515
rect 13163 35451 13182 35515
rect 13246 35451 13264 35515
rect 12587 35431 13264 35451
rect 12587 35367 12598 35431
rect 12662 35367 12682 35431
rect 12746 35367 12766 35431
rect 12830 35367 12850 35431
rect 12914 35367 12933 35431
rect 12997 35367 13016 35431
rect 13080 35367 13099 35431
rect 13163 35367 13182 35431
rect 13246 35367 13264 35431
rect 12587 32613 13264 35367
tri 13957 33764 14399 34206 se
rect 14399 33764 15371 39747
rect 12587 32557 12598 32613
rect 12654 32557 12685 32613
rect 12741 32557 12772 32613
rect 12828 32557 12859 32613
rect 12915 32557 12945 32613
rect 13001 32557 13031 32613
rect 13087 32557 13117 32613
rect 13173 32557 13203 32613
rect 13259 32557 13264 32613
rect 12587 32531 13264 32557
rect 12587 32475 12598 32531
rect 12654 32475 12685 32531
rect 12741 32475 12772 32531
rect 12828 32475 12859 32531
rect 12915 32475 12945 32531
rect 13001 32475 13031 32531
rect 13087 32475 13117 32531
rect 13173 32475 13203 32531
rect 13259 32475 13264 32531
rect 12587 32449 13264 32475
rect 12587 32393 12598 32449
rect 12654 32393 12685 32449
rect 12741 32393 12772 32449
rect 12828 32393 12859 32449
rect 12915 32393 12945 32449
rect 13001 32393 13031 32449
rect 13087 32393 13117 32449
rect 13173 32393 13203 32449
rect 13259 32393 13264 32449
rect 12587 32367 13264 32393
rect 12587 32311 12598 32367
rect 12654 32311 12685 32367
rect 12741 32311 12772 32367
rect 12828 32311 12859 32367
rect 12915 32311 12945 32367
rect 13001 32311 13031 32367
rect 13087 32311 13117 32367
rect 13173 32311 13203 32367
rect 13259 32311 13264 32367
rect 12587 32285 13264 32311
rect 12587 32229 12598 32285
rect 12654 32229 12685 32285
rect 12741 32229 12772 32285
rect 12828 32229 12859 32285
rect 12915 32229 12945 32285
rect 13001 32229 13031 32285
rect 13087 32229 13117 32285
rect 13173 32229 13203 32285
rect 13259 32229 13264 32285
rect 12587 32203 13264 32229
rect 12587 32147 12598 32203
rect 12654 32147 12685 32203
rect 12741 32147 12772 32203
rect 12828 32147 12859 32203
rect 12915 32147 12945 32203
rect 13001 32147 13031 32203
rect 13087 32147 13117 32203
rect 13173 32147 13203 32203
rect 13259 32147 13264 32203
rect 12587 32121 13264 32147
rect 12587 32065 12598 32121
rect 12654 32065 12685 32121
rect 12741 32065 12772 32121
rect 12828 32065 12859 32121
rect 12915 32065 12945 32121
rect 13001 32065 13031 32121
rect 13087 32065 13117 32121
rect 13173 32065 13203 32121
rect 13259 32065 13264 32121
rect 12587 32039 13264 32065
rect 12587 31983 12598 32039
rect 12654 31983 12685 32039
rect 12741 31983 12772 32039
rect 12828 31983 12859 32039
rect 12915 31983 12945 32039
rect 13001 31983 13031 32039
rect 13087 31983 13117 32039
rect 13173 31983 13203 32039
rect 13259 31983 13264 32039
rect 12587 31957 13264 31983
rect 12587 31901 12598 31957
rect 12654 31901 12685 31957
rect 12741 31901 12772 31957
rect 12828 31901 12859 31957
rect 12915 31901 12945 31957
rect 13001 31901 13031 31957
rect 13087 31901 13117 31957
rect 13173 31901 13203 31957
rect 13259 31901 13264 31957
rect 12587 31875 13264 31901
rect 12587 31819 12598 31875
rect 12654 31819 12685 31875
rect 12741 31819 12772 31875
rect 12828 31819 12859 31875
rect 12915 31819 12945 31875
rect 13001 31819 13031 31875
rect 13087 31819 13117 31875
rect 13173 31819 13203 31875
rect 13259 31819 13264 31875
rect 12587 31793 13264 31819
rect 12587 31737 12598 31793
rect 12654 31737 12685 31793
rect 12741 31737 12772 31793
rect 12828 31737 12859 31793
rect 12915 31737 12945 31793
rect 13001 31737 13031 31793
rect 13087 31737 13117 31793
rect 13173 31737 13203 31793
rect 13259 31737 13264 31793
rect 12587 31711 13264 31737
rect 12587 31655 12598 31711
rect 12654 31655 12685 31711
rect 12741 31655 12772 31711
rect 12828 31655 12859 31711
rect 12915 31655 12945 31711
rect 13001 31655 13031 31711
rect 13087 31655 13117 31711
rect 13173 31655 13203 31711
rect 13259 31655 13264 31711
rect 12587 31629 13264 31655
rect 12587 31573 12598 31629
rect 12654 31573 12685 31629
rect 12741 31573 12772 31629
rect 12828 31573 12859 31629
rect 12915 31573 12945 31629
rect 13001 31573 13031 31629
rect 13087 31573 13117 31629
rect 13173 31573 13203 31629
rect 13259 31573 13264 31629
rect 12587 31547 13264 31573
rect 12587 31491 12598 31547
rect 12654 31491 12685 31547
rect 12741 31491 12772 31547
rect 12828 31491 12859 31547
rect 12915 31491 12945 31547
rect 13001 31491 13031 31547
rect 13087 31491 13117 31547
rect 13173 31491 13203 31547
rect 13259 31491 13264 31547
rect 12587 31478 13264 31491
tri 13579 33386 13957 33764 se
rect 13957 33386 14391 33764
rect 5777 31160 13085 31173
rect 5777 31104 6182 31160
rect 6238 31104 6263 31160
rect 6319 31104 6344 31160
rect 6400 31104 6425 31160
rect 6481 31104 6506 31160
rect 6562 31104 6587 31160
rect 6643 31104 6668 31160
rect 6724 31104 6749 31160
rect 6805 31104 6830 31160
rect 6886 31104 6911 31160
rect 6967 31104 6992 31160
rect 7048 31104 7073 31160
rect 7129 31104 7154 31160
rect 7210 31104 7235 31160
rect 7291 31104 7316 31160
rect 7372 31104 7397 31160
rect 7453 31104 7478 31160
rect 7534 31104 7559 31160
rect 7615 31104 7640 31160
rect 7696 31104 7721 31160
rect 7777 31104 7802 31160
rect 7858 31104 7883 31160
rect 7939 31104 7964 31160
rect 8020 31104 8045 31160
rect 8101 31104 8126 31160
rect 8182 31104 8207 31160
rect 8263 31104 8288 31160
rect 8344 31104 8369 31160
rect 8425 31104 8450 31160
rect 8506 31104 8531 31160
rect 8587 31104 8612 31160
rect 8668 31104 8693 31160
rect 8749 31104 8774 31160
rect 8830 31104 8855 31160
rect 8911 31104 8936 31160
rect 8992 31104 9017 31160
rect 9073 31104 9098 31160
rect 9154 31104 9179 31160
rect 9235 31104 9260 31160
rect 9316 31104 9340 31160
rect 9396 31104 9420 31160
rect 9476 31104 9500 31160
rect 9556 31104 9580 31160
rect 9636 31104 9660 31160
rect 9716 31104 9740 31160
rect 9796 31104 9820 31160
rect 9876 31104 9900 31160
rect 9956 31104 9980 31160
rect 10036 31104 10060 31160
rect 10116 31104 10140 31160
rect 10196 31104 10220 31160
rect 10276 31104 10300 31160
rect 10356 31104 10380 31160
rect 10436 31104 10460 31160
rect 10516 31104 10540 31160
rect 10596 31104 10620 31160
rect 10676 31104 10700 31160
rect 10756 31104 10780 31160
rect 10836 31104 10860 31160
rect 10916 31104 10940 31160
rect 10996 31104 11020 31160
rect 11076 31104 11100 31160
rect 11156 31104 11180 31160
rect 11236 31104 11260 31160
rect 11316 31104 11340 31160
rect 11396 31104 11420 31160
rect 11476 31104 11500 31160
rect 11556 31104 11580 31160
rect 11636 31104 11660 31160
rect 11716 31104 11740 31160
rect 11796 31104 11820 31160
rect 11876 31104 11900 31160
rect 11956 31104 11980 31160
rect 12036 31104 12060 31160
rect 12116 31104 12140 31160
rect 12196 31104 12220 31160
rect 12276 31104 12300 31160
rect 12356 31104 12380 31160
rect 12436 31104 12460 31160
rect 12516 31104 12540 31160
rect 12596 31104 12620 31160
rect 12676 31104 12700 31160
rect 12756 31104 12780 31160
rect 12836 31104 12860 31160
rect 12916 31104 12940 31160
rect 12996 31104 13020 31160
rect 13076 31104 13085 31160
rect 5777 31078 13085 31104
rect 5777 31022 6182 31078
rect 6238 31022 6263 31078
rect 6319 31022 6344 31078
rect 6400 31022 6425 31078
rect 6481 31022 6506 31078
rect 6562 31022 6587 31078
rect 6643 31022 6668 31078
rect 6724 31022 6749 31078
rect 6805 31022 6830 31078
rect 6886 31022 6911 31078
rect 6967 31022 6992 31078
rect 7048 31022 7073 31078
rect 7129 31022 7154 31078
rect 7210 31022 7235 31078
rect 7291 31022 7316 31078
rect 7372 31022 7397 31078
rect 7453 31022 7478 31078
rect 7534 31022 7559 31078
rect 7615 31022 7640 31078
rect 7696 31022 7721 31078
rect 7777 31022 7802 31078
rect 7858 31022 7883 31078
rect 7939 31022 7964 31078
rect 8020 31022 8045 31078
rect 8101 31022 8126 31078
rect 8182 31022 8207 31078
rect 8263 31022 8288 31078
rect 8344 31022 8369 31078
rect 8425 31022 8450 31078
rect 8506 31022 8531 31078
rect 8587 31022 8612 31078
rect 8668 31022 8693 31078
rect 8749 31022 8774 31078
rect 8830 31022 8855 31078
rect 8911 31022 8936 31078
rect 8992 31022 9017 31078
rect 9073 31022 9098 31078
rect 9154 31022 9179 31078
rect 9235 31022 9260 31078
rect 9316 31022 9340 31078
rect 9396 31022 9420 31078
rect 9476 31022 9500 31078
rect 9556 31022 9580 31078
rect 9636 31022 9660 31078
rect 9716 31022 9740 31078
rect 9796 31022 9820 31078
rect 9876 31022 9900 31078
rect 9956 31022 9980 31078
rect 10036 31022 10060 31078
rect 10116 31022 10140 31078
rect 10196 31022 10220 31078
rect 10276 31022 10300 31078
rect 10356 31022 10380 31078
rect 10436 31022 10460 31078
rect 10516 31022 10540 31078
rect 10596 31022 10620 31078
rect 10676 31022 10700 31078
rect 10756 31022 10780 31078
rect 10836 31022 10860 31078
rect 10916 31022 10940 31078
rect 10996 31022 11020 31078
rect 11076 31022 11100 31078
rect 11156 31022 11180 31078
rect 11236 31022 11260 31078
rect 11316 31022 11340 31078
rect 11396 31022 11420 31078
rect 11476 31022 11500 31078
rect 11556 31022 11580 31078
rect 11636 31022 11660 31078
rect 11716 31022 11740 31078
rect 11796 31022 11820 31078
rect 11876 31022 11900 31078
rect 11956 31022 11980 31078
rect 12036 31022 12060 31078
rect 12116 31022 12140 31078
rect 12196 31022 12220 31078
rect 12276 31022 12300 31078
rect 12356 31022 12380 31078
rect 12436 31022 12460 31078
rect 12516 31022 12540 31078
rect 12596 31022 12620 31078
rect 12676 31022 12700 31078
rect 12756 31022 12780 31078
rect 12836 31022 12860 31078
rect 12916 31022 12940 31078
rect 12996 31022 13020 31078
rect 13076 31022 13085 31078
rect 5777 30996 13085 31022
rect 5777 30993 6182 30996
rect 5777 30937 5803 30993
rect 5859 30937 5895 30993
rect 5951 30937 5987 30993
rect 6043 30937 6079 30993
rect 6135 30940 6182 30993
rect 6238 30940 6263 30996
rect 6319 30940 6344 30996
rect 6400 30940 6425 30996
rect 6481 30940 6506 30996
rect 6562 30940 6587 30996
rect 6643 30940 6668 30996
rect 6724 30940 6749 30996
rect 6805 30940 6830 30996
rect 6886 30940 6911 30996
rect 6967 30940 6992 30996
rect 7048 30940 7073 30996
rect 7129 30940 7154 30996
rect 7210 30940 7235 30996
rect 7291 30940 7316 30996
rect 7372 30940 7397 30996
rect 7453 30940 7478 30996
rect 7534 30940 7559 30996
rect 7615 30940 7640 30996
rect 7696 30940 7721 30996
rect 7777 30940 7802 30996
rect 7858 30940 7883 30996
rect 7939 30940 7964 30996
rect 8020 30940 8045 30996
rect 8101 30940 8126 30996
rect 8182 30940 8207 30996
rect 8263 30940 8288 30996
rect 8344 30940 8369 30996
rect 8425 30940 8450 30996
rect 8506 30940 8531 30996
rect 8587 30940 8612 30996
rect 8668 30940 8693 30996
rect 8749 30940 8774 30996
rect 8830 30940 8855 30996
rect 8911 30940 8936 30996
rect 8992 30940 9017 30996
rect 9073 30940 9098 30996
rect 9154 30940 9179 30996
rect 9235 30940 9260 30996
rect 9316 30940 9340 30996
rect 9396 30940 9420 30996
rect 9476 30940 9500 30996
rect 9556 30940 9580 30996
rect 9636 30940 9660 30996
rect 9716 30940 9740 30996
rect 9796 30940 9820 30996
rect 9876 30940 9900 30996
rect 9956 30940 9980 30996
rect 10036 30940 10060 30996
rect 10116 30940 10140 30996
rect 10196 30940 10220 30996
rect 10276 30940 10300 30996
rect 10356 30940 10380 30996
rect 10436 30940 10460 30996
rect 10516 30940 10540 30996
rect 10596 30940 10620 30996
rect 10676 30940 10700 30996
rect 10756 30940 10780 30996
rect 10836 30940 10860 30996
rect 10916 30940 10940 30996
rect 10996 30940 11020 30996
rect 11076 30940 11100 30996
rect 11156 30940 11180 30996
rect 11236 30940 11260 30996
rect 11316 30940 11340 30996
rect 11396 30940 11420 30996
rect 11476 30940 11500 30996
rect 11556 30940 11580 30996
rect 11636 30940 11660 30996
rect 11716 30940 11740 30996
rect 11796 30940 11820 30996
rect 11876 30940 11900 30996
rect 11956 30940 11980 30996
rect 12036 30940 12060 30996
rect 12116 30940 12140 30996
rect 12196 30940 12220 30996
rect 12276 30940 12300 30996
rect 12356 30940 12380 30996
rect 12436 30940 12460 30996
rect 12516 30940 12540 30996
rect 12596 30940 12620 30996
rect 12676 30940 12700 30996
rect 12756 30940 12780 30996
rect 12836 30940 12860 30996
rect 12916 30940 12940 30996
rect 12996 30940 13020 30996
rect 13076 30940 13085 30996
rect 6135 30937 13085 30940
rect 5777 30914 13085 30937
rect 5777 30910 6182 30914
rect 5777 30854 5803 30910
rect 5859 30854 5895 30910
rect 5951 30854 5987 30910
rect 6043 30854 6079 30910
rect 6135 30858 6182 30910
rect 6238 30858 6263 30914
rect 6319 30858 6344 30914
rect 6400 30858 6425 30914
rect 6481 30858 6506 30914
rect 6562 30858 6587 30914
rect 6643 30858 6668 30914
rect 6724 30858 6749 30914
rect 6805 30858 6830 30914
rect 6886 30858 6911 30914
rect 6967 30858 6992 30914
rect 7048 30858 7073 30914
rect 7129 30858 7154 30914
rect 7210 30858 7235 30914
rect 7291 30858 7316 30914
rect 7372 30858 7397 30914
rect 7453 30858 7478 30914
rect 7534 30858 7559 30914
rect 7615 30858 7640 30914
rect 7696 30858 7721 30914
rect 7777 30858 7802 30914
rect 7858 30858 7883 30914
rect 7939 30858 7964 30914
rect 8020 30858 8045 30914
rect 8101 30858 8126 30914
rect 8182 30858 8207 30914
rect 8263 30858 8288 30914
rect 8344 30858 8369 30914
rect 8425 30858 8450 30914
rect 8506 30858 8531 30914
rect 8587 30858 8612 30914
rect 8668 30858 8693 30914
rect 8749 30858 8774 30914
rect 8830 30858 8855 30914
rect 8911 30858 8936 30914
rect 8992 30858 9017 30914
rect 9073 30858 9098 30914
rect 9154 30858 9179 30914
rect 9235 30858 9260 30914
rect 9316 30858 9340 30914
rect 9396 30858 9420 30914
rect 9476 30858 9500 30914
rect 9556 30858 9580 30914
rect 9636 30858 9660 30914
rect 9716 30858 9740 30914
rect 9796 30858 9820 30914
rect 9876 30858 9900 30914
rect 9956 30858 9980 30914
rect 10036 30858 10060 30914
rect 10116 30858 10140 30914
rect 10196 30858 10220 30914
rect 10276 30858 10300 30914
rect 10356 30858 10380 30914
rect 10436 30858 10460 30914
rect 10516 30858 10540 30914
rect 10596 30858 10620 30914
rect 10676 30858 10700 30914
rect 10756 30858 10780 30914
rect 10836 30858 10860 30914
rect 10916 30858 10940 30914
rect 10996 30858 11020 30914
rect 11076 30858 11100 30914
rect 11156 30858 11180 30914
rect 11236 30858 11260 30914
rect 11316 30858 11340 30914
rect 11396 30858 11420 30914
rect 11476 30858 11500 30914
rect 11556 30858 11580 30914
rect 11636 30858 11660 30914
rect 11716 30858 11740 30914
rect 11796 30858 11820 30914
rect 11876 30858 11900 30914
rect 11956 30858 11980 30914
rect 12036 30858 12060 30914
rect 12116 30858 12140 30914
rect 12196 30858 12220 30914
rect 12276 30858 12300 30914
rect 12356 30858 12380 30914
rect 12436 30858 12460 30914
rect 12516 30858 12540 30914
rect 12596 30858 12620 30914
rect 12676 30858 12700 30914
rect 12756 30858 12780 30914
rect 12836 30858 12860 30914
rect 12916 30858 12940 30914
rect 12996 30858 13020 30914
rect 13076 30858 13085 30914
rect 6135 30854 13085 30858
rect 5777 30832 13085 30854
rect 5777 30827 6182 30832
rect 5777 30771 5803 30827
rect 5859 30771 5895 30827
rect 5951 30771 5987 30827
rect 6043 30771 6079 30827
rect 6135 30776 6182 30827
rect 6238 30776 6263 30832
rect 6319 30776 6344 30832
rect 6400 30776 6425 30832
rect 6481 30776 6506 30832
rect 6562 30776 6587 30832
rect 6643 30776 6668 30832
rect 6724 30776 6749 30832
rect 6805 30776 6830 30832
rect 6886 30776 6911 30832
rect 6967 30776 6992 30832
rect 7048 30776 7073 30832
rect 7129 30776 7154 30832
rect 7210 30776 7235 30832
rect 7291 30776 7316 30832
rect 7372 30776 7397 30832
rect 7453 30776 7478 30832
rect 7534 30776 7559 30832
rect 7615 30776 7640 30832
rect 7696 30776 7721 30832
rect 7777 30776 7802 30832
rect 7858 30776 7883 30832
rect 7939 30776 7964 30832
rect 8020 30776 8045 30832
rect 8101 30776 8126 30832
rect 8182 30776 8207 30832
rect 8263 30776 8288 30832
rect 8344 30776 8369 30832
rect 8425 30776 8450 30832
rect 8506 30776 8531 30832
rect 8587 30776 8612 30832
rect 8668 30776 8693 30832
rect 8749 30776 8774 30832
rect 8830 30776 8855 30832
rect 8911 30776 8936 30832
rect 8992 30776 9017 30832
rect 9073 30776 9098 30832
rect 9154 30776 9179 30832
rect 9235 30776 9260 30832
rect 9316 30776 9340 30832
rect 9396 30776 9420 30832
rect 9476 30776 9500 30832
rect 9556 30776 9580 30832
rect 9636 30776 9660 30832
rect 9716 30776 9740 30832
rect 9796 30776 9820 30832
rect 9876 30776 9900 30832
rect 9956 30776 9980 30832
rect 10036 30776 10060 30832
rect 10116 30776 10140 30832
rect 10196 30776 10220 30832
rect 10276 30776 10300 30832
rect 10356 30776 10380 30832
rect 10436 30776 10460 30832
rect 10516 30776 10540 30832
rect 10596 30776 10620 30832
rect 10676 30776 10700 30832
rect 10756 30776 10780 30832
rect 10836 30776 10860 30832
rect 10916 30776 10940 30832
rect 10996 30776 11020 30832
rect 11076 30776 11100 30832
rect 11156 30776 11180 30832
rect 11236 30776 11260 30832
rect 11316 30776 11340 30832
rect 11396 30776 11420 30832
rect 11476 30776 11500 30832
rect 11556 30776 11580 30832
rect 11636 30776 11660 30832
rect 11716 30776 11740 30832
rect 11796 30776 11820 30832
rect 11876 30776 11900 30832
rect 11956 30776 11980 30832
rect 12036 30776 12060 30832
rect 12116 30776 12140 30832
rect 12196 30776 12220 30832
rect 12276 30776 12300 30832
rect 12356 30776 12380 30832
rect 12436 30776 12460 30832
rect 12516 30776 12540 30832
rect 12596 30776 12620 30832
rect 12676 30776 12700 30832
rect 12756 30776 12780 30832
rect 12836 30776 12860 30832
rect 12916 30776 12940 30832
rect 12996 30776 13020 30832
rect 13076 30776 13085 30832
rect 6135 30771 13085 30776
rect 5777 30750 13085 30771
rect 5777 30744 6182 30750
rect 5777 30688 5803 30744
rect 5859 30688 5895 30744
rect 5951 30688 5987 30744
rect 6043 30688 6079 30744
rect 6135 30694 6182 30744
rect 6238 30694 6263 30750
rect 6319 30694 6344 30750
rect 6400 30694 6425 30750
rect 6481 30694 6506 30750
rect 6562 30694 6587 30750
rect 6643 30694 6668 30750
rect 6724 30694 6749 30750
rect 6805 30694 6830 30750
rect 6886 30694 6911 30750
rect 6967 30694 6992 30750
rect 7048 30694 7073 30750
rect 7129 30694 7154 30750
rect 7210 30694 7235 30750
rect 7291 30694 7316 30750
rect 7372 30694 7397 30750
rect 7453 30694 7478 30750
rect 7534 30694 7559 30750
rect 7615 30694 7640 30750
rect 7696 30694 7721 30750
rect 7777 30694 7802 30750
rect 7858 30694 7883 30750
rect 7939 30694 7964 30750
rect 8020 30694 8045 30750
rect 8101 30694 8126 30750
rect 8182 30694 8207 30750
rect 8263 30694 8288 30750
rect 8344 30694 8369 30750
rect 8425 30694 8450 30750
rect 8506 30694 8531 30750
rect 8587 30694 8612 30750
rect 8668 30694 8693 30750
rect 8749 30694 8774 30750
rect 8830 30694 8855 30750
rect 8911 30694 8936 30750
rect 8992 30694 9017 30750
rect 9073 30694 9098 30750
rect 9154 30694 9179 30750
rect 9235 30694 9260 30750
rect 9316 30694 9340 30750
rect 9396 30694 9420 30750
rect 9476 30694 9500 30750
rect 9556 30694 9580 30750
rect 9636 30694 9660 30750
rect 9716 30694 9740 30750
rect 9796 30694 9820 30750
rect 9876 30694 9900 30750
rect 9956 30694 9980 30750
rect 10036 30694 10060 30750
rect 10116 30694 10140 30750
rect 10196 30694 10220 30750
rect 10276 30694 10300 30750
rect 10356 30694 10380 30750
rect 10436 30694 10460 30750
rect 10516 30694 10540 30750
rect 10596 30694 10620 30750
rect 10676 30694 10700 30750
rect 10756 30694 10780 30750
rect 10836 30694 10860 30750
rect 10916 30694 10940 30750
rect 10996 30694 11020 30750
rect 11076 30694 11100 30750
rect 11156 30694 11180 30750
rect 11236 30694 11260 30750
rect 11316 30694 11340 30750
rect 11396 30694 11420 30750
rect 11476 30694 11500 30750
rect 11556 30694 11580 30750
rect 11636 30694 11660 30750
rect 11716 30694 11740 30750
rect 11796 30694 11820 30750
rect 11876 30694 11900 30750
rect 11956 30694 11980 30750
rect 12036 30694 12060 30750
rect 12116 30694 12140 30750
rect 12196 30694 12220 30750
rect 12276 30694 12300 30750
rect 12356 30694 12380 30750
rect 12436 30694 12460 30750
rect 12516 30694 12540 30750
rect 12596 30694 12620 30750
rect 12676 30694 12700 30750
rect 12756 30694 12780 30750
rect 12836 30694 12860 30750
rect 12916 30694 12940 30750
rect 12996 30694 13020 30750
rect 13076 30694 13085 30750
rect 6135 30688 13085 30694
rect 5777 30668 13085 30688
rect 5777 30661 6182 30668
rect 5777 30605 5803 30661
rect 5859 30605 5895 30661
rect 5951 30605 5987 30661
rect 6043 30605 6079 30661
rect 6135 30612 6182 30661
rect 6238 30612 6263 30668
rect 6319 30612 6344 30668
rect 6400 30612 6425 30668
rect 6481 30612 6506 30668
rect 6562 30612 6587 30668
rect 6643 30612 6668 30668
rect 6724 30612 6749 30668
rect 6805 30612 6830 30668
rect 6886 30612 6911 30668
rect 6967 30612 6992 30668
rect 7048 30612 7073 30668
rect 7129 30612 7154 30668
rect 7210 30612 7235 30668
rect 7291 30612 7316 30668
rect 7372 30612 7397 30668
rect 7453 30612 7478 30668
rect 7534 30612 7559 30668
rect 7615 30612 7640 30668
rect 7696 30612 7721 30668
rect 7777 30612 7802 30668
rect 7858 30612 7883 30668
rect 7939 30612 7964 30668
rect 8020 30612 8045 30668
rect 8101 30612 8126 30668
rect 8182 30612 8207 30668
rect 8263 30612 8288 30668
rect 8344 30612 8369 30668
rect 8425 30612 8450 30668
rect 8506 30612 8531 30668
rect 8587 30612 8612 30668
rect 8668 30612 8693 30668
rect 8749 30612 8774 30668
rect 8830 30612 8855 30668
rect 8911 30612 8936 30668
rect 8992 30612 9017 30668
rect 9073 30612 9098 30668
rect 9154 30612 9179 30668
rect 9235 30612 9260 30668
rect 9316 30612 9340 30668
rect 9396 30612 9420 30668
rect 9476 30612 9500 30668
rect 9556 30612 9580 30668
rect 9636 30612 9660 30668
rect 9716 30612 9740 30668
rect 9796 30612 9820 30668
rect 9876 30612 9900 30668
rect 9956 30612 9980 30668
rect 10036 30612 10060 30668
rect 10116 30612 10140 30668
rect 10196 30612 10220 30668
rect 10276 30612 10300 30668
rect 10356 30612 10380 30668
rect 10436 30612 10460 30668
rect 10516 30612 10540 30668
rect 10596 30612 10620 30668
rect 10676 30612 10700 30668
rect 10756 30612 10780 30668
rect 10836 30612 10860 30668
rect 10916 30612 10940 30668
rect 10996 30612 11020 30668
rect 11076 30612 11100 30668
rect 11156 30612 11180 30668
rect 11236 30612 11260 30668
rect 11316 30612 11340 30668
rect 11396 30612 11420 30668
rect 11476 30612 11500 30668
rect 11556 30612 11580 30668
rect 11636 30612 11660 30668
rect 11716 30612 11740 30668
rect 11796 30612 11820 30668
rect 11876 30612 11900 30668
rect 11956 30612 11980 30668
rect 12036 30612 12060 30668
rect 12116 30612 12140 30668
rect 12196 30612 12220 30668
rect 12276 30612 12300 30668
rect 12356 30612 12380 30668
rect 12436 30612 12460 30668
rect 12516 30612 12540 30668
rect 12596 30612 12620 30668
rect 12676 30612 12700 30668
rect 12756 30612 12780 30668
rect 12836 30612 12860 30668
rect 12916 30612 12940 30668
rect 12996 30612 13020 30668
rect 13076 30612 13085 30668
rect 6135 30605 13085 30612
rect 5777 30586 13085 30605
rect 5777 30578 6182 30586
rect 5777 30522 5803 30578
rect 5859 30522 5895 30578
rect 5951 30522 5987 30578
rect 6043 30522 6079 30578
rect 6135 30530 6182 30578
rect 6238 30530 6263 30586
rect 6319 30530 6344 30586
rect 6400 30530 6425 30586
rect 6481 30530 6506 30586
rect 6562 30530 6587 30586
rect 6643 30530 6668 30586
rect 6724 30530 6749 30586
rect 6805 30530 6830 30586
rect 6886 30530 6911 30586
rect 6967 30530 6992 30586
rect 7048 30530 7073 30586
rect 7129 30530 7154 30586
rect 7210 30530 7235 30586
rect 7291 30530 7316 30586
rect 7372 30530 7397 30586
rect 7453 30530 7478 30586
rect 7534 30530 7559 30586
rect 7615 30530 7640 30586
rect 7696 30530 7721 30586
rect 7777 30530 7802 30586
rect 7858 30530 7883 30586
rect 7939 30530 7964 30586
rect 8020 30530 8045 30586
rect 8101 30530 8126 30586
rect 8182 30530 8207 30586
rect 8263 30530 8288 30586
rect 8344 30530 8369 30586
rect 8425 30530 8450 30586
rect 8506 30530 8531 30586
rect 8587 30530 8612 30586
rect 8668 30530 8693 30586
rect 8749 30530 8774 30586
rect 8830 30530 8855 30586
rect 8911 30530 8936 30586
rect 8992 30530 9017 30586
rect 9073 30530 9098 30586
rect 9154 30530 9179 30586
rect 9235 30530 9260 30586
rect 9316 30530 9340 30586
rect 9396 30530 9420 30586
rect 9476 30530 9500 30586
rect 9556 30530 9580 30586
rect 9636 30530 9660 30586
rect 9716 30530 9740 30586
rect 9796 30530 9820 30586
rect 9876 30530 9900 30586
rect 9956 30530 9980 30586
rect 10036 30530 10060 30586
rect 10116 30530 10140 30586
rect 10196 30530 10220 30586
rect 10276 30530 10300 30586
rect 10356 30530 10380 30586
rect 10436 30530 10460 30586
rect 10516 30530 10540 30586
rect 10596 30530 10620 30586
rect 10676 30530 10700 30586
rect 10756 30530 10780 30586
rect 10836 30530 10860 30586
rect 10916 30530 10940 30586
rect 10996 30530 11020 30586
rect 11076 30530 11100 30586
rect 11156 30530 11180 30586
rect 11236 30530 11260 30586
rect 11316 30530 11340 30586
rect 11396 30530 11420 30586
rect 11476 30530 11500 30586
rect 11556 30530 11580 30586
rect 11636 30530 11660 30586
rect 11716 30530 11740 30586
rect 11796 30530 11820 30586
rect 11876 30530 11900 30586
rect 11956 30530 11980 30586
rect 12036 30530 12060 30586
rect 12116 30530 12140 30586
rect 12196 30530 12220 30586
rect 12276 30530 12300 30586
rect 12356 30530 12380 30586
rect 12436 30530 12460 30586
rect 12516 30530 12540 30586
rect 12596 30530 12620 30586
rect 12676 30530 12700 30586
rect 12756 30530 12780 30586
rect 12836 30530 12860 30586
rect 12916 30530 12940 30586
rect 12996 30530 13020 30586
rect 13076 30530 13085 30586
rect 6135 30522 13085 30530
rect 5777 30504 13085 30522
rect 5777 30496 6182 30504
rect 5777 30440 5803 30496
rect 5859 30440 5895 30496
rect 5951 30440 5987 30496
rect 6043 30440 6079 30496
rect 6135 30448 6182 30496
rect 6238 30448 6263 30504
rect 6319 30448 6344 30504
rect 6400 30448 6425 30504
rect 6481 30448 6506 30504
rect 6562 30448 6587 30504
rect 6643 30448 6668 30504
rect 6724 30448 6749 30504
rect 6805 30448 6830 30504
rect 6886 30448 6911 30504
rect 6967 30448 6992 30504
rect 7048 30448 7073 30504
rect 7129 30448 7154 30504
rect 7210 30448 7235 30504
rect 7291 30448 7316 30504
rect 7372 30448 7397 30504
rect 7453 30448 7478 30504
rect 7534 30448 7559 30504
rect 7615 30448 7640 30504
rect 7696 30448 7721 30504
rect 7777 30448 7802 30504
rect 7858 30448 7883 30504
rect 7939 30448 7964 30504
rect 8020 30448 8045 30504
rect 8101 30448 8126 30504
rect 8182 30448 8207 30504
rect 8263 30448 8288 30504
rect 8344 30448 8369 30504
rect 8425 30448 8450 30504
rect 8506 30448 8531 30504
rect 8587 30448 8612 30504
rect 8668 30448 8693 30504
rect 8749 30448 8774 30504
rect 8830 30448 8855 30504
rect 8911 30448 8936 30504
rect 8992 30448 9017 30504
rect 9073 30448 9098 30504
rect 9154 30448 9179 30504
rect 9235 30448 9260 30504
rect 9316 30448 9340 30504
rect 9396 30448 9420 30504
rect 9476 30448 9500 30504
rect 9556 30448 9580 30504
rect 9636 30448 9660 30504
rect 9716 30448 9740 30504
rect 9796 30448 9820 30504
rect 9876 30448 9900 30504
rect 9956 30448 9980 30504
rect 10036 30448 10060 30504
rect 10116 30448 10140 30504
rect 10196 30448 10220 30504
rect 10276 30448 10300 30504
rect 10356 30448 10380 30504
rect 10436 30448 10460 30504
rect 10516 30448 10540 30504
rect 10596 30448 10620 30504
rect 10676 30448 10700 30504
rect 10756 30448 10780 30504
rect 10836 30448 10860 30504
rect 10916 30448 10940 30504
rect 10996 30448 11020 30504
rect 11076 30448 11100 30504
rect 11156 30448 11180 30504
rect 11236 30448 11260 30504
rect 11316 30448 11340 30504
rect 11396 30448 11420 30504
rect 11476 30448 11500 30504
rect 11556 30448 11580 30504
rect 11636 30448 11660 30504
rect 11716 30448 11740 30504
rect 11796 30448 11820 30504
rect 11876 30448 11900 30504
rect 11956 30448 11980 30504
rect 12036 30448 12060 30504
rect 12116 30448 12140 30504
rect 12196 30448 12220 30504
rect 12276 30448 12300 30504
rect 12356 30448 12380 30504
rect 12436 30448 12460 30504
rect 12516 30448 12540 30504
rect 12596 30448 12620 30504
rect 12676 30448 12700 30504
rect 12756 30448 12780 30504
rect 12836 30448 12860 30504
rect 12916 30448 12940 30504
rect 12996 30448 13020 30504
rect 13076 30448 13085 30504
rect 6135 30440 13085 30448
rect 5777 30422 13085 30440
rect 5777 30414 6182 30422
rect 5777 30358 5803 30414
rect 5859 30358 5895 30414
rect 5951 30358 5987 30414
rect 6043 30358 6079 30414
rect 6135 30366 6182 30414
rect 6238 30366 6263 30422
rect 6319 30366 6344 30422
rect 6400 30366 6425 30422
rect 6481 30366 6506 30422
rect 6562 30366 6587 30422
rect 6643 30366 6668 30422
rect 6724 30366 6749 30422
rect 6805 30366 6830 30422
rect 6886 30366 6911 30422
rect 6967 30366 6992 30422
rect 7048 30366 7073 30422
rect 7129 30366 7154 30422
rect 7210 30366 7235 30422
rect 7291 30366 7316 30422
rect 7372 30366 7397 30422
rect 7453 30366 7478 30422
rect 7534 30366 7559 30422
rect 7615 30366 7640 30422
rect 7696 30366 7721 30422
rect 7777 30366 7802 30422
rect 7858 30366 7883 30422
rect 7939 30366 7964 30422
rect 8020 30366 8045 30422
rect 8101 30366 8126 30422
rect 8182 30366 8207 30422
rect 8263 30366 8288 30422
rect 8344 30366 8369 30422
rect 8425 30366 8450 30422
rect 8506 30366 8531 30422
rect 8587 30366 8612 30422
rect 8668 30366 8693 30422
rect 8749 30366 8774 30422
rect 8830 30366 8855 30422
rect 8911 30366 8936 30422
rect 8992 30366 9017 30422
rect 9073 30366 9098 30422
rect 9154 30366 9179 30422
rect 9235 30366 9260 30422
rect 9316 30366 9340 30422
rect 9396 30366 9420 30422
rect 9476 30366 9500 30422
rect 9556 30366 9580 30422
rect 9636 30366 9660 30422
rect 9716 30366 9740 30422
rect 9796 30366 9820 30422
rect 9876 30366 9900 30422
rect 9956 30366 9980 30422
rect 10036 30366 10060 30422
rect 10116 30366 10140 30422
rect 10196 30366 10220 30422
rect 10276 30366 10300 30422
rect 10356 30366 10380 30422
rect 10436 30366 10460 30422
rect 10516 30366 10540 30422
rect 10596 30366 10620 30422
rect 10676 30366 10700 30422
rect 10756 30366 10780 30422
rect 10836 30366 10860 30422
rect 10916 30366 10940 30422
rect 10996 30366 11020 30422
rect 11076 30366 11100 30422
rect 11156 30366 11180 30422
rect 11236 30366 11260 30422
rect 11316 30366 11340 30422
rect 11396 30366 11420 30422
rect 11476 30366 11500 30422
rect 11556 30366 11580 30422
rect 11636 30366 11660 30422
rect 11716 30366 11740 30422
rect 11796 30366 11820 30422
rect 11876 30366 11900 30422
rect 11956 30366 11980 30422
rect 12036 30366 12060 30422
rect 12116 30366 12140 30422
rect 12196 30366 12220 30422
rect 12276 30366 12300 30422
rect 12356 30366 12380 30422
rect 12436 30366 12460 30422
rect 12516 30366 12540 30422
rect 12596 30366 12620 30422
rect 12676 30366 12700 30422
rect 12756 30366 12780 30422
rect 12836 30366 12860 30422
rect 12916 30366 12940 30422
rect 12996 30366 13020 30422
rect 13076 30366 13085 30422
rect 6135 30358 13085 30366
rect 5777 30340 13085 30358
rect 5777 30332 6182 30340
rect 5777 30276 5803 30332
rect 5859 30276 5895 30332
rect 5951 30276 5987 30332
rect 6043 30276 6079 30332
rect 6135 30284 6182 30332
rect 6238 30284 6263 30340
rect 6319 30284 6344 30340
rect 6400 30284 6425 30340
rect 6481 30284 6506 30340
rect 6562 30284 6587 30340
rect 6643 30284 6668 30340
rect 6724 30284 6749 30340
rect 6805 30284 6830 30340
rect 6886 30284 6911 30340
rect 6967 30284 6992 30340
rect 7048 30284 7073 30340
rect 7129 30284 7154 30340
rect 7210 30284 7235 30340
rect 7291 30284 7316 30340
rect 7372 30284 7397 30340
rect 7453 30284 7478 30340
rect 7534 30284 7559 30340
rect 7615 30284 7640 30340
rect 7696 30284 7721 30340
rect 7777 30284 7802 30340
rect 7858 30284 7883 30340
rect 7939 30284 7964 30340
rect 8020 30284 8045 30340
rect 8101 30284 8126 30340
rect 8182 30284 8207 30340
rect 8263 30284 8288 30340
rect 8344 30284 8369 30340
rect 8425 30284 8450 30340
rect 8506 30284 8531 30340
rect 8587 30284 8612 30340
rect 8668 30284 8693 30340
rect 8749 30284 8774 30340
rect 8830 30284 8855 30340
rect 8911 30284 8936 30340
rect 8992 30284 9017 30340
rect 9073 30284 9098 30340
rect 9154 30284 9179 30340
rect 9235 30284 9260 30340
rect 9316 30284 9340 30340
rect 9396 30284 9420 30340
rect 9476 30284 9500 30340
rect 9556 30284 9580 30340
rect 9636 30284 9660 30340
rect 9716 30284 9740 30340
rect 9796 30284 9820 30340
rect 9876 30284 9900 30340
rect 9956 30284 9980 30340
rect 10036 30284 10060 30340
rect 10116 30284 10140 30340
rect 10196 30284 10220 30340
rect 10276 30284 10300 30340
rect 10356 30284 10380 30340
rect 10436 30284 10460 30340
rect 10516 30284 10540 30340
rect 10596 30284 10620 30340
rect 10676 30284 10700 30340
rect 10756 30284 10780 30340
rect 10836 30284 10860 30340
rect 10916 30284 10940 30340
rect 10996 30284 11020 30340
rect 11076 30284 11100 30340
rect 11156 30284 11180 30340
rect 11236 30284 11260 30340
rect 11316 30284 11340 30340
rect 11396 30284 11420 30340
rect 11476 30284 11500 30340
rect 11556 30284 11580 30340
rect 11636 30284 11660 30340
rect 11716 30284 11740 30340
rect 11796 30284 11820 30340
rect 11876 30284 11900 30340
rect 11956 30284 11980 30340
rect 12036 30284 12060 30340
rect 12116 30284 12140 30340
rect 12196 30284 12220 30340
rect 12276 30284 12300 30340
rect 12356 30284 12380 30340
rect 12436 30284 12460 30340
rect 12516 30284 12540 30340
rect 12596 30284 12620 30340
rect 12676 30284 12700 30340
rect 12756 30284 12780 30340
rect 12836 30284 12860 30340
rect 12916 30284 12940 30340
rect 12996 30284 13020 30340
rect 13076 30284 13085 30340
rect 6135 30276 13085 30284
rect 5777 30258 13085 30276
rect 5777 30250 6182 30258
rect 5777 30194 5803 30250
rect 5859 30194 5895 30250
rect 5951 30194 5987 30250
rect 6043 30194 6079 30250
rect 6135 30202 6182 30250
rect 6238 30202 6263 30258
rect 6319 30202 6344 30258
rect 6400 30202 6425 30258
rect 6481 30202 6506 30258
rect 6562 30202 6587 30258
rect 6643 30202 6668 30258
rect 6724 30202 6749 30258
rect 6805 30202 6830 30258
rect 6886 30202 6911 30258
rect 6967 30202 6992 30258
rect 7048 30202 7073 30258
rect 7129 30202 7154 30258
rect 7210 30202 7235 30258
rect 7291 30202 7316 30258
rect 7372 30202 7397 30258
rect 7453 30202 7478 30258
rect 7534 30202 7559 30258
rect 7615 30202 7640 30258
rect 7696 30202 7721 30258
rect 7777 30202 7802 30258
rect 7858 30202 7883 30258
rect 7939 30202 7964 30258
rect 8020 30202 8045 30258
rect 8101 30202 8126 30258
rect 8182 30202 8207 30258
rect 8263 30202 8288 30258
rect 8344 30202 8369 30258
rect 8425 30202 8450 30258
rect 8506 30202 8531 30258
rect 8587 30202 8612 30258
rect 8668 30202 8693 30258
rect 8749 30202 8774 30258
rect 8830 30202 8855 30258
rect 8911 30202 8936 30258
rect 8992 30202 9017 30258
rect 9073 30202 9098 30258
rect 9154 30202 9179 30258
rect 9235 30202 9260 30258
rect 9316 30202 9340 30258
rect 9396 30202 9420 30258
rect 9476 30202 9500 30258
rect 9556 30202 9580 30258
rect 9636 30202 9660 30258
rect 9716 30202 9740 30258
rect 9796 30202 9820 30258
rect 9876 30202 9900 30258
rect 9956 30202 9980 30258
rect 10036 30202 10060 30258
rect 10116 30202 10140 30258
rect 10196 30202 10220 30258
rect 10276 30202 10300 30258
rect 10356 30202 10380 30258
rect 10436 30202 10460 30258
rect 10516 30202 10540 30258
rect 10596 30202 10620 30258
rect 10676 30202 10700 30258
rect 10756 30202 10780 30258
rect 10836 30202 10860 30258
rect 10916 30202 10940 30258
rect 10996 30202 11020 30258
rect 11076 30202 11100 30258
rect 11156 30202 11180 30258
rect 11236 30202 11260 30258
rect 11316 30202 11340 30258
rect 11396 30202 11420 30258
rect 11476 30202 11500 30258
rect 11556 30202 11580 30258
rect 11636 30202 11660 30258
rect 11716 30202 11740 30258
rect 11796 30202 11820 30258
rect 11876 30202 11900 30258
rect 11956 30202 11980 30258
rect 12036 30202 12060 30258
rect 12116 30202 12140 30258
rect 12196 30202 12220 30258
rect 12276 30202 12300 30258
rect 12356 30202 12380 30258
rect 12436 30202 12460 30258
rect 12516 30202 12540 30258
rect 12596 30202 12620 30258
rect 12676 30202 12700 30258
rect 12756 30202 12780 30258
rect 12836 30202 12860 30258
rect 12916 30202 12940 30258
rect 12996 30202 13020 30258
rect 13076 30202 13085 30258
rect 6135 30194 13085 30202
rect 5777 30189 13085 30194
rect 5777 29883 13085 29888
rect 5777 29827 5803 29883
rect 5859 29827 5895 29883
rect 5951 29827 5987 29883
rect 6043 29827 6079 29883
rect 6135 29880 13085 29883
rect 6135 29827 6182 29880
rect 5777 29824 6182 29827
rect 6238 29824 6263 29880
rect 6319 29824 6344 29880
rect 6400 29824 6425 29880
rect 6481 29824 6506 29880
rect 6562 29824 6587 29880
rect 6643 29824 6668 29880
rect 6724 29824 6749 29880
rect 6805 29824 6830 29880
rect 6886 29824 6911 29880
rect 6967 29824 6992 29880
rect 7048 29824 7073 29880
rect 7129 29824 7154 29880
rect 7210 29824 7235 29880
rect 7291 29824 7316 29880
rect 7372 29824 7397 29880
rect 7453 29824 7478 29880
rect 7534 29824 7559 29880
rect 7615 29824 7640 29880
rect 7696 29824 7721 29880
rect 7777 29824 7802 29880
rect 7858 29824 7883 29880
rect 7939 29824 7964 29880
rect 8020 29824 8045 29880
rect 8101 29824 8126 29880
rect 8182 29824 8207 29880
rect 8263 29824 8288 29880
rect 8344 29824 8369 29880
rect 8425 29824 8450 29880
rect 8506 29824 8531 29880
rect 8587 29824 8612 29880
rect 8668 29824 8693 29880
rect 8749 29824 8774 29880
rect 8830 29824 8855 29880
rect 8911 29824 8936 29880
rect 8992 29824 9017 29880
rect 9073 29824 9098 29880
rect 9154 29824 9179 29880
rect 9235 29824 9260 29880
rect 5777 29801 9260 29824
rect 5777 29745 5803 29801
rect 5859 29745 5895 29801
rect 5951 29745 5987 29801
rect 6043 29745 6079 29801
rect 6135 29800 9260 29801
rect 6135 29745 6182 29800
rect 5777 29744 6182 29745
rect 6238 29744 6263 29800
rect 6319 29744 6344 29800
rect 6400 29744 6425 29800
rect 6481 29744 6506 29800
rect 6562 29744 6587 29800
rect 6643 29744 6668 29800
rect 6724 29744 6749 29800
rect 6805 29744 6830 29800
rect 6886 29744 6911 29800
rect 6967 29744 6992 29800
rect 7048 29744 7073 29800
rect 7129 29744 7154 29800
rect 7210 29744 7235 29800
rect 7291 29744 7316 29800
rect 7372 29744 7397 29800
rect 7453 29744 7478 29800
rect 7534 29744 7559 29800
rect 7615 29744 7640 29800
rect 7696 29744 7721 29800
rect 7777 29744 7802 29800
rect 7858 29744 7883 29800
rect 7939 29744 7964 29800
rect 8020 29744 8045 29800
rect 8101 29744 8126 29800
rect 8182 29744 8207 29800
rect 8263 29744 8288 29800
rect 8344 29744 8369 29800
rect 8425 29744 8450 29800
rect 8506 29744 8531 29800
rect 8587 29744 8612 29800
rect 8668 29744 8693 29800
rect 8749 29744 8774 29800
rect 8830 29744 8855 29800
rect 8911 29744 8936 29800
rect 8992 29744 9017 29800
rect 9073 29744 9098 29800
rect 9154 29744 9179 29800
rect 9235 29744 9260 29800
rect 5777 29720 9260 29744
rect 5777 29719 6182 29720
rect 5777 29663 5803 29719
rect 5859 29663 5895 29719
rect 5951 29663 5987 29719
rect 6043 29663 6079 29719
rect 6135 29664 6182 29719
rect 6238 29664 6263 29720
rect 6319 29664 6344 29720
rect 6400 29664 6425 29720
rect 6481 29664 6506 29720
rect 6562 29664 6587 29720
rect 6643 29664 6668 29720
rect 6724 29664 6749 29720
rect 6805 29664 6830 29720
rect 6886 29664 6911 29720
rect 6967 29664 6992 29720
rect 7048 29664 7073 29720
rect 7129 29664 7154 29720
rect 7210 29664 7235 29720
rect 7291 29664 7316 29720
rect 7372 29664 7397 29720
rect 7453 29664 7478 29720
rect 7534 29664 7559 29720
rect 7615 29664 7640 29720
rect 7696 29664 7721 29720
rect 7777 29664 7802 29720
rect 7858 29664 7883 29720
rect 7939 29664 7964 29720
rect 8020 29664 8045 29720
rect 8101 29664 8126 29720
rect 8182 29664 8207 29720
rect 8263 29664 8288 29720
rect 8344 29664 8369 29720
rect 8425 29664 8450 29720
rect 8506 29664 8531 29720
rect 8587 29664 8612 29720
rect 8668 29664 8693 29720
rect 8749 29664 8774 29720
rect 8830 29664 8855 29720
rect 8911 29664 8936 29720
rect 8992 29664 9017 29720
rect 9073 29664 9098 29720
rect 9154 29664 9179 29720
rect 9235 29664 9260 29720
rect 6135 29663 9260 29664
rect 5777 29640 9260 29663
rect 5777 29637 6182 29640
rect 5777 29581 5803 29637
rect 5859 29581 5895 29637
rect 5951 29581 5987 29637
rect 6043 29581 6079 29637
rect 6135 29584 6182 29637
rect 6238 29584 6263 29640
rect 6319 29584 6344 29640
rect 6400 29584 6425 29640
rect 6481 29584 6506 29640
rect 6562 29584 6587 29640
rect 6643 29584 6668 29640
rect 6724 29584 6749 29640
rect 6805 29584 6830 29640
rect 6886 29584 6911 29640
rect 6967 29584 6992 29640
rect 7048 29584 7073 29640
rect 7129 29584 7154 29640
rect 7210 29584 7235 29640
rect 7291 29584 7316 29640
rect 7372 29584 7397 29640
rect 7453 29584 7478 29640
rect 7534 29584 7559 29640
rect 7615 29584 7640 29640
rect 7696 29584 7721 29640
rect 7777 29584 7802 29640
rect 7858 29584 7883 29640
rect 7939 29584 7964 29640
rect 8020 29584 8045 29640
rect 8101 29584 8126 29640
rect 8182 29584 8207 29640
rect 8263 29584 8288 29640
rect 8344 29584 8369 29640
rect 8425 29584 8450 29640
rect 8506 29584 8531 29640
rect 8587 29584 8612 29640
rect 8668 29584 8693 29640
rect 8749 29584 8774 29640
rect 8830 29584 8855 29640
rect 8911 29584 8936 29640
rect 8992 29584 9017 29640
rect 9073 29584 9098 29640
rect 9154 29584 9179 29640
rect 9235 29584 9260 29640
rect 6135 29581 9260 29584
rect 5777 29560 9260 29581
rect 5777 29555 6182 29560
rect 5777 29499 5803 29555
rect 5859 29499 5895 29555
rect 5951 29499 5987 29555
rect 6043 29499 6079 29555
rect 6135 29504 6182 29555
rect 6238 29504 6263 29560
rect 6319 29504 6344 29560
rect 6400 29504 6425 29560
rect 6481 29504 6506 29560
rect 6562 29504 6587 29560
rect 6643 29504 6668 29560
rect 6724 29504 6749 29560
rect 6805 29504 6830 29560
rect 6886 29504 6911 29560
rect 6967 29504 6992 29560
rect 7048 29504 7073 29560
rect 7129 29504 7154 29560
rect 7210 29504 7235 29560
rect 7291 29504 7316 29560
rect 7372 29504 7397 29560
rect 7453 29504 7478 29560
rect 7534 29504 7559 29560
rect 7615 29504 7640 29560
rect 7696 29504 7721 29560
rect 7777 29504 7802 29560
rect 7858 29504 7883 29560
rect 7939 29504 7964 29560
rect 8020 29504 8045 29560
rect 8101 29504 8126 29560
rect 8182 29504 8207 29560
rect 8263 29504 8288 29560
rect 8344 29504 8369 29560
rect 8425 29504 8450 29560
rect 8506 29504 8531 29560
rect 8587 29504 8612 29560
rect 8668 29504 8693 29560
rect 8749 29504 8774 29560
rect 8830 29504 8855 29560
rect 8911 29504 8936 29560
rect 8992 29504 9017 29560
rect 9073 29504 9098 29560
rect 9154 29504 9179 29560
rect 9235 29504 9260 29560
rect 6135 29499 9260 29504
rect 5777 29480 9260 29499
rect 5777 29472 6182 29480
rect 5777 29416 5803 29472
rect 5859 29416 5895 29472
rect 5951 29416 5987 29472
rect 6043 29416 6079 29472
rect 6135 29424 6182 29472
rect 6238 29424 6263 29480
rect 6319 29424 6344 29480
rect 6400 29424 6425 29480
rect 6481 29424 6506 29480
rect 6562 29424 6587 29480
rect 6643 29424 6668 29480
rect 6724 29424 6749 29480
rect 6805 29424 6830 29480
rect 6886 29424 6911 29480
rect 6967 29424 6992 29480
rect 7048 29424 7073 29480
rect 7129 29424 7154 29480
rect 7210 29424 7235 29480
rect 7291 29424 7316 29480
rect 7372 29424 7397 29480
rect 7453 29424 7478 29480
rect 7534 29424 7559 29480
rect 7615 29424 7640 29480
rect 7696 29424 7721 29480
rect 7777 29424 7802 29480
rect 7858 29424 7883 29480
rect 7939 29424 7964 29480
rect 8020 29424 8045 29480
rect 8101 29424 8126 29480
rect 8182 29424 8207 29480
rect 8263 29424 8288 29480
rect 8344 29424 8369 29480
rect 8425 29424 8450 29480
rect 8506 29424 8531 29480
rect 8587 29424 8612 29480
rect 8668 29424 8693 29480
rect 8749 29424 8774 29480
rect 8830 29424 8855 29480
rect 8911 29424 8936 29480
rect 8992 29424 9017 29480
rect 9073 29424 9098 29480
rect 9154 29424 9179 29480
rect 9235 29424 9260 29480
rect 6135 29416 9260 29424
rect 5777 29400 9260 29416
rect 5777 29389 6182 29400
rect 5777 29333 5803 29389
rect 5859 29333 5895 29389
rect 5951 29333 5987 29389
rect 6043 29333 6079 29389
rect 6135 29344 6182 29389
rect 6238 29344 6263 29400
rect 6319 29344 6344 29400
rect 6400 29344 6425 29400
rect 6481 29344 6506 29400
rect 6562 29344 6587 29400
rect 6643 29344 6668 29400
rect 6724 29344 6749 29400
rect 6805 29344 6830 29400
rect 6886 29344 6911 29400
rect 6967 29344 6992 29400
rect 7048 29344 7073 29400
rect 7129 29344 7154 29400
rect 7210 29344 7235 29400
rect 7291 29344 7316 29400
rect 7372 29344 7397 29400
rect 7453 29344 7478 29400
rect 7534 29344 7559 29400
rect 7615 29344 7640 29400
rect 7696 29344 7721 29400
rect 7777 29344 7802 29400
rect 7858 29344 7883 29400
rect 7939 29344 7964 29400
rect 8020 29344 8045 29400
rect 8101 29344 8126 29400
rect 8182 29344 8207 29400
rect 8263 29344 8288 29400
rect 8344 29344 8369 29400
rect 8425 29344 8450 29400
rect 8506 29344 8531 29400
rect 8587 29344 8612 29400
rect 8668 29344 8693 29400
rect 8749 29344 8774 29400
rect 8830 29344 8855 29400
rect 8911 29344 8936 29400
rect 8992 29344 9017 29400
rect 9073 29344 9098 29400
rect 9154 29344 9179 29400
rect 9235 29344 9260 29400
rect 6135 29333 9260 29344
rect 5777 29320 9260 29333
rect 5777 29306 6182 29320
rect 5777 29250 5803 29306
rect 5859 29250 5895 29306
rect 5951 29250 5987 29306
rect 6043 29250 6079 29306
rect 6135 29264 6182 29306
rect 6238 29264 6263 29320
rect 6319 29264 6344 29320
rect 6400 29264 6425 29320
rect 6481 29264 6506 29320
rect 6562 29264 6587 29320
rect 6643 29264 6668 29320
rect 6724 29264 6749 29320
rect 6805 29264 6830 29320
rect 6886 29264 6911 29320
rect 6967 29264 6992 29320
rect 7048 29264 7073 29320
rect 7129 29264 7154 29320
rect 7210 29264 7235 29320
rect 7291 29264 7316 29320
rect 7372 29264 7397 29320
rect 7453 29264 7478 29320
rect 7534 29264 7559 29320
rect 7615 29264 7640 29320
rect 7696 29264 7721 29320
rect 7777 29264 7802 29320
rect 7858 29264 7883 29320
rect 7939 29264 7964 29320
rect 8020 29264 8045 29320
rect 8101 29264 8126 29320
rect 8182 29264 8207 29320
rect 8263 29264 8288 29320
rect 8344 29264 8369 29320
rect 8425 29264 8450 29320
rect 8506 29264 8531 29320
rect 8587 29264 8612 29320
rect 8668 29264 8693 29320
rect 8749 29264 8774 29320
rect 8830 29264 8855 29320
rect 8911 29264 8936 29320
rect 8992 29264 9017 29320
rect 9073 29264 9098 29320
rect 9154 29264 9179 29320
rect 9235 29264 9260 29320
rect 6135 29250 9260 29264
rect 5777 29240 9260 29250
rect 5777 29223 6182 29240
rect 5777 29167 5803 29223
rect 5859 29167 5895 29223
rect 5951 29167 5987 29223
rect 6043 29167 6079 29223
rect 6135 29184 6182 29223
rect 6238 29184 6263 29240
rect 6319 29184 6344 29240
rect 6400 29184 6425 29240
rect 6481 29184 6506 29240
rect 6562 29184 6587 29240
rect 6643 29184 6668 29240
rect 6724 29184 6749 29240
rect 6805 29184 6830 29240
rect 6886 29184 6911 29240
rect 6967 29184 6992 29240
rect 7048 29184 7073 29240
rect 7129 29184 7154 29240
rect 7210 29184 7235 29240
rect 7291 29184 7316 29240
rect 7372 29184 7397 29240
rect 7453 29184 7478 29240
rect 7534 29184 7559 29240
rect 7615 29184 7640 29240
rect 7696 29184 7721 29240
rect 7777 29184 7802 29240
rect 7858 29184 7883 29240
rect 7939 29184 7964 29240
rect 8020 29184 8045 29240
rect 8101 29184 8126 29240
rect 8182 29184 8207 29240
rect 8263 29184 8288 29240
rect 8344 29184 8369 29240
rect 8425 29184 8450 29240
rect 8506 29184 8531 29240
rect 8587 29184 8612 29240
rect 8668 29184 8693 29240
rect 8749 29184 8774 29240
rect 8830 29184 8855 29240
rect 8911 29184 8936 29240
rect 8992 29184 9017 29240
rect 9073 29184 9098 29240
rect 9154 29184 9179 29240
rect 9235 29184 9260 29240
rect 6135 29167 9260 29184
rect 5777 29160 9260 29167
rect 5777 29140 6182 29160
rect 5777 29084 5803 29140
rect 5859 29084 5895 29140
rect 5951 29084 5987 29140
rect 6043 29084 6079 29140
rect 6135 29104 6182 29140
rect 6238 29104 6263 29160
rect 6319 29104 6344 29160
rect 6400 29104 6425 29160
rect 6481 29104 6506 29160
rect 6562 29104 6587 29160
rect 6643 29104 6668 29160
rect 6724 29104 6749 29160
rect 6805 29104 6830 29160
rect 6886 29104 6911 29160
rect 6967 29104 6992 29160
rect 7048 29104 7073 29160
rect 7129 29104 7154 29160
rect 7210 29104 7235 29160
rect 7291 29104 7316 29160
rect 7372 29104 7397 29160
rect 7453 29104 7478 29160
rect 7534 29104 7559 29160
rect 7615 29104 7640 29160
rect 7696 29104 7721 29160
rect 7777 29104 7802 29160
rect 7858 29104 7883 29160
rect 7939 29104 7964 29160
rect 8020 29104 8045 29160
rect 8101 29104 8126 29160
rect 8182 29104 8207 29160
rect 8263 29104 8288 29160
rect 8344 29104 8369 29160
rect 8425 29104 8450 29160
rect 8506 29104 8531 29160
rect 8587 29104 8612 29160
rect 8668 29104 8693 29160
rect 8749 29104 8774 29160
rect 8830 29104 8855 29160
rect 8911 29104 8936 29160
rect 8992 29104 9017 29160
rect 9073 29104 9098 29160
rect 9154 29104 9179 29160
rect 9235 29104 9260 29160
rect 6135 29084 9260 29104
rect 5777 29080 9260 29084
rect 5777 29078 6182 29080
tri 5777 29024 5831 29078 ne
rect 5831 29024 6182 29078
rect 6238 29024 6263 29080
rect 6319 29024 6344 29080
rect 6400 29024 6425 29080
rect 6481 29024 6506 29080
rect 6562 29024 6587 29080
rect 6643 29024 6668 29080
rect 6724 29024 6749 29080
rect 6805 29024 6830 29080
rect 6886 29024 6911 29080
rect 6967 29024 6992 29080
rect 7048 29024 7073 29080
rect 7129 29024 7154 29080
rect 7210 29024 7235 29080
rect 7291 29024 7316 29080
rect 7372 29024 7397 29080
rect 7453 29024 7478 29080
rect 7534 29024 7559 29080
rect 7615 29024 7640 29080
rect 7696 29024 7721 29080
rect 7777 29024 7802 29080
rect 7858 29024 7883 29080
rect 7939 29024 7964 29080
rect 8020 29024 8045 29080
rect 8101 29024 8126 29080
rect 8182 29024 8207 29080
rect 8263 29024 8288 29080
rect 8344 29024 8369 29080
rect 8425 29024 8450 29080
rect 8506 29024 8531 29080
rect 8587 29024 8612 29080
rect 8668 29024 8693 29080
rect 8749 29024 8774 29080
rect 8830 29024 8855 29080
rect 8911 29024 8936 29080
rect 8992 29024 9017 29080
rect 9073 29024 9098 29080
rect 9154 29024 9179 29080
rect 9235 29024 9260 29080
tri 5831 29000 5855 29024 ne
rect 5855 29000 9260 29024
tri 5855 28944 5911 29000 ne
rect 5911 28944 6182 29000
rect 6238 28944 6263 29000
rect 6319 28944 6344 29000
rect 6400 28944 6425 29000
rect 6481 28944 6506 29000
rect 6562 28944 6587 29000
rect 6643 28944 6668 29000
rect 6724 28944 6749 29000
rect 6805 28944 6830 29000
rect 6886 28944 6911 29000
rect 6967 28944 6992 29000
rect 7048 28944 7073 29000
rect 7129 28944 7154 29000
rect 7210 28944 7235 29000
rect 7291 28944 7316 29000
rect 7372 28944 7397 29000
rect 7453 28944 7478 29000
rect 7534 28944 7559 29000
rect 7615 28944 7640 29000
rect 7696 28944 7721 29000
rect 7777 28944 7802 29000
rect 7858 28944 7883 29000
rect 7939 28944 7964 29000
rect 8020 28944 8045 29000
rect 8101 28944 8126 29000
rect 8182 28944 8207 29000
rect 8263 28944 8288 29000
rect 8344 28944 8369 29000
rect 8425 28944 8450 29000
rect 8506 28944 8531 29000
rect 8587 28944 8612 29000
rect 8668 28944 8693 29000
rect 8749 28944 8774 29000
rect 8830 28944 8855 29000
rect 8911 28944 8936 29000
rect 8992 28944 9017 29000
rect 9073 28944 9098 29000
rect 9154 28944 9179 29000
rect 9235 28944 9260 29000
tri 5911 28920 5935 28944 ne
rect 5935 28920 9260 28944
tri 5935 28866 5989 28920 ne
rect 5989 28866 6182 28920
tri 5989 28864 5991 28866 ne
rect 5991 28864 6182 28866
rect 6238 28864 6263 28920
rect 6319 28864 6344 28920
rect 6400 28864 6425 28920
rect 6481 28864 6506 28920
rect 6562 28864 6587 28920
rect 6643 28864 6668 28920
rect 6724 28864 6749 28920
rect 6805 28864 6830 28920
rect 6886 28864 6911 28920
rect 6967 28864 6992 28920
rect 7048 28864 7073 28920
rect 7129 28864 7154 28920
rect 7210 28864 7235 28920
rect 7291 28864 7316 28920
rect 7372 28864 7397 28920
rect 7453 28864 7478 28920
rect 7534 28864 7559 28920
rect 7615 28864 7640 28920
rect 7696 28864 7721 28920
rect 7777 28864 7802 28920
rect 7858 28864 7883 28920
rect 7939 28864 7964 28920
rect 8020 28864 8045 28920
rect 8101 28864 8126 28920
rect 8182 28864 8207 28920
rect 8263 28864 8288 28920
rect 8344 28864 8369 28920
rect 8425 28864 8450 28920
rect 8506 28864 8531 28920
rect 8587 28864 8612 28920
rect 8668 28864 8693 28920
rect 8749 28864 8774 28920
rect 8830 28864 8855 28920
rect 8911 28864 8936 28920
rect 8992 28864 9017 28920
rect 9073 28864 9098 28920
rect 9154 28864 9179 28920
rect 9235 28864 9260 28920
rect 13076 28864 13085 29880
tri 5991 28857 5998 28864 ne
rect 5998 28857 13085 28864
tri 5998 28690 6165 28857 ne
rect 6165 28690 13085 28857
tri 2024 28506 2058 28540 sw
rect 2781 28506 2790 28562
rect 2846 28506 2874 28562
rect 2930 28506 2958 28562
rect 3014 28506 3042 28562
rect 3098 28506 3126 28562
rect 3182 28506 3210 28562
rect 3266 28506 3294 28562
rect 3350 28506 3378 28562
rect 3434 28506 3462 28562
rect 3518 28506 3545 28562
rect 3601 28506 3628 28562
rect 3684 28506 3711 28562
rect 3767 28506 3778 28562
rect 1054 28424 2058 28506
tri 2058 28424 2140 28506 sw
rect 2781 28424 3778 28506
rect 1054 28368 2140 28424
tri 2140 28368 2196 28424 sw
rect 2781 28368 2790 28424
rect 2846 28368 2874 28424
rect 2930 28368 2958 28424
rect 3014 28368 3042 28424
rect 3098 28368 3126 28424
rect 3182 28368 3210 28424
rect 3266 28368 3294 28424
rect 3350 28368 3378 28424
rect 3434 28368 3462 28424
rect 3518 28368 3545 28424
rect 3601 28368 3628 28424
rect 3684 28368 3711 28424
rect 3767 28368 3778 28424
rect 1054 28363 2196 28368
tri 2196 28363 2201 28368 sw
rect 1054 28067 2201 28363
tri 2201 28067 2497 28363 sw
rect 1054 28057 2497 28067
rect 1054 28001 2165 28057
rect 2221 28001 2255 28057
rect 2311 28001 2345 28057
rect 2401 28001 2435 28057
rect 2491 28001 2497 28057
rect 1054 27977 2497 28001
rect 1054 27921 2165 27977
rect 2221 27921 2255 27977
rect 2311 27921 2345 27977
rect 2401 27921 2435 27977
rect 2491 27921 2497 27977
rect 1054 27897 2497 27921
rect 1054 27841 2165 27897
rect 2221 27841 2255 27897
rect 2311 27841 2345 27897
rect 2401 27841 2435 27897
rect 2491 27841 2497 27897
rect 1054 27817 2497 27841
rect 1054 27761 2165 27817
rect 2221 27761 2255 27817
rect 2311 27761 2345 27817
rect 2401 27761 2435 27817
rect 2491 27761 2497 27817
rect 1054 27737 2497 27761
rect 1054 27681 2165 27737
rect 2221 27681 2255 27737
rect 2311 27681 2345 27737
rect 2401 27681 2435 27737
rect 2491 27681 2497 27737
rect 1054 27657 2497 27681
rect 1054 27601 2165 27657
rect 2221 27601 2255 27657
rect 2311 27601 2345 27657
rect 2401 27601 2435 27657
rect 2491 27601 2497 27657
rect 1054 27577 2497 27601
rect 1054 27521 2165 27577
rect 2221 27521 2255 27577
rect 2311 27521 2345 27577
rect 2401 27521 2435 27577
rect 2491 27521 2497 27577
rect 1054 27497 2497 27521
rect 1054 27441 2165 27497
rect 2221 27441 2255 27497
rect 2311 27441 2345 27497
rect 2401 27441 2435 27497
rect 2491 27441 2497 27497
rect 1054 27417 2497 27441
rect 1054 27361 2165 27417
rect 2221 27361 2255 27417
rect 2311 27361 2345 27417
rect 2401 27361 2435 27417
rect 2491 27361 2497 27417
rect 1054 27337 2497 27361
rect 1054 27281 2165 27337
rect 2221 27281 2255 27337
rect 2311 27281 2345 27337
rect 2401 27281 2435 27337
rect 2491 27281 2497 27337
rect 1054 27257 2497 27281
rect 1054 27201 2165 27257
rect 2221 27201 2255 27257
rect 2311 27201 2345 27257
rect 2401 27201 2435 27257
rect 2491 27201 2497 27257
rect 1054 27177 2497 27201
rect 1054 27121 2165 27177
rect 2221 27121 2255 27177
rect 2311 27121 2345 27177
rect 2401 27121 2435 27177
rect 2491 27121 2497 27177
rect 1054 27097 2497 27121
rect 1054 27041 2165 27097
rect 2221 27041 2255 27097
rect 2311 27041 2345 27097
rect 2401 27041 2435 27097
rect 2491 27041 2497 27097
rect 1054 27017 2497 27041
rect 1054 26961 2165 27017
rect 2221 26961 2255 27017
rect 2311 26961 2345 27017
rect 2401 26961 2435 27017
rect 2491 26961 2497 27017
rect 1054 26936 2497 26961
rect 1054 26880 2165 26936
rect 2221 26880 2255 26936
rect 2311 26880 2345 26936
rect 2401 26880 2435 26936
rect 2491 26880 2497 26936
rect 1054 26855 2497 26880
rect 1054 26799 2165 26855
rect 2221 26799 2255 26855
rect 2311 26799 2345 26855
rect 2401 26799 2435 26855
rect 2491 26799 2497 26855
rect 1054 26774 2497 26799
rect 1054 26718 2165 26774
rect 2221 26718 2255 26774
rect 2311 26718 2345 26774
rect 2401 26718 2435 26774
rect 2491 26718 2497 26774
rect 1054 26693 2497 26718
rect 1054 26637 2165 26693
rect 2221 26637 2255 26693
rect 2311 26637 2345 26693
rect 2401 26637 2435 26693
rect 2491 26637 2497 26693
rect 1054 26612 2497 26637
rect 1054 26556 2165 26612
rect 2221 26556 2255 26612
rect 2311 26556 2345 26612
rect 2401 26556 2435 26612
rect 2491 26556 2497 26612
rect 1054 26531 2497 26556
rect 1054 26475 2165 26531
rect 2221 26475 2255 26531
rect 2311 26475 2345 26531
rect 2401 26475 2435 26531
rect 2491 26475 2497 26531
rect 1054 26450 2497 26475
rect 1054 26394 2165 26450
rect 2221 26394 2255 26450
rect 2311 26394 2345 26450
rect 2401 26394 2435 26450
rect 2491 26394 2497 26450
rect 1054 26385 2497 26394
rect 292 26309 299 26365
rect 355 26309 393 26365
rect 449 26309 487 26365
rect 543 26309 581 26365
rect 637 26309 656 26365
rect 292 26282 656 26309
rect 292 26226 299 26282
rect 355 26226 393 26282
rect 449 26226 487 26282
rect 543 26226 581 26282
rect 637 26226 656 26282
rect 292 21258 656 26226
rect 1960 25853 2500 25880
rect 1960 25789 1977 25853
rect 2041 25789 2067 25853
rect 2131 25789 2157 25853
rect 2221 25820 2247 25853
rect 2311 25820 2337 25853
rect 2401 25820 2427 25853
rect 2226 25789 2247 25820
rect 2311 25789 2334 25820
rect 2401 25789 2416 25820
rect 2491 25789 2500 25853
rect 1960 25770 2170 25789
rect 2226 25770 2252 25789
rect 2308 25770 2334 25789
rect 2390 25770 2416 25789
rect 2472 25770 2500 25789
rect 1960 25706 1977 25770
rect 2041 25706 2067 25770
rect 2131 25706 2157 25770
rect 2226 25764 2247 25770
rect 2311 25764 2334 25770
rect 2401 25764 2416 25770
rect 2221 25739 2247 25764
rect 2311 25739 2337 25764
rect 2401 25739 2427 25764
rect 2226 25706 2247 25739
rect 2311 25706 2334 25739
rect 2401 25706 2416 25739
rect 2491 25706 2500 25770
rect 1960 25687 2170 25706
rect 2226 25687 2252 25706
rect 2308 25687 2334 25706
rect 2390 25687 2416 25706
rect 2472 25687 2500 25706
rect 1960 25623 1977 25687
rect 2041 25623 2067 25687
rect 2131 25623 2157 25687
rect 2226 25683 2247 25687
rect 2311 25683 2334 25687
rect 2401 25683 2416 25687
rect 2221 25658 2247 25683
rect 2311 25658 2337 25683
rect 2401 25658 2427 25683
rect 2226 25623 2247 25658
rect 2311 25623 2334 25658
rect 2401 25623 2416 25658
rect 2491 25623 2500 25687
rect 1960 25604 2170 25623
rect 2226 25604 2252 25623
rect 2308 25604 2334 25623
rect 2390 25604 2416 25623
rect 2472 25604 2500 25623
rect 1960 25540 1977 25604
rect 2041 25540 2067 25604
rect 2131 25540 2157 25604
rect 2226 25602 2247 25604
rect 2311 25602 2334 25604
rect 2401 25602 2416 25604
rect 2221 25577 2247 25602
rect 2311 25577 2337 25602
rect 2401 25577 2427 25602
rect 2226 25540 2247 25577
rect 2311 25540 2334 25577
rect 2401 25540 2416 25577
rect 2491 25540 2500 25604
rect 1960 25521 2170 25540
rect 2226 25521 2252 25540
rect 2308 25521 2334 25540
rect 2390 25521 2416 25540
rect 2472 25521 2500 25540
rect 1960 25457 1977 25521
rect 2041 25457 2067 25521
rect 2131 25457 2157 25521
rect 2221 25496 2247 25521
rect 2311 25496 2337 25521
rect 2401 25496 2427 25521
rect 2226 25457 2247 25496
rect 2311 25457 2334 25496
rect 2401 25457 2416 25496
rect 2491 25457 2500 25521
rect 1960 25440 2170 25457
rect 2226 25440 2252 25457
rect 2308 25440 2334 25457
rect 2390 25440 2416 25457
rect 2472 25440 2500 25457
rect 1960 25437 2500 25440
rect 1960 25373 1977 25437
rect 2041 25373 2067 25437
rect 2131 25373 2157 25437
rect 2221 25415 2247 25437
rect 2311 25415 2337 25437
rect 2401 25415 2427 25437
rect 2226 25373 2247 25415
rect 2311 25373 2334 25415
rect 2401 25373 2416 25415
rect 2491 25373 2500 25437
rect 1960 25359 2170 25373
rect 2226 25359 2252 25373
rect 2308 25359 2334 25373
rect 2390 25359 2416 25373
rect 2472 25359 2500 25373
rect 1960 25353 2500 25359
rect 1960 25289 1977 25353
rect 2041 25289 2067 25353
rect 2131 25289 2157 25353
rect 2221 25334 2247 25353
rect 2311 25334 2337 25353
rect 2401 25334 2427 25353
rect 2226 25289 2247 25334
rect 2311 25289 2334 25334
rect 2401 25289 2416 25334
rect 2491 25289 2500 25353
rect 1960 25278 2170 25289
rect 2226 25278 2252 25289
rect 2308 25278 2334 25289
rect 2390 25278 2416 25289
rect 2472 25278 2500 25289
rect 1960 25269 2500 25278
rect 1960 25205 1977 25269
rect 2041 25205 2067 25269
rect 2131 25205 2157 25269
rect 2221 25253 2247 25269
rect 2311 25253 2337 25269
rect 2401 25253 2427 25269
rect 2226 25205 2247 25253
rect 2311 25205 2334 25253
rect 2401 25205 2416 25253
rect 2491 25205 2500 25269
rect 1960 25197 2170 25205
rect 2226 25197 2252 25205
rect 2308 25197 2334 25205
rect 2390 25197 2416 25205
rect 2472 25197 2500 25205
rect 1960 25185 2500 25197
rect 1960 25121 1977 25185
rect 2041 25121 2067 25185
rect 2131 25121 2157 25185
rect 2221 25172 2247 25185
rect 2311 25172 2337 25185
rect 2401 25172 2427 25185
rect 2226 25121 2247 25172
rect 2311 25121 2334 25172
rect 2401 25121 2416 25172
rect 2491 25121 2500 25185
rect 1960 25116 2170 25121
rect 2226 25116 2252 25121
rect 2308 25116 2334 25121
rect 2390 25116 2416 25121
rect 2472 25116 2500 25121
rect 1960 25101 2500 25116
rect 1960 25037 1977 25101
rect 2041 25037 2067 25101
rect 2131 25037 2157 25101
rect 2221 25091 2247 25101
rect 2311 25091 2337 25101
rect 2401 25091 2427 25101
rect 2226 25037 2247 25091
rect 2311 25037 2334 25091
rect 2401 25037 2416 25091
rect 2491 25037 2500 25101
rect 1960 25035 2170 25037
rect 2226 25035 2252 25037
rect 2308 25035 2334 25037
rect 2390 25035 2416 25037
rect 2472 25035 2500 25037
rect 1960 25017 2500 25035
rect 1960 24953 1977 25017
rect 2041 24953 2067 25017
rect 2131 24953 2157 25017
rect 2221 25010 2247 25017
rect 2311 25010 2337 25017
rect 2401 25010 2427 25017
rect 2226 24954 2247 25010
rect 2311 24954 2334 25010
rect 2401 24954 2416 25010
rect 2221 24953 2247 24954
rect 2311 24953 2337 24954
rect 2401 24953 2427 24954
rect 2491 24953 2500 25017
rect 1960 24933 2500 24953
rect 1960 24869 1977 24933
rect 2041 24869 2067 24933
rect 2131 24869 2157 24933
rect 2221 24929 2247 24933
rect 2311 24929 2337 24933
rect 2401 24929 2427 24933
rect 2226 24873 2247 24929
rect 2311 24873 2334 24929
rect 2401 24873 2416 24929
rect 2221 24869 2247 24873
rect 2311 24869 2337 24873
rect 2401 24869 2427 24873
rect 2491 24869 2500 24933
rect 1960 24849 2500 24869
rect 1960 24785 1977 24849
rect 2041 24785 2067 24849
rect 2131 24785 2157 24849
rect 2221 24848 2247 24849
rect 2311 24848 2337 24849
rect 2401 24848 2427 24849
rect 2226 24792 2247 24848
rect 2311 24792 2334 24848
rect 2401 24792 2416 24848
rect 2221 24785 2247 24792
rect 2311 24785 2337 24792
rect 2401 24785 2427 24792
rect 2491 24785 2500 24849
rect 1960 24767 2500 24785
rect 1960 24765 2170 24767
rect 2226 24765 2252 24767
rect 2308 24765 2334 24767
rect 2390 24765 2416 24767
rect 2472 24765 2500 24767
rect 1960 24701 1977 24765
rect 2041 24701 2067 24765
rect 2131 24701 2157 24765
rect 2226 24711 2247 24765
rect 2311 24711 2334 24765
rect 2401 24711 2416 24765
rect 2221 24701 2247 24711
rect 2311 24701 2337 24711
rect 2401 24701 2427 24711
rect 2491 24701 2500 24765
rect 1960 24686 2500 24701
rect 1960 24681 2170 24686
rect 2226 24681 2252 24686
rect 2308 24681 2334 24686
rect 2390 24681 2416 24686
rect 2472 24681 2500 24686
rect 1960 24617 1977 24681
rect 2041 24617 2067 24681
rect 2131 24617 2157 24681
rect 2226 24630 2247 24681
rect 2311 24630 2334 24681
rect 2401 24630 2416 24681
rect 2221 24617 2247 24630
rect 2311 24617 2337 24630
rect 2401 24617 2427 24630
rect 2491 24617 2500 24681
rect 1960 24604 2500 24617
rect 1960 24597 2170 24604
rect 2226 24597 2252 24604
rect 2308 24597 2334 24604
rect 2390 24597 2416 24604
rect 2472 24597 2500 24604
rect 1960 24533 1977 24597
rect 2041 24533 2067 24597
rect 2131 24533 2157 24597
rect 2226 24548 2247 24597
rect 2311 24548 2334 24597
rect 2401 24548 2416 24597
rect 2221 24533 2247 24548
rect 2311 24533 2337 24548
rect 2401 24533 2427 24548
rect 2491 24533 2500 24597
rect 1960 24522 2500 24533
rect 1960 24513 2170 24522
rect 2226 24513 2252 24522
rect 2308 24513 2334 24522
rect 2390 24513 2416 24522
rect 2472 24513 2500 24522
rect 1960 24449 1977 24513
rect 2041 24449 2067 24513
rect 2131 24449 2157 24513
rect 2226 24466 2247 24513
rect 2311 24466 2334 24513
rect 2401 24466 2416 24513
rect 2221 24449 2247 24466
rect 2311 24449 2337 24466
rect 2401 24449 2427 24466
rect 2491 24449 2500 24513
rect 1960 24440 2500 24449
rect 1960 24429 2170 24440
rect 2226 24429 2252 24440
rect 2308 24429 2334 24440
rect 2390 24429 2416 24440
rect 2472 24429 2500 24440
rect 1960 24365 1977 24429
rect 2041 24365 2067 24429
rect 2131 24365 2157 24429
rect 2226 24384 2247 24429
rect 2311 24384 2334 24429
rect 2401 24384 2416 24429
rect 2221 24365 2247 24384
rect 2311 24365 2337 24384
rect 2401 24365 2427 24384
rect 2491 24365 2500 24429
rect 1960 24358 2500 24365
rect 1960 24345 2170 24358
rect 2226 24345 2252 24358
rect 2308 24345 2334 24358
rect 2390 24345 2416 24358
rect 2472 24345 2500 24358
rect 1960 24281 1977 24345
rect 2041 24281 2067 24345
rect 2131 24281 2157 24345
rect 2226 24302 2247 24345
rect 2311 24302 2334 24345
rect 2401 24302 2416 24345
rect 2221 24281 2247 24302
rect 2311 24281 2337 24302
rect 2401 24281 2427 24302
rect 2491 24281 2500 24345
rect 1960 24276 2500 24281
tri 1930 24220 1960 24250 se
rect 1960 24240 2170 24276
rect 2226 24240 2252 24276
rect 2308 24240 2334 24276
rect 2390 24240 2416 24276
rect 2472 24240 2500 24276
rect 1960 24220 1977 24240
tri 1904 24194 1930 24220 se
rect 1930 24194 1977 24220
tri 1848 24138 1904 24194 se
rect 1904 24176 1977 24194
rect 2041 24176 2065 24240
rect 2129 24176 2153 24240
rect 2226 24220 2241 24240
rect 2308 24220 2328 24240
rect 2217 24194 2241 24220
rect 2305 24194 2328 24220
rect 2226 24176 2241 24194
rect 2308 24176 2328 24194
rect 2392 24176 2415 24240
rect 2479 24176 2500 24240
rect 1904 24144 2170 24176
rect 2226 24144 2252 24176
rect 2308 24144 2334 24176
rect 2390 24144 2416 24176
rect 2472 24144 2500 24176
rect 1904 24138 1977 24144
tri 1822 24112 1848 24138 se
rect 1848 24112 1977 24138
tri 1766 24056 1822 24112 se
rect 1822 24080 1977 24112
rect 2041 24080 2065 24144
rect 2129 24080 2153 24144
rect 2226 24138 2241 24144
rect 2308 24138 2328 24144
rect 2217 24112 2241 24138
rect 2305 24112 2328 24138
rect 2226 24080 2241 24112
rect 2308 24080 2328 24112
rect 2392 24080 2415 24144
rect 2479 24080 2500 24144
rect 1822 24056 2170 24080
rect 2226 24056 2252 24080
rect 2308 24056 2334 24080
rect 2390 24056 2416 24080
rect 2472 24056 2500 24080
tri 1740 24030 1766 24056 se
rect 1766 24048 2500 24056
rect 1766 24030 1977 24048
tri 1717 24007 1740 24030 se
rect 1740 24007 1977 24030
tri 1684 23974 1717 24007 se
rect 1717 24001 1977 24007
rect 1717 23974 1739 24001
tri 1658 23948 1684 23974 se
rect 1684 23948 1739 23974
tri 1602 23892 1658 23948 se
rect 1658 23937 1739 23948
rect 1803 23937 1875 24001
rect 1939 23984 1977 24001
rect 2041 23984 2065 24048
rect 2129 23984 2153 24048
rect 2217 24030 2241 24048
rect 2305 24030 2328 24048
rect 2226 23984 2241 24030
rect 2308 23984 2328 24030
rect 2392 23984 2415 24048
rect 2479 23984 2500 24048
rect 1939 23974 2170 23984
rect 2226 23974 2252 23984
rect 2308 23974 2334 23984
rect 2390 23974 2416 23984
rect 2472 23974 2500 23984
rect 1939 23952 2500 23974
rect 1939 23937 1977 23952
rect 1658 23892 1977 23937
tri 1577 23867 1602 23892 se
rect 1602 23888 1977 23892
rect 2041 23888 2065 23952
rect 2129 23888 2153 23952
rect 2217 23948 2241 23952
rect 2305 23948 2328 23952
rect 2226 23892 2241 23948
rect 2308 23892 2328 23948
rect 2217 23888 2241 23892
rect 2305 23888 2328 23892
rect 2392 23888 2415 23952
rect 2479 23888 2500 23952
rect 1602 23867 2500 23888
tri 1576 23866 1577 23867 se
rect 1577 23866 2500 23867
tri 1520 23810 1576 23866 se
rect 1576 23865 2170 23866
rect 1576 23810 1739 23865
tri 1501 23791 1520 23810 se
rect 1520 23801 1739 23810
rect 1803 23801 1875 23865
rect 1939 23856 2170 23865
rect 2226 23856 2252 23866
rect 2308 23856 2334 23866
rect 2390 23856 2416 23866
rect 2472 23856 2500 23866
rect 1939 23801 1977 23856
rect 1520 23792 1977 23801
rect 2041 23792 2065 23856
rect 2129 23792 2153 23856
rect 2226 23810 2241 23856
rect 2308 23810 2328 23856
rect 2217 23792 2241 23810
rect 2305 23792 2328 23810
rect 2392 23792 2415 23856
rect 2479 23792 2500 23856
rect 1520 23791 2500 23792
rect 1092 23785 1460 23791
rect 1092 23721 1094 23785
rect 1158 23721 1188 23785
rect 1252 23721 1282 23785
rect 1346 23721 1376 23785
rect 1440 23721 1460 23785
rect 1092 23703 1460 23721
rect 1092 23639 1094 23703
rect 1158 23639 1188 23703
rect 1252 23639 1282 23703
rect 1346 23639 1376 23703
rect 1440 23639 1460 23703
rect 1092 23621 1460 23639
rect 1092 23557 1094 23621
rect 1158 23557 1188 23621
rect 1252 23557 1282 23621
rect 1346 23557 1376 23621
rect 1440 23557 1460 23621
rect 1092 23539 1460 23557
rect 1092 23475 1094 23539
rect 1158 23475 1188 23539
rect 1252 23475 1282 23539
rect 1346 23475 1376 23539
rect 1440 23475 1460 23539
rect 1092 23457 1460 23475
rect 1092 23393 1094 23457
rect 1158 23393 1188 23457
rect 1252 23393 1282 23457
rect 1346 23393 1376 23457
rect 1440 23393 1460 23457
rect 1092 23375 1460 23393
rect 1092 23311 1094 23375
rect 1158 23311 1188 23375
rect 1252 23311 1282 23375
rect 1346 23311 1376 23375
rect 1440 23311 1460 23375
rect 1092 23293 1460 23311
rect 1092 23229 1094 23293
rect 1158 23229 1188 23293
rect 1252 23229 1282 23293
rect 1346 23229 1376 23293
rect 1440 23229 1460 23293
rect 1092 23211 1460 23229
rect 1092 23147 1094 23211
rect 1158 23147 1188 23211
rect 1252 23147 1282 23211
rect 1346 23147 1376 23211
rect 1440 23147 1460 23211
rect 1092 23129 1460 23147
rect 1092 23065 1094 23129
rect 1158 23065 1188 23129
rect 1252 23065 1282 23129
rect 1346 23065 1376 23129
rect 1440 23065 1460 23129
rect 1092 23047 1460 23065
rect 1092 22983 1094 23047
rect 1158 22983 1188 23047
rect 1252 22983 1282 23047
rect 1346 22983 1376 23047
rect 1440 22983 1460 23047
rect 1092 22964 1460 22983
rect 1092 22900 1094 22964
rect 1158 22900 1188 22964
rect 1252 22900 1282 22964
rect 1346 22900 1376 22964
rect 1440 22900 1460 22964
rect 1092 22881 1460 22900
rect 1092 22817 1094 22881
rect 1158 22817 1188 22881
rect 1252 22817 1282 22881
rect 1346 22817 1376 22881
rect 1440 22817 1460 22881
rect 1092 22798 1460 22817
rect 1092 22734 1094 22798
rect 1158 22734 1188 22798
rect 1252 22734 1282 22798
rect 1346 22734 1376 22798
rect 1440 22734 1460 22798
rect 1092 22715 1460 22734
rect 1092 22651 1094 22715
rect 1158 22651 1188 22715
rect 1252 22651 1282 22715
rect 1346 22651 1376 22715
rect 1440 22651 1460 22715
rect 1092 22632 1460 22651
rect 1092 22568 1094 22632
rect 1158 22568 1188 22632
rect 1252 22568 1282 22632
rect 1346 22568 1376 22632
rect 1440 22568 1460 22632
rect 1092 22549 1460 22568
rect 1092 22485 1094 22549
rect 1158 22485 1188 22549
rect 1252 22485 1282 22549
rect 1346 22485 1376 22549
rect 1440 22485 1460 22549
rect 1092 22466 1460 22485
rect 1092 22402 1094 22466
rect 1158 22402 1188 22466
rect 1252 22402 1282 22466
rect 1346 22402 1376 22466
rect 1440 22402 1460 22466
rect 1092 22383 1460 22402
rect 1092 22319 1094 22383
rect 1158 22319 1188 22383
rect 1252 22319 1282 22383
rect 1346 22319 1376 22383
rect 1440 22319 1460 22383
rect 1092 22300 1460 22319
rect 1092 22236 1094 22300
rect 1158 22236 1188 22300
rect 1252 22236 1282 22300
rect 1346 22236 1376 22300
rect 1440 22236 1460 22300
rect 1092 22217 1460 22236
rect 1092 22153 1094 22217
rect 1158 22153 1188 22217
rect 1252 22153 1282 22217
rect 1346 22153 1376 22217
rect 1440 22153 1460 22217
rect 1092 22134 1460 22153
rect 1092 22070 1094 22134
rect 1158 22070 1188 22134
rect 1252 22070 1282 22134
rect 1346 22070 1376 22134
rect 1440 22070 1460 22134
rect 1092 22051 1460 22070
rect 1092 21987 1094 22051
rect 1158 21987 1188 22051
rect 1252 21987 1282 22051
rect 1346 21987 1376 22051
rect 1440 21987 1460 22051
rect 1092 21968 1460 21987
rect 1092 21904 1094 21968
rect 1158 21904 1188 21968
rect 1252 21904 1282 21968
rect 1346 21904 1376 21968
rect 1440 21904 1460 21968
rect 1092 21885 1460 21904
rect 1092 21821 1094 21885
rect 1158 21821 1188 21885
rect 1252 21821 1282 21885
rect 1346 21821 1376 21885
rect 1440 21821 1460 21885
rect 1092 21802 1460 21821
rect 1092 21738 1094 21802
rect 1158 21738 1188 21802
rect 1252 21738 1282 21802
rect 1346 21738 1376 21802
rect 1440 21738 1460 21802
rect 1092 21719 1460 21738
rect 1092 21655 1094 21719
rect 1158 21655 1188 21719
rect 1252 21655 1282 21719
rect 1346 21655 1376 21719
rect 1440 21655 1460 21719
rect 1092 21636 1460 21655
rect 1092 21572 1094 21636
rect 1158 21572 1188 21636
rect 1252 21572 1282 21636
rect 1346 21572 1376 21636
rect 1440 21572 1460 21636
rect 1092 21553 1460 21572
rect 1092 21489 1094 21553
rect 1158 21489 1188 21553
rect 1252 21489 1282 21553
rect 1346 21489 1376 21553
rect 1440 21489 1460 21553
rect 1092 21470 1460 21489
rect 1092 21406 1094 21470
rect 1158 21406 1188 21470
rect 1252 21406 1282 21470
rect 1346 21406 1376 21470
rect 1440 21406 1460 21470
rect 1092 21387 1460 21406
rect 1092 21323 1094 21387
rect 1158 21323 1188 21387
rect 1252 21323 1282 21387
rect 1346 21323 1376 21387
rect 1440 21323 1460 21387
rect 1092 21317 1460 21323
rect 1467 23784 2500 23791
rect 1467 23773 2170 23784
rect 2226 23773 2252 23784
rect 2308 23773 2334 23784
rect 2390 23773 2416 23784
rect 2472 23773 2500 23784
rect 1467 23709 1474 23773
rect 1538 23709 1554 23773
rect 1618 23709 1634 23773
rect 1698 23709 1714 23773
rect 1778 23709 1794 23773
rect 1858 23709 1874 23773
rect 1938 23709 1954 23773
rect 2018 23709 2034 23773
rect 2098 23709 2114 23773
rect 2178 23709 2194 23728
rect 2258 23709 2274 23728
rect 2338 23709 2354 23728
rect 2418 23709 2434 23728
rect 2498 23709 2500 23773
rect 1467 23702 2500 23709
rect 1467 23691 2170 23702
rect 2226 23691 2252 23702
rect 2308 23691 2334 23702
rect 2390 23691 2416 23702
rect 2472 23691 2500 23702
rect 1467 23627 1474 23691
rect 1538 23627 1554 23691
rect 1618 23627 1634 23691
rect 1698 23627 1714 23691
rect 1778 23627 1794 23691
rect 1858 23627 1874 23691
rect 1938 23627 1954 23691
rect 2018 23627 2034 23691
rect 2098 23627 2114 23691
rect 2178 23627 2194 23646
rect 2258 23627 2274 23646
rect 2338 23627 2354 23646
rect 2418 23627 2434 23646
rect 2498 23627 2500 23691
rect 1467 23620 2500 23627
rect 1467 23609 2170 23620
rect 2226 23609 2252 23620
rect 2308 23609 2334 23620
rect 2390 23609 2416 23620
rect 2472 23609 2500 23620
rect 1467 23545 1474 23609
rect 1538 23545 1554 23609
rect 1618 23545 1634 23609
rect 1698 23545 1714 23609
rect 1778 23545 1794 23609
rect 1858 23545 1874 23609
rect 1938 23545 1954 23609
rect 2018 23545 2034 23609
rect 2098 23545 2114 23609
rect 2178 23545 2194 23564
rect 2258 23545 2274 23564
rect 2338 23545 2354 23564
rect 2418 23545 2434 23564
rect 2498 23545 2500 23609
rect 1467 23538 2500 23545
rect 1467 23527 2170 23538
rect 2226 23527 2252 23538
rect 2308 23527 2334 23538
rect 2390 23527 2416 23538
rect 2472 23527 2500 23538
rect 1467 23463 1474 23527
rect 1538 23463 1554 23527
rect 1618 23463 1634 23527
rect 1698 23463 1714 23527
rect 1778 23463 1794 23527
rect 1858 23463 1874 23527
rect 1938 23463 1954 23527
rect 2018 23463 2034 23527
rect 2098 23463 2114 23527
rect 2178 23463 2194 23482
rect 2258 23463 2274 23482
rect 2338 23463 2354 23482
rect 2418 23463 2434 23482
rect 2498 23463 2500 23527
rect 1467 23456 2500 23463
rect 1467 23445 2170 23456
rect 2226 23445 2252 23456
rect 2308 23445 2334 23456
rect 2390 23445 2416 23456
rect 2472 23445 2500 23456
rect 1467 23381 1474 23445
rect 1538 23381 1554 23445
rect 1618 23381 1634 23445
rect 1698 23381 1714 23445
rect 1778 23381 1794 23445
rect 1858 23381 1874 23445
rect 1938 23381 1954 23445
rect 2018 23381 2034 23445
rect 2098 23381 2114 23445
rect 2178 23381 2194 23400
rect 2258 23381 2274 23400
rect 2338 23381 2354 23400
rect 2418 23381 2434 23400
rect 2498 23381 2500 23445
rect 1467 23374 2500 23381
rect 1467 23363 2170 23374
rect 2226 23363 2252 23374
rect 2308 23363 2334 23374
rect 2390 23363 2416 23374
rect 2472 23363 2500 23374
rect 1467 23299 1474 23363
rect 1538 23299 1554 23363
rect 1618 23299 1634 23363
rect 1698 23299 1714 23363
rect 1778 23299 1794 23363
rect 1858 23299 1874 23363
rect 1938 23299 1954 23363
rect 2018 23299 2034 23363
rect 2098 23299 2114 23363
rect 2178 23299 2194 23318
rect 2258 23299 2274 23318
rect 2338 23299 2354 23318
rect 2418 23299 2434 23318
rect 2498 23299 2500 23363
rect 1467 23292 2500 23299
rect 1467 23281 2170 23292
rect 2226 23281 2252 23292
rect 2308 23281 2334 23292
rect 2390 23281 2416 23292
rect 2472 23281 2500 23292
rect 1467 23217 1474 23281
rect 1538 23217 1554 23281
rect 1618 23217 1634 23281
rect 1698 23217 1714 23281
rect 1778 23217 1794 23281
rect 1858 23217 1874 23281
rect 1938 23217 1954 23281
rect 2018 23217 2034 23281
rect 2098 23217 2114 23281
rect 2178 23217 2194 23236
rect 2258 23217 2274 23236
rect 2338 23217 2354 23236
rect 2418 23217 2434 23236
rect 2498 23217 2500 23281
rect 1467 23210 2500 23217
rect 1467 23199 2170 23210
rect 2226 23199 2252 23210
rect 2308 23199 2334 23210
rect 2390 23199 2416 23210
rect 2472 23199 2500 23210
rect 1467 23135 1474 23199
rect 1538 23135 1554 23199
rect 1618 23135 1634 23199
rect 1698 23135 1714 23199
rect 1778 23135 1794 23199
rect 1858 23135 1874 23199
rect 1938 23135 1954 23199
rect 2018 23135 2034 23199
rect 2098 23135 2114 23199
rect 2178 23135 2194 23154
rect 2258 23135 2274 23154
rect 2338 23135 2354 23154
rect 2418 23135 2434 23154
rect 2498 23135 2500 23199
rect 1467 23117 2500 23135
rect 1467 23053 1474 23117
rect 1538 23053 1554 23117
rect 1618 23053 1634 23117
rect 1698 23053 1714 23117
rect 1778 23053 1794 23117
rect 1858 23053 1874 23117
rect 1938 23053 1954 23117
rect 2018 23053 2034 23117
rect 2098 23053 2114 23117
rect 2178 23053 2194 23117
rect 2258 23053 2274 23117
rect 2338 23053 2354 23117
rect 2418 23053 2434 23117
rect 2498 23053 2500 23117
rect 1467 23035 2500 23053
rect 1467 22971 1474 23035
rect 1538 22971 1554 23035
rect 1618 22971 1634 23035
rect 1698 22971 1714 23035
rect 1778 22971 1794 23035
rect 1858 22971 1874 23035
rect 1938 22971 1954 23035
rect 2018 22971 2034 23035
rect 2098 22971 2114 23035
rect 2178 22971 2194 23035
rect 2258 22971 2274 23035
rect 2338 22971 2354 23035
rect 2418 22971 2434 23035
rect 2498 22971 2500 23035
rect 1467 22953 2500 22971
rect 1467 22889 1474 22953
rect 1538 22889 1554 22953
rect 1618 22889 1634 22953
rect 1698 22889 1714 22953
rect 1778 22889 1794 22953
rect 1858 22889 1874 22953
rect 1938 22889 1954 22953
rect 2018 22889 2034 22953
rect 2098 22889 2114 22953
rect 2178 22889 2194 22953
rect 2258 22889 2274 22953
rect 2338 22889 2354 22953
rect 2418 22889 2434 22953
rect 2498 22889 2500 22953
rect 1467 22871 2500 22889
rect 1467 22807 1474 22871
rect 1538 22807 1554 22871
rect 1618 22807 1634 22871
rect 1698 22807 1714 22871
rect 1778 22807 1794 22871
rect 1858 22807 1874 22871
rect 1938 22807 1954 22871
rect 2018 22807 2034 22871
rect 2098 22807 2114 22871
rect 2178 22807 2194 22871
rect 2258 22807 2274 22871
rect 2338 22807 2354 22871
rect 2418 22807 2434 22871
rect 2498 22807 2500 22871
rect 1467 22789 2500 22807
rect 1467 22725 1474 22789
rect 1538 22725 1554 22789
rect 1618 22725 1634 22789
rect 1698 22725 1714 22789
rect 1778 22725 1794 22789
rect 1858 22725 1874 22789
rect 1938 22725 1954 22789
rect 2018 22725 2034 22789
rect 2098 22725 2114 22789
rect 2178 22725 2194 22789
rect 2258 22725 2274 22789
rect 2338 22725 2354 22789
rect 2418 22725 2434 22789
rect 2498 22725 2500 22789
rect 1467 22707 2500 22725
rect 1467 22643 1474 22707
rect 1538 22643 1554 22707
rect 1618 22643 1634 22707
rect 1698 22643 1714 22707
rect 1778 22643 1794 22707
rect 1858 22643 1874 22707
rect 1938 22643 1954 22707
rect 2018 22643 2034 22707
rect 2098 22643 2114 22707
rect 2178 22643 2194 22707
rect 2258 22643 2274 22707
rect 2338 22643 2354 22707
rect 2418 22643 2434 22707
rect 2498 22643 2500 22707
rect 1467 22625 2500 22643
rect 1467 22561 1474 22625
rect 1538 22561 1554 22625
rect 1618 22561 1634 22625
rect 1698 22561 1714 22625
rect 1778 22561 1794 22625
rect 1858 22561 1874 22625
rect 1938 22561 1954 22625
rect 2018 22561 2034 22625
rect 2098 22561 2114 22625
rect 2178 22561 2194 22625
rect 2258 22561 2274 22625
rect 2338 22561 2354 22625
rect 2418 22561 2434 22625
rect 2498 22561 2500 22625
rect 1467 22543 2500 22561
rect 1467 22479 1474 22543
rect 1538 22479 1554 22543
rect 1618 22479 1634 22543
rect 1698 22479 1714 22543
rect 1778 22479 1794 22543
rect 1858 22479 1874 22543
rect 1938 22479 1954 22543
rect 2018 22479 2034 22543
rect 2098 22479 2114 22543
rect 2178 22479 2194 22543
rect 2258 22479 2274 22543
rect 2338 22479 2354 22543
rect 2418 22479 2434 22543
rect 2498 22479 2500 22543
rect 1467 22461 2500 22479
rect 1467 22397 1474 22461
rect 1538 22397 1554 22461
rect 1618 22397 1634 22461
rect 1698 22397 1714 22461
rect 1778 22397 1794 22461
rect 1858 22397 1874 22461
rect 1938 22397 1954 22461
rect 2018 22397 2034 22461
rect 2098 22397 2114 22461
rect 2178 22397 2194 22461
rect 2258 22397 2274 22461
rect 2338 22397 2354 22461
rect 2418 22397 2434 22461
rect 2498 22397 2500 22461
rect 1467 22379 2500 22397
rect 1467 22315 1474 22379
rect 1538 22315 1554 22379
rect 1618 22315 1634 22379
rect 1698 22315 1714 22379
rect 1778 22315 1794 22379
rect 1858 22315 1874 22379
rect 1938 22315 1954 22379
rect 2018 22315 2034 22379
rect 2098 22315 2114 22379
rect 2178 22315 2194 22379
rect 2258 22315 2274 22379
rect 2338 22315 2354 22379
rect 2418 22315 2434 22379
rect 2498 22315 2500 22379
rect 1467 22297 2500 22315
rect 1467 22233 1474 22297
rect 1538 22233 1554 22297
rect 1618 22233 1634 22297
rect 1698 22233 1714 22297
rect 1778 22233 1794 22297
rect 1858 22233 1874 22297
rect 1938 22233 1954 22297
rect 2018 22233 2034 22297
rect 2098 22233 2114 22297
rect 2178 22233 2194 22297
rect 2258 22233 2274 22297
rect 2338 22233 2354 22297
rect 2418 22233 2434 22297
rect 2498 22233 2500 22297
rect 1467 22215 2500 22233
rect 1467 22151 1474 22215
rect 1538 22151 1554 22215
rect 1618 22151 1634 22215
rect 1698 22151 1714 22215
rect 1778 22151 1794 22215
rect 1858 22151 1874 22215
rect 1938 22151 1954 22215
rect 2018 22151 2034 22215
rect 2098 22151 2114 22215
rect 2178 22151 2194 22215
rect 2258 22151 2274 22215
rect 2338 22151 2354 22215
rect 2418 22151 2434 22215
rect 2498 22151 2500 22215
rect 1467 22133 2500 22151
rect 1467 22069 1474 22133
rect 1538 22069 1554 22133
rect 1618 22069 1634 22133
rect 1698 22069 1714 22133
rect 1778 22069 1794 22133
rect 1858 22069 1874 22133
rect 1938 22069 1954 22133
rect 2018 22069 2034 22133
rect 2098 22069 2114 22133
rect 2178 22069 2194 22133
rect 2258 22069 2274 22133
rect 2338 22069 2354 22133
rect 2418 22069 2434 22133
rect 2498 22069 2500 22133
rect 1467 22051 2500 22069
rect 1467 21987 1474 22051
rect 1538 21987 1554 22051
rect 1618 21987 1634 22051
rect 1698 21987 1714 22051
rect 1778 21987 1794 22051
rect 1858 21987 1874 22051
rect 1938 21987 1954 22051
rect 2018 21987 2034 22051
rect 2098 21987 2114 22051
rect 2178 21987 2194 22051
rect 2258 21987 2274 22051
rect 2338 21987 2354 22051
rect 2418 21987 2434 22051
rect 2498 21987 2500 22051
rect 1467 21968 2500 21987
rect 1467 21904 1474 21968
rect 1538 21904 1554 21968
rect 1618 21904 1634 21968
rect 1698 21904 1714 21968
rect 1778 21904 1794 21968
rect 1858 21904 1874 21968
rect 1938 21904 1954 21968
rect 2018 21904 2034 21968
rect 2098 21904 2114 21968
rect 2178 21904 2194 21968
rect 2258 21904 2274 21968
rect 2338 21904 2354 21968
rect 2418 21904 2434 21968
rect 2498 21904 2500 21968
rect 1467 21885 2500 21904
rect 1467 21821 1474 21885
rect 1538 21821 1554 21885
rect 1618 21821 1634 21885
rect 1698 21821 1714 21885
rect 1778 21821 1794 21885
rect 1858 21821 1874 21885
rect 1938 21821 1954 21885
rect 2018 21821 2034 21885
rect 2098 21821 2114 21885
rect 2178 21821 2194 21885
rect 2258 21821 2274 21885
rect 2338 21821 2354 21885
rect 2418 21821 2434 21885
rect 2498 21821 2500 21885
rect 1467 21802 2500 21821
rect 1467 21738 1474 21802
rect 1538 21738 1554 21802
rect 1618 21738 1634 21802
rect 1698 21738 1714 21802
rect 1778 21738 1794 21802
rect 1858 21738 1874 21802
rect 1938 21738 1954 21802
rect 2018 21738 2034 21802
rect 2098 21738 2114 21802
rect 2178 21738 2194 21802
rect 2258 21738 2274 21802
rect 2338 21738 2354 21802
rect 2418 21738 2434 21802
rect 2498 21738 2500 21802
rect 1467 21719 2500 21738
rect 1467 21655 1474 21719
rect 1538 21655 1554 21719
rect 1618 21655 1634 21719
rect 1698 21655 1714 21719
rect 1778 21655 1794 21719
rect 1858 21655 1874 21719
rect 1938 21655 1954 21719
rect 2018 21655 2034 21719
rect 2098 21655 2114 21719
rect 2178 21655 2194 21719
rect 2258 21655 2274 21719
rect 2338 21655 2354 21719
rect 2418 21655 2434 21719
rect 2498 21655 2500 21719
rect 1467 21636 2500 21655
rect 1467 21572 1474 21636
rect 1538 21572 1554 21636
rect 1618 21572 1634 21636
rect 1698 21572 1714 21636
rect 1778 21572 1794 21636
rect 1858 21572 1874 21636
rect 1938 21572 1954 21636
rect 2018 21572 2034 21636
rect 2098 21572 2114 21636
rect 2178 21572 2194 21636
rect 2258 21572 2274 21636
rect 2338 21572 2354 21636
rect 2418 21572 2434 21636
rect 2498 21572 2500 21636
rect 1467 21553 2500 21572
rect 1467 21489 1474 21553
rect 1538 21489 1554 21553
rect 1618 21489 1634 21553
rect 1698 21489 1714 21553
rect 1778 21489 1794 21553
rect 1858 21489 1874 21553
rect 1938 21489 1954 21553
rect 2018 21489 2034 21553
rect 2098 21489 2114 21553
rect 2178 21489 2194 21553
rect 2258 21489 2274 21553
rect 2338 21489 2354 21553
rect 2418 21489 2434 21553
rect 2498 21489 2500 21553
rect 1467 21470 2500 21489
rect 1467 21406 1474 21470
rect 1538 21406 1554 21470
rect 1618 21406 1634 21470
rect 1698 21406 1714 21470
rect 1778 21406 1794 21470
rect 1858 21406 1874 21470
rect 1938 21406 1954 21470
rect 2018 21406 2034 21470
rect 2098 21406 2114 21470
rect 2178 21406 2194 21470
rect 2258 21406 2274 21470
rect 2338 21406 2354 21470
rect 2418 21406 2434 21470
rect 2498 21406 2500 21470
rect 1467 21387 2500 21406
rect 1467 21323 1474 21387
rect 1538 21323 1554 21387
rect 1618 21323 1634 21387
rect 1698 21323 1714 21387
rect 1778 21323 1794 21387
rect 1858 21323 1874 21387
rect 1938 21323 1954 21387
rect 2018 21323 2034 21387
rect 2098 21323 2114 21387
rect 2178 21323 2194 21387
rect 2258 21323 2274 21387
rect 2338 21323 2354 21387
rect 2418 21323 2434 21387
rect 2498 21323 2500 21387
rect 1467 21317 2500 21323
tri 1241 21282 1276 21317 ne
rect 292 20286 574 21258
tri 574 21176 656 21258 nw
rect 1276 21105 1376 21317
tri 1376 21282 1411 21317 nw
tri 1276 21099 1282 21105 ne
rect 1282 21099 1376 21105
tri 1376 21099 1448 21171 sw
tri 1282 21039 1342 21099 ne
rect 1342 21039 2336 21099
tri 2336 21039 2396 21099 sw
tri 1342 21005 1376 21039 ne
rect 1376 21005 2396 21039
tri 1376 20999 1382 21005 ne
rect 1382 20999 2396 21005
tri 2222 20932 2289 20999 ne
rect 2289 20932 2396 20999
rect 665 20923 2130 20932
tri 2289 20931 2290 20932 ne
rect 2290 20931 2396 20932
tri 2290 20925 2296 20931 ne
rect 665 20867 670 20923
rect 726 20867 794 20923
rect 850 20867 1627 20923
rect 1683 20867 1715 20923
rect 1771 20867 1803 20923
rect 1859 20867 1891 20923
rect 1947 20867 1979 20923
rect 2035 20867 2067 20923
rect 2123 20867 2130 20923
rect 665 20832 2130 20867
rect 665 20776 670 20832
rect 726 20776 794 20832
rect 850 20776 1627 20832
rect 1683 20776 1715 20832
rect 1771 20776 1803 20832
rect 1859 20776 1891 20832
rect 1947 20776 1979 20832
rect 2035 20776 2067 20832
rect 2123 20776 2130 20832
rect 665 20741 2130 20776
rect 665 20685 670 20741
rect 726 20685 794 20741
rect 850 20685 1627 20741
rect 1683 20685 1715 20741
rect 1771 20685 1803 20741
rect 1859 20685 1891 20741
rect 1947 20685 1979 20741
rect 2035 20685 2067 20741
rect 2123 20685 2130 20741
rect 665 20650 2130 20685
rect 665 20594 670 20650
rect 726 20594 794 20650
rect 850 20594 1627 20650
rect 1683 20594 1715 20650
rect 1771 20594 1803 20650
rect 1859 20594 1891 20650
rect 1947 20594 1979 20650
rect 2035 20594 2067 20650
rect 2123 20594 2130 20650
rect 665 20559 2130 20594
rect 665 20503 670 20559
rect 726 20503 794 20559
rect 850 20503 1627 20559
rect 1683 20503 1715 20559
rect 1771 20503 1803 20559
rect 1859 20503 1891 20559
rect 1947 20503 1979 20559
rect 2035 20503 2067 20559
rect 2123 20503 2130 20559
rect 665 20468 2130 20503
rect 665 20412 670 20468
rect 726 20412 794 20468
rect 850 20412 1627 20468
rect 1683 20412 1715 20468
rect 1771 20412 1803 20468
rect 1859 20412 1891 20468
rect 1947 20412 1979 20468
rect 2035 20412 2067 20468
rect 2123 20412 2130 20468
rect 665 20403 2130 20412
tri 574 20286 576 20288 sw
rect 292 20206 576 20286
tri 576 20206 656 20286 sw
rect 292 18976 656 20206
tri 2178 20168 2296 20286 se
rect 2296 20200 2396 20931
rect 2296 20168 2364 20200
tri 2364 20168 2396 20200 nw
rect 2781 20931 3778 28368
rect 4099 28057 5099 28066
rect 4099 28001 4105 28057
rect 4161 28001 4189 28057
rect 4245 28001 4273 28057
rect 4329 28001 4357 28057
rect 4413 28001 4441 28057
rect 4497 28001 4525 28057
rect 4581 28001 4609 28057
rect 4665 28001 4693 28057
rect 4749 28001 4777 28057
rect 4833 28001 4861 28057
rect 4917 28001 4945 28057
rect 5001 28001 5029 28057
rect 5085 28001 5099 28057
rect 4099 27977 5099 28001
rect 4099 27921 4105 27977
rect 4161 27921 4189 27977
rect 4245 27921 4273 27977
rect 4329 27921 4357 27977
rect 4413 27921 4441 27977
rect 4497 27921 4525 27977
rect 4581 27921 4609 27977
rect 4665 27921 4693 27977
rect 4749 27921 4777 27977
rect 4833 27921 4861 27977
rect 4917 27921 4945 27977
rect 5001 27921 5029 27977
rect 5085 27921 5099 27977
rect 4099 27897 5099 27921
rect 4099 27841 4105 27897
rect 4161 27841 4189 27897
rect 4245 27841 4273 27897
rect 4329 27841 4357 27897
rect 4413 27841 4441 27897
rect 4497 27841 4525 27897
rect 4581 27841 4609 27897
rect 4665 27841 4693 27897
rect 4749 27841 4777 27897
rect 4833 27841 4861 27897
rect 4917 27841 4945 27897
rect 5001 27841 5029 27897
rect 5085 27841 5099 27897
rect 4099 27817 5099 27841
rect 4099 27761 4105 27817
rect 4161 27761 4189 27817
rect 4245 27761 4273 27817
rect 4329 27761 4357 27817
rect 4413 27761 4441 27817
rect 4497 27761 4525 27817
rect 4581 27761 4609 27817
rect 4665 27761 4693 27817
rect 4749 27761 4777 27817
rect 4833 27761 4861 27817
rect 4917 27761 4945 27817
rect 5001 27761 5029 27817
rect 5085 27761 5099 27817
rect 4099 27737 5099 27761
rect 4099 27681 4105 27737
rect 4161 27681 4189 27737
rect 4245 27681 4273 27737
rect 4329 27681 4357 27737
rect 4413 27681 4441 27737
rect 4497 27681 4525 27737
rect 4581 27681 4609 27737
rect 4665 27681 4693 27737
rect 4749 27681 4777 27737
rect 4833 27681 4861 27737
rect 4917 27681 4945 27737
rect 5001 27681 5029 27737
rect 5085 27681 5099 27737
rect 4099 27657 5099 27681
rect 4099 27601 4105 27657
rect 4161 27601 4189 27657
rect 4245 27601 4273 27657
rect 4329 27601 4357 27657
rect 4413 27601 4441 27657
rect 4497 27601 4525 27657
rect 4581 27601 4609 27657
rect 4665 27601 4693 27657
rect 4749 27601 4777 27657
rect 4833 27601 4861 27657
rect 4917 27601 4945 27657
rect 5001 27601 5029 27657
rect 5085 27601 5099 27657
rect 4099 27577 5099 27601
rect 4099 27521 4105 27577
rect 4161 27521 4189 27577
rect 4245 27521 4273 27577
rect 4329 27521 4357 27577
rect 4413 27521 4441 27577
rect 4497 27521 4525 27577
rect 4581 27521 4609 27577
rect 4665 27521 4693 27577
rect 4749 27521 4777 27577
rect 4833 27521 4861 27577
rect 4917 27521 4945 27577
rect 5001 27521 5029 27577
rect 5085 27521 5099 27577
rect 4099 27497 5099 27521
rect 4099 27441 4105 27497
rect 4161 27441 4189 27497
rect 4245 27441 4273 27497
rect 4329 27441 4357 27497
rect 4413 27441 4441 27497
rect 4497 27441 4525 27497
rect 4581 27441 4609 27497
rect 4665 27441 4693 27497
rect 4749 27441 4777 27497
rect 4833 27441 4861 27497
rect 4917 27441 4945 27497
rect 5001 27441 5029 27497
rect 5085 27441 5099 27497
rect 4099 27417 5099 27441
rect 4099 27361 4105 27417
rect 4161 27361 4189 27417
rect 4245 27361 4273 27417
rect 4329 27361 4357 27417
rect 4413 27361 4441 27417
rect 4497 27361 4525 27417
rect 4581 27361 4609 27417
rect 4665 27361 4693 27417
rect 4749 27361 4777 27417
rect 4833 27361 4861 27417
rect 4917 27361 4945 27417
rect 5001 27361 5029 27417
rect 5085 27361 5099 27417
rect 4099 27337 5099 27361
rect 4099 27281 4105 27337
rect 4161 27281 4189 27337
rect 4245 27281 4273 27337
rect 4329 27281 4357 27337
rect 4413 27281 4441 27337
rect 4497 27281 4525 27337
rect 4581 27281 4609 27337
rect 4665 27281 4693 27337
rect 4749 27281 4777 27337
rect 4833 27281 4861 27337
rect 4917 27281 4945 27337
rect 5001 27281 5029 27337
rect 5085 27281 5099 27337
rect 4099 27257 5099 27281
rect 4099 27201 4105 27257
rect 4161 27201 4189 27257
rect 4245 27201 4273 27257
rect 4329 27201 4357 27257
rect 4413 27201 4441 27257
rect 4497 27201 4525 27257
rect 4581 27201 4609 27257
rect 4665 27201 4693 27257
rect 4749 27201 4777 27257
rect 4833 27201 4861 27257
rect 4917 27201 4945 27257
rect 5001 27201 5029 27257
rect 5085 27201 5099 27257
rect 4099 27177 5099 27201
rect 4099 27121 4105 27177
rect 4161 27121 4189 27177
rect 4245 27121 4273 27177
rect 4329 27121 4357 27177
rect 4413 27121 4441 27177
rect 4497 27121 4525 27177
rect 4581 27121 4609 27177
rect 4665 27121 4693 27177
rect 4749 27121 4777 27177
rect 4833 27121 4861 27177
rect 4917 27121 4945 27177
rect 5001 27121 5029 27177
rect 5085 27121 5099 27177
rect 4099 27097 5099 27121
rect 4099 27041 4105 27097
rect 4161 27041 4189 27097
rect 4245 27041 4273 27097
rect 4329 27041 4357 27097
rect 4413 27041 4441 27097
rect 4497 27041 4525 27097
rect 4581 27041 4609 27097
rect 4665 27041 4693 27097
rect 4749 27041 4777 27097
rect 4833 27041 4861 27097
rect 4917 27041 4945 27097
rect 5001 27041 5029 27097
rect 5085 27041 5099 27097
rect 4099 27017 5099 27041
rect 4099 26961 4105 27017
rect 4161 26961 4189 27017
rect 4245 26961 4273 27017
rect 4329 26961 4357 27017
rect 4413 26961 4441 27017
rect 4497 26961 4525 27017
rect 4581 26961 4609 27017
rect 4665 26961 4693 27017
rect 4749 26961 4777 27017
rect 4833 26961 4861 27017
rect 4917 26961 4945 27017
rect 5001 26961 5029 27017
rect 5085 26961 5099 27017
rect 4099 26936 5099 26961
rect 4099 26880 4105 26936
rect 4161 26880 4189 26936
rect 4245 26880 4273 26936
rect 4329 26880 4357 26936
rect 4413 26880 4441 26936
rect 4497 26880 4525 26936
rect 4581 26880 4609 26936
rect 4665 26880 4693 26936
rect 4749 26880 4777 26936
rect 4833 26880 4861 26936
rect 4917 26880 4945 26936
rect 5001 26880 5029 26936
rect 5085 26880 5099 26936
rect 4099 26855 5099 26880
rect 4099 26799 4105 26855
rect 4161 26799 4189 26855
rect 4245 26799 4273 26855
rect 4329 26799 4357 26855
rect 4413 26799 4441 26855
rect 4497 26799 4525 26855
rect 4581 26799 4609 26855
rect 4665 26799 4693 26855
rect 4749 26799 4777 26855
rect 4833 26799 4861 26855
rect 4917 26799 4945 26855
rect 5001 26799 5029 26855
rect 5085 26799 5099 26855
rect 4099 26774 5099 26799
rect 4099 26718 4105 26774
rect 4161 26718 4189 26774
rect 4245 26718 4273 26774
rect 4329 26718 4357 26774
rect 4413 26718 4441 26774
rect 4497 26718 4525 26774
rect 4581 26718 4609 26774
rect 4665 26718 4693 26774
rect 4749 26718 4777 26774
rect 4833 26718 4861 26774
rect 4917 26718 4945 26774
rect 5001 26718 5029 26774
rect 5085 26718 5099 26774
rect 4099 26693 5099 26718
rect 4099 26637 4105 26693
rect 4161 26637 4189 26693
rect 4245 26637 4273 26693
rect 4329 26637 4357 26693
rect 4413 26637 4441 26693
rect 4497 26637 4525 26693
rect 4581 26637 4609 26693
rect 4665 26637 4693 26693
rect 4749 26637 4777 26693
rect 4833 26637 4861 26693
rect 4917 26637 4945 26693
rect 5001 26637 5029 26693
rect 5085 26637 5099 26693
rect 4099 26612 5099 26637
rect 4099 26556 4105 26612
rect 4161 26556 4189 26612
rect 4245 26556 4273 26612
rect 4329 26556 4357 26612
rect 4413 26556 4441 26612
rect 4497 26556 4525 26612
rect 4581 26556 4609 26612
rect 4665 26556 4693 26612
rect 4749 26556 4777 26612
rect 4833 26556 4861 26612
rect 4917 26556 4945 26612
rect 5001 26556 5029 26612
rect 5085 26556 5099 26612
rect 4099 26531 5099 26556
rect 4099 26475 4105 26531
rect 4161 26475 4189 26531
rect 4245 26475 4273 26531
rect 4329 26475 4357 26531
rect 4413 26475 4441 26531
rect 4497 26475 4525 26531
rect 4581 26475 4609 26531
rect 4665 26475 4693 26531
rect 4749 26475 4777 26531
rect 4833 26475 4861 26531
rect 4917 26475 4945 26531
rect 5001 26475 5029 26531
rect 5085 26475 5099 26531
rect 4099 26450 5099 26475
rect 4099 26394 4105 26450
rect 4161 26394 4189 26450
rect 4245 26394 4273 26450
rect 4329 26394 4357 26450
rect 4413 26394 4441 26450
rect 4497 26394 4525 26450
rect 4581 26394 4609 26450
rect 4665 26394 4693 26450
rect 4749 26394 4777 26450
rect 4833 26394 4861 26450
rect 4917 26394 4945 26450
rect 5001 26394 5029 26450
rect 5085 26394 5099 26450
rect 4099 21433 5099 26394
rect 5416 25828 13085 25839
rect 5416 25772 5425 25828
rect 5481 25772 5506 25828
rect 5562 25772 5587 25828
rect 5643 25772 5668 25828
rect 5724 25772 5749 25828
rect 5805 25772 5830 25828
rect 5886 25772 5911 25828
rect 5967 25772 5992 25828
rect 6048 25772 6073 25828
rect 6129 25772 6154 25828
rect 6210 25772 6235 25828
rect 6291 25772 6316 25828
rect 6372 25772 6397 25828
rect 6453 25772 6478 25828
rect 6534 25772 6559 25828
rect 6615 25772 6640 25828
rect 6696 25772 6721 25828
rect 6777 25772 6802 25828
rect 6858 25772 6883 25828
rect 6939 25772 6964 25828
rect 7020 25772 7045 25828
rect 7101 25772 7126 25828
rect 7182 25772 7207 25828
rect 7263 25772 7288 25828
rect 7344 25772 7369 25828
rect 7425 25772 7450 25828
rect 7506 25772 7531 25828
rect 7587 25772 7612 25828
rect 7668 25772 7693 25828
rect 7749 25772 7774 25828
rect 7830 25772 7855 25828
rect 7911 25772 7936 25828
rect 7992 25772 8017 25828
rect 8073 25772 8098 25828
rect 8154 25772 8179 25828
rect 8235 25772 8260 25828
rect 8316 25772 8341 25828
rect 8397 25772 8422 25828
rect 8478 25772 8503 25828
rect 8559 25772 8584 25828
rect 8640 25772 8665 25828
rect 8721 25772 8746 25828
rect 8802 25772 8827 25828
rect 8883 25772 8908 25828
rect 8964 25772 8989 25828
rect 9045 25772 9070 25828
rect 9126 25772 9151 25828
rect 9207 25772 9232 25828
rect 9288 25772 9313 25828
rect 9369 25772 9394 25828
rect 9450 25772 9475 25828
rect 9531 25772 9556 25828
rect 9612 25772 9637 25828
rect 9693 25772 9718 25828
rect 9774 25772 9799 25828
rect 9855 25772 9880 25828
rect 9936 25772 9961 25828
rect 10017 25772 10042 25828
rect 10098 25772 10123 25828
rect 10179 25772 10204 25828
rect 10260 25772 10285 25828
rect 10341 25772 10366 25828
rect 10422 25772 10447 25828
rect 10503 25772 10528 25828
rect 10584 25772 10609 25828
rect 10665 25772 10690 25828
rect 10746 25772 10771 25828
rect 10827 25772 10852 25828
rect 10908 25772 10933 25828
rect 10989 25772 11014 25828
rect 11070 25772 11095 25828
rect 11151 25772 11176 25828
rect 11232 25772 11257 25828
rect 11313 25772 11338 25828
rect 11394 25772 11419 25828
rect 11475 25772 11500 25828
rect 5416 25748 11500 25772
rect 5416 25692 5425 25748
rect 5481 25692 5506 25748
rect 5562 25692 5587 25748
rect 5643 25692 5668 25748
rect 5724 25692 5749 25748
rect 5805 25692 5830 25748
rect 5886 25692 5911 25748
rect 5967 25692 5992 25748
rect 6048 25692 6073 25748
rect 6129 25692 6154 25748
rect 6210 25692 6235 25748
rect 6291 25692 6316 25748
rect 6372 25692 6397 25748
rect 6453 25692 6478 25748
rect 6534 25692 6559 25748
rect 6615 25692 6640 25748
rect 6696 25692 6721 25748
rect 6777 25692 6802 25748
rect 6858 25692 6883 25748
rect 6939 25692 6964 25748
rect 7020 25692 7045 25748
rect 7101 25692 7126 25748
rect 7182 25692 7207 25748
rect 7263 25692 7288 25748
rect 7344 25692 7369 25748
rect 7425 25692 7450 25748
rect 7506 25692 7531 25748
rect 7587 25692 7612 25748
rect 7668 25692 7693 25748
rect 7749 25692 7774 25748
rect 7830 25692 7855 25748
rect 7911 25692 7936 25748
rect 7992 25692 8017 25748
rect 8073 25692 8098 25748
rect 8154 25692 8179 25748
rect 8235 25692 8260 25748
rect 8316 25692 8341 25748
rect 8397 25692 8422 25748
rect 8478 25692 8503 25748
rect 8559 25692 8584 25748
rect 8640 25692 8665 25748
rect 8721 25692 8746 25748
rect 8802 25692 8827 25748
rect 8883 25692 8908 25748
rect 8964 25692 8989 25748
rect 9045 25692 9070 25748
rect 9126 25692 9151 25748
rect 9207 25692 9232 25748
rect 9288 25692 9313 25748
rect 9369 25692 9394 25748
rect 9450 25692 9475 25748
rect 9531 25692 9556 25748
rect 9612 25692 9637 25748
rect 9693 25692 9718 25748
rect 9774 25692 9799 25748
rect 9855 25692 9880 25748
rect 9936 25692 9961 25748
rect 10017 25692 10042 25748
rect 10098 25692 10123 25748
rect 10179 25692 10204 25748
rect 10260 25692 10285 25748
rect 10341 25692 10366 25748
rect 10422 25692 10447 25748
rect 10503 25692 10528 25748
rect 10584 25692 10609 25748
rect 10665 25692 10690 25748
rect 10746 25692 10771 25748
rect 10827 25692 10852 25748
rect 10908 25692 10933 25748
rect 10989 25692 11014 25748
rect 11070 25692 11095 25748
rect 11151 25692 11176 25748
rect 11232 25692 11257 25748
rect 11313 25692 11338 25748
rect 11394 25692 11419 25748
rect 11475 25692 11500 25748
rect 5416 25668 11500 25692
rect 5416 25612 5425 25668
rect 5481 25612 5506 25668
rect 5562 25612 5587 25668
rect 5643 25612 5668 25668
rect 5724 25612 5749 25668
rect 5805 25612 5830 25668
rect 5886 25612 5911 25668
rect 5967 25612 5992 25668
rect 6048 25612 6073 25668
rect 6129 25612 6154 25668
rect 6210 25612 6235 25668
rect 6291 25612 6316 25668
rect 6372 25612 6397 25668
rect 6453 25612 6478 25668
rect 6534 25612 6559 25668
rect 6615 25612 6640 25668
rect 6696 25612 6721 25668
rect 6777 25612 6802 25668
rect 6858 25612 6883 25668
rect 6939 25612 6964 25668
rect 7020 25612 7045 25668
rect 7101 25612 7126 25668
rect 7182 25612 7207 25668
rect 7263 25612 7288 25668
rect 7344 25612 7369 25668
rect 7425 25612 7450 25668
rect 7506 25612 7531 25668
rect 7587 25612 7612 25668
rect 7668 25612 7693 25668
rect 7749 25612 7774 25668
rect 7830 25612 7855 25668
rect 7911 25612 7936 25668
rect 7992 25612 8017 25668
rect 8073 25612 8098 25668
rect 8154 25612 8179 25668
rect 8235 25612 8260 25668
rect 8316 25612 8341 25668
rect 8397 25612 8422 25668
rect 8478 25612 8503 25668
rect 8559 25612 8584 25668
rect 8640 25612 8665 25668
rect 8721 25612 8746 25668
rect 8802 25612 8827 25668
rect 8883 25612 8908 25668
rect 8964 25612 8989 25668
rect 9045 25612 9070 25668
rect 9126 25612 9151 25668
rect 9207 25612 9232 25668
rect 9288 25612 9313 25668
rect 9369 25612 9394 25668
rect 9450 25612 9475 25668
rect 9531 25612 9556 25668
rect 9612 25612 9637 25668
rect 9693 25612 9718 25668
rect 9774 25612 9799 25668
rect 9855 25612 9880 25668
rect 9936 25612 9961 25668
rect 10017 25612 10042 25668
rect 10098 25612 10123 25668
rect 10179 25612 10204 25668
rect 10260 25612 10285 25668
rect 10341 25612 10366 25668
rect 10422 25612 10447 25668
rect 10503 25612 10528 25668
rect 10584 25612 10609 25668
rect 10665 25612 10690 25668
rect 10746 25612 10771 25668
rect 10827 25612 10852 25668
rect 10908 25612 10933 25668
rect 10989 25612 11014 25668
rect 11070 25612 11095 25668
rect 11151 25612 11176 25668
rect 11232 25612 11257 25668
rect 11313 25612 11338 25668
rect 11394 25612 11419 25668
rect 11475 25612 11500 25668
rect 5416 25588 11500 25612
rect 5416 25532 5425 25588
rect 5481 25532 5506 25588
rect 5562 25532 5587 25588
rect 5643 25532 5668 25588
rect 5724 25532 5749 25588
rect 5805 25532 5830 25588
rect 5886 25532 5911 25588
rect 5967 25532 5992 25588
rect 6048 25532 6073 25588
rect 6129 25532 6154 25588
rect 6210 25532 6235 25588
rect 6291 25532 6316 25588
rect 6372 25532 6397 25588
rect 6453 25532 6478 25588
rect 6534 25532 6559 25588
rect 6615 25532 6640 25588
rect 6696 25532 6721 25588
rect 6777 25532 6802 25588
rect 6858 25532 6883 25588
rect 6939 25532 6964 25588
rect 7020 25532 7045 25588
rect 7101 25532 7126 25588
rect 7182 25532 7207 25588
rect 7263 25532 7288 25588
rect 7344 25532 7369 25588
rect 7425 25532 7450 25588
rect 7506 25532 7531 25588
rect 7587 25532 7612 25588
rect 7668 25532 7693 25588
rect 7749 25532 7774 25588
rect 7830 25532 7855 25588
rect 7911 25532 7936 25588
rect 7992 25532 8017 25588
rect 8073 25532 8098 25588
rect 8154 25532 8179 25588
rect 8235 25532 8260 25588
rect 8316 25532 8341 25588
rect 8397 25532 8422 25588
rect 8478 25532 8503 25588
rect 8559 25532 8584 25588
rect 8640 25532 8665 25588
rect 8721 25532 8746 25588
rect 8802 25532 8827 25588
rect 8883 25532 8908 25588
rect 8964 25532 8989 25588
rect 9045 25532 9070 25588
rect 9126 25532 9151 25588
rect 9207 25532 9232 25588
rect 9288 25532 9313 25588
rect 9369 25532 9394 25588
rect 9450 25532 9475 25588
rect 9531 25532 9556 25588
rect 9612 25532 9637 25588
rect 9693 25532 9718 25588
rect 9774 25532 9799 25588
rect 9855 25532 9880 25588
rect 9936 25532 9961 25588
rect 10017 25532 10042 25588
rect 10098 25532 10123 25588
rect 10179 25532 10204 25588
rect 10260 25532 10285 25588
rect 10341 25532 10366 25588
rect 10422 25532 10447 25588
rect 10503 25532 10528 25588
rect 10584 25532 10609 25588
rect 10665 25532 10690 25588
rect 10746 25532 10771 25588
rect 10827 25532 10852 25588
rect 10908 25532 10933 25588
rect 10989 25532 11014 25588
rect 11070 25532 11095 25588
rect 11151 25532 11176 25588
rect 11232 25532 11257 25588
rect 11313 25532 11338 25588
rect 11394 25532 11419 25588
rect 11475 25532 11500 25588
rect 5416 25508 11500 25532
rect 5416 25452 5425 25508
rect 5481 25452 5506 25508
rect 5562 25452 5587 25508
rect 5643 25452 5668 25508
rect 5724 25452 5749 25508
rect 5805 25452 5830 25508
rect 5886 25452 5911 25508
rect 5967 25452 5992 25508
rect 6048 25452 6073 25508
rect 6129 25452 6154 25508
rect 6210 25452 6235 25508
rect 6291 25452 6316 25508
rect 6372 25452 6397 25508
rect 6453 25452 6478 25508
rect 6534 25452 6559 25508
rect 6615 25452 6640 25508
rect 6696 25452 6721 25508
rect 6777 25452 6802 25508
rect 6858 25452 6883 25508
rect 6939 25452 6964 25508
rect 7020 25452 7045 25508
rect 7101 25452 7126 25508
rect 7182 25452 7207 25508
rect 7263 25452 7288 25508
rect 7344 25452 7369 25508
rect 7425 25452 7450 25508
rect 7506 25452 7531 25508
rect 7587 25452 7612 25508
rect 7668 25452 7693 25508
rect 7749 25452 7774 25508
rect 7830 25452 7855 25508
rect 7911 25452 7936 25508
rect 7992 25452 8017 25508
rect 8073 25452 8098 25508
rect 8154 25452 8179 25508
rect 8235 25452 8260 25508
rect 8316 25452 8341 25508
rect 8397 25452 8422 25508
rect 8478 25452 8503 25508
rect 8559 25452 8584 25508
rect 8640 25452 8665 25508
rect 8721 25452 8746 25508
rect 8802 25452 8827 25508
rect 8883 25452 8908 25508
rect 8964 25452 8989 25508
rect 9045 25452 9070 25508
rect 9126 25452 9151 25508
rect 9207 25452 9232 25508
rect 9288 25452 9313 25508
rect 9369 25452 9394 25508
rect 9450 25452 9475 25508
rect 9531 25452 9556 25508
rect 9612 25452 9637 25508
rect 9693 25452 9718 25508
rect 9774 25452 9799 25508
rect 9855 25452 9880 25508
rect 9936 25452 9961 25508
rect 10017 25452 10042 25508
rect 10098 25452 10123 25508
rect 10179 25452 10204 25508
rect 10260 25452 10285 25508
rect 10341 25452 10366 25508
rect 10422 25452 10447 25508
rect 10503 25452 10528 25508
rect 10584 25452 10609 25508
rect 10665 25452 10690 25508
rect 10746 25452 10771 25508
rect 10827 25452 10852 25508
rect 10908 25452 10933 25508
rect 10989 25452 11014 25508
rect 11070 25452 11095 25508
rect 11151 25452 11176 25508
rect 11232 25452 11257 25508
rect 11313 25452 11338 25508
rect 11394 25452 11419 25508
rect 11475 25452 11500 25508
rect 5416 25428 11500 25452
rect 5416 25372 5425 25428
rect 5481 25372 5506 25428
rect 5562 25372 5587 25428
rect 5643 25372 5668 25428
rect 5724 25372 5749 25428
rect 5805 25372 5830 25428
rect 5886 25372 5911 25428
rect 5967 25372 5992 25428
rect 6048 25372 6073 25428
rect 6129 25372 6154 25428
rect 6210 25372 6235 25428
rect 6291 25372 6316 25428
rect 6372 25372 6397 25428
rect 6453 25372 6478 25428
rect 6534 25372 6559 25428
rect 6615 25372 6640 25428
rect 6696 25372 6721 25428
rect 6777 25372 6802 25428
rect 6858 25372 6883 25428
rect 6939 25372 6964 25428
rect 7020 25372 7045 25428
rect 7101 25372 7126 25428
rect 7182 25372 7207 25428
rect 7263 25372 7288 25428
rect 7344 25372 7369 25428
rect 7425 25372 7450 25428
rect 7506 25372 7531 25428
rect 7587 25372 7612 25428
rect 7668 25372 7693 25428
rect 7749 25372 7774 25428
rect 7830 25372 7855 25428
rect 7911 25372 7936 25428
rect 7992 25372 8017 25428
rect 8073 25372 8098 25428
rect 8154 25372 8179 25428
rect 8235 25372 8260 25428
rect 8316 25372 8341 25428
rect 8397 25372 8422 25428
rect 8478 25372 8503 25428
rect 8559 25372 8584 25428
rect 8640 25372 8665 25428
rect 8721 25372 8746 25428
rect 8802 25372 8827 25428
rect 8883 25372 8908 25428
rect 8964 25372 8989 25428
rect 9045 25372 9070 25428
rect 9126 25372 9151 25428
rect 9207 25372 9232 25428
rect 9288 25372 9313 25428
rect 9369 25372 9394 25428
rect 9450 25372 9475 25428
rect 9531 25372 9556 25428
rect 9612 25372 9637 25428
rect 9693 25372 9718 25428
rect 9774 25372 9799 25428
rect 9855 25372 9880 25428
rect 9936 25372 9961 25428
rect 10017 25372 10042 25428
rect 10098 25372 10123 25428
rect 10179 25372 10204 25428
rect 10260 25372 10285 25428
rect 10341 25372 10366 25428
rect 10422 25372 10447 25428
rect 10503 25372 10528 25428
rect 10584 25372 10609 25428
rect 10665 25372 10690 25428
rect 10746 25372 10771 25428
rect 10827 25372 10852 25428
rect 10908 25372 10933 25428
rect 10989 25372 11014 25428
rect 11070 25372 11095 25428
rect 11151 25372 11176 25428
rect 11232 25372 11257 25428
rect 11313 25372 11338 25428
rect 11394 25372 11419 25428
rect 11475 25372 11500 25428
rect 5416 25348 11500 25372
rect 5416 25292 5425 25348
rect 5481 25292 5506 25348
rect 5562 25292 5587 25348
rect 5643 25292 5668 25348
rect 5724 25292 5749 25348
rect 5805 25292 5830 25348
rect 5886 25292 5911 25348
rect 5967 25292 5992 25348
rect 6048 25292 6073 25348
rect 6129 25292 6154 25348
rect 6210 25292 6235 25348
rect 6291 25292 6316 25348
rect 6372 25292 6397 25348
rect 6453 25292 6478 25348
rect 6534 25292 6559 25348
rect 6615 25292 6640 25348
rect 6696 25292 6721 25348
rect 6777 25292 6802 25348
rect 6858 25292 6883 25348
rect 6939 25292 6964 25348
rect 7020 25292 7045 25348
rect 7101 25292 7126 25348
rect 7182 25292 7207 25348
rect 7263 25292 7288 25348
rect 7344 25292 7369 25348
rect 7425 25292 7450 25348
rect 7506 25292 7531 25348
rect 7587 25292 7612 25348
rect 7668 25292 7693 25348
rect 7749 25292 7774 25348
rect 7830 25292 7855 25348
rect 7911 25292 7936 25348
rect 7992 25292 8017 25348
rect 8073 25292 8098 25348
rect 8154 25292 8179 25348
rect 8235 25292 8260 25348
rect 8316 25292 8341 25348
rect 8397 25292 8422 25348
rect 8478 25292 8503 25348
rect 8559 25292 8584 25348
rect 8640 25292 8665 25348
rect 8721 25292 8746 25348
rect 8802 25292 8827 25348
rect 8883 25292 8908 25348
rect 8964 25292 8989 25348
rect 9045 25292 9070 25348
rect 9126 25292 9151 25348
rect 9207 25292 9232 25348
rect 9288 25292 9313 25348
rect 9369 25292 9394 25348
rect 9450 25292 9475 25348
rect 9531 25292 9556 25348
rect 9612 25292 9637 25348
rect 9693 25292 9718 25348
rect 9774 25292 9799 25348
rect 9855 25292 9880 25348
rect 9936 25292 9961 25348
rect 10017 25292 10042 25348
rect 10098 25292 10123 25348
rect 10179 25292 10204 25348
rect 10260 25292 10285 25348
rect 10341 25292 10366 25348
rect 10422 25292 10447 25348
rect 10503 25292 10528 25348
rect 10584 25292 10609 25348
rect 10665 25292 10690 25348
rect 10746 25292 10771 25348
rect 10827 25292 10852 25348
rect 10908 25292 10933 25348
rect 10989 25292 11014 25348
rect 11070 25292 11095 25348
rect 11151 25292 11176 25348
rect 11232 25292 11257 25348
rect 11313 25292 11338 25348
rect 11394 25292 11419 25348
rect 11475 25292 11500 25348
rect 5416 25268 11500 25292
rect 5416 25212 5425 25268
rect 5481 25212 5506 25268
rect 5562 25212 5587 25268
rect 5643 25212 5668 25268
rect 5724 25212 5749 25268
rect 5805 25212 5830 25268
rect 5886 25212 5911 25268
rect 5967 25212 5992 25268
rect 6048 25212 6073 25268
rect 6129 25212 6154 25268
rect 6210 25212 6235 25268
rect 6291 25212 6316 25268
rect 6372 25212 6397 25268
rect 6453 25212 6478 25268
rect 6534 25212 6559 25268
rect 6615 25212 6640 25268
rect 6696 25212 6721 25268
rect 6777 25212 6802 25268
rect 6858 25212 6883 25268
rect 6939 25212 6964 25268
rect 7020 25212 7045 25268
rect 7101 25212 7126 25268
rect 7182 25212 7207 25268
rect 7263 25212 7288 25268
rect 7344 25212 7369 25268
rect 7425 25212 7450 25268
rect 7506 25212 7531 25268
rect 7587 25212 7612 25268
rect 7668 25212 7693 25268
rect 7749 25212 7774 25268
rect 7830 25212 7855 25268
rect 7911 25212 7936 25268
rect 7992 25212 8017 25268
rect 8073 25212 8098 25268
rect 8154 25212 8179 25268
rect 8235 25212 8260 25268
rect 8316 25212 8341 25268
rect 8397 25212 8422 25268
rect 8478 25212 8503 25268
rect 8559 25212 8584 25268
rect 8640 25212 8665 25268
rect 8721 25212 8746 25268
rect 8802 25212 8827 25268
rect 8883 25212 8908 25268
rect 8964 25212 8989 25268
rect 9045 25212 9070 25268
rect 9126 25212 9151 25268
rect 9207 25212 9232 25268
rect 9288 25212 9313 25268
rect 9369 25212 9394 25268
rect 9450 25212 9475 25268
rect 9531 25212 9556 25268
rect 9612 25212 9637 25268
rect 9693 25212 9718 25268
rect 9774 25212 9799 25268
rect 9855 25212 9880 25268
rect 9936 25212 9961 25268
rect 10017 25212 10042 25268
rect 10098 25212 10123 25268
rect 10179 25212 10204 25268
rect 10260 25212 10285 25268
rect 10341 25212 10366 25268
rect 10422 25212 10447 25268
rect 10503 25212 10528 25268
rect 10584 25212 10609 25268
rect 10665 25212 10690 25268
rect 10746 25212 10771 25268
rect 10827 25212 10852 25268
rect 10908 25212 10933 25268
rect 10989 25212 11014 25268
rect 11070 25212 11095 25268
rect 11151 25212 11176 25268
rect 11232 25212 11257 25268
rect 11313 25212 11338 25268
rect 11394 25212 11419 25268
rect 11475 25212 11500 25268
rect 5416 25188 11500 25212
rect 5416 25132 5425 25188
rect 5481 25132 5506 25188
rect 5562 25132 5587 25188
rect 5643 25132 5668 25188
rect 5724 25132 5749 25188
rect 5805 25132 5830 25188
rect 5886 25132 5911 25188
rect 5967 25132 5992 25188
rect 6048 25132 6073 25188
rect 6129 25132 6154 25188
rect 6210 25132 6235 25188
rect 6291 25132 6316 25188
rect 6372 25132 6397 25188
rect 6453 25132 6478 25188
rect 6534 25132 6559 25188
rect 6615 25132 6640 25188
rect 6696 25132 6721 25188
rect 6777 25132 6802 25188
rect 6858 25132 6883 25188
rect 6939 25132 6964 25188
rect 7020 25132 7045 25188
rect 7101 25132 7126 25188
rect 7182 25132 7207 25188
rect 7263 25132 7288 25188
rect 7344 25132 7369 25188
rect 7425 25132 7450 25188
rect 7506 25132 7531 25188
rect 7587 25132 7612 25188
rect 7668 25132 7693 25188
rect 7749 25132 7774 25188
rect 7830 25132 7855 25188
rect 7911 25132 7936 25188
rect 7992 25132 8017 25188
rect 8073 25132 8098 25188
rect 8154 25132 8179 25188
rect 8235 25132 8260 25188
rect 8316 25132 8341 25188
rect 8397 25132 8422 25188
rect 8478 25132 8503 25188
rect 8559 25132 8584 25188
rect 8640 25132 8665 25188
rect 8721 25132 8746 25188
rect 8802 25132 8827 25188
rect 8883 25132 8908 25188
rect 8964 25132 8989 25188
rect 9045 25132 9070 25188
rect 9126 25132 9151 25188
rect 9207 25132 9232 25188
rect 9288 25132 9313 25188
rect 9369 25132 9394 25188
rect 9450 25132 9475 25188
rect 9531 25132 9556 25188
rect 9612 25132 9637 25188
rect 9693 25132 9718 25188
rect 9774 25132 9799 25188
rect 9855 25132 9880 25188
rect 9936 25132 9961 25188
rect 10017 25132 10042 25188
rect 10098 25132 10123 25188
rect 10179 25132 10204 25188
rect 10260 25132 10285 25188
rect 10341 25132 10366 25188
rect 10422 25132 10447 25188
rect 10503 25132 10528 25188
rect 10584 25132 10609 25188
rect 10665 25132 10690 25188
rect 10746 25132 10771 25188
rect 10827 25132 10852 25188
rect 10908 25132 10933 25188
rect 10989 25132 11014 25188
rect 11070 25132 11095 25188
rect 11151 25132 11176 25188
rect 11232 25132 11257 25188
rect 11313 25132 11338 25188
rect 11394 25132 11419 25188
rect 11475 25132 11500 25188
rect 5416 25108 11500 25132
rect 5416 25052 5425 25108
rect 5481 25052 5506 25108
rect 5562 25052 5587 25108
rect 5643 25052 5668 25108
rect 5724 25052 5749 25108
rect 5805 25052 5830 25108
rect 5886 25052 5911 25108
rect 5967 25052 5992 25108
rect 6048 25052 6073 25108
rect 6129 25052 6154 25108
rect 6210 25052 6235 25108
rect 6291 25052 6316 25108
rect 6372 25052 6397 25108
rect 6453 25052 6478 25108
rect 6534 25052 6559 25108
rect 6615 25052 6640 25108
rect 6696 25052 6721 25108
rect 6777 25052 6802 25108
rect 6858 25052 6883 25108
rect 6939 25052 6964 25108
rect 7020 25052 7045 25108
rect 7101 25052 7126 25108
rect 7182 25052 7207 25108
rect 7263 25052 7288 25108
rect 7344 25052 7369 25108
rect 7425 25052 7450 25108
rect 7506 25052 7531 25108
rect 7587 25052 7612 25108
rect 7668 25052 7693 25108
rect 7749 25052 7774 25108
rect 7830 25052 7855 25108
rect 7911 25052 7936 25108
rect 7992 25052 8017 25108
rect 8073 25052 8098 25108
rect 8154 25052 8179 25108
rect 8235 25052 8260 25108
rect 8316 25052 8341 25108
rect 8397 25052 8422 25108
rect 8478 25052 8503 25108
rect 8559 25052 8584 25108
rect 8640 25052 8665 25108
rect 8721 25052 8746 25108
rect 8802 25052 8827 25108
rect 8883 25052 8908 25108
rect 8964 25052 8989 25108
rect 9045 25052 9070 25108
rect 9126 25052 9151 25108
rect 9207 25052 9232 25108
rect 9288 25052 9313 25108
rect 9369 25052 9394 25108
rect 9450 25052 9475 25108
rect 9531 25052 9556 25108
rect 9612 25052 9637 25108
rect 9693 25052 9718 25108
rect 9774 25052 9799 25108
rect 9855 25052 9880 25108
rect 9936 25052 9961 25108
rect 10017 25052 10042 25108
rect 10098 25052 10123 25108
rect 10179 25052 10204 25108
rect 10260 25052 10285 25108
rect 10341 25052 10366 25108
rect 10422 25052 10447 25108
rect 10503 25052 10528 25108
rect 10584 25052 10609 25108
rect 10665 25052 10690 25108
rect 10746 25052 10771 25108
rect 10827 25052 10852 25108
rect 10908 25052 10933 25108
rect 10989 25052 11014 25108
rect 11070 25052 11095 25108
rect 11151 25052 11176 25108
rect 11232 25052 11257 25108
rect 11313 25052 11338 25108
rect 11394 25052 11419 25108
rect 11475 25052 11500 25108
rect 5416 25028 11500 25052
rect 5416 24972 5425 25028
rect 5481 24972 5506 25028
rect 5562 24972 5587 25028
rect 5643 24972 5668 25028
rect 5724 24972 5749 25028
rect 5805 24972 5830 25028
rect 5886 24972 5911 25028
rect 5967 24972 5992 25028
rect 6048 24972 6073 25028
rect 6129 24972 6154 25028
rect 6210 24972 6235 25028
rect 6291 24972 6316 25028
rect 6372 24972 6397 25028
rect 6453 24972 6478 25028
rect 6534 24972 6559 25028
rect 6615 24972 6640 25028
rect 6696 24972 6721 25028
rect 6777 24972 6802 25028
rect 6858 24972 6883 25028
rect 6939 24972 6964 25028
rect 7020 24972 7045 25028
rect 7101 24972 7126 25028
rect 7182 24972 7207 25028
rect 7263 24972 7288 25028
rect 7344 24972 7369 25028
rect 7425 24972 7450 25028
rect 7506 24972 7531 25028
rect 7587 24972 7612 25028
rect 7668 24972 7693 25028
rect 7749 24972 7774 25028
rect 7830 24972 7855 25028
rect 7911 24972 7936 25028
rect 7992 24972 8017 25028
rect 8073 24972 8098 25028
rect 8154 24972 8179 25028
rect 8235 24972 8260 25028
rect 8316 24972 8341 25028
rect 8397 24972 8422 25028
rect 8478 24972 8503 25028
rect 8559 24972 8584 25028
rect 8640 24972 8665 25028
rect 8721 24972 8746 25028
rect 8802 24972 8827 25028
rect 8883 24972 8908 25028
rect 8964 24972 8989 25028
rect 9045 24972 9070 25028
rect 9126 24972 9151 25028
rect 9207 24972 9232 25028
rect 9288 24972 9313 25028
rect 9369 24972 9394 25028
rect 9450 24972 9475 25028
rect 9531 24972 9556 25028
rect 9612 24972 9637 25028
rect 9693 24972 9718 25028
rect 9774 24972 9799 25028
rect 9855 24972 9880 25028
rect 9936 24972 9961 25028
rect 10017 24972 10042 25028
rect 10098 24972 10123 25028
rect 10179 24972 10204 25028
rect 10260 24972 10285 25028
rect 10341 24972 10366 25028
rect 10422 24972 10447 25028
rect 10503 24972 10528 25028
rect 10584 24972 10609 25028
rect 10665 24972 10690 25028
rect 10746 24972 10771 25028
rect 10827 24972 10852 25028
rect 10908 24972 10933 25028
rect 10989 24972 11014 25028
rect 11070 24972 11095 25028
rect 11151 24972 11176 25028
rect 11232 24972 11257 25028
rect 11313 24972 11338 25028
rect 11394 24972 11419 25028
rect 11475 24972 11500 25028
rect 5416 24948 11500 24972
rect 5416 24892 5425 24948
rect 5481 24892 5506 24948
rect 5562 24892 5587 24948
rect 5643 24892 5668 24948
rect 5724 24892 5749 24948
rect 5805 24892 5830 24948
rect 5886 24892 5911 24948
rect 5967 24892 5992 24948
rect 6048 24892 6073 24948
rect 6129 24892 6154 24948
rect 6210 24892 6235 24948
rect 6291 24892 6316 24948
rect 6372 24892 6397 24948
rect 6453 24892 6478 24948
rect 6534 24892 6559 24948
rect 6615 24892 6640 24948
rect 6696 24892 6721 24948
rect 6777 24892 6802 24948
rect 6858 24892 6883 24948
rect 6939 24892 6964 24948
rect 7020 24892 7045 24948
rect 7101 24892 7126 24948
rect 7182 24892 7207 24948
rect 7263 24892 7288 24948
rect 7344 24892 7369 24948
rect 7425 24892 7450 24948
rect 7506 24892 7531 24948
rect 7587 24892 7612 24948
rect 7668 24892 7693 24948
rect 7749 24892 7774 24948
rect 7830 24892 7855 24948
rect 7911 24892 7936 24948
rect 7992 24892 8017 24948
rect 8073 24892 8098 24948
rect 8154 24892 8179 24948
rect 8235 24892 8260 24948
rect 8316 24892 8341 24948
rect 8397 24892 8422 24948
rect 8478 24892 8503 24948
rect 8559 24892 8584 24948
rect 8640 24892 8665 24948
rect 8721 24892 8746 24948
rect 8802 24892 8827 24948
rect 8883 24892 8908 24948
rect 8964 24892 8989 24948
rect 9045 24892 9070 24948
rect 9126 24892 9151 24948
rect 9207 24892 9232 24948
rect 9288 24892 9313 24948
rect 9369 24892 9394 24948
rect 9450 24892 9475 24948
rect 9531 24892 9556 24948
rect 9612 24892 9637 24948
rect 9693 24892 9718 24948
rect 9774 24892 9799 24948
rect 9855 24892 9880 24948
rect 9936 24892 9961 24948
rect 10017 24892 10042 24948
rect 10098 24892 10123 24948
rect 10179 24892 10204 24948
rect 10260 24892 10285 24948
rect 10341 24892 10366 24948
rect 10422 24892 10447 24948
rect 10503 24892 10528 24948
rect 10584 24892 10609 24948
rect 10665 24892 10690 24948
rect 10746 24892 10771 24948
rect 10827 24892 10852 24948
rect 10908 24892 10933 24948
rect 10989 24892 11014 24948
rect 11070 24892 11095 24948
rect 11151 24892 11176 24948
rect 11232 24892 11257 24948
rect 11313 24892 11338 24948
rect 11394 24892 11419 24948
rect 11475 24892 11500 24948
rect 5416 24868 11500 24892
rect 5416 24812 5425 24868
rect 5481 24812 5506 24868
rect 5562 24812 5587 24868
rect 5643 24812 5668 24868
rect 5724 24812 5749 24868
rect 5805 24812 5830 24868
rect 5886 24812 5911 24868
rect 5967 24812 5992 24868
rect 6048 24812 6073 24868
rect 6129 24812 6154 24868
rect 6210 24812 6235 24868
rect 6291 24812 6316 24868
rect 6372 24812 6397 24868
rect 6453 24812 6478 24868
rect 6534 24812 6559 24868
rect 6615 24812 6640 24868
rect 6696 24812 6721 24868
rect 6777 24812 6802 24868
rect 6858 24812 6883 24868
rect 6939 24812 6964 24868
rect 7020 24812 7045 24868
rect 7101 24812 7126 24868
rect 7182 24812 7207 24868
rect 7263 24812 7288 24868
rect 7344 24812 7369 24868
rect 7425 24812 7450 24868
rect 7506 24812 7531 24868
rect 7587 24812 7612 24868
rect 7668 24812 7693 24868
rect 7749 24812 7774 24868
rect 7830 24812 7855 24868
rect 7911 24812 7936 24868
rect 7992 24812 8017 24868
rect 8073 24812 8098 24868
rect 8154 24812 8179 24868
rect 8235 24812 8260 24868
rect 8316 24812 8341 24868
rect 8397 24812 8422 24868
rect 8478 24812 8503 24868
rect 8559 24812 8584 24868
rect 8640 24812 8665 24868
rect 8721 24812 8746 24868
rect 8802 24812 8827 24868
rect 8883 24812 8908 24868
rect 8964 24812 8989 24868
rect 9045 24812 9070 24868
rect 9126 24812 9151 24868
rect 9207 24812 9232 24868
rect 9288 24812 9313 24868
rect 9369 24812 9394 24868
rect 9450 24812 9475 24868
rect 9531 24812 9556 24868
rect 9612 24812 9637 24868
rect 9693 24812 9718 24868
rect 9774 24812 9799 24868
rect 9855 24812 9880 24868
rect 9936 24812 9961 24868
rect 10017 24812 10042 24868
rect 10098 24812 10123 24868
rect 10179 24812 10204 24868
rect 10260 24812 10285 24868
rect 10341 24812 10366 24868
rect 10422 24812 10447 24868
rect 10503 24812 10528 24868
rect 10584 24812 10609 24868
rect 10665 24812 10690 24868
rect 10746 24812 10771 24868
rect 10827 24812 10852 24868
rect 10908 24812 10933 24868
rect 10989 24812 11014 24868
rect 11070 24812 11095 24868
rect 11151 24812 11176 24868
rect 11232 24812 11257 24868
rect 11313 24812 11338 24868
rect 11394 24812 11419 24868
rect 11475 24812 11500 24868
rect 5416 24788 11500 24812
rect 5416 24732 5425 24788
rect 5481 24732 5506 24788
rect 5562 24732 5587 24788
rect 5643 24732 5668 24788
rect 5724 24732 5749 24788
rect 5805 24732 5830 24788
rect 5886 24732 5911 24788
rect 5967 24732 5992 24788
rect 6048 24732 6073 24788
rect 6129 24732 6154 24788
rect 6210 24732 6235 24788
rect 6291 24732 6316 24788
rect 6372 24732 6397 24788
rect 6453 24732 6478 24788
rect 6534 24732 6559 24788
rect 6615 24732 6640 24788
rect 6696 24732 6721 24788
rect 6777 24732 6802 24788
rect 6858 24732 6883 24788
rect 6939 24732 6964 24788
rect 7020 24732 7045 24788
rect 7101 24732 7126 24788
rect 7182 24732 7207 24788
rect 7263 24732 7288 24788
rect 7344 24732 7369 24788
rect 7425 24732 7450 24788
rect 7506 24732 7531 24788
rect 7587 24732 7612 24788
rect 7668 24732 7693 24788
rect 7749 24732 7774 24788
rect 7830 24732 7855 24788
rect 7911 24732 7936 24788
rect 7992 24732 8017 24788
rect 8073 24732 8098 24788
rect 8154 24732 8179 24788
rect 8235 24732 8260 24788
rect 8316 24732 8341 24788
rect 8397 24732 8422 24788
rect 8478 24732 8503 24788
rect 8559 24732 8584 24788
rect 8640 24732 8665 24788
rect 8721 24732 8746 24788
rect 8802 24732 8827 24788
rect 8883 24732 8908 24788
rect 8964 24732 8989 24788
rect 9045 24732 9070 24788
rect 9126 24732 9151 24788
rect 9207 24732 9232 24788
rect 9288 24732 9313 24788
rect 9369 24732 9394 24788
rect 9450 24732 9475 24788
rect 9531 24732 9556 24788
rect 9612 24732 9637 24788
rect 9693 24732 9718 24788
rect 9774 24732 9799 24788
rect 9855 24732 9880 24788
rect 9936 24732 9961 24788
rect 10017 24732 10042 24788
rect 10098 24732 10123 24788
rect 10179 24732 10204 24788
rect 10260 24732 10285 24788
rect 10341 24732 10366 24788
rect 10422 24732 10447 24788
rect 10503 24732 10528 24788
rect 10584 24732 10609 24788
rect 10665 24732 10690 24788
rect 10746 24732 10771 24788
rect 10827 24732 10852 24788
rect 10908 24732 10933 24788
rect 10989 24732 11014 24788
rect 11070 24732 11095 24788
rect 11151 24732 11176 24788
rect 11232 24732 11257 24788
rect 11313 24732 11338 24788
rect 11394 24732 11419 24788
rect 11475 24732 11500 24788
rect 5416 24708 11500 24732
rect 5416 24652 5425 24708
rect 5481 24652 5506 24708
rect 5562 24652 5587 24708
rect 5643 24652 5668 24708
rect 5724 24652 5749 24708
rect 5805 24652 5830 24708
rect 5886 24652 5911 24708
rect 5967 24652 5992 24708
rect 6048 24652 6073 24708
rect 6129 24652 6154 24708
rect 6210 24652 6235 24708
rect 6291 24652 6316 24708
rect 6372 24652 6397 24708
rect 6453 24652 6478 24708
rect 6534 24652 6559 24708
rect 6615 24652 6640 24708
rect 6696 24652 6721 24708
rect 6777 24652 6802 24708
rect 6858 24652 6883 24708
rect 6939 24652 6964 24708
rect 7020 24652 7045 24708
rect 7101 24652 7126 24708
rect 7182 24652 7207 24708
rect 7263 24652 7288 24708
rect 7344 24652 7369 24708
rect 7425 24652 7450 24708
rect 7506 24652 7531 24708
rect 7587 24652 7612 24708
rect 7668 24652 7693 24708
rect 7749 24652 7774 24708
rect 7830 24652 7855 24708
rect 7911 24652 7936 24708
rect 7992 24652 8017 24708
rect 8073 24652 8098 24708
rect 8154 24652 8179 24708
rect 8235 24652 8260 24708
rect 8316 24652 8341 24708
rect 8397 24652 8422 24708
rect 8478 24652 8503 24708
rect 8559 24652 8584 24708
rect 8640 24652 8665 24708
rect 8721 24652 8746 24708
rect 8802 24652 8827 24708
rect 8883 24652 8908 24708
rect 8964 24652 8989 24708
rect 9045 24652 9070 24708
rect 9126 24652 9151 24708
rect 9207 24652 9232 24708
rect 9288 24652 9313 24708
rect 9369 24652 9394 24708
rect 9450 24652 9475 24708
rect 9531 24652 9556 24708
rect 9612 24652 9637 24708
rect 9693 24652 9718 24708
rect 9774 24652 9799 24708
rect 9855 24652 9880 24708
rect 9936 24652 9961 24708
rect 10017 24652 10042 24708
rect 10098 24652 10123 24708
rect 10179 24652 10204 24708
rect 10260 24652 10285 24708
rect 10341 24652 10366 24708
rect 10422 24652 10447 24708
rect 10503 24652 10528 24708
rect 10584 24652 10609 24708
rect 10665 24652 10690 24708
rect 10746 24652 10771 24708
rect 10827 24652 10852 24708
rect 10908 24652 10933 24708
rect 10989 24652 11014 24708
rect 11070 24652 11095 24708
rect 11151 24652 11176 24708
rect 11232 24652 11257 24708
rect 11313 24652 11338 24708
rect 11394 24652 11419 24708
rect 11475 24652 11500 24708
rect 13076 24652 13085 25828
rect 5416 24641 13085 24652
rect 5416 24323 13085 24334
rect 5416 24267 5425 24323
rect 5481 24267 5506 24323
rect 5562 24267 5587 24323
rect 5643 24267 5668 24323
rect 5724 24267 5749 24323
rect 5805 24267 5830 24323
rect 5886 24267 5911 24323
rect 5967 24267 5992 24323
rect 6048 24267 6073 24323
rect 6129 24267 6154 24323
rect 6210 24267 6235 24323
rect 6291 24267 6316 24323
rect 6372 24267 6397 24323
rect 6453 24267 6478 24323
rect 6534 24267 6559 24323
rect 6615 24267 6640 24323
rect 6696 24267 6721 24323
rect 6777 24267 6802 24323
rect 6858 24267 6883 24323
rect 6939 24267 6964 24323
rect 7020 24267 7045 24323
rect 7101 24267 7126 24323
rect 7182 24267 7207 24323
rect 7263 24267 7288 24323
rect 7344 24267 7369 24323
rect 7425 24267 7450 24323
rect 7506 24267 7531 24323
rect 7587 24267 7612 24323
rect 7668 24267 7693 24323
rect 7749 24267 7774 24323
rect 7830 24267 7855 24323
rect 7911 24267 7936 24323
rect 7992 24267 8017 24323
rect 8073 24267 8098 24323
rect 8154 24267 8179 24323
rect 8235 24267 8260 24323
rect 8316 24267 8341 24323
rect 8397 24267 8422 24323
rect 8478 24267 8503 24323
rect 8559 24267 8584 24323
rect 8640 24267 8665 24323
rect 8721 24267 8746 24323
rect 8802 24267 8827 24323
rect 8883 24267 8908 24323
rect 8964 24267 8989 24323
rect 9045 24267 9070 24323
rect 9126 24267 9151 24323
rect 9207 24267 9232 24323
rect 9288 24267 9313 24323
rect 9369 24267 9394 24323
rect 9450 24267 9475 24323
rect 9531 24267 9556 24323
rect 9612 24267 9637 24323
rect 9693 24267 9718 24323
rect 9774 24267 9799 24323
rect 9855 24267 9880 24323
rect 9936 24267 9961 24323
rect 10017 24267 10042 24323
rect 10098 24267 10123 24323
rect 10179 24267 10204 24323
rect 10260 24267 10285 24323
rect 10341 24267 10366 24323
rect 10422 24267 10447 24323
rect 10503 24267 10528 24323
rect 10584 24267 10609 24323
rect 10665 24267 10690 24323
rect 10746 24267 10771 24323
rect 10827 24267 10852 24323
rect 10908 24267 10933 24323
rect 10989 24267 11014 24323
rect 11070 24267 11095 24323
rect 11151 24267 11176 24323
rect 11232 24267 11257 24323
rect 11313 24267 11338 24323
rect 11394 24267 11419 24323
rect 11475 24267 11500 24323
rect 5416 24243 11500 24267
rect 5416 24187 5425 24243
rect 5481 24187 5506 24243
rect 5562 24187 5587 24243
rect 5643 24187 5668 24243
rect 5724 24187 5749 24243
rect 5805 24187 5830 24243
rect 5886 24187 5911 24243
rect 5967 24187 5992 24243
rect 6048 24187 6073 24243
rect 6129 24187 6154 24243
rect 6210 24187 6235 24243
rect 6291 24187 6316 24243
rect 6372 24187 6397 24243
rect 6453 24187 6478 24243
rect 6534 24187 6559 24243
rect 6615 24187 6640 24243
rect 6696 24187 6721 24243
rect 6777 24187 6802 24243
rect 6858 24187 6883 24243
rect 6939 24187 6964 24243
rect 7020 24187 7045 24243
rect 7101 24187 7126 24243
rect 7182 24187 7207 24243
rect 7263 24187 7288 24243
rect 7344 24187 7369 24243
rect 7425 24187 7450 24243
rect 7506 24187 7531 24243
rect 7587 24187 7612 24243
rect 7668 24187 7693 24243
rect 7749 24187 7774 24243
rect 7830 24187 7855 24243
rect 7911 24187 7936 24243
rect 7992 24187 8017 24243
rect 8073 24187 8098 24243
rect 8154 24187 8179 24243
rect 8235 24187 8260 24243
rect 8316 24187 8341 24243
rect 8397 24187 8422 24243
rect 8478 24187 8503 24243
rect 8559 24187 8584 24243
rect 8640 24187 8665 24243
rect 8721 24187 8746 24243
rect 8802 24187 8827 24243
rect 8883 24187 8908 24243
rect 8964 24187 8989 24243
rect 9045 24187 9070 24243
rect 9126 24187 9151 24243
rect 9207 24187 9232 24243
rect 9288 24187 9313 24243
rect 9369 24187 9394 24243
rect 9450 24187 9475 24243
rect 9531 24187 9556 24243
rect 9612 24187 9637 24243
rect 9693 24187 9718 24243
rect 9774 24187 9799 24243
rect 9855 24187 9880 24243
rect 9936 24187 9961 24243
rect 10017 24187 10042 24243
rect 10098 24187 10123 24243
rect 10179 24187 10204 24243
rect 10260 24187 10285 24243
rect 10341 24187 10366 24243
rect 10422 24187 10447 24243
rect 10503 24187 10528 24243
rect 10584 24187 10609 24243
rect 10665 24187 10690 24243
rect 10746 24187 10771 24243
rect 10827 24187 10852 24243
rect 10908 24187 10933 24243
rect 10989 24187 11014 24243
rect 11070 24187 11095 24243
rect 11151 24187 11176 24243
rect 11232 24187 11257 24243
rect 11313 24187 11338 24243
rect 11394 24187 11419 24243
rect 11475 24187 11500 24243
rect 5416 24163 11500 24187
rect 5416 24107 5425 24163
rect 5481 24107 5506 24163
rect 5562 24107 5587 24163
rect 5643 24107 5668 24163
rect 5724 24107 5749 24163
rect 5805 24107 5830 24163
rect 5886 24107 5911 24163
rect 5967 24107 5992 24163
rect 6048 24107 6073 24163
rect 6129 24107 6154 24163
rect 6210 24107 6235 24163
rect 6291 24107 6316 24163
rect 6372 24107 6397 24163
rect 6453 24107 6478 24163
rect 6534 24107 6559 24163
rect 6615 24107 6640 24163
rect 6696 24107 6721 24163
rect 6777 24107 6802 24163
rect 6858 24107 6883 24163
rect 6939 24107 6964 24163
rect 7020 24107 7045 24163
rect 7101 24107 7126 24163
rect 7182 24107 7207 24163
rect 7263 24107 7288 24163
rect 7344 24107 7369 24163
rect 7425 24107 7450 24163
rect 7506 24107 7531 24163
rect 7587 24107 7612 24163
rect 7668 24107 7693 24163
rect 7749 24107 7774 24163
rect 7830 24107 7855 24163
rect 7911 24107 7936 24163
rect 7992 24107 8017 24163
rect 8073 24107 8098 24163
rect 8154 24107 8179 24163
rect 8235 24107 8260 24163
rect 8316 24107 8341 24163
rect 8397 24107 8422 24163
rect 8478 24107 8503 24163
rect 8559 24107 8584 24163
rect 8640 24107 8665 24163
rect 8721 24107 8746 24163
rect 8802 24107 8827 24163
rect 8883 24107 8908 24163
rect 8964 24107 8989 24163
rect 9045 24107 9070 24163
rect 9126 24107 9151 24163
rect 9207 24107 9232 24163
rect 9288 24107 9313 24163
rect 9369 24107 9394 24163
rect 9450 24107 9475 24163
rect 9531 24107 9556 24163
rect 9612 24107 9637 24163
rect 9693 24107 9718 24163
rect 9774 24107 9799 24163
rect 9855 24107 9880 24163
rect 9936 24107 9961 24163
rect 10017 24107 10042 24163
rect 10098 24107 10123 24163
rect 10179 24107 10204 24163
rect 10260 24107 10285 24163
rect 10341 24107 10366 24163
rect 10422 24107 10447 24163
rect 10503 24107 10528 24163
rect 10584 24107 10609 24163
rect 10665 24107 10690 24163
rect 10746 24107 10771 24163
rect 10827 24107 10852 24163
rect 10908 24107 10933 24163
rect 10989 24107 11014 24163
rect 11070 24107 11095 24163
rect 11151 24107 11176 24163
rect 11232 24107 11257 24163
rect 11313 24107 11338 24163
rect 11394 24107 11419 24163
rect 11475 24107 11500 24163
rect 5416 24083 11500 24107
rect 5416 24027 5425 24083
rect 5481 24027 5506 24083
rect 5562 24027 5587 24083
rect 5643 24027 5668 24083
rect 5724 24027 5749 24083
rect 5805 24027 5830 24083
rect 5886 24027 5911 24083
rect 5967 24027 5992 24083
rect 6048 24027 6073 24083
rect 6129 24027 6154 24083
rect 6210 24027 6235 24083
rect 6291 24027 6316 24083
rect 6372 24027 6397 24083
rect 6453 24027 6478 24083
rect 6534 24027 6559 24083
rect 6615 24027 6640 24083
rect 6696 24027 6721 24083
rect 6777 24027 6802 24083
rect 6858 24027 6883 24083
rect 6939 24027 6964 24083
rect 7020 24027 7045 24083
rect 7101 24027 7126 24083
rect 7182 24027 7207 24083
rect 7263 24027 7288 24083
rect 7344 24027 7369 24083
rect 7425 24027 7450 24083
rect 7506 24027 7531 24083
rect 7587 24027 7612 24083
rect 7668 24027 7693 24083
rect 7749 24027 7774 24083
rect 7830 24027 7855 24083
rect 7911 24027 7936 24083
rect 7992 24027 8017 24083
rect 8073 24027 8098 24083
rect 8154 24027 8179 24083
rect 8235 24027 8260 24083
rect 8316 24027 8341 24083
rect 8397 24027 8422 24083
rect 8478 24027 8503 24083
rect 8559 24027 8584 24083
rect 8640 24027 8665 24083
rect 8721 24027 8746 24083
rect 8802 24027 8827 24083
rect 8883 24027 8908 24083
rect 8964 24027 8989 24083
rect 9045 24027 9070 24083
rect 9126 24027 9151 24083
rect 9207 24027 9232 24083
rect 9288 24027 9313 24083
rect 9369 24027 9394 24083
rect 9450 24027 9475 24083
rect 9531 24027 9556 24083
rect 9612 24027 9637 24083
rect 9693 24027 9718 24083
rect 9774 24027 9799 24083
rect 9855 24027 9880 24083
rect 9936 24027 9961 24083
rect 10017 24027 10042 24083
rect 10098 24027 10123 24083
rect 10179 24027 10204 24083
rect 10260 24027 10285 24083
rect 10341 24027 10366 24083
rect 10422 24027 10447 24083
rect 10503 24027 10528 24083
rect 10584 24027 10609 24083
rect 10665 24027 10690 24083
rect 10746 24027 10771 24083
rect 10827 24027 10852 24083
rect 10908 24027 10933 24083
rect 10989 24027 11014 24083
rect 11070 24027 11095 24083
rect 11151 24027 11176 24083
rect 11232 24027 11257 24083
rect 11313 24027 11338 24083
rect 11394 24027 11419 24083
rect 11475 24027 11500 24083
rect 5416 24003 11500 24027
rect 5416 23947 5425 24003
rect 5481 23947 5506 24003
rect 5562 23947 5587 24003
rect 5643 23947 5668 24003
rect 5724 23947 5749 24003
rect 5805 23947 5830 24003
rect 5886 23947 5911 24003
rect 5967 23947 5992 24003
rect 6048 23947 6073 24003
rect 6129 23947 6154 24003
rect 6210 23947 6235 24003
rect 6291 23947 6316 24003
rect 6372 23947 6397 24003
rect 6453 23947 6478 24003
rect 6534 23947 6559 24003
rect 6615 23947 6640 24003
rect 6696 23947 6721 24003
rect 6777 23947 6802 24003
rect 6858 23947 6883 24003
rect 6939 23947 6964 24003
rect 7020 23947 7045 24003
rect 7101 23947 7126 24003
rect 7182 23947 7207 24003
rect 7263 23947 7288 24003
rect 7344 23947 7369 24003
rect 7425 23947 7450 24003
rect 7506 23947 7531 24003
rect 7587 23947 7612 24003
rect 7668 23947 7693 24003
rect 7749 23947 7774 24003
rect 7830 23947 7855 24003
rect 7911 23947 7936 24003
rect 7992 23947 8017 24003
rect 8073 23947 8098 24003
rect 8154 23947 8179 24003
rect 8235 23947 8260 24003
rect 8316 23947 8341 24003
rect 8397 23947 8422 24003
rect 8478 23947 8503 24003
rect 8559 23947 8584 24003
rect 8640 23947 8665 24003
rect 8721 23947 8746 24003
rect 8802 23947 8827 24003
rect 8883 23947 8908 24003
rect 8964 23947 8989 24003
rect 9045 23947 9070 24003
rect 9126 23947 9151 24003
rect 9207 23947 9232 24003
rect 9288 23947 9313 24003
rect 9369 23947 9394 24003
rect 9450 23947 9475 24003
rect 9531 23947 9556 24003
rect 9612 23947 9637 24003
rect 9693 23947 9718 24003
rect 9774 23947 9799 24003
rect 9855 23947 9880 24003
rect 9936 23947 9961 24003
rect 10017 23947 10042 24003
rect 10098 23947 10123 24003
rect 10179 23947 10204 24003
rect 10260 23947 10285 24003
rect 10341 23947 10366 24003
rect 10422 23947 10447 24003
rect 10503 23947 10528 24003
rect 10584 23947 10609 24003
rect 10665 23947 10690 24003
rect 10746 23947 10771 24003
rect 10827 23947 10852 24003
rect 10908 23947 10933 24003
rect 10989 23947 11014 24003
rect 11070 23947 11095 24003
rect 11151 23947 11176 24003
rect 11232 23947 11257 24003
rect 11313 23947 11338 24003
rect 11394 23947 11419 24003
rect 11475 23947 11500 24003
rect 5416 23923 11500 23947
rect 5416 23867 5425 23923
rect 5481 23867 5506 23923
rect 5562 23867 5587 23923
rect 5643 23867 5668 23923
rect 5724 23867 5749 23923
rect 5805 23867 5830 23923
rect 5886 23867 5911 23923
rect 5967 23867 5992 23923
rect 6048 23867 6073 23923
rect 6129 23867 6154 23923
rect 6210 23867 6235 23923
rect 6291 23867 6316 23923
rect 6372 23867 6397 23923
rect 6453 23867 6478 23923
rect 6534 23867 6559 23923
rect 6615 23867 6640 23923
rect 6696 23867 6721 23923
rect 6777 23867 6802 23923
rect 6858 23867 6883 23923
rect 6939 23867 6964 23923
rect 7020 23867 7045 23923
rect 7101 23867 7126 23923
rect 7182 23867 7207 23923
rect 7263 23867 7288 23923
rect 7344 23867 7369 23923
rect 7425 23867 7450 23923
rect 7506 23867 7531 23923
rect 7587 23867 7612 23923
rect 7668 23867 7693 23923
rect 7749 23867 7774 23923
rect 7830 23867 7855 23923
rect 7911 23867 7936 23923
rect 7992 23867 8017 23923
rect 8073 23867 8098 23923
rect 8154 23867 8179 23923
rect 8235 23867 8260 23923
rect 8316 23867 8341 23923
rect 8397 23867 8422 23923
rect 8478 23867 8503 23923
rect 8559 23867 8584 23923
rect 8640 23867 8665 23923
rect 8721 23867 8746 23923
rect 8802 23867 8827 23923
rect 8883 23867 8908 23923
rect 8964 23867 8989 23923
rect 9045 23867 9070 23923
rect 9126 23867 9151 23923
rect 9207 23867 9232 23923
rect 9288 23867 9313 23923
rect 9369 23867 9394 23923
rect 9450 23867 9475 23923
rect 9531 23867 9556 23923
rect 9612 23867 9637 23923
rect 9693 23867 9718 23923
rect 9774 23867 9799 23923
rect 9855 23867 9880 23923
rect 9936 23867 9961 23923
rect 10017 23867 10042 23923
rect 10098 23867 10123 23923
rect 10179 23867 10204 23923
rect 10260 23867 10285 23923
rect 10341 23867 10366 23923
rect 10422 23867 10447 23923
rect 10503 23867 10528 23923
rect 10584 23867 10609 23923
rect 10665 23867 10690 23923
rect 10746 23867 10771 23923
rect 10827 23867 10852 23923
rect 10908 23867 10933 23923
rect 10989 23867 11014 23923
rect 11070 23867 11095 23923
rect 11151 23867 11176 23923
rect 11232 23867 11257 23923
rect 11313 23867 11338 23923
rect 11394 23867 11419 23923
rect 11475 23867 11500 23923
rect 5416 23843 11500 23867
rect 5416 23787 5425 23843
rect 5481 23787 5506 23843
rect 5562 23787 5587 23843
rect 5643 23787 5668 23843
rect 5724 23787 5749 23843
rect 5805 23787 5830 23843
rect 5886 23787 5911 23843
rect 5967 23787 5992 23843
rect 6048 23787 6073 23843
rect 6129 23787 6154 23843
rect 6210 23787 6235 23843
rect 6291 23787 6316 23843
rect 6372 23787 6397 23843
rect 6453 23787 6478 23843
rect 6534 23787 6559 23843
rect 6615 23787 6640 23843
rect 6696 23787 6721 23843
rect 6777 23787 6802 23843
rect 6858 23787 6883 23843
rect 6939 23787 6964 23843
rect 7020 23787 7045 23843
rect 7101 23787 7126 23843
rect 7182 23787 7207 23843
rect 7263 23787 7288 23843
rect 7344 23787 7369 23843
rect 7425 23787 7450 23843
rect 7506 23787 7531 23843
rect 7587 23787 7612 23843
rect 7668 23787 7693 23843
rect 7749 23787 7774 23843
rect 7830 23787 7855 23843
rect 7911 23787 7936 23843
rect 7992 23787 8017 23843
rect 8073 23787 8098 23843
rect 8154 23787 8179 23843
rect 8235 23787 8260 23843
rect 8316 23787 8341 23843
rect 8397 23787 8422 23843
rect 8478 23787 8503 23843
rect 8559 23787 8584 23843
rect 8640 23787 8665 23843
rect 8721 23787 8746 23843
rect 8802 23787 8827 23843
rect 8883 23787 8908 23843
rect 8964 23787 8989 23843
rect 9045 23787 9070 23843
rect 9126 23787 9151 23843
rect 9207 23787 9232 23843
rect 9288 23787 9313 23843
rect 9369 23787 9394 23843
rect 9450 23787 9475 23843
rect 9531 23787 9556 23843
rect 9612 23787 9637 23843
rect 9693 23787 9718 23843
rect 9774 23787 9799 23843
rect 9855 23787 9880 23843
rect 9936 23787 9961 23843
rect 10017 23787 10042 23843
rect 10098 23787 10123 23843
rect 10179 23787 10204 23843
rect 10260 23787 10285 23843
rect 10341 23787 10366 23843
rect 10422 23787 10447 23843
rect 10503 23787 10528 23843
rect 10584 23787 10609 23843
rect 10665 23787 10690 23843
rect 10746 23787 10771 23843
rect 10827 23787 10852 23843
rect 10908 23787 10933 23843
rect 10989 23787 11014 23843
rect 11070 23787 11095 23843
rect 11151 23787 11176 23843
rect 11232 23787 11257 23843
rect 11313 23787 11338 23843
rect 11394 23787 11419 23843
rect 11475 23787 11500 23843
rect 5416 23763 11500 23787
rect 5416 23707 5425 23763
rect 5481 23707 5506 23763
rect 5562 23707 5587 23763
rect 5643 23707 5668 23763
rect 5724 23707 5749 23763
rect 5805 23707 5830 23763
rect 5886 23707 5911 23763
rect 5967 23707 5992 23763
rect 6048 23707 6073 23763
rect 6129 23707 6154 23763
rect 6210 23707 6235 23763
rect 6291 23707 6316 23763
rect 6372 23707 6397 23763
rect 6453 23707 6478 23763
rect 6534 23707 6559 23763
rect 6615 23707 6640 23763
rect 6696 23707 6721 23763
rect 6777 23707 6802 23763
rect 6858 23707 6883 23763
rect 6939 23707 6964 23763
rect 7020 23707 7045 23763
rect 7101 23707 7126 23763
rect 7182 23707 7207 23763
rect 7263 23707 7288 23763
rect 7344 23707 7369 23763
rect 7425 23707 7450 23763
rect 7506 23707 7531 23763
rect 7587 23707 7612 23763
rect 7668 23707 7693 23763
rect 7749 23707 7774 23763
rect 7830 23707 7855 23763
rect 7911 23707 7936 23763
rect 7992 23707 8017 23763
rect 8073 23707 8098 23763
rect 8154 23707 8179 23763
rect 8235 23707 8260 23763
rect 8316 23707 8341 23763
rect 8397 23707 8422 23763
rect 8478 23707 8503 23763
rect 8559 23707 8584 23763
rect 8640 23707 8665 23763
rect 8721 23707 8746 23763
rect 8802 23707 8827 23763
rect 8883 23707 8908 23763
rect 8964 23707 8989 23763
rect 9045 23707 9070 23763
rect 9126 23707 9151 23763
rect 9207 23707 9232 23763
rect 9288 23707 9313 23763
rect 9369 23707 9394 23763
rect 9450 23707 9475 23763
rect 9531 23707 9556 23763
rect 9612 23707 9637 23763
rect 9693 23707 9718 23763
rect 9774 23707 9799 23763
rect 9855 23707 9880 23763
rect 9936 23707 9961 23763
rect 10017 23707 10042 23763
rect 10098 23707 10123 23763
rect 10179 23707 10204 23763
rect 10260 23707 10285 23763
rect 10341 23707 10366 23763
rect 10422 23707 10447 23763
rect 10503 23707 10528 23763
rect 10584 23707 10609 23763
rect 10665 23707 10690 23763
rect 10746 23707 10771 23763
rect 10827 23707 10852 23763
rect 10908 23707 10933 23763
rect 10989 23707 11014 23763
rect 11070 23707 11095 23763
rect 11151 23707 11176 23763
rect 11232 23707 11257 23763
rect 11313 23707 11338 23763
rect 11394 23707 11419 23763
rect 11475 23707 11500 23763
rect 5416 23683 11500 23707
rect 5416 23627 5425 23683
rect 5481 23627 5506 23683
rect 5562 23627 5587 23683
rect 5643 23627 5668 23683
rect 5724 23627 5749 23683
rect 5805 23627 5830 23683
rect 5886 23627 5911 23683
rect 5967 23627 5992 23683
rect 6048 23627 6073 23683
rect 6129 23627 6154 23683
rect 6210 23627 6235 23683
rect 6291 23627 6316 23683
rect 6372 23627 6397 23683
rect 6453 23627 6478 23683
rect 6534 23627 6559 23683
rect 6615 23627 6640 23683
rect 6696 23627 6721 23683
rect 6777 23627 6802 23683
rect 6858 23627 6883 23683
rect 6939 23627 6964 23683
rect 7020 23627 7045 23683
rect 7101 23627 7126 23683
rect 7182 23627 7207 23683
rect 7263 23627 7288 23683
rect 7344 23627 7369 23683
rect 7425 23627 7450 23683
rect 7506 23627 7531 23683
rect 7587 23627 7612 23683
rect 7668 23627 7693 23683
rect 7749 23627 7774 23683
rect 7830 23627 7855 23683
rect 7911 23627 7936 23683
rect 7992 23627 8017 23683
rect 8073 23627 8098 23683
rect 8154 23627 8179 23683
rect 8235 23627 8260 23683
rect 8316 23627 8341 23683
rect 8397 23627 8422 23683
rect 8478 23627 8503 23683
rect 8559 23627 8584 23683
rect 8640 23627 8665 23683
rect 8721 23627 8746 23683
rect 8802 23627 8827 23683
rect 8883 23627 8908 23683
rect 8964 23627 8989 23683
rect 9045 23627 9070 23683
rect 9126 23627 9151 23683
rect 9207 23627 9232 23683
rect 9288 23627 9313 23683
rect 9369 23627 9394 23683
rect 9450 23627 9475 23683
rect 9531 23627 9556 23683
rect 9612 23627 9637 23683
rect 9693 23627 9718 23683
rect 9774 23627 9799 23683
rect 9855 23627 9880 23683
rect 9936 23627 9961 23683
rect 10017 23627 10042 23683
rect 10098 23627 10123 23683
rect 10179 23627 10204 23683
rect 10260 23627 10285 23683
rect 10341 23627 10366 23683
rect 10422 23627 10447 23683
rect 10503 23627 10528 23683
rect 10584 23627 10609 23683
rect 10665 23627 10690 23683
rect 10746 23627 10771 23683
rect 10827 23627 10852 23683
rect 10908 23627 10933 23683
rect 10989 23627 11014 23683
rect 11070 23627 11095 23683
rect 11151 23627 11176 23683
rect 11232 23627 11257 23683
rect 11313 23627 11338 23683
rect 11394 23627 11419 23683
rect 11475 23627 11500 23683
rect 5416 23603 11500 23627
rect 5416 23547 5425 23603
rect 5481 23547 5506 23603
rect 5562 23547 5587 23603
rect 5643 23547 5668 23603
rect 5724 23547 5749 23603
rect 5805 23547 5830 23603
rect 5886 23547 5911 23603
rect 5967 23547 5992 23603
rect 6048 23547 6073 23603
rect 6129 23547 6154 23603
rect 6210 23547 6235 23603
rect 6291 23547 6316 23603
rect 6372 23547 6397 23603
rect 6453 23547 6478 23603
rect 6534 23547 6559 23603
rect 6615 23547 6640 23603
rect 6696 23547 6721 23603
rect 6777 23547 6802 23603
rect 6858 23547 6883 23603
rect 6939 23547 6964 23603
rect 7020 23547 7045 23603
rect 7101 23547 7126 23603
rect 7182 23547 7207 23603
rect 7263 23547 7288 23603
rect 7344 23547 7369 23603
rect 7425 23547 7450 23603
rect 7506 23547 7531 23603
rect 7587 23547 7612 23603
rect 7668 23547 7693 23603
rect 7749 23547 7774 23603
rect 7830 23547 7855 23603
rect 7911 23547 7936 23603
rect 7992 23547 8017 23603
rect 8073 23547 8098 23603
rect 8154 23547 8179 23603
rect 8235 23547 8260 23603
rect 8316 23547 8341 23603
rect 8397 23547 8422 23603
rect 8478 23547 8503 23603
rect 8559 23547 8584 23603
rect 8640 23547 8665 23603
rect 8721 23547 8746 23603
rect 8802 23547 8827 23603
rect 8883 23547 8908 23603
rect 8964 23547 8989 23603
rect 9045 23547 9070 23603
rect 9126 23547 9151 23603
rect 9207 23547 9232 23603
rect 9288 23547 9313 23603
rect 9369 23547 9394 23603
rect 9450 23547 9475 23603
rect 9531 23547 9556 23603
rect 9612 23547 9637 23603
rect 9693 23547 9718 23603
rect 9774 23547 9799 23603
rect 9855 23547 9880 23603
rect 9936 23547 9961 23603
rect 10017 23547 10042 23603
rect 10098 23547 10123 23603
rect 10179 23547 10204 23603
rect 10260 23547 10285 23603
rect 10341 23547 10366 23603
rect 10422 23547 10447 23603
rect 10503 23547 10528 23603
rect 10584 23547 10609 23603
rect 10665 23547 10690 23603
rect 10746 23547 10771 23603
rect 10827 23547 10852 23603
rect 10908 23547 10933 23603
rect 10989 23547 11014 23603
rect 11070 23547 11095 23603
rect 11151 23547 11176 23603
rect 11232 23547 11257 23603
rect 11313 23547 11338 23603
rect 11394 23547 11419 23603
rect 11475 23547 11500 23603
rect 5416 23523 11500 23547
rect 5416 23467 5425 23523
rect 5481 23467 5506 23523
rect 5562 23467 5587 23523
rect 5643 23467 5668 23523
rect 5724 23467 5749 23523
rect 5805 23467 5830 23523
rect 5886 23467 5911 23523
rect 5967 23467 5992 23523
rect 6048 23467 6073 23523
rect 6129 23467 6154 23523
rect 6210 23467 6235 23523
rect 6291 23467 6316 23523
rect 6372 23467 6397 23523
rect 6453 23467 6478 23523
rect 6534 23467 6559 23523
rect 6615 23467 6640 23523
rect 6696 23467 6721 23523
rect 6777 23467 6802 23523
rect 6858 23467 6883 23523
rect 6939 23467 6964 23523
rect 7020 23467 7045 23523
rect 7101 23467 7126 23523
rect 7182 23467 7207 23523
rect 7263 23467 7288 23523
rect 7344 23467 7369 23523
rect 7425 23467 7450 23523
rect 7506 23467 7531 23523
rect 7587 23467 7612 23523
rect 7668 23467 7693 23523
rect 7749 23467 7774 23523
rect 7830 23467 7855 23523
rect 7911 23467 7936 23523
rect 7992 23467 8017 23523
rect 8073 23467 8098 23523
rect 8154 23467 8179 23523
rect 8235 23467 8260 23523
rect 8316 23467 8341 23523
rect 8397 23467 8422 23523
rect 8478 23467 8503 23523
rect 8559 23467 8584 23523
rect 8640 23467 8665 23523
rect 8721 23467 8746 23523
rect 8802 23467 8827 23523
rect 8883 23467 8908 23523
rect 8964 23467 8989 23523
rect 9045 23467 9070 23523
rect 9126 23467 9151 23523
rect 9207 23467 9232 23523
rect 9288 23467 9313 23523
rect 9369 23467 9394 23523
rect 9450 23467 9475 23523
rect 9531 23467 9556 23523
rect 9612 23467 9637 23523
rect 9693 23467 9718 23523
rect 9774 23467 9799 23523
rect 9855 23467 9880 23523
rect 9936 23467 9961 23523
rect 10017 23467 10042 23523
rect 10098 23467 10123 23523
rect 10179 23467 10204 23523
rect 10260 23467 10285 23523
rect 10341 23467 10366 23523
rect 10422 23467 10447 23523
rect 10503 23467 10528 23523
rect 10584 23467 10609 23523
rect 10665 23467 10690 23523
rect 10746 23467 10771 23523
rect 10827 23467 10852 23523
rect 10908 23467 10933 23523
rect 10989 23467 11014 23523
rect 11070 23467 11095 23523
rect 11151 23467 11176 23523
rect 11232 23467 11257 23523
rect 11313 23467 11338 23523
rect 11394 23467 11419 23523
rect 11475 23467 11500 23523
rect 5416 23443 11500 23467
rect 5416 23387 5425 23443
rect 5481 23387 5506 23443
rect 5562 23387 5587 23443
rect 5643 23387 5668 23443
rect 5724 23387 5749 23443
rect 5805 23387 5830 23443
rect 5886 23387 5911 23443
rect 5967 23387 5992 23443
rect 6048 23387 6073 23443
rect 6129 23387 6154 23443
rect 6210 23387 6235 23443
rect 6291 23387 6316 23443
rect 6372 23387 6397 23443
rect 6453 23387 6478 23443
rect 6534 23387 6559 23443
rect 6615 23387 6640 23443
rect 6696 23387 6721 23443
rect 6777 23387 6802 23443
rect 6858 23387 6883 23443
rect 6939 23387 6964 23443
rect 7020 23387 7045 23443
rect 7101 23387 7126 23443
rect 7182 23387 7207 23443
rect 7263 23387 7288 23443
rect 7344 23387 7369 23443
rect 7425 23387 7450 23443
rect 7506 23387 7531 23443
rect 7587 23387 7612 23443
rect 7668 23387 7693 23443
rect 7749 23387 7774 23443
rect 7830 23387 7855 23443
rect 7911 23387 7936 23443
rect 7992 23387 8017 23443
rect 8073 23387 8098 23443
rect 8154 23387 8179 23443
rect 8235 23387 8260 23443
rect 8316 23387 8341 23443
rect 8397 23387 8422 23443
rect 8478 23387 8503 23443
rect 8559 23387 8584 23443
rect 8640 23387 8665 23443
rect 8721 23387 8746 23443
rect 8802 23387 8827 23443
rect 8883 23387 8908 23443
rect 8964 23387 8989 23443
rect 9045 23387 9070 23443
rect 9126 23387 9151 23443
rect 9207 23387 9232 23443
rect 9288 23387 9313 23443
rect 9369 23387 9394 23443
rect 9450 23387 9475 23443
rect 9531 23387 9556 23443
rect 9612 23387 9637 23443
rect 9693 23387 9718 23443
rect 9774 23387 9799 23443
rect 9855 23387 9880 23443
rect 9936 23387 9961 23443
rect 10017 23387 10042 23443
rect 10098 23387 10123 23443
rect 10179 23387 10204 23443
rect 10260 23387 10285 23443
rect 10341 23387 10366 23443
rect 10422 23387 10447 23443
rect 10503 23387 10528 23443
rect 10584 23387 10609 23443
rect 10665 23387 10690 23443
rect 10746 23387 10771 23443
rect 10827 23387 10852 23443
rect 10908 23387 10933 23443
rect 10989 23387 11014 23443
rect 11070 23387 11095 23443
rect 11151 23387 11176 23443
rect 11232 23387 11257 23443
rect 11313 23387 11338 23443
rect 11394 23387 11419 23443
rect 11475 23387 11500 23443
rect 5416 23363 11500 23387
rect 5416 23307 5425 23363
rect 5481 23307 5506 23363
rect 5562 23307 5587 23363
rect 5643 23307 5668 23363
rect 5724 23307 5749 23363
rect 5805 23307 5830 23363
rect 5886 23307 5911 23363
rect 5967 23307 5992 23363
rect 6048 23307 6073 23363
rect 6129 23307 6154 23363
rect 6210 23307 6235 23363
rect 6291 23307 6316 23363
rect 6372 23307 6397 23363
rect 6453 23307 6478 23363
rect 6534 23307 6559 23363
rect 6615 23307 6640 23363
rect 6696 23307 6721 23363
rect 6777 23307 6802 23363
rect 6858 23307 6883 23363
rect 6939 23307 6964 23363
rect 7020 23307 7045 23363
rect 7101 23307 7126 23363
rect 7182 23307 7207 23363
rect 7263 23307 7288 23363
rect 7344 23307 7369 23363
rect 7425 23307 7450 23363
rect 7506 23307 7531 23363
rect 7587 23307 7612 23363
rect 7668 23307 7693 23363
rect 7749 23307 7774 23363
rect 7830 23307 7855 23363
rect 7911 23307 7936 23363
rect 7992 23307 8017 23363
rect 8073 23307 8098 23363
rect 8154 23307 8179 23363
rect 8235 23307 8260 23363
rect 8316 23307 8341 23363
rect 8397 23307 8422 23363
rect 8478 23307 8503 23363
rect 8559 23307 8584 23363
rect 8640 23307 8665 23363
rect 8721 23307 8746 23363
rect 8802 23307 8827 23363
rect 8883 23307 8908 23363
rect 8964 23307 8989 23363
rect 9045 23307 9070 23363
rect 9126 23307 9151 23363
rect 9207 23307 9232 23363
rect 9288 23307 9313 23363
rect 9369 23307 9394 23363
rect 9450 23307 9475 23363
rect 9531 23307 9556 23363
rect 9612 23307 9637 23363
rect 9693 23307 9718 23363
rect 9774 23307 9799 23363
rect 9855 23307 9880 23363
rect 9936 23307 9961 23363
rect 10017 23307 10042 23363
rect 10098 23307 10123 23363
rect 10179 23307 10204 23363
rect 10260 23307 10285 23363
rect 10341 23307 10366 23363
rect 10422 23307 10447 23363
rect 10503 23307 10528 23363
rect 10584 23307 10609 23363
rect 10665 23307 10690 23363
rect 10746 23307 10771 23363
rect 10827 23307 10852 23363
rect 10908 23307 10933 23363
rect 10989 23307 11014 23363
rect 11070 23307 11095 23363
rect 11151 23307 11176 23363
rect 11232 23307 11257 23363
rect 11313 23307 11338 23363
rect 11394 23307 11419 23363
rect 11475 23307 11500 23363
rect 5416 23283 11500 23307
rect 5416 23227 5425 23283
rect 5481 23227 5506 23283
rect 5562 23227 5587 23283
rect 5643 23227 5668 23283
rect 5724 23227 5749 23283
rect 5805 23227 5830 23283
rect 5886 23227 5911 23283
rect 5967 23227 5992 23283
rect 6048 23227 6073 23283
rect 6129 23227 6154 23283
rect 6210 23227 6235 23283
rect 6291 23227 6316 23283
rect 6372 23227 6397 23283
rect 6453 23227 6478 23283
rect 6534 23227 6559 23283
rect 6615 23227 6640 23283
rect 6696 23227 6721 23283
rect 6777 23227 6802 23283
rect 6858 23227 6883 23283
rect 6939 23227 6964 23283
rect 7020 23227 7045 23283
rect 7101 23227 7126 23283
rect 7182 23227 7207 23283
rect 7263 23227 7288 23283
rect 7344 23227 7369 23283
rect 7425 23227 7450 23283
rect 7506 23227 7531 23283
rect 7587 23227 7612 23283
rect 7668 23227 7693 23283
rect 7749 23227 7774 23283
rect 7830 23227 7855 23283
rect 7911 23227 7936 23283
rect 7992 23227 8017 23283
rect 8073 23227 8098 23283
rect 8154 23227 8179 23283
rect 8235 23227 8260 23283
rect 8316 23227 8341 23283
rect 8397 23227 8422 23283
rect 8478 23227 8503 23283
rect 8559 23227 8584 23283
rect 8640 23227 8665 23283
rect 8721 23227 8746 23283
rect 8802 23227 8827 23283
rect 8883 23227 8908 23283
rect 8964 23227 8989 23283
rect 9045 23227 9070 23283
rect 9126 23227 9151 23283
rect 9207 23227 9232 23283
rect 9288 23227 9313 23283
rect 9369 23227 9394 23283
rect 9450 23227 9475 23283
rect 9531 23227 9556 23283
rect 9612 23227 9637 23283
rect 9693 23227 9718 23283
rect 9774 23227 9799 23283
rect 9855 23227 9880 23283
rect 9936 23227 9961 23283
rect 10017 23227 10042 23283
rect 10098 23227 10123 23283
rect 10179 23227 10204 23283
rect 10260 23227 10285 23283
rect 10341 23227 10366 23283
rect 10422 23227 10447 23283
rect 10503 23227 10528 23283
rect 10584 23227 10609 23283
rect 10665 23227 10690 23283
rect 10746 23227 10771 23283
rect 10827 23227 10852 23283
rect 10908 23227 10933 23283
rect 10989 23227 11014 23283
rect 11070 23227 11095 23283
rect 11151 23227 11176 23283
rect 11232 23227 11257 23283
rect 11313 23227 11338 23283
rect 11394 23227 11419 23283
rect 11475 23227 11500 23283
rect 5416 23203 11500 23227
rect 5416 23147 5425 23203
rect 5481 23147 5506 23203
rect 5562 23147 5587 23203
rect 5643 23147 5668 23203
rect 5724 23147 5749 23203
rect 5805 23147 5830 23203
rect 5886 23147 5911 23203
rect 5967 23147 5992 23203
rect 6048 23147 6073 23203
rect 6129 23147 6154 23203
rect 6210 23147 6235 23203
rect 6291 23147 6316 23203
rect 6372 23147 6397 23203
rect 6453 23147 6478 23203
rect 6534 23147 6559 23203
rect 6615 23147 6640 23203
rect 6696 23147 6721 23203
rect 6777 23147 6802 23203
rect 6858 23147 6883 23203
rect 6939 23147 6964 23203
rect 7020 23147 7045 23203
rect 7101 23147 7126 23203
rect 7182 23147 7207 23203
rect 7263 23147 7288 23203
rect 7344 23147 7369 23203
rect 7425 23147 7450 23203
rect 7506 23147 7531 23203
rect 7587 23147 7612 23203
rect 7668 23147 7693 23203
rect 7749 23147 7774 23203
rect 7830 23147 7855 23203
rect 7911 23147 7936 23203
rect 7992 23147 8017 23203
rect 8073 23147 8098 23203
rect 8154 23147 8179 23203
rect 8235 23147 8260 23203
rect 8316 23147 8341 23203
rect 8397 23147 8422 23203
rect 8478 23147 8503 23203
rect 8559 23147 8584 23203
rect 8640 23147 8665 23203
rect 8721 23147 8746 23203
rect 8802 23147 8827 23203
rect 8883 23147 8908 23203
rect 8964 23147 8989 23203
rect 9045 23147 9070 23203
rect 9126 23147 9151 23203
rect 9207 23147 9232 23203
rect 9288 23147 9313 23203
rect 9369 23147 9394 23203
rect 9450 23147 9475 23203
rect 9531 23147 9556 23203
rect 9612 23147 9637 23203
rect 9693 23147 9718 23203
rect 9774 23147 9799 23203
rect 9855 23147 9880 23203
rect 9936 23147 9961 23203
rect 10017 23147 10042 23203
rect 10098 23147 10123 23203
rect 10179 23147 10204 23203
rect 10260 23147 10285 23203
rect 10341 23147 10366 23203
rect 10422 23147 10447 23203
rect 10503 23147 10528 23203
rect 10584 23147 10609 23203
rect 10665 23147 10690 23203
rect 10746 23147 10771 23203
rect 10827 23147 10852 23203
rect 10908 23147 10933 23203
rect 10989 23147 11014 23203
rect 11070 23147 11095 23203
rect 11151 23147 11176 23203
rect 11232 23147 11257 23203
rect 11313 23147 11338 23203
rect 11394 23147 11419 23203
rect 11475 23147 11500 23203
rect 13076 23147 13085 24323
rect 5416 23136 13085 23147
rect 13579 21961 14391 33386
tri 14391 32784 15371 33764 nw
rect 14502 31178 15298 31184
rect 14502 29034 14508 31178
rect 15292 29034 15298 31178
rect 14502 29017 15298 29034
rect 14502 28953 14508 29017
rect 14572 28953 14588 29017
rect 14652 28953 14668 29017
rect 14732 28953 14748 29017
rect 14812 28953 14828 29017
rect 14892 28953 14908 29017
rect 14972 28953 14988 29017
rect 15052 28953 15068 29017
rect 15132 28953 15148 29017
rect 15212 28953 15228 29017
rect 15292 28953 15298 29017
rect 14502 28936 15298 28953
rect 14502 28872 14508 28936
rect 14572 28872 14588 28936
rect 14652 28872 14668 28936
rect 14732 28872 14748 28936
rect 14812 28872 14828 28936
rect 14892 28872 14908 28936
rect 14972 28872 14988 28936
rect 15052 28872 15068 28936
rect 15132 28872 15148 28936
rect 15212 28872 15228 28936
rect 15292 28872 15298 28936
rect 14502 28871 14514 28872
rect 14570 28871 14594 28872
rect 14650 28871 14674 28872
rect 14730 28871 14754 28872
rect 14810 28871 14834 28872
rect 14890 28871 14914 28872
rect 14970 28871 14994 28872
rect 15050 28871 15074 28872
rect 15130 28871 15154 28872
rect 15210 28871 15234 28872
rect 15290 28871 15298 28872
rect 14502 28866 15298 28871
rect 14517 27593 15039 27599
rect 14517 27529 14521 27593
rect 14585 27529 14611 27593
rect 14675 27529 14701 27593
rect 14765 27529 14791 27593
rect 14855 27574 14881 27593
rect 14945 27574 14971 27593
rect 14855 27529 14880 27574
rect 14945 27529 14969 27574
rect 15035 27529 15039 27593
rect 14517 27518 14522 27529
rect 14578 27518 14612 27529
rect 14668 27518 14702 27529
rect 14758 27518 14791 27529
rect 14847 27518 14880 27529
rect 14936 27518 14969 27529
rect 15025 27518 15039 27529
rect 14517 27512 15039 27518
rect 14517 27448 14521 27512
rect 14585 27448 14611 27512
rect 14675 27448 14701 27512
rect 14765 27448 14791 27512
rect 14855 27488 14881 27512
rect 14945 27488 14971 27512
rect 14855 27448 14880 27488
rect 14945 27448 14969 27488
rect 15035 27448 15039 27512
rect 14517 27432 14522 27448
rect 14578 27432 14612 27448
rect 14668 27432 14702 27448
rect 14758 27432 14791 27448
rect 14847 27432 14880 27448
rect 14936 27432 14969 27448
rect 15025 27432 15039 27448
rect 14517 27431 15039 27432
rect 14517 27367 14521 27431
rect 14585 27367 14611 27431
rect 14675 27367 14701 27431
rect 14765 27367 14791 27431
rect 14855 27402 14881 27431
rect 14945 27402 14971 27431
rect 14855 27367 14880 27402
rect 14945 27367 14969 27402
rect 15035 27367 15039 27431
rect 14517 27350 14522 27367
rect 14578 27350 14612 27367
rect 14668 27350 14702 27367
rect 14758 27350 14791 27367
rect 14847 27350 14880 27367
rect 14936 27350 14969 27367
rect 15025 27350 15039 27367
rect 14517 27286 14521 27350
rect 14585 27286 14611 27350
rect 14675 27286 14701 27350
rect 14765 27286 14791 27350
rect 14855 27346 14880 27350
rect 14945 27346 14969 27350
rect 14855 27316 14881 27346
rect 14945 27316 14971 27346
rect 14855 27286 14880 27316
rect 14945 27286 14969 27316
rect 15035 27286 15039 27350
rect 14517 27268 14522 27286
rect 14578 27268 14612 27286
rect 14668 27268 14702 27286
rect 14758 27268 14791 27286
rect 14847 27268 14880 27286
rect 14936 27268 14969 27286
rect 15025 27268 15039 27286
rect 14517 27204 14521 27268
rect 14585 27204 14611 27268
rect 14675 27204 14701 27268
rect 14765 27204 14791 27268
rect 14855 27260 14880 27268
rect 14945 27260 14969 27268
rect 14855 27230 14881 27260
rect 14945 27230 14971 27260
rect 14855 27204 14880 27230
rect 14945 27204 14969 27230
rect 15035 27204 15039 27268
rect 14517 27186 14522 27204
rect 14578 27186 14612 27204
rect 14668 27186 14702 27204
rect 14758 27186 14791 27204
rect 14847 27186 14880 27204
rect 14936 27186 14969 27204
rect 15025 27186 15039 27204
rect 14517 27122 14521 27186
rect 14585 27122 14611 27186
rect 14675 27122 14701 27186
rect 14765 27122 14791 27186
rect 14855 27174 14880 27186
rect 14945 27174 14969 27186
rect 14855 27144 14881 27174
rect 14945 27144 14971 27174
rect 14855 27122 14880 27144
rect 14945 27122 14969 27144
rect 15035 27122 15039 27186
rect 14517 27104 14522 27122
rect 14578 27104 14612 27122
rect 14668 27104 14702 27122
rect 14758 27104 14791 27122
rect 14847 27104 14880 27122
rect 14936 27104 14969 27122
rect 15025 27104 15039 27122
rect 14517 27040 14521 27104
rect 14585 27040 14611 27104
rect 14675 27040 14701 27104
rect 14765 27040 14791 27104
rect 14855 27088 14880 27104
rect 14945 27088 14969 27104
rect 14855 27040 14881 27088
rect 14945 27040 14971 27088
rect 15035 27040 15039 27104
rect 14517 27034 15039 27040
rect 14504 25822 15040 25827
rect 14504 25766 14509 25822
rect 14565 25809 14603 25822
rect 14659 25809 14697 25822
rect 14753 25809 14791 25822
rect 14847 25809 14885 25822
rect 14941 25809 14979 25822
rect 14504 25745 14510 25766
rect 14574 25745 14602 25809
rect 14666 25745 14694 25809
rect 14758 25745 14786 25809
rect 14850 25745 14878 25809
rect 14942 25745 14970 25809
rect 15035 25766 15040 25822
rect 15034 25745 15040 25766
rect 14504 25741 15040 25745
rect 14504 25685 14509 25741
rect 14565 25729 14603 25741
rect 14659 25729 14697 25741
rect 14753 25729 14791 25741
rect 14847 25729 14885 25741
rect 14941 25729 14979 25741
rect 14504 25665 14510 25685
rect 14574 25665 14602 25729
rect 14666 25665 14694 25729
rect 14758 25665 14786 25729
rect 14850 25665 14878 25729
rect 14942 25665 14970 25729
rect 15035 25685 15040 25741
rect 15034 25665 15040 25685
rect 14504 25660 15040 25665
rect 14504 25604 14509 25660
rect 14565 25648 14603 25660
rect 14659 25648 14697 25660
rect 14753 25648 14791 25660
rect 14847 25648 14885 25660
rect 14941 25648 14979 25660
rect 14504 25584 14510 25604
rect 14574 25584 14602 25648
rect 14666 25584 14694 25648
rect 14758 25584 14786 25648
rect 14850 25584 14878 25648
rect 14942 25584 14970 25648
rect 15035 25604 15040 25660
rect 15034 25584 15040 25604
rect 14504 25579 15040 25584
rect 14504 25523 14509 25579
rect 14565 25567 14603 25579
rect 14659 25567 14697 25579
rect 14753 25567 14791 25579
rect 14847 25567 14885 25579
rect 14941 25567 14979 25579
rect 14504 25503 14510 25523
rect 14574 25503 14602 25567
rect 14666 25503 14694 25567
rect 14758 25503 14786 25567
rect 14850 25503 14878 25567
rect 14942 25503 14970 25567
rect 15035 25523 15040 25579
rect 15034 25503 15040 25523
rect 14504 25498 15040 25503
rect 14504 25442 14509 25498
rect 14565 25486 14603 25498
rect 14659 25486 14697 25498
rect 14753 25486 14791 25498
rect 14847 25486 14885 25498
rect 14941 25486 14979 25498
rect 14504 25422 14510 25442
rect 14574 25422 14602 25486
rect 14666 25422 14694 25486
rect 14758 25422 14786 25486
rect 14850 25422 14878 25486
rect 14942 25422 14970 25486
rect 15035 25442 15040 25498
rect 15034 25422 15040 25442
rect 14504 25417 15040 25422
rect 14504 25361 14509 25417
rect 14565 25405 14603 25417
rect 14659 25405 14697 25417
rect 14753 25405 14791 25417
rect 14847 25405 14885 25417
rect 14941 25405 14979 25417
rect 14504 25341 14510 25361
rect 14574 25341 14602 25405
rect 14666 25341 14694 25405
rect 14758 25341 14786 25405
rect 14850 25341 14878 25405
rect 14942 25341 14970 25405
rect 15035 25361 15040 25417
rect 15034 25341 15040 25361
rect 14504 25336 15040 25341
rect 14504 25280 14509 25336
rect 14565 25324 14603 25336
rect 14659 25324 14697 25336
rect 14753 25324 14791 25336
rect 14847 25324 14885 25336
rect 14941 25324 14979 25336
rect 14504 25260 14510 25280
rect 14574 25260 14602 25324
rect 14666 25260 14694 25324
rect 14758 25260 14786 25324
rect 14850 25260 14878 25324
rect 14942 25260 14970 25324
rect 15035 25280 15040 25336
rect 15034 25260 15040 25280
rect 14504 25255 15040 25260
rect 14504 25199 14509 25255
rect 14565 25243 14603 25255
rect 14659 25243 14697 25255
rect 14753 25243 14791 25255
rect 14847 25243 14885 25255
rect 14941 25243 14979 25255
rect 14504 25179 14510 25199
rect 14574 25179 14602 25243
rect 14666 25179 14694 25243
rect 14758 25179 14786 25243
rect 14850 25179 14878 25243
rect 14942 25179 14970 25243
rect 15035 25199 15040 25255
rect 15034 25179 15040 25199
rect 14504 25174 15040 25179
rect 14504 25118 14509 25174
rect 14565 25162 14603 25174
rect 14659 25162 14697 25174
rect 14753 25162 14791 25174
rect 14847 25162 14885 25174
rect 14941 25162 14979 25174
rect 14504 25098 14510 25118
rect 14574 25098 14602 25162
rect 14666 25098 14694 25162
rect 14758 25098 14786 25162
rect 14850 25098 14878 25162
rect 14942 25098 14970 25162
rect 15035 25118 15040 25174
rect 15034 25098 15040 25118
rect 14504 25093 15040 25098
rect 14504 25037 14509 25093
rect 14565 25081 14603 25093
rect 14659 25081 14697 25093
rect 14753 25081 14791 25093
rect 14847 25081 14885 25093
rect 14941 25081 14979 25093
rect 14504 25017 14510 25037
rect 14574 25017 14602 25081
rect 14666 25017 14694 25081
rect 14758 25017 14786 25081
rect 14850 25017 14878 25081
rect 14942 25017 14970 25081
rect 15035 25037 15040 25093
rect 15034 25017 15040 25037
rect 14504 25011 15040 25017
rect 14504 24955 14509 25011
rect 14565 25000 14603 25011
rect 14659 25000 14697 25011
rect 14753 25000 14791 25011
rect 14847 25000 14885 25011
rect 14941 25000 14979 25011
rect 14504 24936 14510 24955
rect 14574 24936 14602 25000
rect 14666 24936 14694 25000
rect 14758 24936 14786 25000
rect 14850 24936 14878 25000
rect 14942 24936 14970 25000
rect 15035 24955 15040 25011
rect 15034 24936 15040 24955
rect 14504 24929 15040 24936
rect 14504 24873 14509 24929
rect 14565 24919 14603 24929
rect 14659 24919 14697 24929
rect 14753 24919 14791 24929
rect 14847 24919 14885 24929
rect 14941 24919 14979 24929
rect 14504 24855 14510 24873
rect 14574 24855 14602 24919
rect 14666 24855 14694 24919
rect 14758 24855 14786 24919
rect 14850 24855 14878 24919
rect 14942 24855 14970 24919
rect 15035 24873 15040 24929
rect 15034 24855 15040 24873
rect 14504 24847 15040 24855
rect 14504 24791 14509 24847
rect 14565 24838 14603 24847
rect 14659 24838 14697 24847
rect 14753 24838 14791 24847
rect 14847 24838 14885 24847
rect 14941 24838 14979 24847
rect 14504 24774 14510 24791
rect 14574 24774 14602 24838
rect 14666 24774 14694 24838
rect 14758 24774 14786 24838
rect 14850 24774 14878 24838
rect 14942 24774 14970 24838
rect 15035 24791 15040 24847
rect 15034 24774 15040 24791
rect 14504 24765 15040 24774
rect 14504 24709 14509 24765
rect 14565 24757 14603 24765
rect 14659 24757 14697 24765
rect 14753 24757 14791 24765
rect 14847 24757 14885 24765
rect 14941 24757 14979 24765
rect 14504 24693 14510 24709
rect 14574 24693 14602 24757
rect 14666 24693 14694 24757
rect 14758 24693 14786 24757
rect 14850 24693 14878 24757
rect 14942 24693 14970 24757
rect 15035 24709 15040 24765
rect 15034 24693 15040 24709
rect 14504 24683 15040 24693
rect 14504 24627 14509 24683
rect 14565 24676 14603 24683
rect 14659 24676 14697 24683
rect 14753 24676 14791 24683
rect 14847 24676 14885 24683
rect 14941 24676 14979 24683
rect 14504 24612 14510 24627
rect 14574 24612 14602 24676
rect 14666 24612 14694 24676
rect 14758 24612 14786 24676
rect 14850 24612 14878 24676
rect 14942 24612 14970 24676
rect 15035 24627 15040 24683
rect 15034 24612 15040 24627
rect 14504 24601 15040 24612
rect 14504 24545 14509 24601
rect 14565 24595 14603 24601
rect 14659 24595 14697 24601
rect 14753 24595 14791 24601
rect 14847 24595 14885 24601
rect 14941 24595 14979 24601
rect 14504 24531 14510 24545
rect 14574 24531 14602 24595
rect 14666 24531 14694 24595
rect 14758 24531 14786 24595
rect 14850 24531 14878 24595
rect 14942 24531 14970 24595
rect 15035 24545 15040 24601
rect 15034 24531 15040 24545
rect 14504 24519 15040 24531
rect 14504 24463 14509 24519
rect 14565 24514 14603 24519
rect 14659 24514 14697 24519
rect 14753 24514 14791 24519
rect 14847 24514 14885 24519
rect 14941 24514 14979 24519
rect 14504 24450 14510 24463
rect 14574 24450 14602 24514
rect 14666 24450 14694 24514
rect 14758 24450 14786 24514
rect 14850 24450 14878 24514
rect 14942 24450 14970 24514
rect 15035 24463 15040 24519
rect 15034 24450 15040 24463
rect 14504 24437 15040 24450
rect 14504 24381 14509 24437
rect 14565 24433 14603 24437
rect 14659 24433 14697 24437
rect 14753 24433 14791 24437
rect 14847 24433 14885 24437
rect 14941 24433 14979 24437
rect 14504 24369 14510 24381
rect 14574 24369 14602 24433
rect 14666 24369 14694 24433
rect 14758 24369 14786 24433
rect 14850 24369 14878 24433
rect 14942 24369 14970 24433
rect 15035 24381 15040 24437
rect 15034 24369 15040 24381
rect 14504 24355 15040 24369
rect 14504 24299 14509 24355
rect 14565 24352 14603 24355
rect 14659 24352 14697 24355
rect 14753 24352 14791 24355
rect 14847 24352 14885 24355
rect 14941 24352 14979 24355
rect 14504 24288 14510 24299
rect 14574 24288 14602 24352
rect 14666 24288 14694 24352
rect 14758 24288 14786 24352
rect 14850 24288 14878 24352
rect 14942 24288 14970 24352
rect 15035 24299 15040 24355
rect 15034 24288 15040 24299
rect 14504 24273 15040 24288
rect 14504 24217 14509 24273
rect 14565 24271 14603 24273
rect 14659 24271 14697 24273
rect 14753 24271 14791 24273
rect 14847 24271 14885 24273
rect 14941 24271 14979 24273
rect 14504 24207 14510 24217
rect 14574 24207 14602 24271
rect 14666 24207 14694 24271
rect 14758 24207 14786 24271
rect 14850 24207 14878 24271
rect 14942 24207 14970 24271
rect 15035 24217 15040 24273
rect 15034 24207 15040 24217
rect 14504 24191 15040 24207
rect 14504 24135 14509 24191
rect 14565 24190 14603 24191
rect 14659 24190 14697 24191
rect 14753 24190 14791 24191
rect 14847 24190 14885 24191
rect 14941 24190 14979 24191
rect 14504 24126 14510 24135
rect 14574 24126 14602 24190
rect 14666 24126 14694 24190
rect 14758 24126 14786 24190
rect 14850 24126 14878 24190
rect 14942 24126 14970 24190
rect 15035 24135 15040 24191
rect 15034 24126 15040 24135
rect 14504 24109 15040 24126
rect 14504 24053 14509 24109
rect 14504 24045 14510 24053
rect 14574 24045 14602 24109
rect 14666 24045 14694 24109
rect 14758 24045 14786 24109
rect 14850 24045 14878 24109
rect 14942 24045 14970 24109
rect 15035 24053 15040 24109
rect 15034 24045 15040 24053
rect 14504 24028 15040 24045
rect 14504 24027 14510 24028
rect 14504 23971 14509 24027
rect 14504 23964 14510 23971
rect 14574 23964 14602 24028
rect 14666 23964 14694 24028
rect 14758 23964 14786 24028
rect 14850 23964 14878 24028
rect 14942 23964 14970 24028
rect 15034 24027 15040 24028
rect 15035 23971 15040 24027
rect 15034 23964 15040 23971
rect 14504 23947 15040 23964
rect 14504 23945 14510 23947
rect 14504 23889 14509 23945
rect 14504 23883 14510 23889
rect 14574 23883 14602 23947
rect 14666 23883 14694 23947
rect 14758 23883 14786 23947
rect 14850 23883 14878 23947
rect 14942 23883 14970 23947
rect 15034 23945 15040 23947
rect 15035 23889 15040 23945
rect 15034 23883 15040 23889
rect 14504 23866 15040 23883
rect 14504 23863 14510 23866
rect 14504 23807 14509 23863
rect 14504 23802 14510 23807
rect 14574 23802 14602 23866
rect 14666 23802 14694 23866
rect 14758 23802 14786 23866
rect 14850 23802 14878 23866
rect 14942 23802 14970 23866
rect 15034 23863 15040 23866
rect 15035 23807 15040 23863
rect 15034 23802 15040 23807
rect 14504 23785 15040 23802
rect 14504 23781 14510 23785
rect 14504 23725 14509 23781
rect 14504 23721 14510 23725
rect 14574 23721 14602 23785
rect 14666 23721 14694 23785
rect 14758 23721 14786 23785
rect 14850 23721 14878 23785
rect 14942 23721 14970 23785
rect 15034 23781 15040 23785
rect 15035 23725 15040 23781
rect 15034 23721 15040 23725
rect 14504 23704 15040 23721
rect 14504 23699 14510 23704
rect 14504 23643 14509 23699
rect 14504 23640 14510 23643
rect 14574 23640 14602 23704
rect 14666 23640 14694 23704
rect 14758 23640 14786 23704
rect 14850 23640 14878 23704
rect 14942 23640 14970 23704
rect 15034 23699 15040 23704
rect 15035 23643 15040 23699
rect 15034 23640 15040 23643
rect 14504 23623 15040 23640
rect 14504 23617 14510 23623
rect 14504 23561 14509 23617
rect 14504 23559 14510 23561
rect 14574 23559 14602 23623
rect 14666 23559 14694 23623
rect 14758 23559 14786 23623
rect 14850 23559 14878 23623
rect 14942 23559 14970 23623
rect 15034 23617 15040 23623
rect 15035 23561 15040 23617
rect 15034 23559 15040 23561
rect 14504 23542 15040 23559
rect 14504 23535 14510 23542
rect 14504 23479 14509 23535
rect 14504 23478 14510 23479
rect 14574 23478 14602 23542
rect 14666 23478 14694 23542
rect 14758 23478 14786 23542
rect 14850 23478 14878 23542
rect 14942 23478 14970 23542
rect 15034 23535 15040 23542
rect 15035 23479 15040 23535
rect 15034 23478 15040 23479
rect 14504 23461 15040 23478
rect 14504 23453 14510 23461
rect 14504 23397 14509 23453
rect 14574 23397 14602 23461
rect 14666 23397 14694 23461
rect 14758 23397 14786 23461
rect 14850 23397 14878 23461
rect 14942 23397 14970 23461
rect 15034 23453 15040 23461
rect 15035 23397 15040 23453
rect 14504 23380 15040 23397
rect 14504 23371 14510 23380
rect 14504 23315 14509 23371
rect 14574 23316 14602 23380
rect 14666 23316 14694 23380
rect 14758 23316 14786 23380
rect 14850 23316 14878 23380
rect 14942 23316 14970 23380
rect 15034 23371 15040 23380
rect 14565 23315 14603 23316
rect 14659 23315 14697 23316
rect 14753 23315 14791 23316
rect 14847 23315 14885 23316
rect 14941 23315 14979 23316
rect 15035 23315 15040 23371
rect 14504 23299 15040 23315
rect 14504 23289 14510 23299
rect 14504 23233 14509 23289
rect 14574 23235 14602 23299
rect 14666 23235 14694 23299
rect 14758 23235 14786 23299
rect 14850 23235 14878 23299
rect 14942 23235 14970 23299
rect 15034 23289 15040 23299
rect 14565 23233 14603 23235
rect 14659 23233 14697 23235
rect 14753 23233 14791 23235
rect 14847 23233 14885 23235
rect 14941 23233 14979 23235
rect 15035 23233 15040 23289
rect 14504 23218 15040 23233
rect 14504 23207 14510 23218
rect 14504 23151 14509 23207
rect 14574 23154 14602 23218
rect 14666 23154 14694 23218
rect 14758 23154 14786 23218
rect 14850 23154 14878 23218
rect 14942 23154 14970 23218
rect 15034 23207 15040 23218
rect 14565 23151 14603 23154
rect 14659 23151 14697 23154
rect 14753 23151 14791 23154
rect 14847 23151 14885 23154
rect 14941 23151 14979 23154
rect 15035 23151 15040 23207
rect 14504 23146 15040 23151
tri 13579 21847 13693 21961 ne
rect 13693 21847 14391 21961
tri 14391 21847 15107 22563 sw
tri 4099 21317 4215 21433 ne
rect 4215 21317 5099 21433
tri 5099 21317 5629 21847 sw
tri 13693 21583 13957 21847 ne
rect 13957 21583 15107 21847
tri 15107 21583 15371 21847 sw
tri 13957 21317 14223 21583 ne
rect 14223 21317 15371 21583
tri 4215 21282 4250 21317 ne
rect 4250 21282 5629 21317
tri 5629 21282 5664 21317 sw
tri 14223 21282 14258 21317 ne
rect 14258 21282 15371 21317
tri 4250 21171 4361 21282 ne
rect 4361 21171 5664 21282
tri 5664 21171 5775 21282 sw
tri 14258 21171 14369 21282 ne
rect 14369 21171 15371 21282
tri 4361 21099 4433 21171 ne
rect 4433 21099 5775 21171
tri 5775 21099 5847 21171 sw
tri 14369 21149 14391 21171 ne
rect 14391 21149 15371 21171
tri 14391 21112 14428 21149 ne
tri 4433 20955 4577 21099 ne
rect 4577 20955 5847 21099
tri 5847 20955 5991 21099 sw
rect 2781 20875 2790 20931
rect 2846 20875 2873 20931
rect 2929 20875 2956 20931
rect 3012 20875 3039 20931
rect 3095 20875 3122 20931
rect 3178 20875 3205 20931
rect 3261 20875 3288 20931
rect 3344 20875 3371 20931
rect 3427 20875 3454 20931
rect 3510 20875 3537 20931
rect 3593 20875 3620 20931
rect 3676 20875 3703 20931
rect 3759 20875 3778 20931
rect 2781 20837 3778 20875
rect 2781 20781 2790 20837
rect 2846 20781 2873 20837
rect 2929 20781 2956 20837
rect 3012 20781 3039 20837
rect 3095 20781 3122 20837
rect 3178 20781 3205 20837
rect 3261 20781 3288 20837
rect 3344 20781 3371 20837
rect 3427 20781 3454 20837
rect 3510 20781 3537 20837
rect 3593 20781 3620 20837
rect 3676 20781 3703 20837
rect 3759 20781 3778 20837
rect 2781 20743 3778 20781
rect 2781 20687 2790 20743
rect 2846 20687 2873 20743
rect 2929 20687 2956 20743
rect 3012 20687 3039 20743
rect 3095 20687 3122 20743
rect 3178 20687 3205 20743
rect 3261 20687 3288 20743
rect 3344 20687 3371 20743
rect 3427 20687 3454 20743
rect 3510 20687 3537 20743
rect 3593 20687 3620 20743
rect 3676 20687 3703 20743
rect 3759 20687 3778 20743
rect 2781 20649 3778 20687
rect 2781 20593 2790 20649
rect 2846 20593 2873 20649
rect 2929 20593 2956 20649
rect 3012 20593 3039 20649
rect 3095 20593 3122 20649
rect 3178 20593 3205 20649
rect 3261 20593 3288 20649
rect 3344 20593 3371 20649
rect 3427 20593 3454 20649
rect 3510 20593 3537 20649
rect 3593 20593 3620 20649
rect 3676 20593 3703 20649
rect 3759 20593 3778 20649
rect 2781 20555 3778 20593
rect 2781 20499 2790 20555
rect 2846 20499 2873 20555
rect 2929 20499 2956 20555
rect 3012 20499 3039 20555
rect 3095 20499 3122 20555
rect 3178 20499 3205 20555
rect 3261 20499 3288 20555
rect 3344 20499 3371 20555
rect 3427 20499 3454 20555
rect 3510 20499 3537 20555
rect 3593 20499 3620 20555
rect 3676 20499 3703 20555
rect 3759 20499 3778 20555
tri 4577 20541 4991 20955 ne
rect 2781 20461 3778 20499
rect 2781 20405 2790 20461
rect 2846 20405 2873 20461
rect 2929 20405 2956 20461
rect 3012 20405 3039 20461
rect 3095 20405 3122 20461
rect 3178 20405 3205 20461
rect 3261 20405 3288 20461
rect 3344 20405 3371 20461
rect 3427 20405 3454 20461
rect 3510 20405 3537 20461
rect 3593 20405 3620 20461
rect 3676 20405 3703 20461
rect 3759 20405 3778 20461
rect 356 18912 392 18976
rect 456 18912 492 18976
rect 556 18912 592 18976
rect 292 18896 656 18912
rect 356 18832 392 18896
rect 456 18832 492 18896
rect 556 18832 592 18896
rect 292 18816 656 18832
rect 356 18752 392 18816
rect 456 18752 492 18816
rect 556 18752 592 18816
rect 292 18736 656 18752
rect 356 18672 392 18736
rect 456 18672 492 18736
rect 556 18672 592 18736
rect 292 18656 656 18672
rect 356 18592 392 18656
rect 456 18592 492 18656
rect 556 18592 592 18656
rect 292 18576 656 18592
rect 356 18512 392 18576
rect 456 18512 492 18576
rect 556 18512 592 18576
rect 292 18496 656 18512
rect 356 18432 392 18496
rect 456 18432 492 18496
rect 556 18432 592 18496
rect 292 18416 656 18432
rect 356 18352 392 18416
rect 456 18352 492 18416
rect 556 18352 592 18416
rect 292 18336 656 18352
rect 356 18272 392 18336
rect 456 18272 492 18336
rect 556 18272 592 18336
rect 292 18256 656 18272
rect 356 18192 392 18256
rect 456 18192 492 18256
rect 556 18192 592 18256
rect 292 18176 656 18192
rect 356 18112 392 18176
rect 456 18112 492 18176
rect 556 18112 592 18176
tri 1276 20079 1365 20168 se
rect 1365 20079 2275 20168
tri 2275 20079 2364 20168 nw
rect 1276 20068 2264 20079
tri 2264 20068 2275 20079 nw
rect 1276 18312 1376 20068
tri 1376 19950 1494 20068 nw
rect 2781 19243 3778 20405
rect 2781 19187 2790 19243
rect 2846 19187 2874 19243
rect 2930 19187 2958 19243
rect 3014 19187 3042 19243
rect 3098 19187 3126 19243
rect 3182 19187 3210 19243
rect 3266 19187 3294 19243
rect 3350 19187 3378 19243
rect 3434 19187 3462 19243
rect 3518 19187 3546 19243
rect 3602 19187 3630 19243
rect 3686 19187 3713 19243
rect 3769 19187 3778 19243
rect 2781 19073 3778 19187
rect 2781 19017 3025 19073
rect 3081 19017 3111 19073
rect 3167 19017 3197 19073
rect 3253 19017 3283 19073
rect 3339 19017 3369 19073
rect 3425 19017 3455 19073
rect 3511 19017 3541 19073
rect 3597 19017 3627 19073
rect 3683 19017 3713 19073
rect 3769 19017 3778 19073
tri 1376 18312 1384 18320 sw
rect 1276 18278 1384 18312
tri 1384 18278 1418 18312 sw
tri 1276 18170 1384 18278 ne
rect 1384 18212 1418 18278
tri 1418 18212 1484 18278 sw
rect 292 18096 656 18112
rect 356 18032 392 18096
rect 456 18032 492 18096
rect 556 18032 592 18096
rect 292 18015 656 18032
rect 356 17951 392 18015
rect 456 17951 492 18015
rect 556 17951 592 18015
rect 292 17934 656 17951
rect 356 17870 392 17934
rect 456 17870 492 17934
rect 556 17870 592 17934
rect 292 17853 656 17870
rect 356 17789 392 17853
rect 456 17789 492 17853
rect 556 17789 592 17853
rect 292 17772 656 17789
rect 356 17708 392 17772
rect 456 17708 492 17772
rect 556 17708 592 17772
rect 292 17691 656 17708
rect 356 17627 392 17691
rect 456 17627 492 17691
rect 556 17627 592 17691
rect 292 17610 656 17627
rect 356 17546 392 17610
rect 456 17546 492 17610
rect 556 17546 592 17610
rect 292 17529 656 17546
rect 356 17465 392 17529
rect 456 17465 492 17529
rect 556 17465 592 17529
rect 292 17448 656 17465
rect 356 17384 392 17448
rect 456 17384 492 17448
rect 556 17384 592 17448
rect 292 17367 656 17384
rect 356 17303 392 17367
rect 456 17303 492 17367
rect 556 17303 592 17367
rect 292 17286 656 17303
rect 356 17222 392 17286
rect 456 17222 492 17286
rect 556 17222 592 17286
rect 292 17205 656 17222
rect 356 17141 392 17205
rect 456 17141 492 17205
rect 556 17141 592 17205
rect 292 17124 656 17141
rect 356 17060 392 17124
rect 456 17060 492 17124
rect 556 17060 592 17124
rect 292 17043 656 17060
rect 356 16979 392 17043
rect 456 16979 492 17043
rect 556 16979 592 17043
rect 292 16962 656 16979
rect 356 16898 392 16962
rect 456 16898 492 16962
rect 556 16898 592 16962
rect 292 16881 656 16898
rect 356 16817 392 16881
rect 456 16817 492 16881
rect 556 16817 592 16881
rect 292 16800 656 16817
rect 356 16736 392 16800
rect 456 16736 492 16800
rect 556 16736 592 16800
rect 292 16719 656 16736
rect 356 16655 392 16719
rect 456 16655 492 16719
rect 556 16655 592 16719
rect 292 16638 656 16655
rect 356 16574 392 16638
rect 456 16574 492 16638
rect 556 16574 592 16638
rect 292 16557 656 16574
rect 356 16493 392 16557
rect 456 16493 492 16557
rect 556 16493 592 16557
rect 292 16476 656 16493
rect 356 16412 392 16476
rect 456 16412 492 16476
rect 556 16412 592 16476
rect 292 16395 656 16412
rect 356 16331 392 16395
rect 456 16331 492 16395
rect 556 16331 592 16395
rect 292 16314 656 16331
rect 356 16250 392 16314
rect 456 16250 492 16314
rect 556 16250 592 16314
rect 292 16233 656 16250
rect 356 16169 392 16233
rect 456 16169 492 16233
rect 556 16169 592 16233
rect 292 16152 656 16169
rect 356 16088 392 16152
rect 456 16088 492 16152
rect 556 16088 592 16152
rect 292 16071 656 16088
rect 356 16007 392 16071
rect 456 16007 492 16071
rect 556 16007 592 16071
rect 292 15990 656 16007
rect 356 15926 392 15990
rect 456 15926 492 15990
rect 556 15926 592 15990
rect 292 15909 656 15926
rect 356 15845 392 15909
rect 456 15845 492 15909
rect 556 15845 592 15909
rect 292 15828 656 15845
rect 356 15764 392 15828
rect 456 15764 492 15828
rect 556 15764 592 15828
rect 292 15747 656 15764
rect 356 15683 392 15747
rect 456 15683 492 15747
rect 556 15683 592 15747
rect 292 15666 656 15683
rect 356 15602 392 15666
rect 456 15602 492 15666
rect 556 15602 592 15666
rect 292 15585 656 15602
rect 356 15521 392 15585
rect 456 15521 492 15585
rect 556 15521 592 15585
rect 292 15504 656 15521
rect 356 15440 392 15504
rect 456 15440 492 15504
rect 556 15440 592 15504
rect 292 15423 656 15440
rect 356 15359 392 15423
rect 456 15359 492 15423
rect 556 15359 592 15423
rect 292 15342 656 15359
rect 356 15278 392 15342
rect 456 15278 492 15342
rect 556 15278 592 15342
rect 292 15261 656 15278
rect 356 15197 392 15261
rect 456 15197 492 15261
rect 556 15197 592 15261
rect 292 15180 656 15197
rect 356 15116 392 15180
rect 456 15116 492 15180
rect 556 15116 592 15180
rect 292 15099 656 15116
rect 356 15035 392 15099
rect 456 15035 492 15099
rect 556 15035 592 15099
rect 292 15018 656 15035
rect 356 14954 392 15018
rect 456 14954 492 15018
rect 556 14954 592 15018
tri 1242 14988 1384 15130 se
rect 1384 15088 1484 18212
tri 1384 14988 1484 15088 nw
rect 2781 17353 3778 19017
rect 2781 17297 3207 17353
rect 3263 17297 3289 17353
rect 3345 17297 3778 17353
rect 292 14937 656 14954
rect 356 14873 392 14937
rect 456 14873 492 14937
rect 556 14873 592 14937
rect 292 14856 656 14873
rect 356 14792 392 14856
rect 456 14792 492 14856
rect 556 14792 592 14856
rect 292 14775 656 14792
rect 356 14711 392 14775
rect 456 14711 492 14775
rect 556 14711 592 14775
rect 292 14694 656 14711
rect 356 14630 392 14694
rect 456 14630 492 14694
rect 556 14630 592 14694
rect 292 14613 656 14630
rect 356 14549 392 14613
rect 456 14549 492 14613
rect 556 14549 592 14613
rect 292 14532 656 14549
rect 356 14468 392 14532
rect 456 14468 492 14532
rect 556 14468 592 14532
rect 292 14451 656 14468
rect 356 14387 392 14451
rect 456 14387 492 14451
rect 556 14387 592 14451
rect 292 14370 656 14387
rect 356 14306 392 14370
rect 456 14306 492 14370
rect 556 14306 592 14370
rect 292 14289 656 14306
rect 356 14225 392 14289
rect 456 14225 492 14289
rect 556 14225 592 14289
rect 292 14208 656 14225
rect 356 14144 392 14208
rect 456 14144 492 14208
rect 556 14144 592 14208
rect 292 14127 656 14144
rect 356 14063 392 14127
rect 456 14063 492 14127
rect 556 14063 592 14127
rect 292 14057 656 14063
tri 1188 14934 1242 14988 se
rect 1242 14934 1330 14988
tri 1330 14934 1384 14988 nw
rect 516 11282 522 11346
rect 586 11282 606 11346
rect 670 11282 690 11346
rect 754 11282 760 11346
rect 516 10563 760 11282
rect 516 10499 522 10563
rect 586 10499 606 10563
rect 670 10499 690 10563
rect 754 10499 760 10563
rect 516 10479 760 10499
rect 516 10415 522 10479
rect 586 10415 606 10479
rect 670 10415 690 10479
rect 754 10415 760 10479
rect 516 10395 760 10415
rect 516 10331 522 10395
rect 586 10331 606 10395
rect 670 10331 690 10395
rect 754 10331 760 10395
rect 516 9612 760 10331
rect 516 9548 522 9612
rect 586 9548 606 9612
rect 670 9548 690 9612
rect 754 9548 760 9612
tri 1132 9472 1188 9528 se
rect 1188 9472 1288 14934
tri 1288 14892 1330 14934 nw
rect 1370 13596 1570 13605
rect 1370 13532 1372 13596
rect 1436 13532 1502 13596
rect 1566 13532 1570 13596
rect 1370 13509 1570 13532
rect 1370 13445 1372 13509
rect 1436 13445 1502 13509
rect 1566 13445 1570 13509
rect 1370 13422 1570 13445
rect 1370 13358 1372 13422
rect 1436 13358 1502 13422
rect 1566 13358 1570 13422
rect 1370 13335 1570 13358
rect 1370 13271 1372 13335
rect 1436 13271 1502 13335
rect 1566 13271 1570 13335
rect 1370 13248 1570 13271
rect 1370 13184 1372 13248
rect 1436 13184 1502 13248
rect 1566 13184 1570 13248
rect 1370 13161 1570 13184
rect 1370 13097 1372 13161
rect 1436 13097 1502 13161
rect 1566 13097 1570 13161
rect 1370 13074 1570 13097
rect 1370 13010 1372 13074
rect 1436 13010 1502 13074
rect 1566 13010 1570 13074
rect 1370 12986 1570 13010
rect 1370 12922 1372 12986
rect 1436 12922 1502 12986
rect 1566 12922 1570 12986
rect 1370 12898 1570 12922
rect 1370 12834 1372 12898
rect 1436 12834 1502 12898
rect 1566 12834 1570 12898
rect 1370 9923 1570 12834
rect 2781 10398 3778 17297
rect 4991 18320 5991 20955
rect 13738 20376 13952 20382
rect 13802 20312 13888 20376
rect 13738 20282 13952 20312
rect 13802 20218 13888 20282
rect 13738 20188 13952 20218
rect 13802 20124 13888 20188
rect 13738 20094 13952 20124
rect 13802 20030 13888 20094
rect 13738 19999 13952 20030
rect 13802 19935 13888 19999
rect 13738 19904 13952 19935
rect 13802 19840 13888 19904
tri 5991 18457 6039 18505 sw
tri 5991 18320 6001 18330 sw
rect 4991 18312 6001 18320
tri 6001 18312 6009 18320 sw
rect 4991 18282 6009 18312
tri 6009 18282 6039 18312 sw
rect 3889 16383 4620 16388
rect 3889 16327 3894 16383
rect 3950 16327 4019 16383
rect 4075 16327 4144 16383
rect 4200 16327 4269 16383
rect 4325 16363 4620 16383
tri 4620 16363 4645 16388 sw
rect 4325 16327 4645 16363
rect 3889 16307 4645 16327
tri 4645 16307 4701 16363 sw
rect 3889 16303 4701 16307
rect 3889 16247 3894 16303
rect 3950 16247 4019 16303
rect 4075 16247 4144 16303
rect 4200 16247 4269 16303
rect 4325 16275 4701 16303
tri 4701 16275 4733 16307 sw
rect 4325 16247 4733 16275
rect 3889 16223 4733 16247
rect 3889 16167 3894 16223
rect 3950 16167 4019 16223
rect 4075 16167 4144 16223
rect 4200 16167 4269 16223
rect 4325 16219 4733 16223
tri 4733 16219 4789 16275 sw
rect 4325 16167 4789 16219
rect 3889 16162 4789 16167
tri 4789 16162 4846 16219 sw
tri 3957 16125 3994 16162 ne
rect 3994 16125 4846 16162
tri 4846 16125 4883 16162 sw
tri 3994 15832 4287 16125 ne
rect 2781 10342 2999 10398
rect 3055 10342 3088 10398
rect 3144 10342 3177 10398
rect 3233 10342 3265 10398
rect 3321 10342 3353 10398
rect 3409 10342 3441 10398
rect 3497 10342 3529 10398
rect 3585 10342 3617 10398
rect 3673 10342 3705 10398
rect 3761 10342 3778 10398
rect 2781 10318 3778 10342
rect 2781 10262 2999 10318
rect 3055 10262 3088 10318
rect 3144 10262 3177 10318
rect 3233 10262 3265 10318
rect 3321 10262 3353 10318
rect 3409 10262 3441 10318
rect 3497 10262 3529 10318
rect 3585 10262 3617 10318
rect 3673 10262 3705 10318
rect 3761 10262 3778 10318
rect 2225 10044 2699 10051
rect 2225 9988 2234 10044
rect 2290 9988 2333 10044
rect 2389 9988 2431 10044
rect 2487 9988 2529 10044
rect 2585 9988 2627 10044
rect 2683 9988 2699 10044
rect 2225 9950 2699 9988
rect 1132 9408 1138 9472
rect 1202 9408 1218 9472
rect 1282 9408 1288 9472
rect 2225 9894 2234 9950
rect 2290 9894 2333 9950
rect 2389 9894 2431 9950
rect 2487 9894 2529 9950
rect 2585 9894 2627 9950
rect 2683 9894 2699 9950
rect 2225 9856 2699 9894
rect 2225 9800 2234 9856
rect 2290 9800 2333 9856
rect 2389 9800 2431 9856
rect 2487 9800 2529 9856
rect 2585 9800 2627 9856
rect 2683 9800 2699 9856
rect 2225 9762 2699 9800
rect 2225 9706 2234 9762
rect 2290 9706 2333 9762
rect 2389 9706 2431 9762
rect 2487 9706 2529 9762
rect 2585 9706 2627 9762
rect 2683 9706 2699 9762
rect 1485 8077 2143 8082
rect 1485 8021 1536 8077
rect 1592 8021 1626 8077
rect 1682 8021 1716 8077
rect 1772 8021 1806 8077
rect 1862 8021 1896 8077
rect 1952 8021 1986 8077
rect 2042 8021 2076 8077
rect 2132 8021 2143 8077
rect 1485 7993 2143 8021
rect 1485 7937 1536 7993
rect 1592 7937 1626 7993
rect 1682 7937 1716 7993
rect 1772 7937 1806 7993
rect 1862 7937 1896 7993
rect 1952 7937 1986 7993
rect 2042 7937 2076 7993
rect 2132 7937 2143 7993
rect 1485 7909 2143 7937
rect 1485 7853 1536 7909
rect 1592 7853 1626 7909
rect 1682 7853 1716 7909
rect 1772 7853 1806 7909
rect 1862 7853 1896 7909
rect 1952 7853 1986 7909
rect 2042 7853 2076 7909
rect 2132 7853 2143 7909
rect 1485 7825 2143 7853
rect 1485 7769 1536 7825
rect 1592 7769 1626 7825
rect 1682 7769 1716 7825
rect 1772 7769 1806 7825
rect 1862 7769 1896 7825
rect 1952 7769 1986 7825
rect 2042 7769 2076 7825
rect 2132 7769 2143 7825
rect 1485 7741 2143 7769
rect 1485 7685 1536 7741
rect 1592 7685 1626 7741
rect 1682 7685 1716 7741
rect 1772 7685 1806 7741
rect 1862 7685 1896 7741
rect 1952 7685 1986 7741
rect 2042 7685 2076 7741
rect 2132 7685 2143 7741
rect 1485 7657 2143 7685
rect 1485 7601 1536 7657
rect 1592 7601 1626 7657
rect 1682 7601 1716 7657
rect 1772 7601 1806 7657
rect 1862 7601 1896 7657
rect 1952 7601 1986 7657
rect 2042 7601 2076 7657
rect 2132 7601 2143 7657
rect 1485 7573 2143 7601
rect 1485 7517 1536 7573
rect 1592 7517 1626 7573
rect 1682 7517 1716 7573
rect 1772 7517 1806 7573
rect 1862 7517 1896 7573
rect 1952 7517 1986 7573
rect 2042 7517 2076 7573
rect 2132 7517 2143 7573
rect 1485 7489 2143 7517
rect 1485 7433 1536 7489
rect 1592 7433 1626 7489
rect 1682 7433 1716 7489
rect 1772 7433 1806 7489
rect 1862 7433 1896 7489
rect 1952 7433 1986 7489
rect 2042 7433 2076 7489
rect 2132 7433 2143 7489
rect 1485 7405 2143 7433
rect 1485 7349 1536 7405
rect 1592 7349 1626 7405
rect 1682 7349 1716 7405
rect 1772 7349 1806 7405
rect 1862 7349 1896 7405
rect 1952 7349 1986 7405
rect 2042 7349 2076 7405
rect 2132 7349 2143 7405
rect 1485 7321 2143 7349
rect 1485 7265 1536 7321
rect 1592 7265 1626 7321
rect 1682 7265 1716 7321
rect 1772 7265 1806 7321
rect 1862 7265 1896 7321
rect 1952 7265 1986 7321
rect 2042 7265 2076 7321
rect 2132 7265 2143 7321
rect 905 7174 911 7238
rect 975 7174 991 7238
rect 1055 7174 1061 7238
tri 905 7153 926 7174 ne
rect 926 7153 1041 7174
tri 1041 7154 1061 7174 nw
rect 1485 7237 2143 7265
rect 1485 7181 1536 7237
rect 1592 7181 1626 7237
rect 1682 7181 1716 7237
rect 1772 7181 1806 7237
rect 1862 7181 1896 7237
rect 1952 7181 1986 7237
rect 2042 7181 2076 7237
rect 2132 7181 2143 7237
tri 926 7152 927 7153 ne
rect 927 7152 1041 7153
tri 927 7102 977 7152 ne
tri 976 4852 977 4853 se
rect 977 4852 1041 7152
tri 952 4828 976 4852 se
rect 976 4828 1041 4852
tri 896 4772 952 4828 se
rect 952 4827 1041 4828
rect 952 4772 986 4827
tri 986 4772 1041 4827 nw
rect 1485 7152 2143 7181
rect 1485 7096 1536 7152
rect 1592 7096 1626 7152
rect 1682 7096 1716 7152
rect 1772 7096 1806 7152
rect 1862 7096 1896 7152
rect 1952 7096 1986 7152
rect 2042 7096 2076 7152
rect 2132 7096 2143 7152
rect 1485 7067 2143 7096
rect 1485 7011 1536 7067
rect 1592 7011 1626 7067
rect 1682 7011 1716 7067
rect 1772 7011 1806 7067
rect 1862 7011 1896 7067
rect 1952 7011 1986 7067
rect 2042 7011 2076 7067
rect 2132 7011 2143 7067
rect 1485 6982 2143 7011
rect 1485 6926 1536 6982
rect 1592 6926 1626 6982
rect 1682 6926 1716 6982
rect 1772 6926 1806 6982
rect 1862 6926 1896 6982
rect 1952 6926 1986 6982
rect 2042 6926 2076 6982
rect 2132 6926 2143 6982
rect 1485 6897 2143 6926
rect 1485 6841 1536 6897
rect 1592 6841 1626 6897
rect 1682 6841 1716 6897
rect 1772 6841 1806 6897
rect 1862 6841 1896 6897
rect 1952 6841 1986 6897
rect 2042 6841 2076 6897
rect 2132 6841 2143 6897
rect 1485 6812 2143 6841
rect 1485 6756 1536 6812
rect 1592 6756 1626 6812
rect 1682 6756 1716 6812
rect 1772 6756 1806 6812
rect 1862 6756 1896 6812
rect 1952 6756 1986 6812
rect 2042 6756 2076 6812
rect 2132 6756 2143 6812
rect 1485 6727 2143 6756
rect 1485 6671 1536 6727
rect 1592 6671 1626 6727
rect 1682 6671 1716 6727
rect 1772 6671 1806 6727
rect 1862 6671 1896 6727
rect 1952 6671 1986 6727
rect 2042 6671 2076 6727
rect 2132 6671 2143 6727
rect 1485 6635 2143 6671
rect 1485 6579 1709 6635
rect 1765 6579 1797 6635
rect 1853 6579 1885 6635
rect 1941 6579 1973 6635
rect 2029 6579 2061 6635
rect 2117 6579 2143 6635
rect 1485 6551 2143 6579
rect 1485 6495 1709 6551
rect 1765 6495 1797 6551
rect 1853 6495 1885 6551
rect 1941 6495 1973 6551
rect 2029 6495 2061 6551
rect 2117 6495 2143 6551
rect 1485 6467 2143 6495
rect 1485 6411 1709 6467
rect 1765 6411 1797 6467
rect 1853 6411 1885 6467
rect 1941 6411 1973 6467
rect 2029 6411 2061 6467
rect 2117 6411 2143 6467
rect 1485 6383 2143 6411
rect 1485 6327 1709 6383
rect 1765 6327 1797 6383
rect 1853 6327 1885 6383
rect 1941 6327 1973 6383
rect 2029 6327 2061 6383
rect 2117 6327 2143 6383
rect 1485 6299 2143 6327
rect 1485 6243 1709 6299
rect 1765 6243 1797 6299
rect 1853 6243 1885 6299
rect 1941 6243 1973 6299
rect 2029 6243 2061 6299
rect 2117 6243 2143 6299
rect 1485 6215 2143 6243
rect 1485 6159 1709 6215
rect 1765 6159 1797 6215
rect 1853 6159 1885 6215
rect 1941 6159 1973 6215
rect 2029 6159 2061 6215
rect 2117 6159 2143 6215
rect 1485 6131 2143 6159
rect 1485 6075 1709 6131
rect 1765 6075 1797 6131
rect 1853 6075 1885 6131
rect 1941 6075 1973 6131
rect 2029 6075 2061 6131
rect 2117 6075 2143 6131
rect 1485 6046 2143 6075
rect 1485 5990 1709 6046
rect 1765 5990 1797 6046
rect 1853 5990 1885 6046
rect 1941 5990 1973 6046
rect 2029 5990 2061 6046
rect 2117 5990 2143 6046
rect 1485 5961 2143 5990
rect 1485 5905 1709 5961
rect 1765 5905 1797 5961
rect 1853 5905 1885 5961
rect 1941 5905 1973 5961
rect 2029 5905 2061 5961
rect 2117 5905 2143 5961
rect 1485 5836 2143 5905
rect 1485 5780 1708 5836
rect 1764 5780 1814 5836
rect 1870 5780 1920 5836
rect 1976 5780 2143 5836
rect 1485 5754 2143 5780
rect 1485 5698 1708 5754
rect 1764 5698 1814 5754
rect 1870 5698 1920 5754
rect 1976 5698 2143 5754
rect 1485 5672 2143 5698
rect 1485 5616 1708 5672
rect 1764 5616 1814 5672
rect 1870 5616 1920 5672
rect 1976 5616 2143 5672
rect 1485 5590 2143 5616
rect 1485 5534 1708 5590
rect 1764 5534 1814 5590
rect 1870 5534 1920 5590
rect 1976 5534 2143 5590
rect 1485 5508 2143 5534
rect 1485 5452 1708 5508
rect 1764 5452 1814 5508
rect 1870 5452 1920 5508
rect 1976 5452 2143 5508
rect 1485 5426 2143 5452
rect 1485 5370 1708 5426
rect 1764 5370 1814 5426
rect 1870 5370 1920 5426
rect 1976 5370 2143 5426
rect 1485 5343 2143 5370
rect 1485 5287 1708 5343
rect 1764 5287 1814 5343
rect 1870 5287 1920 5343
rect 1976 5287 2143 5343
rect 1485 5228 2143 5287
rect 1485 5172 1709 5228
rect 1765 5172 1797 5228
rect 1853 5172 1885 5228
rect 1941 5172 1973 5228
rect 2029 5172 2061 5228
rect 2117 5172 2143 5228
rect 1485 5148 2143 5172
rect 1485 5092 1709 5148
rect 1765 5092 1797 5148
rect 1853 5092 1885 5148
rect 1941 5092 1973 5148
rect 2029 5092 2061 5148
rect 2117 5092 2143 5148
rect 1485 5068 2143 5092
rect 1485 5012 1709 5068
rect 1765 5012 1797 5068
rect 1853 5012 1885 5068
rect 1941 5012 1973 5068
rect 2029 5012 2061 5068
rect 2117 5012 2143 5068
rect 1485 4988 2143 5012
rect 1485 4932 1709 4988
rect 1765 4932 1797 4988
rect 1853 4932 1885 4988
rect 1941 4932 1973 4988
rect 2029 4932 2061 4988
rect 2117 4932 2143 4988
rect 1485 4908 2143 4932
rect 1485 4886 1709 4908
rect 1765 4886 1797 4908
rect 1853 4886 1885 4908
rect 1941 4886 1973 4908
rect 2029 4886 2061 4908
rect 2117 4886 2143 4908
rect 1485 4822 1486 4886
rect 1550 4822 1570 4886
rect 1634 4822 1654 4886
rect 1970 4852 1973 4886
rect 2054 4852 2061 4886
rect 1718 4828 1738 4852
rect 1802 4828 1822 4852
rect 1886 4828 1906 4852
rect 1970 4828 1990 4852
rect 2054 4828 2074 4852
rect 1970 4822 1973 4828
rect 2054 4822 2061 4828
rect 2138 4822 2143 4886
rect 1485 4800 1709 4822
rect 1765 4800 1797 4822
rect 1853 4800 1885 4822
rect 1941 4800 1973 4822
rect 2029 4800 2061 4822
rect 2117 4800 2143 4822
tri 887 4763 896 4772 se
rect 896 4763 977 4772
tri 977 4763 986 4772 nw
tri 871 4747 887 4763 se
rect 887 4747 961 4763
tri 961 4747 977 4763 nw
tri 852 4728 871 4747 se
rect 871 4728 942 4747
tri 942 4728 961 4747 nw
rect 1485 4736 1486 4800
rect 1550 4736 1570 4800
rect 1634 4736 1654 4800
rect 1970 4772 1973 4800
rect 2054 4772 2061 4800
rect 1718 4747 1738 4772
rect 1802 4747 1822 4772
rect 1886 4747 1906 4772
rect 1970 4747 1990 4772
rect 2054 4747 2074 4772
rect 1970 4736 1973 4747
rect 2054 4736 2061 4747
rect 2138 4736 2143 4800
rect 852 3811 916 4728
tri 916 4702 942 4728 nw
rect 1485 4714 1709 4736
rect 1765 4714 1797 4736
rect 1853 4714 1885 4736
rect 1941 4714 1973 4736
rect 2029 4714 2061 4736
rect 2117 4714 2143 4736
rect 1485 4650 1486 4714
rect 1550 4650 1570 4714
rect 1634 4650 1654 4714
rect 1970 4691 1973 4714
rect 2054 4691 2061 4714
rect 1718 4666 1738 4691
rect 1802 4666 1822 4691
rect 1886 4666 1906 4691
rect 1970 4666 1990 4691
rect 2054 4666 2074 4691
rect 1970 4650 1973 4666
rect 2054 4650 2061 4666
rect 2138 4650 2143 4714
rect 1485 4628 1709 4650
rect 1765 4628 1797 4650
rect 1853 4628 1885 4650
rect 1941 4628 1973 4650
rect 2029 4628 2061 4650
rect 2117 4628 2143 4650
rect 1485 4564 1486 4628
rect 1550 4564 1570 4628
rect 1634 4564 1654 4628
rect 1970 4610 1973 4628
rect 2054 4610 2061 4628
rect 1718 4585 1738 4610
rect 1802 4585 1822 4610
rect 1886 4585 1906 4610
rect 1970 4585 1990 4610
rect 2054 4585 2074 4610
rect 1970 4564 1973 4585
rect 2054 4564 2061 4585
rect 2138 4564 2143 4628
rect 1485 4542 1709 4564
rect 1765 4542 1797 4564
rect 1853 4542 1885 4564
rect 1941 4542 1973 4564
rect 2029 4542 2061 4564
rect 2117 4542 2143 4564
rect 1485 4478 1486 4542
rect 1550 4478 1570 4542
rect 1634 4478 1654 4542
rect 1970 4529 1973 4542
rect 2054 4529 2061 4542
rect 1718 4504 1738 4529
rect 1802 4504 1822 4529
rect 1886 4504 1906 4529
rect 1970 4504 1990 4529
rect 2054 4504 2074 4529
rect 1970 4478 1973 4504
rect 2054 4478 2061 4504
rect 2138 4478 2143 4542
rect 1485 4456 1709 4478
rect 1765 4456 1797 4478
rect 1853 4456 1885 4478
rect 1941 4456 1973 4478
rect 2029 4456 2061 4478
rect 2117 4456 2143 4478
rect 1485 4392 1486 4456
rect 1550 4392 1570 4456
rect 1634 4392 1654 4456
rect 1970 4448 1973 4456
rect 2054 4448 2061 4456
rect 1718 4423 1738 4448
rect 1802 4423 1822 4448
rect 1886 4423 1906 4448
rect 1970 4423 1990 4448
rect 2054 4423 2074 4448
rect 1970 4392 1973 4423
rect 2054 4392 2061 4423
rect 2138 4392 2143 4456
rect 1485 4370 1709 4392
rect 1765 4370 1797 4392
rect 1853 4370 1885 4392
rect 1941 4370 1973 4392
rect 2029 4370 2061 4392
rect 2117 4370 2143 4392
rect 1485 4306 1486 4370
rect 1550 4306 1570 4370
rect 1634 4306 1654 4370
rect 1970 4367 1973 4370
rect 2054 4367 2061 4370
rect 1718 4342 1738 4367
rect 1802 4342 1822 4367
rect 1886 4342 1906 4367
rect 1970 4342 1990 4367
rect 2054 4342 2074 4367
rect 1970 4306 1973 4342
rect 2054 4306 2061 4342
rect 2138 4306 2143 4370
rect 1485 4286 1709 4306
rect 1765 4286 1797 4306
rect 1853 4286 1885 4306
rect 1941 4286 1973 4306
rect 2029 4286 2061 4306
rect 2117 4286 2143 4306
rect 1485 4283 2143 4286
rect 1485 4219 1486 4283
rect 1550 4219 1570 4283
rect 1634 4219 1654 4283
rect 1718 4261 1738 4283
rect 1802 4261 1822 4283
rect 1886 4261 1906 4283
rect 1970 4261 1990 4283
rect 2054 4261 2074 4283
rect 1970 4219 1973 4261
rect 2054 4219 2061 4261
rect 2138 4219 2143 4283
rect 1485 4205 1709 4219
rect 1765 4205 1797 4219
rect 1853 4205 1885 4219
rect 1941 4205 1973 4219
rect 2029 4205 2061 4219
rect 2117 4205 2143 4219
rect 1485 4196 2143 4205
rect 1485 4132 1486 4196
rect 1550 4132 1570 4196
rect 1634 4132 1654 4196
rect 1718 4180 1738 4196
rect 1802 4180 1822 4196
rect 1886 4180 1906 4196
rect 1970 4180 1990 4196
rect 2054 4180 2074 4196
rect 1970 4132 1973 4180
rect 2054 4132 2061 4180
rect 2138 4132 2143 4196
rect 1485 4124 1709 4132
rect 1765 4124 1797 4132
rect 1853 4124 1885 4132
rect 1941 4124 1973 4132
rect 2029 4124 2061 4132
rect 2117 4124 2143 4132
rect 1485 4109 2143 4124
rect 1485 4045 1486 4109
rect 1550 4045 1570 4109
rect 1634 4045 1654 4109
rect 1718 4099 1738 4109
rect 1802 4099 1822 4109
rect 1886 4099 1906 4109
rect 1970 4099 1990 4109
rect 2054 4099 2074 4109
rect 1970 4045 1973 4099
rect 2054 4045 2061 4099
rect 2138 4045 2143 4109
rect 1485 4043 1709 4045
rect 1765 4043 1797 4045
rect 1853 4043 1885 4045
rect 1941 4043 1973 4045
rect 2029 4043 2061 4045
rect 2117 4043 2143 4045
rect 1485 4022 2143 4043
rect 1485 3958 1486 4022
rect 1550 3958 1570 4022
rect 1634 3958 1654 4022
rect 1718 4018 1738 4022
rect 1802 4018 1822 4022
rect 1886 4018 1906 4022
rect 1970 4018 1990 4022
rect 2054 4018 2074 4022
rect 1970 3962 1973 4018
rect 2054 3962 2061 4018
rect 1718 3958 1738 3962
rect 1802 3958 1822 3962
rect 1886 3958 1906 3962
rect 1970 3958 1990 3962
rect 2054 3958 2074 3962
rect 2138 3958 2143 4022
rect 1485 3937 2143 3958
rect 1485 3881 1709 3937
rect 1765 3881 1797 3937
rect 1853 3881 1885 3937
rect 1941 3881 1973 3937
rect 2029 3881 2061 3937
rect 2117 3881 2143 3937
rect 1485 3863 2143 3881
tri 916 3811 936 3831 sw
rect 852 3805 936 3811
tri 936 3805 942 3811 sw
tri 852 3721 936 3805 ne
rect 936 3745 942 3805
tri 942 3745 1002 3805 sw
rect 936 2813 1002 3745
rect 936 2757 941 2813
rect 997 2757 1002 2813
rect 936 2733 1002 2757
rect 936 2677 941 2733
rect 997 2677 1002 2733
rect 936 2672 1002 2677
rect 1472 1653 2143 1663
rect 1472 1652 1789 1653
rect 1472 1596 1507 1652
rect 1563 1596 1590 1652
rect 1646 1597 1789 1652
rect 1845 1597 2143 1653
rect 1646 1596 2143 1597
rect 1472 1507 2143 1596
rect 1472 1506 1789 1507
rect 1472 1450 1507 1506
rect 1563 1450 1590 1506
rect 1646 1451 1789 1506
rect 1845 1451 2143 1507
rect 1646 1450 2143 1451
tri 1466 1409 1472 1415 se
rect 1472 1409 2143 1450
tri 1291 1234 1466 1409 se
rect 1466 1234 2143 1409
rect 283 330 441 335
rect 283 274 288 330
rect 344 298 441 330
rect 283 250 291 274
rect 283 194 288 250
rect 355 234 371 298
rect 435 234 441 298
rect 344 194 441 234
rect 283 189 441 194
rect 1291 256 2143 1234
rect 2225 1496 2699 9706
rect 2225 1432 2230 1496
rect 2294 1432 2310 1496
rect 2374 1432 2390 1496
rect 2454 1432 2470 1496
rect 2534 1432 2550 1496
rect 2614 1432 2630 1496
rect 2694 1432 2699 1496
rect 2225 1412 2699 1432
rect 2225 1348 2230 1412
rect 2294 1348 2310 1412
rect 2374 1348 2390 1412
rect 2454 1348 2470 1412
rect 2534 1348 2550 1412
rect 2614 1348 2630 1412
rect 2694 1348 2699 1412
rect 2225 1328 2699 1348
rect 2225 1264 2230 1328
rect 2294 1264 2310 1328
rect 2374 1264 2390 1328
rect 2454 1264 2470 1328
rect 2534 1264 2550 1328
rect 2614 1264 2630 1328
rect 2694 1264 2699 1328
rect 2225 1244 2699 1264
rect 2225 1180 2230 1244
rect 2294 1180 2310 1244
rect 2374 1180 2390 1244
rect 2454 1180 2470 1244
rect 2534 1180 2550 1244
rect 2614 1180 2630 1244
rect 2694 1180 2699 1244
rect 2225 1160 2699 1180
rect 2225 1096 2230 1160
rect 2294 1096 2310 1160
rect 2374 1096 2390 1160
rect 2454 1096 2470 1160
rect 2534 1096 2550 1160
rect 2614 1096 2630 1160
rect 2694 1096 2699 1160
rect 2225 1076 2699 1096
rect 2225 1012 2230 1076
rect 2294 1012 2310 1076
rect 2374 1012 2390 1076
rect 2454 1012 2470 1076
rect 2534 1012 2550 1076
rect 2614 1012 2630 1076
rect 2694 1012 2699 1076
rect 2225 992 2699 1012
rect 2225 928 2230 992
rect 2294 928 2310 992
rect 2374 928 2390 992
rect 2454 928 2470 992
rect 2534 928 2550 992
rect 2614 928 2630 992
rect 2694 928 2699 992
rect 2225 908 2699 928
rect 2225 844 2230 908
rect 2294 844 2310 908
rect 2374 844 2390 908
rect 2454 844 2470 908
rect 2534 844 2550 908
rect 2614 844 2630 908
rect 2694 844 2699 908
rect 2225 823 2699 844
rect 2225 759 2230 823
rect 2294 759 2310 823
rect 2374 759 2390 823
rect 2454 759 2470 823
rect 2534 759 2550 823
rect 2614 759 2630 823
rect 2694 759 2699 823
rect 2225 738 2699 759
rect 2225 674 2230 738
rect 2294 674 2310 738
rect 2374 674 2390 738
rect 2454 674 2470 738
rect 2534 674 2550 738
rect 2614 674 2630 738
rect 2694 674 2699 738
rect 2225 653 2699 674
rect 2225 589 2230 653
rect 2294 589 2310 653
rect 2374 589 2390 653
rect 2454 589 2470 653
rect 2534 589 2550 653
rect 2614 589 2630 653
rect 2694 589 2699 653
rect 2781 9260 3778 10262
rect 2781 9246 2789 9260
rect 2845 9246 2921 9260
rect 2977 9246 3053 9260
rect 3109 9246 3185 9260
rect 3241 9246 3317 9260
rect 3373 9246 3449 9260
rect 3505 9246 3581 9260
rect 3637 9246 3713 9260
rect 3769 9246 3778 9260
rect 2781 9182 2782 9246
rect 2846 9182 2866 9246
rect 2930 9182 2950 9204
rect 3014 9182 3034 9246
rect 3109 9204 3118 9246
rect 3098 9182 3118 9204
rect 3182 9204 3185 9246
rect 3182 9182 3202 9204
rect 3266 9182 3286 9246
rect 3434 9204 3449 9246
rect 3350 9182 3370 9204
rect 3434 9182 3454 9204
rect 3518 9182 3538 9246
rect 3602 9182 3622 9204
rect 3686 9182 3706 9246
rect 3770 9182 3778 9246
rect 2781 9160 3778 9182
rect 2781 9096 2782 9160
rect 2846 9096 2866 9160
rect 2930 9120 2950 9160
rect 3014 9096 3034 9160
rect 3098 9120 3118 9160
rect 3109 9096 3118 9120
rect 3182 9120 3202 9160
rect 3182 9096 3185 9120
rect 3266 9096 3286 9160
rect 3350 9120 3370 9160
rect 3434 9120 3454 9160
rect 3434 9096 3449 9120
rect 3518 9096 3538 9160
rect 3602 9120 3622 9160
rect 3686 9096 3706 9160
rect 3770 9096 3778 9160
rect 2781 9074 2789 9096
rect 2845 9074 2921 9096
rect 2977 9074 3053 9096
rect 3109 9074 3185 9096
rect 3241 9074 3317 9096
rect 3373 9074 3449 9096
rect 3505 9074 3581 9096
rect 3637 9074 3713 9096
rect 3769 9074 3778 9096
rect 2781 9010 2782 9074
rect 2846 9010 2866 9074
rect 2930 9010 2950 9064
rect 3014 9010 3034 9074
rect 3109 9064 3118 9074
rect 3098 9010 3118 9064
rect 3182 9064 3185 9074
rect 3182 9010 3202 9064
rect 3266 9010 3286 9074
rect 3434 9064 3449 9074
rect 3350 9010 3370 9064
rect 3434 9010 3454 9064
rect 3518 9010 3538 9074
rect 3602 9010 3622 9064
rect 3686 9010 3706 9074
rect 3770 9010 3778 9074
rect 2781 8988 3778 9010
rect 2781 8924 2782 8988
rect 2846 8924 2866 8988
rect 2930 8924 2950 8988
rect 3014 8924 3034 8988
rect 3098 8924 3118 8988
rect 3182 8924 3202 8988
rect 3266 8924 3286 8988
rect 3350 8924 3370 8988
rect 3434 8924 3454 8988
rect 3518 8924 3538 8988
rect 3602 8924 3622 8988
rect 3686 8924 3706 8988
rect 3770 8924 3778 8988
rect 2781 8902 3778 8924
rect 2781 8838 2782 8902
rect 2846 8838 2866 8902
rect 2930 8838 2950 8902
rect 3014 8838 3034 8902
rect 3098 8838 3118 8902
rect 3182 8838 3202 8902
rect 3266 8838 3286 8902
rect 3350 8838 3370 8902
rect 3434 8838 3454 8902
rect 3518 8838 3538 8902
rect 3602 8838 3622 8902
rect 3686 8838 3706 8902
rect 3770 8838 3778 8902
rect 2781 8816 3778 8838
rect 2781 8752 2782 8816
rect 2846 8752 2866 8816
rect 2930 8752 2950 8816
rect 3014 8752 3034 8816
rect 3098 8752 3118 8816
rect 3182 8752 3202 8816
rect 3266 8752 3286 8816
rect 3350 8752 3370 8816
rect 3434 8752 3454 8816
rect 3518 8752 3538 8816
rect 3602 8752 3622 8816
rect 3686 8752 3706 8816
rect 3770 8752 3778 8816
rect 2781 8730 3778 8752
rect 2781 8666 2782 8730
rect 2846 8666 2866 8730
rect 2930 8666 2950 8730
rect 3014 8666 3034 8730
rect 3098 8666 3118 8730
rect 3182 8666 3202 8730
rect 3266 8666 3286 8730
rect 3350 8666 3370 8730
rect 3434 8666 3454 8730
rect 3518 8666 3538 8730
rect 3602 8666 3622 8730
rect 3686 8666 3706 8730
rect 3770 8666 3778 8730
rect 2781 8643 3778 8666
rect 2781 8579 2782 8643
rect 2846 8579 2866 8643
rect 2930 8579 2950 8643
rect 3014 8579 3034 8643
rect 3098 8579 3118 8643
rect 3182 8579 3202 8643
rect 3266 8579 3286 8643
rect 3350 8579 3370 8643
rect 3434 8579 3454 8643
rect 3518 8579 3538 8643
rect 3602 8579 3622 8643
rect 3686 8579 3706 8643
rect 3770 8579 3778 8643
rect 2781 8556 3778 8579
rect 2781 8492 2782 8556
rect 2846 8492 2866 8556
rect 2930 8492 2950 8556
rect 3014 8492 3034 8556
rect 3098 8492 3118 8556
rect 3182 8492 3202 8556
rect 3266 8492 3286 8556
rect 3350 8492 3370 8556
rect 3434 8492 3454 8556
rect 3518 8492 3538 8556
rect 3602 8492 3622 8556
rect 3686 8492 3706 8556
rect 3770 8492 3778 8556
rect 2781 8469 3778 8492
rect 2781 8405 2782 8469
rect 2846 8405 2866 8469
rect 2930 8405 2950 8469
rect 3014 8405 3034 8469
rect 3098 8405 3118 8469
rect 3182 8405 3202 8469
rect 3266 8405 3286 8469
rect 3350 8405 3370 8469
rect 3434 8405 3454 8469
rect 3518 8405 3538 8469
rect 3602 8405 3622 8469
rect 3686 8405 3706 8469
rect 3770 8405 3778 8469
rect 2781 8382 3778 8405
rect 2781 8318 2782 8382
rect 2846 8318 2866 8382
rect 2930 8318 2950 8382
rect 3014 8318 3034 8382
rect 3098 8318 3118 8382
rect 3182 8318 3202 8382
rect 3266 8318 3286 8382
rect 3350 8318 3370 8382
rect 3434 8318 3454 8382
rect 3518 8318 3538 8382
rect 3602 8318 3622 8382
rect 3686 8318 3706 8382
rect 3770 8318 3778 8382
rect 2781 8232 3778 8318
rect 2781 8176 2850 8232
rect 2906 8176 2974 8232
rect 3030 8176 3098 8232
rect 3154 8176 3221 8232
rect 3277 8176 3344 8232
rect 3400 8176 3467 8232
rect 3523 8176 3590 8232
rect 3646 8176 3713 8232
rect 3769 8176 3778 8232
rect 2781 3150 3778 8176
rect 3858 7884 4178 14686
rect 4287 14332 4883 16125
rect 4991 14988 5991 18282
rect 8266 17283 9136 17289
rect 8266 17227 8454 17283
rect 8510 17227 8604 17283
rect 8660 17227 8754 17283
rect 8810 17227 8903 17283
rect 8959 17227 9052 17283
rect 9108 17227 9136 17283
rect 8266 17195 9136 17227
rect 8266 17139 8454 17195
rect 8510 17139 8604 17195
rect 8660 17139 8754 17195
rect 8810 17139 8903 17195
rect 8959 17139 9052 17195
rect 9108 17139 9136 17195
rect 8266 17107 9136 17139
rect 8266 17051 8454 17107
rect 8510 17051 8604 17107
rect 8660 17051 8754 17107
rect 8810 17051 8903 17107
rect 8959 17051 9052 17107
rect 9108 17051 9136 17107
rect 7036 16795 7182 16803
rect 7036 16739 7041 16795
rect 7097 16739 7121 16795
rect 7177 16739 7182 16795
tri 6915 15706 7036 15827 se
rect 7036 15706 7182 16739
tri 8213 16456 8266 16509 se
rect 8266 16456 9136 17051
tri 8208 16451 8213 16456 se
rect 8213 16451 9136 16456
tri 5991 14988 6251 15248 sw
rect 4991 14934 6251 14988
tri 6251 14934 6305 14988 sw
rect 4991 14892 6305 14934
tri 6305 14892 6347 14934 sw
rect 4991 14873 6347 14892
tri 4991 14604 5260 14873 ne
rect 5260 14604 6347 14873
tri 6347 14604 6635 14892 sw
tri 5260 14411 5453 14604 ne
rect 5453 14411 6635 14604
rect 6915 14578 7182 15706
tri 8156 16399 8208 16451 se
rect 8208 16399 8454 16451
rect 8156 16395 8454 16399
rect 8510 16395 8604 16451
rect 8660 16395 8754 16451
rect 8810 16395 8903 16451
rect 8959 16395 9052 16451
rect 9108 16395 9136 16451
rect 8156 16363 9136 16395
rect 8156 16307 8454 16363
rect 8510 16307 8604 16363
rect 8660 16307 8754 16363
rect 8810 16307 8903 16363
rect 8959 16307 9052 16363
rect 9108 16307 9136 16363
rect 8156 16275 9136 16307
rect 8156 16219 8454 16275
rect 8510 16219 8604 16275
rect 8660 16219 8754 16275
rect 8810 16219 8903 16275
rect 8959 16219 9052 16275
rect 9108 16219 9136 16275
rect 8156 15947 9136 16219
rect 8156 14988 8468 15947
tri 8468 15688 8727 15947 nw
tri 13561 15067 13738 15244 se
rect 13738 15094 13952 19840
rect 13738 15067 13925 15094
tri 13925 15067 13952 15094 nw
tri 12529 15024 12572 15067 se
rect 12572 15024 13711 15067
tri 8468 14988 8504 15024 sw
tri 12493 14988 12529 15024 se
rect 12529 14988 13711 15024
rect 8156 14934 8504 14988
tri 8504 14934 8558 14988 sw
tri 12439 14934 12493 14988 se
rect 12493 14934 13711 14988
rect 8156 14892 8558 14934
tri 8558 14892 8600 14934 sw
tri 12397 14892 12439 14934 se
rect 12439 14892 13711 14934
rect 8156 14780 8600 14892
tri 8600 14780 8712 14892 sw
tri 12342 14837 12397 14892 se
rect 12397 14853 13711 14892
tri 13711 14853 13925 15067 nw
rect 12397 14837 12792 14853
tri 12792 14837 12808 14853 nw
rect 12342 14780 12735 14837
tri 12735 14780 12792 14837 nw
rect 8156 14660 9484 14780
tri 9484 14660 9604 14780 sw
rect 12342 14660 12615 14780
tri 12615 14660 12735 14780 nw
rect 8156 14490 9604 14660
tri 4883 14332 4962 14411 sw
tri 5453 14332 5532 14411 ne
rect 5532 14332 6635 14411
rect 4287 14224 4962 14332
tri 4962 14224 5070 14332 sw
tri 5532 14224 5640 14332 ne
rect 4287 14129 5070 14224
tri 4287 13900 4516 14129 ne
rect 4516 13900 5070 14129
tri 5070 13900 5394 14224 sw
tri 4516 13844 4572 13900 ne
rect 4572 13844 5394 13900
tri 5394 13844 5450 13900 sw
tri 4572 13762 4654 13844 ne
rect 4654 13762 5450 13844
tri 5450 13762 5532 13844 sw
tri 4654 13533 4883 13762 ne
rect 4883 13533 5532 13762
tri 4883 13504 4912 13533 ne
rect 4264 8422 4446 11564
rect 4620 11528 4626 11533
rect 4620 11472 4625 11528
rect 4620 11469 4626 11472
rect 4690 11469 4706 11533
rect 4770 11528 4776 11533
rect 4771 11472 4776 11528
rect 4770 11469 4776 11472
rect 4620 11467 4776 11469
rect 4544 11282 4550 11346
rect 4614 11282 4634 11346
rect 4698 11282 4718 11346
rect 4782 11282 4788 11346
rect 4544 10563 4788 11282
rect 4544 10499 4550 10563
rect 4614 10499 4634 10563
rect 4698 10499 4718 10563
rect 4782 10499 4788 10563
rect 4544 10479 4788 10499
rect 4544 10415 4550 10479
rect 4614 10415 4634 10479
rect 4698 10415 4718 10479
rect 4782 10415 4788 10479
rect 4544 10395 4788 10415
rect 4544 10331 4550 10395
rect 4614 10331 4634 10395
rect 4698 10331 4718 10395
rect 4782 10331 4788 10395
rect 4544 9612 4788 10331
rect 4544 9548 4550 9612
rect 4614 9548 4634 9612
rect 4698 9548 4718 9612
rect 4782 9548 4788 9612
tri 4446 8422 4448 8424 sw
rect 4264 8390 4448 8422
tri 4448 8390 4480 8422 sw
rect 4264 8334 4480 8390
tri 4480 8334 4536 8390 sw
rect 4264 8313 4536 8334
tri 4536 8313 4557 8334 sw
rect 4264 8257 4557 8313
tri 4557 8257 4613 8313 sw
rect 4264 8235 4613 8257
tri 4613 8235 4635 8257 sw
rect 4264 8179 4635 8235
tri 4635 8179 4691 8235 sw
rect 4264 8127 4691 8179
tri 4691 8127 4743 8179 sw
rect 4264 8120 4743 8127
tri 4743 8120 4750 8127 sw
rect 4264 7989 4750 8120
rect 4264 7964 4332 7989
tri 4264 7940 4288 7964 ne
rect 4288 7940 4332 7964
tri 4288 7923 4305 7940 ne
rect 4305 7925 4332 7940
rect 4396 7925 4416 7989
rect 4480 7925 4499 7989
rect 4563 7925 4582 7989
rect 4646 7925 4665 7989
rect 4729 7925 4750 7989
rect 4305 7923 4750 7925
tri 4305 7906 4322 7923 ne
rect 4322 7906 4750 7923
tri 4178 7884 4200 7906 sw
tri 4322 7884 4344 7906 ne
rect 4344 7904 4750 7906
rect 4344 7884 4415 7904
rect 3858 7859 4200 7884
tri 4200 7859 4225 7884 sw
tri 4344 7859 4369 7884 ne
rect 4369 7859 4415 7884
rect 3858 7820 4225 7859
tri 4225 7820 4264 7859 sw
tri 4369 7838 4390 7859 ne
rect 4390 7840 4415 7859
rect 4479 7840 4499 7904
rect 4563 7840 4582 7904
rect 4646 7840 4665 7904
rect 4729 7840 4750 7904
rect 4390 7838 4750 7840
tri 4390 7820 4408 7838 ne
rect 4408 7820 4750 7838
rect 3858 7803 4264 7820
tri 4264 7803 4281 7820 sw
tri 4408 7803 4425 7820 ne
rect 4425 7818 4750 7820
rect 4425 7803 4496 7818
rect 3858 7778 4281 7803
tri 4281 7778 4306 7803 sw
tri 4425 7778 4450 7803 ne
rect 4450 7778 4496 7803
rect 3858 7772 4306 7778
tri 3858 7766 3864 7772 ne
rect 3864 7766 4306 7772
tri 4306 7766 4318 7778 sw
tri 4450 7766 4462 7778 ne
rect 4462 7766 4496 7778
tri 3864 7722 3908 7766 ne
rect 3908 7722 4318 7766
tri 4318 7722 4362 7766 sw
tri 4462 7752 4476 7766 ne
rect 4476 7754 4496 7766
rect 4560 7754 4581 7818
rect 4645 7754 4665 7818
rect 4729 7754 4750 7818
rect 4476 7752 4750 7754
tri 4476 7722 4506 7752 ne
rect 4506 7722 4750 7752
tri 3908 7697 3933 7722 ne
rect 3933 7700 4362 7722
tri 4362 7700 4384 7722 sw
tri 4506 7700 4528 7722 ne
rect 4528 7700 4750 7722
rect 3933 7697 4384 7700
tri 4384 7697 4387 7700 sw
tri 4528 7697 4531 7700 ne
rect 4531 7698 4750 7700
rect 4531 7697 4578 7698
tri 3933 7641 3989 7697 ne
rect 3989 7660 4387 7697
tri 4387 7660 4424 7697 sw
tri 4531 7660 4568 7697 ne
rect 3989 7641 4424 7660
tri 4424 7641 4443 7660 sw
tri 3989 7616 4014 7641 ne
rect 4014 7632 4443 7641
tri 4443 7632 4452 7641 sw
rect 4568 7634 4578 7697
rect 4642 7634 4665 7698
rect 4729 7634 4750 7698
rect 4014 7617 4452 7632
tri 4452 7617 4467 7632 sw
rect 4568 7617 4750 7634
rect 4014 7616 4467 7617
tri 4467 7616 4468 7617 sw
tri 4014 7560 4070 7616 ne
rect 4070 7560 4468 7616
tri 4468 7560 4524 7616 sw
tri 4070 7535 4095 7560 ne
rect 4095 7535 4524 7560
tri 4524 7535 4549 7560 sw
tri 4095 7479 4151 7535 ne
rect 4151 7479 4549 7535
tri 4549 7479 4605 7535 sw
tri 4151 7454 4176 7479 ne
rect 4176 7454 4605 7479
tri 4605 7454 4630 7479 sw
tri 4176 7452 4178 7454 ne
rect 4178 7452 4630 7454
tri 4178 7398 4232 7452 ne
rect 4232 7398 4630 7452
tri 4630 7398 4686 7454 sw
tri 4232 7373 4257 7398 ne
rect 4257 7373 4686 7398
tri 4686 7373 4711 7398 sw
tri 4257 7317 4313 7373 ne
rect 4313 7317 4711 7373
tri 4711 7317 4767 7373 sw
tri 4313 7312 4318 7317 ne
rect 4318 7312 4767 7317
tri 4767 7312 4772 7317 sw
tri 4318 7291 4339 7312 ne
rect 4339 7291 4772 7312
tri 4339 7235 4395 7291 ne
rect 4395 7235 4772 7291
tri 4395 7209 4421 7235 ne
rect 4421 7066 4772 7235
rect 4421 7002 4454 7066
rect 4518 7002 4538 7066
rect 4602 7002 4622 7066
rect 4686 7002 4706 7066
rect 4770 7002 4772 7066
rect 4421 6980 4772 7002
rect 4421 6916 4454 6980
rect 4518 6916 4538 6980
rect 4602 6916 4622 6980
rect 4686 6916 4706 6980
rect 4770 6916 4772 6980
rect 4421 6894 4772 6916
rect 4421 6830 4454 6894
rect 4518 6830 4538 6894
rect 4602 6830 4622 6894
rect 4686 6830 4706 6894
rect 4770 6830 4772 6894
rect 4421 6807 4772 6830
rect 4421 6743 4454 6807
rect 4518 6743 4538 6807
rect 4602 6743 4622 6807
rect 4686 6743 4706 6807
rect 4770 6743 4772 6807
rect 4421 6720 4772 6743
rect 4421 6656 4454 6720
rect 4518 6656 4538 6720
rect 4602 6656 4622 6720
rect 4686 6656 4706 6720
rect 4770 6656 4772 6720
rect 4421 6633 4772 6656
rect 4421 6569 4454 6633
rect 4518 6569 4538 6633
rect 4602 6569 4622 6633
rect 4686 6569 4706 6633
rect 4770 6569 4772 6633
rect 4421 6546 4772 6569
rect 4421 6482 4454 6546
rect 4518 6482 4538 6546
rect 4602 6482 4622 6546
rect 4686 6482 4706 6546
rect 4770 6482 4772 6546
rect 4421 6459 4772 6482
rect 4421 6395 4454 6459
rect 4518 6395 4538 6459
rect 4602 6395 4622 6459
rect 4686 6395 4706 6459
rect 4770 6395 4772 6459
rect 4421 6377 4772 6395
rect 4912 3676 5532 13533
rect 4912 3612 4918 3676
rect 4982 3612 5008 3676
rect 5072 3612 5098 3676
rect 5162 3612 5188 3676
rect 5252 3612 5278 3676
rect 5342 3612 5368 3676
rect 5432 3612 5458 3676
rect 5522 3612 5532 3676
rect 4912 3590 5532 3612
rect 4912 3526 4918 3590
rect 4982 3526 5008 3590
rect 5072 3526 5098 3590
rect 5162 3526 5188 3590
rect 5252 3526 5278 3590
rect 5342 3526 5368 3590
rect 5432 3526 5458 3590
rect 5522 3526 5532 3590
rect 4912 3503 5532 3526
rect 4912 3439 4918 3503
rect 4982 3439 5008 3503
rect 5072 3439 5098 3503
rect 5162 3439 5188 3503
rect 5252 3439 5278 3503
rect 5342 3439 5368 3503
rect 5432 3439 5458 3503
rect 5522 3439 5532 3503
rect 4912 3416 5532 3439
rect 4912 3352 4918 3416
rect 4982 3352 5008 3416
rect 5072 3352 5098 3416
rect 5162 3352 5188 3416
rect 5252 3352 5278 3416
rect 5342 3352 5368 3416
rect 5432 3352 5458 3416
rect 5522 3352 5532 3416
rect 4912 3329 5532 3352
tri 3778 3150 3912 3284 sw
rect 4912 3265 4918 3329
rect 4982 3265 5008 3329
rect 5072 3265 5098 3329
rect 5162 3265 5188 3329
rect 5252 3265 5278 3329
rect 5342 3265 5368 3329
rect 5432 3265 5458 3329
rect 5522 3265 5532 3329
rect 4912 3242 5532 3265
rect 4912 3178 4918 3242
rect 4982 3178 5008 3242
rect 5072 3178 5098 3242
rect 5162 3178 5188 3242
rect 5252 3178 5278 3242
rect 5342 3178 5368 3242
rect 5432 3178 5458 3242
rect 5522 3178 5532 3242
rect 4912 3155 5532 3178
rect 2781 3145 3912 3150
tri 3912 3145 3917 3150 sw
rect 2781 3089 3917 3145
tri 3917 3089 3973 3145 sw
rect 4912 3091 4918 3155
rect 4982 3091 5008 3155
rect 5072 3091 5098 3155
rect 5162 3091 5188 3155
rect 5252 3091 5278 3155
rect 5342 3091 5368 3155
rect 5432 3091 5458 3155
rect 5522 3091 5532 3155
rect 2781 3023 3973 3089
tri 3973 3023 4039 3089 sw
rect 4912 3068 5532 3091
rect 2781 3022 4039 3023
tri 4039 3022 4040 3023 sw
rect 2781 2966 4040 3022
tri 4040 2966 4096 3022 sw
rect 4912 3004 4918 3068
rect 4982 3004 5008 3068
rect 5072 3004 5098 3068
rect 5162 3004 5188 3068
rect 5252 3004 5278 3068
rect 5342 3004 5368 3068
rect 5432 3004 5458 3068
rect 5522 3004 5532 3068
rect 4912 2988 5532 3004
rect 5640 13698 6635 14332
tri 9364 14250 9604 14490 ne
tri 9604 14250 10014 14660 sw
tri 9604 14130 9724 14250 ne
rect 5640 13634 5648 13698
rect 5712 13634 5731 13698
rect 5795 13634 5814 13698
rect 5878 13634 5897 13698
rect 5961 13634 5980 13698
rect 6044 13634 6063 13698
rect 6127 13634 6146 13698
rect 6210 13634 6229 13698
rect 6293 13634 6312 13698
rect 6376 13634 6395 13698
rect 6459 13634 6478 13698
rect 6542 13634 6561 13698
rect 6625 13634 6635 13698
rect 5640 13618 6635 13634
rect 5640 13554 5648 13618
rect 5712 13554 5731 13618
rect 5795 13554 5814 13618
rect 5878 13554 5897 13618
rect 5961 13554 5980 13618
rect 6044 13554 6063 13618
rect 6127 13554 6146 13618
rect 6210 13554 6229 13618
rect 6293 13554 6312 13618
rect 6376 13554 6395 13618
rect 6459 13554 6478 13618
rect 6542 13554 6561 13618
rect 6625 13554 6635 13618
rect 5640 13538 6635 13554
rect 5640 13474 5648 13538
rect 5712 13474 5731 13538
rect 5795 13474 5814 13538
rect 5878 13474 5897 13538
rect 5961 13474 5980 13538
rect 6044 13474 6063 13538
rect 6127 13474 6146 13538
rect 6210 13474 6229 13538
rect 6293 13474 6312 13538
rect 6376 13474 6395 13538
rect 6459 13474 6478 13538
rect 6542 13474 6561 13538
rect 6625 13474 6635 13538
rect 5640 13458 6635 13474
rect 5640 13394 5648 13458
rect 5712 13394 5731 13458
rect 5795 13394 5814 13458
rect 5878 13394 5897 13458
rect 5961 13394 5980 13458
rect 6044 13394 6063 13458
rect 6127 13394 6146 13458
rect 6210 13394 6229 13458
rect 6293 13394 6312 13458
rect 6376 13394 6395 13458
rect 6459 13394 6478 13458
rect 6542 13394 6561 13458
rect 6625 13394 6635 13458
rect 5640 13378 6635 13394
rect 5640 13314 5648 13378
rect 5712 13314 5731 13378
rect 5795 13314 5814 13378
rect 5878 13314 5897 13378
rect 5961 13314 5980 13378
rect 6044 13314 6063 13378
rect 6127 13314 6146 13378
rect 6210 13314 6229 13378
rect 6293 13314 6312 13378
rect 6376 13314 6395 13378
rect 6459 13314 6478 13378
rect 6542 13314 6561 13378
rect 6625 13314 6635 13378
rect 5640 13298 6635 13314
rect 5640 13234 5648 13298
rect 5712 13234 5731 13298
rect 5795 13234 5814 13298
rect 5878 13234 5897 13298
rect 5961 13234 5980 13298
rect 6044 13234 6063 13298
rect 6127 13234 6146 13298
rect 6210 13234 6229 13298
rect 6293 13234 6312 13298
rect 6376 13234 6395 13298
rect 6459 13234 6478 13298
rect 6542 13234 6561 13298
rect 6625 13234 6635 13298
rect 5640 13218 6635 13234
rect 5640 13154 5648 13218
rect 5712 13154 5731 13218
rect 5795 13154 5814 13218
rect 5878 13154 5897 13218
rect 5961 13154 5980 13218
rect 6044 13154 6063 13218
rect 6127 13154 6146 13218
rect 6210 13154 6229 13218
rect 6293 13154 6312 13218
rect 6376 13154 6395 13218
rect 6459 13154 6478 13218
rect 6542 13154 6561 13218
rect 6625 13154 6635 13218
rect 5640 13138 6635 13154
rect 5640 13074 5648 13138
rect 5712 13074 5731 13138
rect 5795 13074 5814 13138
rect 5878 13074 5897 13138
rect 5961 13074 5980 13138
rect 6044 13074 6063 13138
rect 6127 13074 6146 13138
rect 6210 13074 6229 13138
rect 6293 13074 6312 13138
rect 6376 13074 6395 13138
rect 6459 13074 6478 13138
rect 6542 13074 6561 13138
rect 6625 13074 6635 13138
rect 5640 13058 6635 13074
rect 5640 12994 5648 13058
rect 5712 12994 5731 13058
rect 5795 12994 5814 13058
rect 5878 12994 5897 13058
rect 5961 12994 5980 13058
rect 6044 12994 6063 13058
rect 6127 12994 6146 13058
rect 6210 12994 6229 13058
rect 6293 12994 6312 13058
rect 6376 12994 6395 13058
rect 6459 12994 6478 13058
rect 6542 12994 6561 13058
rect 6625 12994 6635 13058
rect 5640 12978 6635 12994
rect 5640 12914 5648 12978
rect 5712 12914 5731 12978
rect 5795 12914 5814 12978
rect 5878 12914 5897 12978
rect 5961 12914 5980 12978
rect 6044 12914 6063 12978
rect 6127 12914 6146 12978
rect 6210 12914 6229 12978
rect 6293 12914 6312 12978
rect 6376 12914 6395 12978
rect 6459 12914 6478 12978
rect 6542 12914 6561 12978
rect 6625 12914 6635 12978
rect 5640 12898 6635 12914
rect 5640 12834 5648 12898
rect 5712 12834 5731 12898
rect 5795 12834 5814 12898
rect 5878 12834 5897 12898
rect 5961 12834 5980 12898
rect 6044 12834 6063 12898
rect 6127 12834 6146 12898
rect 6210 12834 6229 12898
rect 6293 12834 6312 12898
rect 6376 12834 6395 12898
rect 6459 12834 6478 12898
rect 6542 12834 6561 12898
rect 6625 12834 6635 12898
rect 5640 11721 6635 12834
rect 5640 11373 6619 11721
tri 6619 11705 6635 11721 nw
rect 6699 11586 6855 11591
rect 6699 11530 6704 11586
rect 6760 11533 6855 11586
rect 6699 11506 6705 11530
rect 6699 11450 6704 11506
rect 6769 11469 6785 11533
rect 6849 11469 6855 11533
rect 6760 11450 6855 11469
rect 6699 11445 6855 11450
tri 6619 11373 6635 11389 sw
rect 2781 2901 4096 2966
tri 4096 2901 4161 2966 sw
rect 2781 2899 4161 2901
tri 4161 2899 4163 2901 sw
rect 2781 2843 4163 2899
tri 4163 2843 4219 2899 sw
rect 2781 2779 4219 2843
tri 4219 2779 4283 2843 sw
tri 5596 2779 5640 2823 se
rect 5640 2779 6635 11373
rect 6915 9238 7182 13498
rect 9341 13077 9407 13082
rect 9341 13021 9346 13077
rect 9402 13021 9407 13077
rect 9341 12997 9407 13021
rect 9341 12941 9346 12997
rect 9402 12941 9407 12997
rect 8018 11840 8084 11845
rect 8018 11784 8023 11840
rect 8079 11784 8084 11840
rect 8018 11760 8084 11784
rect 8018 11704 8023 11760
rect 8079 11704 8084 11760
tri 7924 11608 8018 11702 se
rect 8018 11674 8084 11704
tri 8018 11608 8084 11674 nw
tri 7867 11551 7924 11608 se
rect 7924 11551 7961 11608
tri 7961 11551 8018 11608 nw
rect 7867 10030 7933 11551
tri 7933 11523 7961 11551 nw
rect 9341 11526 9407 12941
rect 9470 13080 9536 13085
rect 9470 13024 9475 13080
rect 9531 13024 9536 13080
rect 9470 13000 9536 13024
rect 9470 12944 9475 13000
rect 9531 12944 9536 13000
rect 9470 11594 9536 12944
rect 9724 12066 10014 14250
rect 11001 13900 11287 13939
rect 11001 13844 11011 13900
rect 11067 13844 11111 13900
rect 11167 13844 11211 13900
rect 11267 13844 11287 13900
tri 9724 11885 9905 12066 ne
rect 9905 11885 10014 12066
tri 10014 11885 10315 12186 sw
tri 9905 11776 10014 11885 ne
rect 10014 11776 10315 11885
tri 10014 11765 10025 11776 ne
tri 9470 11554 9510 11594 ne
rect 9510 11554 9536 11594
tri 9536 11554 9604 11622 sw
tri 9407 11526 9435 11554 sw
tri 9510 11541 9523 11554 ne
rect 9523 11541 9604 11554
tri 9604 11541 9617 11554 sw
tri 9523 11528 9536 11541 ne
rect 9536 11528 9617 11541
tri 9536 11526 9538 11528 ne
rect 9538 11526 9617 11528
tri 9617 11526 9632 11541 sw
tri 9341 11523 9344 11526 ne
rect 9344 11523 9435 11526
tri 9344 11432 9435 11523 ne
tri 9435 11432 9529 11526 sw
tri 9538 11447 9617 11526 ne
rect 9617 11447 9632 11526
tri 9632 11447 9711 11526 sw
tri 9617 11432 9632 11447 ne
rect 9632 11432 9711 11447
tri 9711 11432 9726 11447 sw
tri 9435 11346 9521 11432 ne
rect 9521 11353 9529 11432
tri 9529 11353 9608 11432 sw
tri 9632 11353 9711 11432 ne
rect 9711 11353 9726 11432
tri 9726 11353 9805 11432 sw
rect 9521 11346 9608 11353
rect 7867 9974 7872 10030
rect 7928 9974 7933 10030
rect 7867 9950 7933 9974
rect 7867 9894 7872 9950
rect 7928 9894 7933 9950
rect 7867 9889 7933 9894
rect 8165 11282 8171 11346
rect 8235 11282 8255 11346
rect 8319 11282 8339 11346
rect 8403 11282 8409 11346
rect 8165 10563 8409 11282
rect 9180 11282 9186 11346
rect 9250 11282 9270 11346
rect 9334 11282 9354 11346
rect 9418 11282 9424 11346
tri 9521 11338 9529 11346 ne
rect 9529 11338 9608 11346
tri 9608 11338 9623 11353 sw
tri 9711 11338 9726 11353 ne
rect 9726 11338 9805 11353
tri 9805 11338 9820 11353 sw
rect 8165 10499 8171 10563
rect 8235 10499 8255 10563
rect 8319 10499 8339 10563
rect 8403 10499 8409 10563
rect 8165 10479 8409 10499
rect 8165 10415 8171 10479
rect 8235 10415 8255 10479
rect 8319 10415 8339 10479
rect 8403 10415 8409 10479
rect 8165 10395 8409 10415
rect 8165 10331 8171 10395
rect 8235 10331 8255 10395
rect 8319 10331 8339 10395
rect 8403 10331 8409 10395
rect 8165 9612 8409 10331
rect 8165 9548 8171 9612
rect 8235 9548 8255 9612
rect 8319 9548 8339 9612
rect 8403 9548 8409 9612
rect 6915 9174 6916 9238
rect 6980 9174 7014 9238
rect 7078 9174 7112 9238
rect 7176 9174 7182 9238
rect 6915 9153 7182 9174
rect 6915 9089 6916 9153
rect 6980 9089 7014 9153
rect 7078 9089 7112 9153
rect 7176 9089 7182 9153
rect 6915 9068 7182 9089
rect 6915 9004 6916 9068
rect 6980 9004 7014 9068
rect 7078 9004 7112 9068
rect 7176 9004 7182 9068
rect 6915 8983 7182 9004
rect 6915 8919 6916 8983
rect 6980 8919 7014 8983
rect 7078 8919 7112 8983
rect 7176 8919 7182 8983
rect 6915 8898 7182 8919
rect 6915 8834 6916 8898
rect 6980 8834 7014 8898
rect 7078 8834 7112 8898
rect 7176 8834 7182 8898
rect 6915 8813 7182 8834
rect 6915 8749 6916 8813
rect 6980 8749 7014 8813
rect 7078 8749 7112 8813
rect 7176 8749 7182 8813
rect 6915 8728 7182 8749
rect 6915 8664 6916 8728
rect 6980 8664 7014 8728
rect 7078 8664 7112 8728
rect 7176 8664 7182 8728
rect 6915 8643 7182 8664
rect 6915 8579 6916 8643
rect 6980 8579 7014 8643
rect 7078 8579 7112 8643
rect 7176 8579 7182 8643
rect 6915 8558 7182 8579
rect 6915 8494 6916 8558
rect 6980 8494 7014 8558
rect 7078 8494 7112 8558
rect 7176 8494 7182 8558
rect 6915 8472 7182 8494
rect 6915 8408 6916 8472
rect 6980 8408 7014 8472
rect 7078 8408 7112 8472
rect 7176 8408 7182 8472
rect 6915 8386 7182 8408
rect 6915 8322 6916 8386
rect 6980 8322 7014 8386
rect 7078 8322 7112 8386
rect 7176 8322 7182 8386
rect 6915 8315 7182 8322
rect 8595 9241 8862 11188
rect 9180 10563 9424 11282
tri 9529 11244 9623 11338 ne
tri 9623 11284 9677 11338 sw
tri 9726 11284 9780 11338 ne
rect 9780 11284 9820 11338
tri 9820 11284 9874 11338 sw
rect 9623 11259 9677 11284
tri 9677 11259 9702 11284 sw
tri 9780 11259 9805 11284 ne
rect 9805 11259 9874 11284
tri 9874 11259 9899 11284 sw
rect 9623 11244 9702 11259
tri 9702 11244 9717 11259 sw
tri 9805 11244 9820 11259 ne
rect 9820 11244 9899 11259
tri 9623 11190 9677 11244 ne
rect 9677 11218 9717 11244
tri 9717 11218 9743 11244 sw
tri 9820 11231 9833 11244 ne
rect 9180 10499 9186 10563
rect 9250 10499 9270 10563
rect 9334 10499 9354 10563
rect 9418 10499 9424 10563
rect 9180 10479 9424 10499
rect 9180 10415 9186 10479
rect 9250 10415 9270 10479
rect 9334 10415 9354 10479
rect 9418 10415 9424 10479
rect 9180 10395 9424 10415
rect 9180 10331 9186 10395
rect 9250 10331 9270 10395
rect 9334 10331 9354 10395
rect 9418 10331 9424 10395
rect 9180 9612 9424 10331
rect 9677 9988 9743 11218
rect 9677 9932 9682 9988
rect 9738 9932 9743 9988
rect 9677 9908 9743 9932
rect 9677 9852 9682 9908
rect 9738 9852 9743 9908
rect 9677 9847 9743 9852
rect 9180 9548 9186 9612
rect 9250 9548 9270 9612
rect 9334 9548 9354 9612
rect 9418 9548 9424 9612
rect 8595 9177 8601 9241
rect 8665 9177 8699 9241
rect 8763 9177 8797 9241
rect 8861 9177 8862 9241
rect 8595 9156 8862 9177
rect 8595 9092 8601 9156
rect 8665 9092 8699 9156
rect 8763 9092 8797 9156
rect 8861 9092 8862 9156
rect 8595 9070 8862 9092
rect 8595 9006 8601 9070
rect 8665 9006 8699 9070
rect 8763 9006 8797 9070
rect 8861 9006 8862 9070
rect 8595 8984 8862 9006
rect 8595 8920 8601 8984
rect 8665 8920 8699 8984
rect 8763 8920 8797 8984
rect 8861 8920 8862 8984
rect 8595 8898 8862 8920
rect 8595 8834 8601 8898
rect 8665 8834 8699 8898
rect 8763 8834 8797 8898
rect 8861 8834 8862 8898
rect 8595 8812 8862 8834
rect 8595 8748 8601 8812
rect 8665 8748 8699 8812
rect 8763 8748 8797 8812
rect 8861 8748 8862 8812
rect 8595 8726 8862 8748
rect 8595 8662 8601 8726
rect 8665 8662 8699 8726
rect 8763 8662 8797 8726
rect 8861 8662 8862 8726
rect 8595 8640 8862 8662
rect 8595 8576 8601 8640
rect 8665 8576 8699 8640
rect 8763 8576 8797 8640
rect 8861 8576 8862 8640
rect 8595 8554 8862 8576
rect 8595 8490 8601 8554
rect 8665 8490 8699 8554
rect 8763 8490 8797 8554
rect 8861 8490 8862 8554
rect 8595 8468 8862 8490
rect 8595 8404 8601 8468
rect 8665 8404 8699 8468
rect 8763 8404 8797 8468
rect 8861 8404 8862 8468
rect 8595 8382 8862 8404
rect 8595 8318 8601 8382
rect 8665 8318 8699 8382
rect 8763 8318 8797 8382
rect 8861 8318 8862 8382
rect 8595 8312 8862 8318
rect 9106 9265 9687 9445
rect 9106 9241 9121 9265
rect 9177 9241 9217 9265
rect 9273 9241 9313 9265
rect 9369 9241 9409 9265
rect 9465 9241 9505 9265
rect 9561 9241 9687 9265
rect 9106 9177 9114 9241
rect 9178 9177 9198 9241
rect 9273 9209 9282 9241
rect 9262 9178 9282 9209
rect 9346 9178 9366 9209
rect 9430 9178 9450 9209
rect 9514 9178 9534 9209
rect 9273 9177 9282 9178
rect 9598 9177 9618 9241
rect 9682 9177 9687 9241
rect 9106 9156 9121 9177
rect 9177 9156 9217 9177
rect 9273 9156 9313 9177
rect 9369 9156 9409 9177
rect 9465 9156 9505 9177
rect 9561 9156 9687 9177
rect 9106 9092 9114 9156
rect 9178 9092 9198 9156
rect 9273 9122 9282 9156
rect 9262 9092 9282 9122
rect 9346 9092 9366 9122
rect 9430 9092 9450 9122
rect 9514 9092 9534 9122
rect 9598 9092 9618 9156
rect 9682 9092 9687 9156
rect 9106 9091 9687 9092
rect 9106 9071 9121 9091
rect 9177 9071 9217 9091
rect 9273 9071 9313 9091
rect 9369 9071 9409 9091
rect 9465 9071 9505 9091
rect 9561 9071 9687 9091
rect 9106 9007 9114 9071
rect 9178 9007 9198 9071
rect 9273 9035 9282 9071
rect 9262 9007 9282 9035
rect 9346 9007 9366 9035
rect 9430 9007 9450 9035
rect 9514 9007 9534 9035
rect 9598 9007 9618 9071
rect 9682 9007 9687 9071
rect 9106 9004 9687 9007
rect 9106 8986 9121 9004
rect 9177 8986 9217 9004
rect 9273 8986 9313 9004
rect 9369 8986 9409 9004
rect 9465 8986 9505 9004
rect 9561 8986 9687 9004
rect 9106 8922 9114 8986
rect 9178 8922 9198 8986
rect 9273 8948 9282 8986
rect 9262 8922 9282 8948
rect 9346 8922 9366 8948
rect 9430 8922 9450 8948
rect 9514 8922 9534 8948
rect 9598 8922 9618 8986
rect 9682 8922 9687 8986
rect 9106 8917 9687 8922
rect 9106 8901 9121 8917
rect 9177 8901 9217 8917
rect 9273 8901 9313 8917
rect 9369 8901 9409 8917
rect 9465 8901 9505 8917
rect 9561 8901 9687 8917
rect 9106 8837 9114 8901
rect 9178 8837 9198 8901
rect 9273 8861 9282 8901
rect 9262 8837 9282 8861
rect 9346 8837 9366 8861
rect 9430 8837 9450 8861
rect 9514 8837 9534 8861
rect 9598 8837 9618 8901
rect 9682 8837 9687 8901
rect 9106 8830 9687 8837
rect 9106 8816 9121 8830
rect 9177 8816 9217 8830
rect 9273 8816 9313 8830
rect 9369 8816 9409 8830
rect 9465 8816 9505 8830
rect 9561 8816 9687 8830
rect 9106 8752 9114 8816
rect 9178 8752 9198 8816
rect 9273 8774 9282 8816
rect 9262 8752 9282 8774
rect 9346 8752 9366 8774
rect 9430 8752 9450 8774
rect 9514 8752 9534 8774
rect 9598 8752 9618 8816
rect 9682 8752 9687 8816
rect 9106 8742 9687 8752
rect 9106 8731 9121 8742
rect 9177 8731 9217 8742
rect 9273 8731 9313 8742
rect 9369 8731 9409 8742
rect 9465 8731 9505 8742
rect 9561 8731 9687 8742
rect 9106 8667 9114 8731
rect 9178 8667 9198 8731
rect 9273 8686 9282 8731
rect 9262 8667 9282 8686
rect 9346 8667 9366 8686
rect 9430 8667 9450 8686
rect 9514 8667 9534 8686
rect 9598 8667 9618 8731
rect 9682 8667 9687 8731
rect 9106 8654 9687 8667
rect 9106 8645 9121 8654
rect 9177 8645 9217 8654
rect 9273 8645 9313 8654
rect 9369 8645 9409 8654
rect 9465 8645 9505 8654
rect 9561 8645 9687 8654
rect 9106 8581 9114 8645
rect 9178 8581 9198 8645
rect 9273 8598 9282 8645
rect 9262 8581 9282 8598
rect 9346 8581 9366 8598
rect 9430 8581 9450 8598
rect 9514 8581 9534 8598
rect 9598 8581 9618 8645
rect 9682 8581 9687 8645
rect 9106 8566 9687 8581
rect 9106 8559 9121 8566
rect 9177 8559 9217 8566
rect 9273 8559 9313 8566
rect 9369 8559 9409 8566
rect 9465 8559 9505 8566
rect 9561 8559 9687 8566
rect 9106 8495 9114 8559
rect 9178 8495 9198 8559
rect 9273 8510 9282 8559
rect 9262 8495 9282 8510
rect 9346 8495 9366 8510
rect 9430 8495 9450 8510
rect 9514 8495 9534 8510
rect 9598 8495 9618 8559
rect 9682 8495 9687 8559
rect 9106 8478 9687 8495
rect 9106 8473 9121 8478
rect 9177 8473 9217 8478
rect 9273 8473 9313 8478
rect 9369 8473 9409 8478
rect 9465 8473 9505 8478
rect 9561 8473 9687 8478
rect 9106 8409 9114 8473
rect 9178 8409 9198 8473
rect 9273 8422 9282 8473
rect 9262 8409 9282 8422
rect 9346 8409 9366 8422
rect 9430 8409 9450 8422
rect 9514 8409 9534 8422
rect 9598 8409 9618 8473
rect 9682 8409 9687 8473
rect 9106 8390 9687 8409
rect 9106 8387 9121 8390
rect 9177 8387 9217 8390
rect 9273 8387 9313 8390
rect 9369 8387 9409 8390
rect 9465 8387 9505 8390
rect 9561 8387 9687 8390
rect 9106 8323 9114 8387
rect 9178 8323 9198 8387
rect 9273 8334 9282 8387
rect 9262 8323 9282 8334
rect 9346 8323 9366 8334
rect 9430 8323 9450 8334
rect 9514 8323 9534 8334
rect 9598 8323 9618 8387
rect 9682 8323 9687 8387
rect 9106 8134 9687 8323
tri 9266 7454 9280 7468 se
rect 9280 7454 9609 7468
tri 9609 7454 9623 7468 sw
tri 9210 7398 9266 7454 se
rect 9266 7402 9623 7454
rect 9266 7398 9304 7402
tri 9304 7398 9308 7402 nw
tri 9581 7398 9585 7402 ne
rect 9585 7398 9623 7402
tri 9623 7398 9679 7454 sw
tri 9187 7375 9210 7398 se
rect 9210 7375 9281 7398
tri 9281 7375 9304 7398 nw
tri 9585 7375 9608 7398 ne
rect 9608 7375 9679 7398
tri 9679 7375 9702 7398 sw
tri 9186 7374 9187 7375 se
rect 9187 7374 9280 7375
tri 9280 7374 9281 7375 nw
tri 9608 7374 9609 7375 ne
rect 9609 7374 9702 7375
tri 9185 7373 9186 7374 se
rect 9186 7373 9279 7374
tri 9279 7373 9280 7374 nw
tri 9609 7373 9610 7374 ne
rect 9610 7373 9702 7374
tri 9173 7361 9185 7373 se
rect 9185 7361 9267 7373
tri 9267 7361 9279 7373 nw
tri 9610 7361 9622 7373 ne
rect 9622 7361 9702 7373
rect 2781 2776 4283 2779
tri 4283 2776 4286 2779 sw
tri 5593 2776 5596 2779 se
rect 5596 2776 6635 2779
rect 2781 2750 4286 2776
tri 4286 2750 4312 2776 sw
rect 2781 2639 4312 2750
tri 5537 2720 5593 2776 se
rect 5593 2720 6635 2776
tri 5474 2657 5537 2720 se
rect 5537 2657 6635 2720
tri 5470 2653 5474 2657 se
rect 5474 2653 6635 2657
rect 2781 2583 3674 2639
rect 3730 2583 3756 2639
rect 3812 2583 3837 2639
rect 3893 2583 3918 2639
rect 3974 2583 3999 2639
rect 4055 2583 4080 2639
rect 4136 2583 4161 2639
rect 4217 2583 4242 2639
rect 4298 2583 4312 2639
tri 5414 2597 5470 2653 se
rect 5470 2597 6635 2653
rect 2781 2509 4312 2583
tri 5398 2581 5414 2597 se
rect 5414 2581 6635 2597
tri 5352 2535 5398 2581 se
rect 5398 2535 6635 2581
tri 5347 2530 5352 2535 se
rect 5352 2530 6635 2535
rect 2781 2453 3674 2509
rect 3730 2453 3756 2509
rect 3812 2453 3837 2509
rect 3893 2453 3918 2509
rect 3974 2453 3999 2509
rect 4055 2453 4080 2509
rect 4136 2453 4161 2509
rect 4217 2453 4242 2509
rect 4298 2453 4312 2509
tri 5291 2474 5347 2530 se
rect 5347 2474 6635 2530
tri 5276 2459 5291 2474 se
rect 5291 2459 6635 2474
rect 2781 2405 4312 2453
tri 5229 2412 5276 2459 se
rect 5276 2412 6635 2459
tri 5224 2407 5229 2412 se
rect 5229 2407 6635 2412
rect 2781 2351 4258 2405
tri 4258 2351 4312 2405 nw
tri 5168 2351 5224 2407 se
rect 5224 2404 6635 2407
rect 5224 2351 6582 2404
tri 6582 2351 6635 2404 nw
rect 6842 3145 7076 3150
rect 6842 3089 6847 3145
rect 6903 3089 6931 3145
rect 6987 3089 7015 3145
rect 7071 3089 7076 3145
rect 6842 3022 7076 3089
rect 6842 2966 6847 3022
rect 6903 2966 6931 3022
rect 6987 2966 7015 3022
rect 7071 2966 7076 3022
rect 6842 2899 7076 2966
rect 6842 2843 6847 2899
rect 6903 2843 6931 2899
rect 6987 2843 7015 2899
rect 7071 2843 7076 2899
rect 6842 2776 7076 2843
rect 6842 2720 6847 2776
rect 6903 2720 6931 2776
rect 6987 2720 7015 2776
rect 7071 2720 7076 2776
rect 6842 2706 7076 2720
rect 6842 2556 6847 2706
rect 6911 2642 6927 2706
rect 6991 2642 7007 2706
rect 6903 2620 6931 2642
rect 6987 2620 7015 2642
rect 6911 2556 6927 2620
rect 6991 2556 7007 2620
rect 7071 2556 7076 2706
rect 6842 2534 7076 2556
rect 6842 2470 6847 2534
rect 6911 2470 6927 2534
rect 6991 2470 7007 2534
rect 7071 2470 7076 2534
rect 6842 2448 7076 2470
rect 2781 2289 4196 2351
tri 4196 2289 4258 2351 nw
tri 5106 2289 5168 2351 se
rect 5168 2289 6520 2351
tri 6520 2289 6582 2351 nw
rect 6842 2298 6847 2448
rect 6911 2384 6927 2448
rect 6991 2384 7007 2448
rect 6903 2362 6931 2384
rect 6987 2362 7015 2384
rect 6911 2298 6927 2362
rect 6991 2298 7007 2362
rect 7071 2298 7076 2448
rect 2781 2284 4191 2289
tri 4191 2284 4196 2289 nw
tri 5101 2284 5106 2289 se
rect 5106 2284 6515 2289
tri 6515 2284 6520 2289 nw
rect 6842 2284 7076 2298
rect 2781 2228 4135 2284
tri 4135 2228 4191 2284 nw
tri 5045 2228 5101 2284 se
rect 5101 2228 6459 2284
tri 6459 2228 6515 2284 nw
rect 2781 2166 4073 2228
tri 4073 2166 4135 2228 nw
tri 4983 2166 5045 2228 se
rect 5045 2166 6397 2228
tri 6397 2166 6459 2228 nw
rect 6842 2212 6847 2284
rect 6903 2276 6931 2284
rect 6987 2276 7015 2284
rect 6911 2212 6927 2276
rect 6991 2212 7007 2276
rect 7071 2212 7076 2284
rect 6842 2190 7076 2212
rect 2781 2161 4068 2166
tri 4068 2161 4073 2166 nw
tri 4978 2161 4983 2166 se
rect 4983 2161 6392 2166
tri 6392 2161 6397 2166 nw
rect 2781 2105 4012 2161
tri 4012 2105 4068 2161 nw
tri 4922 2105 4978 2161 se
rect 4978 2105 6336 2161
tri 6336 2105 6392 2161 nw
rect 6842 2105 6847 2190
rect 6911 2126 6927 2190
rect 6991 2126 7007 2190
rect 6903 2105 6931 2126
rect 6987 2105 7015 2126
rect 7071 2105 7076 2190
rect 2781 2043 3950 2105
tri 3950 2043 4012 2105 nw
tri 4860 2043 4922 2105 se
rect 4922 2043 6274 2105
tri 6274 2043 6336 2105 nw
rect 6842 2103 7076 2105
rect 2781 2038 3945 2043
tri 3945 2038 3950 2043 nw
tri 4855 2038 4860 2043 se
rect 4860 2038 6269 2043
tri 6269 2038 6274 2043 nw
rect 6842 2039 6847 2103
rect 6911 2039 6927 2103
rect 6991 2039 7007 2103
rect 7071 2039 7076 2103
rect 6842 2038 7076 2039
rect 2781 1982 3889 2038
tri 3889 1982 3945 2038 nw
tri 4799 1982 4855 2038 se
rect 4855 1982 6213 2038
tri 6213 1982 6269 2038 nw
rect 2781 1915 3822 1982
tri 3822 1915 3889 1982 nw
tri 4732 1915 4799 1982 se
rect 4799 1915 6146 1982
tri 6146 1915 6213 1982 nw
rect 6842 1952 6847 2038
rect 6903 2016 6931 2038
rect 6987 2016 7015 2038
rect 6911 1952 6927 2016
rect 6991 1952 7007 2016
rect 7071 1952 7076 2038
rect 6842 1929 7076 1952
rect 2781 1087 3778 1915
tri 3778 1871 3822 1915 nw
tri 4688 1871 4732 1915 se
rect 4732 1871 6090 1915
tri 4676 1859 4688 1871 se
rect 4688 1859 6090 1871
tri 6090 1859 6146 1915 nw
rect 6842 1859 6847 1929
rect 6911 1865 6927 1929
rect 6991 1865 7007 1929
rect 6903 1859 6931 1865
rect 6987 1859 7015 1865
rect 7071 1859 7076 1929
tri 4671 1854 4676 1859 se
rect 4676 1854 6003 1859
tri 4666 1849 4671 1854 se
rect 4671 1849 6003 1854
tri 4589 1772 4666 1849 se
rect 4666 1772 6003 1849
tri 6003 1772 6090 1859 nw
rect 6842 1842 7076 1859
rect 6842 1778 6847 1842
rect 6911 1778 6927 1842
rect 6991 1778 7007 1842
rect 7071 1778 7076 1842
rect 8610 3145 8780 3150
rect 8610 3089 8615 3145
rect 8671 3089 8719 3145
rect 8775 3089 8780 3145
rect 8610 3023 8780 3089
rect 8610 2967 8615 3023
rect 8671 2967 8719 3023
rect 8775 2967 8780 3023
rect 8610 2901 8780 2967
rect 8610 2845 8615 2901
rect 8671 2845 8719 2901
rect 8775 2845 8780 2901
rect 8610 2779 8780 2845
rect 8610 2723 8615 2779
rect 8671 2723 8719 2779
rect 8775 2723 8780 2779
rect 8610 2706 8780 2723
rect 8674 2642 8716 2706
rect 8610 2621 8615 2642
rect 8671 2621 8719 2642
rect 8775 2621 8780 2642
rect 8674 2557 8716 2621
rect 8610 2536 8780 2557
rect 8674 2472 8716 2536
rect 8610 2450 8780 2472
rect 8674 2386 8716 2450
rect 8610 2364 8615 2386
rect 8671 2364 8719 2386
rect 8775 2364 8780 2386
rect 8674 2300 8716 2364
rect 8610 2289 8780 2300
rect 8610 2278 8615 2289
rect 8671 2278 8719 2289
rect 8775 2278 8780 2289
rect 8674 2214 8716 2278
rect 8610 2192 8780 2214
rect 8674 2128 8716 2192
rect 8610 2110 8615 2128
rect 8671 2110 8719 2128
rect 8775 2110 8780 2128
rect 8610 2106 8780 2110
rect 8674 2042 8716 2106
rect 8610 2020 8615 2042
rect 8671 2020 8719 2042
rect 8775 2020 8780 2042
rect 8674 1956 8716 2020
rect 8610 1934 8780 1956
rect 8674 1870 8716 1934
rect 8610 1848 8780 1870
rect 8674 1784 8716 1848
rect 8610 1778 8780 1784
rect 6842 1772 7076 1778
rect 2781 1031 2788 1087
rect 2844 1031 2889 1087
rect 2945 1031 2990 1087
rect 3046 1031 3091 1087
rect 3147 1031 3192 1087
rect 3248 1031 3293 1087
rect 3349 1031 3778 1087
rect 2781 937 3778 1031
rect 2781 881 2788 937
rect 2844 881 2889 937
rect 2945 881 2990 937
rect 3046 881 3091 937
rect 3147 881 3192 937
rect 3248 881 3293 937
rect 3349 881 3778 937
rect 2781 632 3778 881
tri 4527 1710 4589 1772 se
rect 4589 1710 5941 1772
tri 5941 1710 6003 1772 nw
rect 4527 1658 5889 1710
tri 5889 1658 5941 1710 nw
rect 4527 1653 5723 1658
rect 4527 1597 4857 1653
rect 4913 1597 4940 1653
rect 4996 1597 5023 1653
rect 5079 1597 5106 1653
rect 5162 1597 5188 1653
rect 5244 1597 5723 1653
rect 4527 1507 5723 1597
rect 4527 1451 4857 1507
rect 4913 1451 4940 1507
rect 4996 1451 5023 1507
rect 5079 1451 5106 1507
rect 5162 1451 5188 1507
rect 5244 1492 5723 1507
tri 5723 1492 5889 1658 nw
rect 5244 1486 5717 1492
tri 5717 1486 5723 1492 nw
rect 5244 1451 5677 1486
rect 4527 1446 5677 1451
tri 5677 1446 5717 1486 nw
rect 4527 1445 5676 1446
tri 5676 1445 5677 1446 nw
rect 4527 1430 5661 1445
tri 5661 1430 5676 1445 nw
rect 4527 1409 5635 1430
rect 4527 713 4862 1409
rect 5238 1404 5635 1409
tri 5635 1404 5661 1430 nw
rect 5238 1348 5579 1404
tri 5579 1348 5635 1404 nw
rect 5238 1322 5553 1348
tri 5553 1322 5579 1348 nw
rect 5238 713 5527 1322
tri 5527 1296 5553 1322 nw
rect 4527 688 5527 713
rect 4527 632 4862 688
rect 4918 632 4942 688
rect 4998 632 5022 688
rect 5078 632 5102 688
rect 5158 632 5182 688
rect 5238 632 5527 688
rect 2225 568 2699 589
rect 2225 504 2230 568
rect 2294 504 2310 568
rect 2374 504 2390 568
rect 2454 504 2470 568
rect 2534 504 2550 568
rect 2614 504 2630 568
rect 2694 504 2699 568
rect 2225 483 2699 504
rect 2225 419 2230 483
rect 2294 419 2310 483
rect 2374 419 2390 483
rect 2454 419 2470 483
rect 2534 419 2550 483
rect 2614 419 2630 483
rect 2694 419 2699 483
rect 2225 407 2699 419
rect 4527 607 5527 632
rect 4527 551 4862 607
rect 4918 551 4942 607
rect 4998 551 5022 607
rect 5078 551 5102 607
rect 5158 551 5182 607
rect 5238 551 5527 607
rect 4527 526 5527 551
rect 4527 470 4862 526
rect 4918 470 4942 526
rect 4998 470 5022 526
rect 5078 470 5102 526
rect 5158 470 5182 526
rect 5238 470 5527 526
rect 4527 445 5527 470
rect 1291 200 1388 256
rect 1444 200 1475 256
rect 1531 200 1562 256
rect 1618 200 1648 256
rect 1704 200 1734 256
rect 1790 200 1820 256
rect 1876 200 1906 256
rect 1962 200 1992 256
rect 2048 200 2078 256
rect 2134 200 2143 256
rect 1291 110 2143 200
rect 1291 54 1388 110
rect 1444 54 1475 110
rect 1531 54 1562 110
rect 1618 54 1648 110
rect 1704 54 1734 110
rect 1790 54 1820 110
rect 1876 54 1906 110
rect 1962 54 1992 110
rect 2048 54 2078 110
rect 2134 54 2143 110
rect 1291 49 2143 54
rect 4527 389 4862 445
rect 4918 389 4942 445
rect 4998 389 5022 445
rect 5078 389 5102 445
rect 5158 389 5182 445
rect 5238 389 5527 445
rect 4527 364 5527 389
rect 4527 308 4862 364
rect 4918 308 4942 364
rect 4998 308 5022 364
rect 5078 308 5102 364
rect 5158 308 5182 364
rect 5238 308 5527 364
rect 4527 257 5527 308
rect 4527 201 4608 257
rect 4664 201 4691 257
rect 4747 201 4774 257
rect 4830 201 4857 257
rect 4913 201 4940 257
rect 4996 201 5023 257
rect 5079 201 5106 257
rect 5162 201 5188 257
rect 5244 201 5527 257
rect 4527 111 5527 201
rect 4527 55 4608 111
rect 4664 55 4691 111
rect 4747 55 4774 111
rect 4830 55 4857 111
rect 4913 55 4940 111
rect 4996 55 5023 111
rect 5079 55 5106 111
rect 5162 55 5188 111
rect 5244 55 5527 111
rect 4527 50 5527 55
rect 9173 0 9239 7361
tri 9239 7333 9267 7361 nw
tri 9622 7347 9636 7361 ne
tri 9592 7238 9636 7282 se
rect 9636 7262 9702 7361
rect 9833 7291 9899 11244
tri 9899 7291 9912 7304 sw
tri 9702 7262 9724 7284 sw
rect 9636 7238 9724 7262
tri 9724 7238 9748 7262 sw
rect 9376 7174 9382 7238
rect 9446 7174 9462 7238
rect 9526 7174 9532 7238
rect 9592 7174 9598 7238
rect 9662 7174 9678 7238
rect 9742 7174 9748 7238
tri 9809 7238 9833 7262 se
rect 9833 7238 9912 7291
tri 9912 7238 9965 7291 sw
rect 9809 7174 9815 7238
rect 9879 7174 9895 7238
rect 9959 7174 9965 7238
tri 9382 7153 9403 7174 ne
rect 9403 7153 9511 7174
tri 9511 7153 9532 7174 nw
tri 9403 7132 9424 7153 ne
rect 9424 5949 9490 7153
tri 9490 7132 9511 7153 nw
tri 9424 5912 9461 5949 ne
rect 9461 5912 9490 5949
tri 9490 5912 9555 5977 sw
tri 9461 5883 9490 5912 ne
rect 9490 5883 9555 5912
tri 9490 5818 9555 5883 ne
tri 9555 5818 9649 5912 sw
tri 9555 5724 9649 5818 ne
tri 9649 5724 9743 5818 sw
tri 9649 5630 9743 5724 ne
tri 9743 5630 9837 5724 sw
tri 9743 5602 9771 5630 ne
rect 9771 758 9837 5630
rect 10025 3676 10315 11776
rect 11001 11604 11287 13844
rect 11010 10326 11277 10331
rect 11010 10270 11015 10326
rect 11071 10270 11116 10326
rect 11172 10270 11216 10326
rect 11272 10270 11277 10326
rect 11010 10216 11277 10270
rect 11010 10160 11015 10216
rect 11071 10160 11116 10216
rect 11172 10160 11216 10216
rect 11272 10160 11277 10216
rect 11010 10155 11277 10160
rect 10951 9471 11183 9476
rect 10951 9415 10956 9471
rect 11012 9415 11039 9471
rect 11095 9415 11122 9471
rect 11178 9415 11183 9471
rect 10951 9387 11183 9415
rect 10951 9331 10956 9387
rect 11012 9331 11039 9387
rect 11095 9331 11122 9387
rect 11178 9331 11183 9387
rect 10951 9326 11183 9331
rect 12122 9408 12128 9472
rect 12192 9408 12209 9472
rect 12273 9408 12279 9472
rect 10025 3612 10026 3676
rect 10090 3612 10138 3676
rect 10202 3612 10250 3676
rect 10314 3612 10315 3676
rect 10025 3590 10315 3612
rect 10025 3526 10026 3590
rect 10090 3526 10138 3590
rect 10202 3526 10250 3590
rect 10314 3526 10315 3590
rect 10025 3503 10315 3526
rect 10025 3439 10026 3503
rect 10090 3439 10138 3503
rect 10202 3439 10250 3503
rect 10314 3439 10315 3503
rect 10025 3416 10315 3439
rect 10025 3352 10026 3416
rect 10090 3352 10138 3416
rect 10202 3352 10250 3416
rect 10314 3352 10315 3416
rect 10025 3329 10315 3352
rect 10025 3265 10026 3329
rect 10090 3265 10138 3329
rect 10202 3265 10250 3329
rect 10314 3265 10315 3329
rect 10025 3242 10315 3265
rect 10025 3178 10026 3242
rect 10090 3178 10138 3242
rect 10202 3178 10250 3242
rect 10314 3178 10315 3242
rect 10025 3155 10315 3178
rect 10025 3091 10026 3155
rect 10090 3091 10138 3155
rect 10202 3091 10250 3155
rect 10314 3091 10315 3155
rect 10025 3068 10315 3091
rect 10025 3004 10026 3068
rect 10090 3004 10138 3068
rect 10202 3004 10250 3068
rect 10314 3004 10315 3068
rect 10025 2998 10315 3004
rect 10496 9238 11163 9246
rect 10496 9174 10503 9238
rect 10567 9174 10585 9238
rect 10649 9174 10667 9238
rect 10731 9174 10749 9238
rect 10813 9174 10831 9238
rect 10895 9174 10913 9238
rect 10977 9174 10995 9238
rect 11059 9174 11077 9238
rect 11141 9174 11163 9238
rect 10496 9154 11163 9174
rect 10496 9090 10503 9154
rect 10567 9090 10585 9154
rect 10649 9090 10667 9154
rect 10731 9090 10749 9154
rect 10813 9090 10831 9154
rect 10895 9090 10913 9154
rect 10977 9090 10995 9154
rect 11059 9090 11077 9154
rect 11141 9090 11163 9154
rect 10496 9070 11163 9090
rect 10496 9006 10503 9070
rect 10567 9006 10585 9070
rect 10649 9006 10667 9070
rect 10731 9006 10749 9070
rect 10813 9006 10831 9070
rect 10895 9006 10913 9070
rect 10977 9006 10995 9070
rect 11059 9006 11077 9070
rect 11141 9006 11163 9070
rect 10496 8986 11163 9006
rect 10496 8922 10503 8986
rect 10567 8922 10585 8986
rect 10649 8922 10667 8986
rect 10731 8922 10749 8986
rect 10813 8922 10831 8986
rect 10895 8922 10913 8986
rect 10977 8922 10995 8986
rect 11059 8922 11077 8986
rect 11141 8922 11163 8986
rect 10496 8902 11163 8922
rect 10496 8838 10503 8902
rect 10567 8838 10585 8902
rect 10649 8838 10667 8902
rect 10731 8838 10749 8902
rect 10813 8838 10831 8902
rect 10895 8838 10913 8902
rect 10977 8838 10995 8902
rect 11059 8838 11077 8902
rect 11141 8838 11163 8902
rect 10496 8818 11163 8838
rect 10496 8754 10503 8818
rect 10567 8754 10585 8818
rect 10649 8754 10667 8818
rect 10731 8754 10749 8818
rect 10813 8754 10831 8818
rect 10895 8754 10913 8818
rect 10977 8754 10995 8818
rect 11059 8754 11077 8818
rect 11141 8754 11163 8818
rect 10496 8734 11163 8754
rect 10496 8670 10503 8734
rect 10567 8670 10585 8734
rect 10649 8670 10667 8734
rect 10731 8670 10749 8734
rect 10813 8670 10831 8734
rect 10895 8670 10913 8734
rect 10977 8670 10995 8734
rect 11059 8670 11077 8734
rect 11141 8670 11163 8734
rect 10496 8650 11163 8670
rect 10496 8586 10503 8650
rect 10567 8586 10585 8650
rect 10649 8586 10667 8650
rect 10731 8586 10749 8650
rect 10813 8586 10831 8650
rect 10895 8586 10913 8650
rect 10977 8586 10995 8650
rect 11059 8586 11077 8650
rect 11141 8586 11163 8650
rect 10496 8566 11163 8586
rect 10496 8502 10503 8566
rect 10567 8502 10585 8566
rect 10649 8502 10667 8566
rect 10731 8502 10749 8566
rect 10813 8502 10831 8566
rect 10895 8502 10913 8566
rect 10977 8502 10995 8566
rect 11059 8502 11077 8566
rect 11141 8502 11163 8566
rect 10496 8482 11163 8502
rect 10496 8418 10503 8482
rect 10567 8418 10585 8482
rect 10649 8418 10667 8482
rect 10731 8418 10749 8482
rect 10813 8418 10831 8482
rect 10895 8418 10913 8482
rect 10977 8418 10995 8482
rect 11059 8418 11077 8482
rect 11141 8418 11163 8482
rect 10496 8397 11163 8418
rect 10496 8333 10503 8397
rect 10567 8333 10585 8397
rect 10649 8333 10667 8397
rect 10731 8333 10749 8397
rect 10813 8333 10831 8397
rect 10895 8333 10913 8397
rect 10977 8333 10995 8397
rect 11059 8333 11077 8397
rect 11141 8333 11163 8397
rect 10496 8235 11163 8333
rect 10496 8179 10506 8235
rect 10562 8179 10587 8235
rect 10643 8179 10668 8235
rect 10724 8179 11163 8235
rect 10496 5314 11163 8179
rect 10496 4831 11038 5314
tri 11038 5189 11163 5314 nw
rect 11122 4990 11132 5056
tri 11038 4831 11163 4956 sw
rect 9771 702 9776 758
rect 9832 702 9837 758
rect 9771 678 9837 702
rect 9771 622 9776 678
rect 9832 622 9837 678
rect 9771 617 9837 622
rect 10496 2637 11163 4831
rect 12122 3813 12279 9408
rect 12342 7235 12556 14660
tri 12556 14601 12615 14660 nw
tri 12998 9472 13068 9542 se
rect 13068 9472 13884 11557
tri 12934 9408 12998 9472 se
rect 12998 9408 13884 9472
tri 12772 9246 12934 9408 se
rect 12934 9246 13884 9408
tri 12664 9138 12772 9246 se
rect 12772 9204 13884 9246
rect 12772 9138 13818 9204
tri 13818 9138 13884 9204 nw
rect 14428 9647 15371 21149
rect 14428 9293 15315 9647
tri 15315 9591 15371 9647 nw
tri 15315 9293 15371 9349 sw
rect 12664 8030 13480 9138
tri 13480 8800 13818 9138 nw
rect 14428 8467 15371 9293
rect 12664 7966 12674 8030
rect 12738 7966 12755 8030
rect 12819 7966 12836 8030
rect 12900 7966 12917 8030
rect 12981 7966 12998 8030
rect 13062 7966 13078 8030
rect 13142 7966 13158 8030
rect 13222 7966 13238 8030
rect 13302 7966 13318 8030
rect 13382 7966 13398 8030
rect 13462 7966 13480 8030
rect 12664 7944 13480 7966
rect 12664 7880 12674 7944
rect 12738 7880 12755 7944
rect 12819 7880 12836 7944
rect 12900 7880 12917 7944
rect 12981 7880 12998 7944
rect 13062 7880 13078 7944
rect 13142 7880 13158 7944
rect 13222 7880 13238 7944
rect 13302 7880 13318 7944
rect 13382 7880 13398 7944
rect 13462 7880 13480 7944
rect 12664 7858 13480 7880
rect 12664 7794 12674 7858
rect 12738 7794 12755 7858
rect 12819 7794 12836 7858
rect 12900 7794 12917 7858
rect 12981 7794 12998 7858
rect 13062 7794 13078 7858
rect 13142 7794 13158 7858
rect 13222 7794 13238 7858
rect 13302 7794 13318 7858
rect 13382 7794 13398 7858
rect 13462 7794 13480 7858
rect 12664 7772 13480 7794
rect 12664 7708 12674 7772
rect 12738 7708 12755 7772
rect 12819 7708 12836 7772
rect 12900 7708 12917 7772
rect 12981 7708 12998 7772
rect 13062 7708 13078 7772
rect 13142 7708 13158 7772
rect 13222 7708 13238 7772
rect 13302 7708 13318 7772
rect 13382 7708 13398 7772
rect 13462 7708 13480 7772
rect 12664 7686 13480 7708
rect 12664 7622 12674 7686
rect 12738 7622 12755 7686
rect 12819 7622 12836 7686
rect 12900 7622 12917 7686
rect 12981 7622 12998 7686
rect 13062 7622 13078 7686
rect 13142 7622 13158 7686
rect 13222 7622 13238 7686
rect 13302 7622 13318 7686
rect 13382 7622 13398 7686
rect 13462 7622 13480 7686
rect 12664 7600 13480 7622
rect 12664 7536 12674 7600
rect 12738 7536 12755 7600
rect 12819 7536 12836 7600
rect 12900 7536 12917 7600
rect 12981 7536 12998 7600
rect 13062 7536 13078 7600
rect 13142 7536 13158 7600
rect 13222 7536 13238 7600
rect 13302 7536 13318 7600
rect 13382 7536 13398 7600
rect 13462 7536 13480 7600
rect 12664 7514 13480 7536
rect 12664 7450 12674 7514
rect 12738 7450 12755 7514
rect 12819 7450 12836 7514
rect 12900 7450 12917 7514
rect 12981 7450 12998 7514
rect 13062 7450 13078 7514
rect 13142 7450 13158 7514
rect 13222 7450 13238 7514
rect 13302 7450 13318 7514
rect 13382 7450 13398 7514
rect 13462 7450 13480 7514
rect 12664 7428 13480 7450
rect 12664 7364 12674 7428
rect 12738 7364 12755 7428
rect 12819 7364 12836 7428
rect 12900 7364 12917 7428
rect 12981 7364 12998 7428
rect 13062 7364 13078 7428
rect 13142 7364 13158 7428
rect 13222 7364 13238 7428
rect 13302 7364 13318 7428
rect 13382 7364 13398 7428
rect 13462 7364 13480 7428
rect 12664 7347 13480 7364
rect 13566 8313 14056 8355
rect 13566 8257 13577 8313
rect 13633 8257 13661 8313
rect 13717 8257 13745 8313
rect 13801 8257 13829 8313
rect 13885 8257 13912 8313
rect 13968 8257 13995 8313
rect 14051 8257 14056 8313
tri 12556 7235 12561 7240 sw
rect 12342 7209 12561 7235
tri 12561 7209 12587 7235 sw
rect 12342 7153 12587 7209
tri 12587 7153 12643 7209 sw
rect 12342 7152 12643 7153
tri 12643 7152 12644 7153 sw
tri 12342 7127 12367 7152 ne
rect 12367 7127 12644 7152
tri 12644 7127 12669 7152 sw
tri 12367 7071 12423 7127 ne
rect 12423 7071 12669 7127
tri 12669 7071 12725 7127 sw
tri 12423 7045 12449 7071 ne
rect 12449 7057 12725 7071
tri 12725 7057 12739 7071 sw
rect 12449 7045 12739 7057
tri 12449 6989 12505 7045 ne
rect 12505 6989 12739 7045
tri 12505 6969 12525 6989 ne
tri 12122 3707 12228 3813 ne
rect 12228 3707 12279 3813
tri 12279 3707 12450 3878 sw
tri 12228 3656 12279 3707 ne
rect 12279 3656 12450 3707
tri 12279 3641 12294 3656 ne
rect 10496 2581 10522 2637
rect 10578 2581 10614 2637
rect 10670 2581 10706 2637
rect 10762 2581 10798 2637
rect 10854 2581 10890 2637
rect 10946 2581 10982 2637
rect 11038 2581 11163 2637
rect 10496 2515 11163 2581
rect 10496 2459 10522 2515
rect 10578 2459 10614 2515
rect 10670 2459 10706 2515
rect 10762 2459 10798 2515
rect 10854 2459 10890 2515
rect 10946 2459 10982 2515
rect 11038 2459 11163 2515
rect 10496 1076 11163 2459
rect 11341 2706 11707 2712
rect 11341 2642 11342 2706
rect 11406 2642 11442 2706
rect 11506 2642 11542 2706
rect 11606 2642 11642 2706
rect 11706 2642 11707 2706
rect 11341 2621 11707 2642
rect 11341 2557 11342 2621
rect 11406 2557 11442 2621
rect 11506 2557 11542 2621
rect 11606 2557 11642 2621
rect 11706 2557 11707 2621
rect 11341 2536 11707 2557
rect 11341 2472 11342 2536
rect 11406 2472 11442 2536
rect 11506 2472 11542 2536
rect 11606 2472 11642 2536
rect 11706 2472 11707 2536
tri 12228 2495 12294 2561 se
rect 12294 2495 12450 3656
rect 12525 3614 12739 6989
tri 12739 3614 12778 3653 sw
rect 12525 3565 12778 3614
tri 12525 3526 12564 3565 ne
rect 11341 2451 11707 2472
rect 11341 2387 11342 2451
rect 11406 2387 11442 2451
rect 11506 2387 11542 2451
rect 11606 2387 11642 2451
rect 11706 2387 11707 2451
rect 11341 2366 11707 2387
rect 11341 2302 11342 2366
rect 11406 2302 11442 2366
rect 11506 2302 11542 2366
rect 11606 2302 11642 2366
rect 11706 2302 11707 2366
tri 12077 2344 12228 2495 se
rect 12228 2344 12299 2495
tri 12299 2344 12450 2495 nw
rect 11341 2280 11707 2302
rect 11341 2216 11342 2280
rect 11406 2216 11442 2280
rect 11506 2216 11542 2280
rect 11606 2216 11642 2280
rect 11706 2216 11707 2280
rect 11341 2194 11707 2216
rect 11341 2130 11342 2194
rect 11406 2130 11442 2194
rect 11506 2130 11542 2194
rect 11606 2130 11642 2194
rect 11706 2130 11707 2194
rect 11341 2108 11707 2130
rect 11341 2044 11342 2108
rect 11406 2044 11442 2108
rect 11506 2044 11542 2108
rect 11606 2044 11642 2108
rect 11706 2044 11707 2108
rect 11341 2022 11707 2044
rect 11341 1958 11342 2022
rect 11406 1958 11442 2022
rect 11506 1958 11542 2022
rect 11606 1958 11642 2022
rect 11706 1958 11707 2022
rect 11341 1936 11707 1958
rect 11341 1872 11342 1936
rect 11406 1872 11442 1936
rect 11506 1872 11542 1936
rect 11606 1872 11642 1936
rect 11706 1872 11707 1936
rect 11341 1850 11707 1872
rect 11341 1786 11342 1850
rect 11406 1786 11442 1850
rect 11506 1786 11542 1850
rect 11606 1786 11642 1850
rect 11706 1786 11707 1850
rect 11341 1780 11707 1786
tri 11920 2187 12077 2344 se
rect 11920 1486 12077 2187
tri 12077 2122 12299 2344 nw
rect 12564 1948 12778 3565
tri 12553 1550 12564 1561 se
rect 12564 1550 12778 1941
rect 13566 2706 14056 8257
rect 14136 8183 14348 8192
rect 14136 8127 14141 8183
rect 14197 8127 14285 8183
rect 14341 8127 14348 8183
rect 14136 8102 14348 8127
rect 14136 8046 14141 8102
rect 14197 8046 14285 8102
rect 14341 8046 14348 8102
rect 14136 8021 14348 8046
rect 14136 7965 14141 8021
rect 14197 7965 14285 8021
rect 14341 7965 14348 8021
rect 14136 7940 14348 7965
rect 14136 7884 14141 7940
rect 14197 7884 14285 7940
rect 14341 7884 14348 7940
rect 14136 7859 14348 7884
rect 14136 7803 14141 7859
rect 14197 7803 14285 7859
rect 14341 7803 14348 7859
rect 14136 7778 14348 7803
rect 14136 7722 14141 7778
rect 14197 7722 14285 7778
rect 14341 7722 14348 7778
rect 14136 7697 14348 7722
rect 14136 7641 14141 7697
rect 14197 7641 14285 7697
rect 14341 7641 14348 7697
rect 14136 7616 14348 7641
rect 14136 7560 14141 7616
rect 14197 7560 14285 7616
rect 14341 7560 14348 7616
rect 14136 7535 14348 7560
rect 14136 7479 14141 7535
rect 14197 7479 14285 7535
rect 14341 7479 14348 7535
rect 14136 7454 14348 7479
rect 14136 7398 14141 7454
rect 14197 7398 14285 7454
rect 14341 7398 14348 7454
rect 14136 7373 14348 7398
rect 14136 7317 14141 7373
rect 14197 7317 14285 7373
rect 14341 7317 14348 7373
rect 14136 7291 14348 7317
rect 14136 7235 14141 7291
rect 14197 7235 14285 7291
rect 14341 7235 14348 7291
rect 14136 7209 14348 7235
rect 14136 7153 14141 7209
rect 14197 7153 14285 7209
rect 14341 7153 14348 7209
rect 14136 7127 14348 7153
rect 14136 7071 14141 7127
rect 14197 7071 14285 7127
rect 14341 7071 14348 7127
rect 14136 7045 14348 7071
rect 14136 6989 14141 7045
rect 14197 6989 14285 7045
rect 14341 6989 14348 7045
rect 14136 6963 14348 6989
rect 14136 6907 14141 6963
rect 14197 6907 14285 6963
rect 14341 6907 14348 6963
rect 14136 6881 14348 6907
rect 14136 6825 14141 6881
rect 14197 6825 14285 6881
rect 14341 6825 14348 6881
rect 14136 6799 14348 6825
rect 14136 6743 14141 6799
rect 14197 6743 14285 6799
rect 14341 6743 14348 6799
rect 14136 6717 14348 6743
rect 14136 6661 14141 6717
rect 14197 6661 14285 6717
rect 14341 6661 14348 6717
rect 14136 6635 14348 6661
rect 14136 6579 14141 6635
rect 14197 6579 14285 6635
rect 14341 6579 14348 6635
rect 14136 6553 14348 6579
rect 14136 6497 14141 6553
rect 14197 6497 14285 6553
rect 14341 6497 14348 6553
rect 14136 6471 14348 6497
rect 14136 6415 14141 6471
rect 14197 6415 14285 6471
rect 14341 6415 14348 6471
rect 14136 6389 14348 6415
rect 14136 6333 14141 6389
rect 14197 6333 14285 6389
rect 14341 6333 14348 6389
rect 14136 4881 14348 6333
rect 14136 4817 14139 4881
rect 14203 4817 14283 4881
rect 14347 4817 14348 4881
rect 14136 4796 14348 4817
rect 14136 4732 14139 4796
rect 14203 4732 14283 4796
rect 14347 4732 14348 4796
rect 14136 4711 14348 4732
rect 14136 4647 14139 4711
rect 14203 4647 14283 4711
rect 14347 4647 14348 4711
rect 14136 4626 14348 4647
rect 14136 4562 14139 4626
rect 14203 4562 14283 4626
rect 14347 4562 14348 4626
rect 14136 4541 14348 4562
rect 14136 4477 14139 4541
rect 14203 4477 14283 4541
rect 14347 4477 14348 4541
rect 14136 4456 14348 4477
rect 14136 4392 14139 4456
rect 14203 4392 14283 4456
rect 14347 4392 14348 4456
rect 14136 4371 14348 4392
rect 14136 4307 14139 4371
rect 14203 4307 14283 4371
rect 14347 4307 14348 4371
rect 14136 4286 14348 4307
rect 14136 4222 14139 4286
rect 14203 4222 14283 4286
rect 14347 4222 14348 4286
rect 14136 4201 14348 4222
rect 14136 4137 14139 4201
rect 14203 4137 14283 4201
rect 14347 4137 14348 4201
rect 14136 4115 14348 4137
rect 14136 4051 14139 4115
rect 14203 4051 14283 4115
rect 14347 4051 14348 4115
rect 14136 4029 14348 4051
rect 14136 3965 14139 4029
rect 14203 3965 14283 4029
rect 14347 3965 14348 4029
rect 14136 3958 14348 3965
rect 14428 7930 15361 8467
tri 15361 8457 15371 8467 nw
tri 15361 7930 15371 7940 sw
rect 13566 2642 13569 2706
rect 13633 2642 13653 2706
rect 13717 2642 13737 2706
rect 13801 2642 13821 2706
rect 13885 2642 13905 2706
rect 13969 2642 13989 2706
rect 14053 2642 14056 2706
rect 13566 2621 14056 2642
rect 13566 2557 13569 2621
rect 13633 2557 13653 2621
rect 13717 2557 13737 2621
rect 13801 2557 13821 2621
rect 13885 2557 13905 2621
rect 13969 2557 13989 2621
rect 14053 2557 14056 2621
rect 13566 2535 14056 2557
rect 13566 2471 13569 2535
rect 13633 2471 13653 2535
rect 13717 2471 13737 2535
rect 13801 2471 13821 2535
rect 13885 2471 13905 2535
rect 13969 2471 13989 2535
rect 14053 2471 14056 2535
rect 13566 2449 14056 2471
rect 13566 2385 13569 2449
rect 13633 2385 13653 2449
rect 13717 2385 13737 2449
rect 13801 2385 13821 2449
rect 13885 2385 13905 2449
rect 13969 2385 13989 2449
rect 14053 2385 14056 2449
rect 13566 2363 14056 2385
rect 13566 2299 13569 2363
rect 13633 2299 13653 2363
rect 13717 2299 13737 2363
rect 13801 2299 13821 2363
rect 13885 2299 13905 2363
rect 13969 2299 13989 2363
rect 14053 2299 14056 2363
rect 13566 2277 14056 2299
rect 13566 2213 13569 2277
rect 13633 2213 13653 2277
rect 13717 2213 13737 2277
rect 13801 2213 13821 2277
rect 13885 2213 13905 2277
rect 13969 2213 13989 2277
rect 14053 2213 14056 2277
rect 13566 2191 14056 2213
rect 13566 2127 13569 2191
rect 13633 2127 13653 2191
rect 13717 2127 13737 2191
rect 13801 2127 13821 2191
rect 13885 2127 13905 2191
rect 13969 2127 13989 2191
rect 14053 2127 14056 2191
rect 13566 2105 14056 2127
rect 13566 2041 13569 2105
rect 13633 2041 13653 2105
rect 13717 2041 13737 2105
rect 13801 2041 13821 2105
rect 13885 2041 13905 2105
rect 13969 2041 13989 2105
rect 14053 2041 14056 2105
rect 13566 2019 14056 2041
rect 13566 1955 13569 2019
rect 13633 1955 13653 2019
rect 13717 1955 13737 2019
rect 13801 1955 13821 2019
rect 13885 1955 13905 2019
rect 13969 1955 13989 2019
rect 14053 1955 14056 2019
rect 13566 1933 14056 1955
rect 13566 1869 13569 1933
rect 13633 1869 13653 1933
rect 13717 1869 13737 1933
rect 13801 1869 13821 1933
rect 13885 1869 13905 1933
rect 13969 1869 13989 1933
rect 14053 1869 14056 1933
rect 13566 1847 14056 1869
rect 13566 1783 13569 1847
rect 13633 1783 13653 1847
rect 13717 1783 13737 1847
rect 13801 1783 13821 1847
rect 13885 1783 13905 1847
rect 13969 1783 13989 1847
rect 14053 1783 14056 1847
rect 13566 1777 14056 1783
tri 12077 1486 12141 1550 sw
tri 12489 1486 12553 1550 se
rect 12553 1486 12778 1550
rect 11920 1485 12141 1486
tri 11920 1430 11975 1485 ne
rect 11975 1430 12141 1485
tri 12141 1430 12197 1486 sw
tri 12433 1430 12489 1486 se
rect 12489 1430 12778 1486
tri 11975 1414 11991 1430 ne
rect 11991 1414 12197 1430
tri 12197 1414 12213 1430 sw
tri 12417 1414 12433 1430 se
rect 12433 1414 12778 1430
tri 11991 1404 12001 1414 ne
rect 12001 1404 12778 1414
tri 12001 1348 12057 1404 ne
rect 12057 1348 12778 1404
tri 12057 1328 12077 1348 ne
rect 12077 1328 12778 1348
tri 12077 1322 12083 1328 ne
rect 12083 1322 12778 1328
tri 12083 1266 12139 1322 ne
rect 12139 1266 12778 1322
tri 12139 1258 12147 1266 ne
rect 12147 1258 12778 1266
tri 12417 1111 12564 1258 ne
rect 10496 1020 10519 1076
rect 10575 1020 10600 1076
rect 10656 1020 10681 1076
rect 10737 1020 10763 1076
rect 10819 1020 11163 1076
rect 10496 994 11163 1020
rect 10496 938 10519 994
rect 10575 938 10600 994
rect 10656 938 10681 994
rect 10737 938 10763 994
rect 10819 938 11163 994
rect 10496 912 11163 938
rect 10496 856 10519 912
rect 10575 856 10600 912
rect 10656 856 10681 912
rect 10737 856 10763 912
rect 10819 856 11163 912
rect 10496 830 11163 856
rect 10496 774 10519 830
rect 10575 774 10600 830
rect 10656 774 10681 830
rect 10737 774 10763 830
rect 10819 774 11163 830
rect 10496 748 11163 774
rect 10496 692 10519 748
rect 10575 692 10600 748
rect 10656 692 10681 748
rect 10737 692 10763 748
rect 10819 692 11163 748
rect 10496 666 11163 692
rect 10496 610 10519 666
rect 10575 610 10600 666
rect 10656 610 10681 666
rect 10737 610 10763 666
rect 10819 610 11163 666
rect 10496 584 11163 610
rect 10496 528 10519 584
rect 10575 528 10600 584
rect 10656 528 10681 584
rect 10737 528 10763 584
rect 10819 528 11163 584
rect 10496 515 11163 528
rect 9883 430 10579 435
rect 9883 374 9888 430
rect 9944 374 9968 430
rect 10024 374 10579 430
rect 9883 369 10579 374
tri 10579 369 10645 435 sw
tri 10551 298 10622 369 ne
rect 10622 298 10645 369
tri 10645 298 10716 369 sw
rect 10337 234 10343 298
rect 10407 234 10423 298
rect 10487 234 10493 298
tri 10622 295 10625 298 ne
rect 10625 295 10714 298
tri 10625 275 10645 295 ne
rect 10645 275 10714 295
tri 10645 239 10681 275 ne
rect 10681 239 10714 275
tri 10681 237 10683 239 ne
rect 10683 237 10714 239
tri 10683 234 10686 237 ne
rect 10686 234 10714 237
rect 10778 234 10794 298
rect 10858 234 10864 298
tri 11099 295 11102 298 se
rect 11102 295 11207 298
tri 11043 239 11099 295 se
rect 11099 239 11207 295
tri 11041 237 11043 239 se
rect 11043 237 11207 239
tri 11038 234 11041 237 se
rect 11041 234 11207 237
rect 11271 234 11287 298
rect 11351 234 11357 298
rect 10337 232 10493 234
tri 11036 232 11038 234 se
rect 11038 232 11102 234
tri 11012 208 11036 232 se
rect 11036 208 11102 232
tri 11102 208 11128 234 nw
tri 10974 170 11012 208 se
rect 11012 170 11064 208
tri 11064 170 11102 208 nw
rect 9922 165 11000 170
rect 9922 109 9927 165
rect 9983 109 10007 165
rect 10063 109 11000 165
rect 9922 106 11000 109
tri 11000 106 11064 170 nw
rect 9922 104 10068 106
tri 10068 104 10070 106 nw
rect 12564 0 12778 1258
rect 14428 1486 15371 7930
rect 14428 1422 14438 1486
rect 14502 1422 14524 1486
rect 14588 1422 14610 1486
rect 14674 1422 14696 1486
rect 14760 1422 14782 1486
rect 14846 1422 14868 1486
rect 14932 1422 14954 1486
rect 15018 1422 15040 1486
rect 15104 1422 15126 1486
rect 15190 1422 15212 1486
rect 15276 1422 15298 1486
rect 15362 1422 15371 1486
rect 14428 1401 15371 1422
rect 14428 1337 14438 1401
rect 14502 1337 14524 1401
rect 14588 1337 14610 1401
rect 14674 1337 14696 1401
rect 14760 1337 14782 1401
rect 14846 1337 14868 1401
rect 14932 1337 14954 1401
rect 15018 1337 15040 1401
rect 15104 1337 15126 1401
rect 15190 1337 15212 1401
rect 15276 1337 15298 1401
rect 15362 1337 15371 1401
rect 14428 1316 15371 1337
rect 14428 1252 14438 1316
rect 14502 1252 14524 1316
rect 14588 1252 14610 1316
rect 14674 1252 14696 1316
rect 14760 1252 14782 1316
rect 14846 1252 14868 1316
rect 14932 1252 14954 1316
rect 15018 1252 15040 1316
rect 15104 1252 15126 1316
rect 15190 1252 15212 1316
rect 15276 1252 15298 1316
rect 15362 1252 15371 1316
rect 14428 1230 15371 1252
rect 14428 1166 14438 1230
rect 14502 1166 14524 1230
rect 14588 1166 14610 1230
rect 14674 1166 14696 1230
rect 14760 1166 14782 1230
rect 14846 1166 14868 1230
rect 14932 1166 14954 1230
rect 15018 1166 15040 1230
rect 15104 1166 15126 1230
rect 15190 1166 15212 1230
rect 15276 1166 15298 1230
rect 15362 1166 15371 1230
rect 14428 1144 15371 1166
rect 14428 1080 14438 1144
rect 14502 1080 14524 1144
rect 14588 1080 14610 1144
rect 14674 1080 14696 1144
rect 14760 1080 14782 1144
rect 14846 1080 14868 1144
rect 14932 1080 14954 1144
rect 15018 1080 15040 1144
rect 15104 1080 15126 1144
rect 15190 1080 15212 1144
rect 15276 1080 15298 1144
rect 15362 1080 15371 1144
rect 14428 1058 15371 1080
rect 14428 994 14438 1058
rect 14502 994 14524 1058
rect 14588 994 14610 1058
rect 14674 994 14696 1058
rect 14760 994 14782 1058
rect 14846 994 14868 1058
rect 14932 994 14954 1058
rect 15018 994 15040 1058
rect 15104 994 15126 1058
rect 15190 994 15212 1058
rect 15276 994 15298 1058
rect 15362 994 15371 1058
rect 14428 972 15371 994
rect 14428 908 14438 972
rect 14502 908 14524 972
rect 14588 908 14610 972
rect 14674 908 14696 972
rect 14760 908 14782 972
rect 14846 908 14868 972
rect 14932 908 14954 972
rect 15018 908 15040 972
rect 15104 908 15126 972
rect 15190 908 15212 972
rect 15276 908 15298 972
rect 15362 908 15371 972
rect 14428 886 15371 908
rect 14428 822 14438 886
rect 14502 822 14524 886
rect 14588 822 14610 886
rect 14674 822 14696 886
rect 14760 822 14782 886
rect 14846 822 14868 886
rect 14932 822 14954 886
rect 15018 822 15040 886
rect 15104 822 15126 886
rect 15190 822 15212 886
rect 15276 822 15298 886
rect 15362 822 15371 886
rect 14428 800 15371 822
rect 14428 736 14438 800
rect 14502 736 14524 800
rect 14588 736 14610 800
rect 14674 736 14696 800
rect 14760 736 14782 800
rect 14846 736 14868 800
rect 14932 736 14954 800
rect 15018 736 15040 800
rect 15104 736 15126 800
rect 15190 736 15212 800
rect 15276 736 15298 800
rect 15362 736 15371 800
rect 14428 714 15371 736
rect 14428 650 14438 714
rect 14502 650 14524 714
rect 14588 650 14610 714
rect 14674 650 14696 714
rect 14760 650 14782 714
rect 14846 650 14868 714
rect 14932 650 14954 714
rect 15018 650 15040 714
rect 15104 650 15126 714
rect 15190 650 15212 714
rect 15276 650 15298 714
rect 15362 650 15371 714
rect 14428 628 15371 650
rect 14428 564 14438 628
rect 14502 564 14524 628
rect 14588 564 14610 628
rect 14674 564 14696 628
rect 14760 564 14782 628
rect 14846 564 14868 628
rect 14932 564 14954 628
rect 15018 564 15040 628
rect 15104 564 15126 628
rect 15190 564 15212 628
rect 15276 564 15298 628
rect 15362 564 15371 628
rect 15589 1486 15655 1491
rect 15589 1430 15594 1486
rect 15650 1430 15655 1486
rect 15589 1404 15655 1430
rect 15589 1348 15594 1404
rect 15650 1348 15655 1404
rect 15589 1322 15655 1348
rect 15589 1266 15594 1322
rect 15650 1266 15655 1322
rect 14428 557 15371 564
tri 15565 557 15589 581 se
rect 15589 557 15655 1266
tri 15552 544 15565 557 se
rect 15565 544 15642 557
tri 15642 544 15655 557 nw
rect 13007 539 13163 544
rect 13007 483 13012 539
rect 13068 483 13102 539
rect 13158 483 13163 539
tri 15512 504 15552 544 se
rect 15552 504 15602 544
tri 15602 504 15642 544 nw
rect 13007 478 13163 483
tri 13054 430 13102 478 ne
tri 13055 298 13102 345 se
rect 13102 298 13163 478
tri 15422 414 15512 504 se
tri 15512 414 15602 504 nw
tri 15332 324 15422 414 se
tri 15422 324 15512 414 nw
tri 15308 300 15332 324 se
rect 15332 300 15398 324
tri 15398 300 15422 324 nw
rect 13007 234 13013 298
rect 13077 234 13093 298
rect 13157 234 13163 298
rect 13312 298 13468 300
tri 15306 298 15308 300 se
rect 15308 298 15391 300
rect 13312 295 13318 298
rect 13312 239 13317 295
rect 13312 234 13318 239
rect 13382 234 13398 298
rect 13462 295 13468 298
rect 13463 239 13468 295
rect 13462 234 13468 239
rect 15024 234 15030 298
rect 15094 234 15110 298
rect 15174 293 15391 298
tri 15391 293 15398 300 nw
rect 15482 293 15488 298
rect 15174 237 15335 293
tri 15335 237 15391 293 nw
rect 15482 237 15487 293
rect 15174 234 15332 237
tri 15332 234 15335 237 nw
rect 15482 234 15488 237
rect 15552 234 15568 298
rect 15632 293 15638 298
rect 15633 237 15638 293
rect 15632 234 15638 237
rect 15482 232 15638 234
rect 15716 0 15782 35296
rect 15848 0 15914 35296
<< rmetal3 >>
rect 1460 21317 1467 23791
rect 12564 1941 12778 1948
<< via3 >>
rect 5110 39301 5174 39365
rect 5190 39301 5254 39365
rect 5270 39301 5334 39365
rect 5350 39301 5414 39365
rect 5430 39301 5494 39365
rect 5510 39301 5574 39365
rect 5590 39301 5654 39365
rect 5670 39301 5734 39365
rect 5750 39301 5814 39365
rect 5830 39301 5894 39365
rect 5910 39301 5974 39365
rect 5990 39301 6054 39365
rect 6070 39301 6134 39365
rect 6150 39301 6214 39365
rect 6230 39301 6294 39365
rect 5110 39220 5174 39284
rect 5190 39220 5254 39284
rect 5270 39220 5334 39284
rect 5350 39220 5414 39284
rect 5430 39220 5494 39284
rect 5510 39220 5574 39284
rect 5590 39220 5654 39284
rect 5670 39220 5734 39284
rect 5750 39220 5814 39284
rect 5830 39220 5894 39284
rect 5910 39220 5974 39284
rect 5990 39220 6054 39284
rect 6070 39220 6134 39284
rect 6150 39220 6214 39284
rect 6230 39220 6294 39284
rect 5110 39139 5174 39203
rect 5190 39139 5254 39203
rect 5270 39139 5334 39203
rect 5350 39139 5414 39203
rect 5430 39139 5494 39203
rect 5510 39139 5574 39203
rect 5590 39139 5654 39203
rect 5670 39139 5734 39203
rect 5750 39139 5814 39203
rect 5830 39139 5894 39203
rect 5910 39139 5974 39203
rect 5990 39139 6054 39203
rect 6070 39139 6134 39203
rect 6150 39139 6214 39203
rect 6230 39139 6294 39203
rect 5110 39058 5174 39122
rect 5190 39058 5254 39122
rect 5270 39058 5334 39122
rect 5350 39058 5414 39122
rect 5430 39058 5494 39122
rect 5510 39058 5574 39122
rect 5590 39058 5654 39122
rect 5670 39058 5734 39122
rect 5750 39058 5814 39122
rect 5830 39058 5894 39122
rect 5910 39058 5974 39122
rect 5990 39058 6054 39122
rect 6070 39058 6134 39122
rect 6150 39058 6214 39122
rect 6230 39058 6294 39122
rect 5110 38977 5174 39041
rect 5190 38977 5254 39041
rect 5270 38977 5334 39041
rect 5350 38977 5414 39041
rect 5430 38977 5494 39041
rect 5510 38977 5574 39041
rect 5590 38977 5654 39041
rect 5670 38977 5734 39041
rect 5750 38977 5814 39041
rect 5830 38977 5894 39041
rect 5910 38977 5974 39041
rect 5990 38977 6054 39041
rect 6070 38977 6134 39041
rect 6150 38977 6214 39041
rect 6230 38977 6294 39041
rect 5110 38896 5174 38960
rect 5190 38896 5254 38960
rect 5270 38896 5334 38960
rect 5350 38896 5414 38960
rect 5430 38896 5494 38960
rect 5510 38896 5574 38960
rect 5590 38896 5654 38960
rect 5670 38896 5734 38960
rect 5750 38896 5814 38960
rect 5830 38896 5894 38960
rect 5910 38896 5974 38960
rect 5990 38896 6054 38960
rect 6070 38896 6134 38960
rect 6150 38896 6214 38960
rect 6230 38896 6294 38960
rect 5110 38815 5174 38879
rect 5190 38815 5254 38879
rect 5270 38815 5334 38879
rect 5350 38815 5414 38879
rect 5430 38815 5494 38879
rect 5510 38815 5574 38879
rect 5590 38815 5654 38879
rect 5670 38815 5734 38879
rect 5750 38815 5814 38879
rect 5830 38815 5894 38879
rect 5910 38815 5974 38879
rect 5990 38815 6054 38879
rect 6070 38815 6134 38879
rect 6150 38815 6214 38879
rect 6230 38815 6294 38879
rect 5110 38734 5174 38798
rect 5190 38734 5254 38798
rect 5270 38734 5334 38798
rect 5350 38734 5414 38798
rect 5430 38734 5494 38798
rect 5510 38734 5574 38798
rect 5590 38734 5654 38798
rect 5670 38734 5734 38798
rect 5750 38734 5814 38798
rect 5830 38734 5894 38798
rect 5910 38734 5974 38798
rect 5990 38734 6054 38798
rect 6070 38734 6134 38798
rect 6150 38734 6214 38798
rect 6230 38734 6294 38798
rect 5110 38653 5174 38717
rect 5190 38653 5254 38717
rect 5270 38653 5334 38717
rect 5350 38653 5414 38717
rect 5430 38653 5494 38717
rect 5510 38653 5574 38717
rect 5590 38653 5654 38717
rect 5670 38653 5734 38717
rect 5750 38653 5814 38717
rect 5830 38653 5894 38717
rect 5910 38653 5974 38717
rect 5990 38653 6054 38717
rect 6070 38653 6134 38717
rect 6150 38653 6214 38717
rect 6230 38653 6294 38717
rect 5110 38572 5174 38636
rect 5190 38572 5254 38636
rect 5270 38572 5334 38636
rect 5350 38572 5414 38636
rect 5430 38572 5494 38636
rect 5510 38572 5574 38636
rect 5590 38572 5654 38636
rect 5670 38572 5734 38636
rect 5750 38572 5814 38636
rect 5830 38572 5894 38636
rect 5910 38572 5974 38636
rect 5990 38572 6054 38636
rect 6070 38572 6134 38636
rect 6150 38572 6214 38636
rect 6230 38572 6294 38636
rect 5110 38491 5174 38555
rect 5190 38491 5254 38555
rect 5270 38491 5334 38555
rect 5350 38491 5414 38555
rect 5430 38491 5494 38555
rect 5510 38491 5574 38555
rect 5590 38491 5654 38555
rect 5670 38491 5734 38555
rect 5750 38491 5814 38555
rect 5830 38491 5894 38555
rect 5910 38491 5974 38555
rect 5990 38491 6054 38555
rect 6070 38491 6134 38555
rect 6150 38491 6214 38555
rect 6230 38491 6294 38555
rect 5110 38410 5174 38474
rect 5190 38410 5254 38474
rect 5270 38410 5334 38474
rect 5350 38410 5414 38474
rect 5430 38410 5494 38474
rect 5510 38410 5574 38474
rect 5590 38410 5654 38474
rect 5670 38410 5734 38474
rect 5750 38410 5814 38474
rect 5830 38410 5894 38474
rect 5910 38410 5974 38474
rect 5990 38410 6054 38474
rect 6070 38410 6134 38474
rect 6150 38410 6214 38474
rect 6230 38410 6294 38474
rect 5110 38329 5174 38393
rect 5190 38329 5254 38393
rect 5270 38329 5334 38393
rect 5350 38329 5414 38393
rect 5430 38329 5494 38393
rect 5510 38329 5574 38393
rect 5590 38329 5654 38393
rect 5670 38329 5734 38393
rect 5750 38329 5814 38393
rect 5830 38329 5894 38393
rect 5910 38329 5974 38393
rect 5990 38329 6054 38393
rect 6070 38329 6134 38393
rect 6150 38329 6214 38393
rect 6230 38329 6294 38393
rect 5110 38248 5174 38312
rect 5190 38248 5254 38312
rect 5270 38248 5334 38312
rect 5350 38248 5414 38312
rect 5430 38248 5494 38312
rect 5510 38248 5574 38312
rect 5590 38248 5654 38312
rect 5670 38248 5734 38312
rect 5750 38248 5814 38312
rect 5830 38248 5894 38312
rect 5910 38248 5974 38312
rect 5990 38248 6054 38312
rect 6070 38248 6134 38312
rect 6150 38248 6214 38312
rect 6230 38248 6294 38312
rect 5110 38167 5174 38231
rect 5190 38167 5254 38231
rect 5270 38167 5334 38231
rect 5350 38167 5414 38231
rect 5430 38167 5494 38231
rect 5510 38167 5574 38231
rect 5590 38167 5654 38231
rect 5670 38167 5734 38231
rect 5750 38167 5814 38231
rect 5830 38167 5894 38231
rect 5910 38167 5974 38231
rect 5990 38167 6054 38231
rect 6070 38167 6134 38231
rect 6150 38167 6214 38231
rect 6230 38167 6294 38231
rect 5110 38086 5174 38150
rect 5190 38086 5254 38150
rect 5270 38086 5334 38150
rect 5350 38086 5414 38150
rect 5430 38086 5494 38150
rect 5510 38086 5574 38150
rect 5590 38086 5654 38150
rect 5670 38086 5734 38150
rect 5750 38086 5814 38150
rect 5830 38086 5894 38150
rect 5910 38086 5974 38150
rect 5990 38086 6054 38150
rect 6070 38086 6134 38150
rect 6150 38086 6214 38150
rect 6230 38086 6294 38150
rect 5110 38005 5174 38069
rect 5190 38005 5254 38069
rect 5270 38005 5334 38069
rect 5350 38005 5414 38069
rect 5430 38005 5494 38069
rect 5510 38005 5574 38069
rect 5590 38005 5654 38069
rect 5670 38005 5734 38069
rect 5750 38005 5814 38069
rect 5830 38005 5894 38069
rect 5910 38005 5974 38069
rect 5990 38005 6054 38069
rect 6070 38005 6134 38069
rect 6150 38005 6214 38069
rect 6230 38005 6294 38069
rect 5110 37924 5174 37988
rect 5190 37924 5254 37988
rect 5270 37924 5334 37988
rect 5350 37924 5414 37988
rect 5430 37924 5494 37988
rect 5510 37924 5574 37988
rect 5590 37924 5654 37988
rect 5670 37924 5734 37988
rect 5750 37924 5814 37988
rect 5830 37924 5894 37988
rect 5910 37924 5974 37988
rect 5990 37924 6054 37988
rect 6070 37924 6134 37988
rect 6150 37924 6214 37988
rect 6230 37924 6294 37988
rect 5110 37843 5174 37907
rect 5190 37843 5254 37907
rect 5270 37843 5334 37907
rect 5350 37843 5414 37907
rect 5430 37843 5494 37907
rect 5510 37843 5574 37907
rect 5590 37843 5654 37907
rect 5670 37843 5734 37907
rect 5750 37843 5814 37907
rect 5830 37843 5894 37907
rect 5910 37843 5974 37907
rect 5990 37843 6054 37907
rect 6070 37843 6134 37907
rect 6150 37843 6214 37907
rect 6230 37843 6294 37907
rect 5110 37762 5174 37826
rect 5190 37762 5254 37826
rect 5270 37762 5334 37826
rect 5350 37762 5414 37826
rect 5430 37762 5494 37826
rect 5510 37762 5574 37826
rect 5590 37762 5654 37826
rect 5670 37762 5734 37826
rect 5750 37762 5814 37826
rect 5830 37762 5894 37826
rect 5910 37762 5974 37826
rect 5990 37762 6054 37826
rect 6070 37762 6134 37826
rect 6150 37762 6214 37826
rect 6230 37762 6294 37826
rect 5110 37681 5174 37745
rect 5190 37681 5254 37745
rect 5270 37681 5334 37745
rect 5350 37681 5414 37745
rect 5430 37681 5494 37745
rect 5510 37681 5574 37745
rect 5590 37681 5654 37745
rect 5670 37681 5734 37745
rect 5750 37681 5814 37745
rect 5830 37681 5894 37745
rect 5910 37681 5974 37745
rect 5990 37681 6054 37745
rect 6070 37681 6134 37745
rect 6150 37681 6214 37745
rect 6230 37681 6294 37745
rect 5110 37600 5174 37664
rect 5190 37600 5254 37664
rect 5270 37600 5334 37664
rect 5350 37600 5414 37664
rect 5430 37600 5494 37664
rect 5510 37600 5574 37664
rect 5590 37600 5654 37664
rect 5670 37600 5734 37664
rect 5750 37600 5814 37664
rect 5830 37600 5894 37664
rect 5910 37600 5974 37664
rect 5990 37600 6054 37664
rect 6070 37600 6134 37664
rect 6150 37600 6214 37664
rect 6230 37600 6294 37664
rect 5110 37519 5174 37583
rect 5190 37519 5254 37583
rect 5270 37519 5334 37583
rect 5350 37519 5414 37583
rect 5430 37519 5494 37583
rect 5510 37519 5574 37583
rect 5590 37519 5654 37583
rect 5670 37519 5734 37583
rect 5750 37519 5814 37583
rect 5830 37519 5894 37583
rect 5910 37519 5974 37583
rect 5990 37519 6054 37583
rect 6070 37519 6134 37583
rect 6150 37519 6214 37583
rect 6230 37519 6294 37583
rect 5110 37438 5174 37502
rect 5190 37438 5254 37502
rect 5270 37438 5334 37502
rect 5350 37438 5414 37502
rect 5430 37438 5494 37502
rect 5510 37438 5574 37502
rect 5590 37438 5654 37502
rect 5670 37438 5734 37502
rect 5750 37438 5814 37502
rect 5830 37438 5894 37502
rect 5910 37438 5974 37502
rect 5990 37438 6054 37502
rect 6070 37438 6134 37502
rect 6150 37438 6214 37502
rect 6230 37438 6294 37502
rect 5110 37357 5174 37421
rect 5190 37357 5254 37421
rect 5270 37357 5334 37421
rect 5350 37357 5414 37421
rect 5430 37357 5494 37421
rect 5510 37357 5574 37421
rect 5590 37357 5654 37421
rect 5670 37357 5734 37421
rect 5750 37357 5814 37421
rect 5830 37357 5894 37421
rect 5910 37357 5974 37421
rect 5990 37357 6054 37421
rect 6070 37357 6134 37421
rect 6150 37357 6214 37421
rect 6230 37357 6294 37421
rect 5110 37276 5174 37340
rect 5190 37276 5254 37340
rect 5270 37276 5334 37340
rect 5350 37276 5414 37340
rect 5430 37276 5494 37340
rect 5510 37276 5574 37340
rect 5590 37276 5654 37340
rect 5670 37276 5734 37340
rect 5750 37276 5814 37340
rect 5830 37276 5894 37340
rect 5910 37276 5974 37340
rect 5990 37276 6054 37340
rect 6070 37276 6134 37340
rect 6150 37276 6214 37340
rect 6230 37276 6294 37340
rect 5110 37195 5174 37259
rect 5190 37195 5254 37259
rect 5270 37195 5334 37259
rect 5350 37195 5414 37259
rect 5430 37195 5494 37259
rect 5510 37195 5574 37259
rect 5590 37195 5654 37259
rect 5670 37195 5734 37259
rect 5750 37195 5814 37259
rect 5830 37195 5894 37259
rect 5910 37195 5974 37259
rect 5990 37195 6054 37259
rect 6070 37195 6134 37259
rect 6150 37195 6214 37259
rect 6230 37195 6294 37259
rect 5110 37114 5174 37178
rect 5190 37114 5254 37178
rect 5270 37114 5334 37178
rect 5350 37114 5414 37178
rect 5430 37114 5494 37178
rect 5510 37114 5574 37178
rect 5590 37114 5654 37178
rect 5670 37114 5734 37178
rect 5750 37114 5814 37178
rect 5830 37114 5894 37178
rect 5910 37114 5974 37178
rect 5990 37114 6054 37178
rect 6070 37114 6134 37178
rect 6150 37114 6214 37178
rect 6230 37114 6294 37178
rect 5110 37033 5174 37097
rect 5190 37033 5254 37097
rect 5270 37033 5334 37097
rect 5350 37033 5414 37097
rect 5430 37033 5494 37097
rect 5510 37033 5574 37097
rect 5590 37033 5654 37097
rect 5670 37033 5734 37097
rect 5750 37033 5814 37097
rect 5830 37033 5894 37097
rect 5910 37033 5974 37097
rect 5990 37033 6054 37097
rect 6070 37033 6134 37097
rect 6150 37033 6214 37097
rect 6230 37033 6294 37097
rect 5110 36952 5174 37016
rect 5190 36952 5254 37016
rect 5270 36952 5334 37016
rect 5350 36952 5414 37016
rect 5430 36952 5494 37016
rect 5510 36952 5574 37016
rect 5590 36952 5654 37016
rect 5670 36952 5734 37016
rect 5750 36952 5814 37016
rect 5830 36952 5894 37016
rect 5910 36952 5974 37016
rect 5990 36952 6054 37016
rect 6070 36952 6134 37016
rect 6150 36952 6214 37016
rect 6230 36952 6294 37016
rect 5110 36871 5174 36935
rect 5190 36871 5254 36935
rect 5270 36871 5334 36935
rect 5350 36871 5414 36935
rect 5430 36871 5494 36935
rect 5510 36871 5574 36935
rect 5590 36871 5654 36935
rect 5670 36871 5734 36935
rect 5750 36871 5814 36935
rect 5830 36871 5894 36935
rect 5910 36871 5974 36935
rect 5990 36871 6054 36935
rect 6070 36871 6134 36935
rect 6150 36871 6214 36935
rect 6230 36871 6294 36935
rect 5110 36790 5174 36854
rect 5190 36790 5254 36854
rect 5270 36790 5334 36854
rect 5350 36790 5414 36854
rect 5430 36790 5494 36854
rect 5510 36790 5574 36854
rect 5590 36790 5654 36854
rect 5670 36790 5734 36854
rect 5750 36790 5814 36854
rect 5830 36790 5894 36854
rect 5910 36790 5974 36854
rect 5990 36790 6054 36854
rect 6070 36790 6134 36854
rect 6150 36790 6214 36854
rect 6230 36790 6294 36854
rect 5110 36709 5174 36773
rect 5190 36709 5254 36773
rect 5270 36709 5334 36773
rect 5350 36709 5414 36773
rect 5430 36709 5494 36773
rect 5510 36709 5574 36773
rect 5590 36709 5654 36773
rect 5670 36709 5734 36773
rect 5750 36709 5814 36773
rect 5830 36709 5894 36773
rect 5910 36709 5974 36773
rect 5990 36709 6054 36773
rect 6070 36709 6134 36773
rect 6150 36709 6214 36773
rect 6230 36709 6294 36773
rect 5110 36628 5174 36692
rect 5190 36628 5254 36692
rect 5270 36628 5334 36692
rect 5350 36628 5414 36692
rect 5430 36628 5494 36692
rect 5510 36628 5574 36692
rect 5590 36628 5654 36692
rect 5670 36628 5734 36692
rect 5750 36628 5814 36692
rect 5830 36628 5894 36692
rect 5910 36628 5974 36692
rect 5990 36628 6054 36692
rect 6070 36628 6134 36692
rect 6150 36628 6214 36692
rect 6230 36628 6294 36692
rect 5110 36547 5174 36611
rect 5190 36547 5254 36611
rect 5270 36547 5334 36611
rect 5350 36547 5414 36611
rect 5430 36547 5494 36611
rect 5510 36547 5574 36611
rect 5590 36547 5654 36611
rect 5670 36547 5734 36611
rect 5750 36547 5814 36611
rect 5830 36547 5894 36611
rect 5910 36547 5974 36611
rect 5990 36547 6054 36611
rect 6070 36547 6134 36611
rect 6150 36547 6214 36611
rect 6230 36547 6294 36611
rect 5110 36466 5174 36530
rect 5190 36466 5254 36530
rect 5270 36466 5334 36530
rect 5350 36466 5414 36530
rect 5430 36466 5494 36530
rect 5510 36466 5574 36530
rect 5590 36466 5654 36530
rect 5670 36466 5734 36530
rect 5750 36466 5814 36530
rect 5830 36466 5894 36530
rect 5910 36466 5974 36530
rect 5990 36466 6054 36530
rect 6070 36466 6134 36530
rect 6150 36466 6214 36530
rect 6230 36466 6294 36530
rect 2132 31159 2196 31167
rect 2132 31103 2139 31159
rect 2139 31103 2195 31159
rect 2195 31103 2196 31159
rect 2232 31159 2296 31167
rect 2232 31103 2237 31159
rect 2237 31103 2293 31159
rect 2293 31103 2296 31159
rect 2332 31159 2396 31167
rect 2332 31103 2335 31159
rect 2335 31103 2391 31159
rect 2391 31103 2396 31159
rect 2432 31159 2496 31167
rect 2432 31103 2433 31159
rect 2433 31103 2489 31159
rect 2489 31103 2496 31159
rect 2132 31077 2196 31085
rect 2132 31021 2139 31077
rect 2139 31021 2195 31077
rect 2195 31021 2196 31077
rect 2232 31077 2296 31085
rect 2232 31021 2237 31077
rect 2237 31021 2293 31077
rect 2293 31021 2296 31077
rect 2332 31077 2396 31085
rect 2332 31021 2335 31077
rect 2335 31021 2391 31077
rect 2391 31021 2396 31077
rect 2432 31077 2496 31085
rect 2432 31021 2433 31077
rect 2433 31021 2489 31077
rect 2489 31021 2496 31077
rect 2132 30995 2196 31003
rect 2132 30939 2139 30995
rect 2139 30939 2195 30995
rect 2195 30939 2196 30995
rect 2232 30995 2296 31003
rect 2232 30939 2237 30995
rect 2237 30939 2293 30995
rect 2293 30939 2296 30995
rect 2332 30995 2396 31003
rect 2332 30939 2335 30995
rect 2335 30939 2391 30995
rect 2391 30939 2396 30995
rect 2432 30995 2496 31003
rect 2432 30939 2433 30995
rect 2433 30939 2489 30995
rect 2489 30939 2496 30995
rect 2132 30913 2196 30921
rect 2132 30857 2139 30913
rect 2139 30857 2195 30913
rect 2195 30857 2196 30913
rect 2232 30913 2296 30921
rect 2232 30857 2237 30913
rect 2237 30857 2293 30913
rect 2293 30857 2296 30913
rect 2332 30913 2396 30921
rect 2332 30857 2335 30913
rect 2335 30857 2391 30913
rect 2391 30857 2396 30913
rect 2432 30913 2496 30921
rect 2432 30857 2433 30913
rect 2433 30857 2489 30913
rect 2489 30857 2496 30913
rect 2132 30831 2196 30839
rect 2132 30775 2139 30831
rect 2139 30775 2195 30831
rect 2195 30775 2196 30831
rect 2232 30831 2296 30839
rect 2232 30775 2237 30831
rect 2237 30775 2293 30831
rect 2293 30775 2296 30831
rect 2332 30831 2396 30839
rect 2332 30775 2335 30831
rect 2335 30775 2391 30831
rect 2391 30775 2396 30831
rect 2432 30831 2496 30839
rect 2432 30775 2433 30831
rect 2433 30775 2489 30831
rect 2489 30775 2496 30831
rect 2132 30749 2196 30757
rect 2132 30693 2139 30749
rect 2139 30693 2195 30749
rect 2195 30693 2196 30749
rect 2232 30749 2296 30757
rect 2232 30693 2237 30749
rect 2237 30693 2293 30749
rect 2293 30693 2296 30749
rect 2332 30749 2396 30757
rect 2332 30693 2335 30749
rect 2335 30693 2391 30749
rect 2391 30693 2396 30749
rect 2432 30749 2496 30757
rect 2432 30693 2433 30749
rect 2433 30693 2489 30749
rect 2489 30693 2496 30749
rect 2132 30667 2196 30675
rect 2132 30611 2139 30667
rect 2139 30611 2195 30667
rect 2195 30611 2196 30667
rect 2232 30667 2296 30675
rect 2232 30611 2237 30667
rect 2237 30611 2293 30667
rect 2293 30611 2296 30667
rect 2332 30667 2396 30675
rect 2332 30611 2335 30667
rect 2335 30611 2391 30667
rect 2391 30611 2396 30667
rect 2432 30667 2496 30675
rect 2432 30611 2433 30667
rect 2433 30611 2489 30667
rect 2489 30611 2496 30667
rect 2132 30585 2196 30593
rect 2132 30529 2139 30585
rect 2139 30529 2195 30585
rect 2195 30529 2196 30585
rect 2232 30585 2296 30593
rect 2232 30529 2237 30585
rect 2237 30529 2293 30585
rect 2293 30529 2296 30585
rect 2332 30585 2396 30593
rect 2332 30529 2335 30585
rect 2335 30529 2391 30585
rect 2391 30529 2396 30585
rect 2432 30585 2496 30593
rect 2432 30529 2433 30585
rect 2433 30529 2489 30585
rect 2489 30529 2496 30585
rect 2132 30503 2196 30511
rect 2132 30447 2139 30503
rect 2139 30447 2195 30503
rect 2195 30447 2196 30503
rect 2232 30503 2296 30511
rect 2232 30447 2237 30503
rect 2237 30447 2293 30503
rect 2293 30447 2296 30503
rect 2332 30503 2396 30511
rect 2332 30447 2335 30503
rect 2335 30447 2391 30503
rect 2391 30447 2396 30503
rect 2432 30503 2496 30511
rect 2432 30447 2433 30503
rect 2433 30447 2489 30503
rect 2489 30447 2496 30503
rect 2132 30421 2196 30429
rect 2132 30365 2139 30421
rect 2139 30365 2195 30421
rect 2195 30365 2196 30421
rect 2232 30421 2296 30429
rect 2232 30365 2237 30421
rect 2237 30365 2293 30421
rect 2293 30365 2296 30421
rect 2332 30421 2396 30429
rect 2332 30365 2335 30421
rect 2335 30365 2391 30421
rect 2391 30365 2396 30421
rect 2432 30421 2496 30429
rect 2432 30365 2433 30421
rect 2433 30365 2489 30421
rect 2489 30365 2496 30421
rect 2132 30338 2196 30347
rect 2132 30283 2139 30338
rect 2139 30283 2195 30338
rect 2195 30283 2196 30338
rect 2232 30338 2296 30347
rect 2232 30283 2237 30338
rect 2237 30283 2293 30338
rect 2293 30283 2296 30338
rect 2332 30338 2396 30347
rect 2332 30283 2335 30338
rect 2335 30283 2391 30338
rect 2391 30283 2396 30338
rect 2432 30338 2496 30347
rect 2432 30283 2433 30338
rect 2433 30283 2489 30338
rect 2489 30283 2496 30338
rect 2132 30255 2196 30264
rect 2132 30200 2139 30255
rect 2139 30200 2195 30255
rect 2195 30200 2196 30255
rect 2232 30255 2296 30264
rect 2232 30200 2237 30255
rect 2237 30200 2293 30255
rect 2293 30200 2296 30255
rect 2332 30255 2396 30264
rect 2332 30200 2335 30255
rect 2335 30200 2391 30255
rect 2391 30200 2396 30255
rect 2432 30255 2496 30264
rect 2432 30200 2433 30255
rect 2433 30200 2489 30255
rect 2489 30200 2496 30255
rect 2132 30172 2196 30181
rect 2132 30117 2139 30172
rect 2139 30117 2195 30172
rect 2195 30117 2196 30172
rect 2232 30172 2296 30181
rect 2232 30117 2237 30172
rect 2237 30117 2293 30172
rect 2293 30117 2296 30172
rect 2332 30172 2396 30181
rect 2332 30117 2335 30172
rect 2335 30117 2391 30172
rect 2391 30117 2396 30172
rect 2432 30172 2496 30181
rect 2432 30117 2433 30172
rect 2433 30117 2489 30172
rect 2489 30117 2496 30172
rect 2132 30089 2196 30098
rect 2132 30034 2139 30089
rect 2139 30034 2195 30089
rect 2195 30034 2196 30089
rect 2232 30089 2296 30098
rect 2232 30034 2237 30089
rect 2237 30034 2293 30089
rect 2293 30034 2296 30089
rect 2332 30089 2396 30098
rect 2332 30034 2335 30089
rect 2335 30034 2391 30089
rect 2391 30034 2396 30089
rect 2432 30089 2496 30098
rect 2432 30034 2433 30089
rect 2433 30034 2489 30089
rect 2489 30034 2496 30089
rect 2132 30006 2196 30015
rect 2132 29951 2139 30006
rect 2139 29951 2195 30006
rect 2195 29951 2196 30006
rect 2232 30006 2296 30015
rect 2232 29951 2237 30006
rect 2237 29951 2293 30006
rect 2293 29951 2296 30006
rect 2332 30006 2396 30015
rect 2332 29951 2335 30006
rect 2335 29951 2391 30006
rect 2391 29951 2396 30006
rect 2432 30006 2496 30015
rect 2432 29951 2433 30006
rect 2433 29951 2489 30006
rect 2489 29951 2496 30006
rect 2132 29923 2196 29932
rect 2132 29868 2139 29923
rect 2139 29868 2195 29923
rect 2195 29868 2196 29923
rect 2232 29923 2296 29932
rect 2232 29868 2237 29923
rect 2237 29868 2293 29923
rect 2293 29868 2296 29923
rect 2332 29923 2396 29932
rect 2332 29868 2335 29923
rect 2335 29868 2391 29923
rect 2391 29868 2396 29923
rect 2432 29923 2496 29932
rect 2432 29868 2433 29923
rect 2433 29868 2489 29923
rect 2489 29868 2496 29923
rect 2132 29840 2196 29849
rect 2132 29785 2139 29840
rect 2139 29785 2195 29840
rect 2195 29785 2196 29840
rect 2232 29840 2296 29849
rect 2232 29785 2237 29840
rect 2237 29785 2293 29840
rect 2293 29785 2296 29840
rect 2332 29840 2396 29849
rect 2332 29785 2335 29840
rect 2335 29785 2391 29840
rect 2391 29785 2396 29840
rect 2432 29840 2496 29849
rect 2432 29785 2433 29840
rect 2433 29785 2489 29840
rect 2489 29785 2496 29840
rect 2132 29757 2196 29766
rect 2132 29702 2139 29757
rect 2139 29702 2195 29757
rect 2195 29702 2196 29757
rect 2232 29757 2296 29766
rect 2232 29702 2237 29757
rect 2237 29702 2293 29757
rect 2293 29702 2296 29757
rect 2332 29757 2396 29766
rect 2332 29702 2335 29757
rect 2335 29702 2391 29757
rect 2391 29702 2396 29757
rect 2432 29757 2496 29766
rect 2432 29702 2433 29757
rect 2433 29702 2489 29757
rect 2489 29702 2496 29757
rect 2132 29674 2196 29683
rect 2132 29619 2139 29674
rect 2139 29619 2195 29674
rect 2195 29619 2196 29674
rect 2232 29674 2296 29683
rect 2232 29619 2237 29674
rect 2237 29619 2293 29674
rect 2293 29619 2296 29674
rect 2332 29674 2396 29683
rect 2332 29619 2335 29674
rect 2335 29619 2391 29674
rect 2391 29619 2396 29674
rect 2432 29674 2496 29683
rect 2432 29619 2433 29674
rect 2433 29619 2489 29674
rect 2489 29619 2496 29674
rect 2132 29591 2196 29600
rect 2132 29536 2139 29591
rect 2139 29536 2195 29591
rect 2195 29536 2196 29591
rect 2232 29591 2296 29600
rect 2232 29536 2237 29591
rect 2237 29536 2293 29591
rect 2293 29536 2296 29591
rect 2332 29591 2396 29600
rect 2332 29536 2335 29591
rect 2335 29536 2391 29591
rect 2391 29536 2396 29591
rect 2432 29591 2496 29600
rect 2432 29536 2433 29591
rect 2433 29536 2489 29591
rect 2489 29536 2496 29591
rect 2132 29508 2196 29517
rect 2132 29453 2139 29508
rect 2139 29453 2195 29508
rect 2195 29453 2196 29508
rect 2232 29508 2296 29517
rect 2232 29453 2237 29508
rect 2237 29453 2293 29508
rect 2293 29453 2296 29508
rect 2332 29508 2396 29517
rect 2332 29453 2335 29508
rect 2335 29453 2391 29508
rect 2391 29453 2396 29508
rect 2432 29508 2496 29517
rect 2432 29453 2433 29508
rect 2433 29453 2489 29508
rect 2489 29453 2496 29508
rect 2132 29425 2196 29434
rect 2132 29370 2139 29425
rect 2139 29370 2195 29425
rect 2195 29370 2196 29425
rect 2232 29425 2296 29434
rect 2232 29370 2237 29425
rect 2237 29370 2293 29425
rect 2293 29370 2296 29425
rect 2332 29425 2396 29434
rect 2332 29370 2335 29425
rect 2335 29370 2391 29425
rect 2391 29370 2396 29425
rect 2432 29425 2496 29434
rect 2432 29370 2433 29425
rect 2433 29370 2489 29425
rect 2489 29370 2496 29425
rect 2132 29342 2196 29351
rect 2132 29287 2139 29342
rect 2139 29287 2195 29342
rect 2195 29287 2196 29342
rect 2232 29342 2296 29351
rect 2232 29287 2237 29342
rect 2237 29287 2293 29342
rect 2293 29287 2296 29342
rect 2332 29342 2396 29351
rect 2332 29287 2335 29342
rect 2335 29287 2391 29342
rect 2391 29287 2396 29342
rect 2432 29342 2496 29351
rect 2432 29287 2433 29342
rect 2433 29287 2489 29342
rect 2489 29287 2496 29342
rect 2132 29259 2196 29268
rect 2132 29204 2139 29259
rect 2139 29204 2195 29259
rect 2195 29204 2196 29259
rect 2232 29259 2296 29268
rect 2232 29204 2237 29259
rect 2237 29204 2293 29259
rect 2293 29204 2296 29259
rect 2332 29259 2396 29268
rect 2332 29204 2335 29259
rect 2335 29204 2391 29259
rect 2391 29204 2396 29259
rect 2432 29259 2496 29268
rect 2432 29204 2433 29259
rect 2433 29204 2489 29259
rect 2489 29204 2496 29259
rect 2132 29176 2196 29185
rect 2132 29121 2139 29176
rect 2139 29121 2195 29176
rect 2195 29121 2196 29176
rect 2232 29176 2296 29185
rect 2232 29121 2237 29176
rect 2237 29121 2293 29176
rect 2293 29121 2296 29176
rect 2332 29176 2396 29185
rect 2332 29121 2335 29176
rect 2335 29121 2391 29176
rect 2391 29121 2396 29176
rect 2432 29176 2496 29185
rect 2432 29121 2433 29176
rect 2433 29121 2489 29176
rect 2489 29121 2496 29176
rect 2132 29093 2196 29102
rect 2132 29038 2139 29093
rect 2139 29038 2195 29093
rect 2195 29038 2196 29093
rect 2232 29093 2296 29102
rect 2232 29038 2237 29093
rect 2237 29038 2293 29093
rect 2293 29038 2296 29093
rect 2332 29093 2396 29102
rect 2332 29038 2335 29093
rect 2335 29038 2391 29093
rect 2391 29038 2396 29093
rect 2432 29093 2496 29102
rect 2432 29038 2433 29093
rect 2433 29038 2489 29093
rect 2489 29038 2496 29093
rect 2132 29010 2196 29019
rect 2132 28955 2139 29010
rect 2139 28955 2195 29010
rect 2195 28955 2196 29010
rect 2232 29010 2296 29019
rect 2232 28955 2237 29010
rect 2237 28955 2293 29010
rect 2293 28955 2296 29010
rect 2332 29010 2396 29019
rect 2332 28955 2335 29010
rect 2335 28955 2391 29010
rect 2391 28955 2396 29010
rect 2432 29010 2496 29019
rect 2432 28955 2433 29010
rect 2433 28955 2489 29010
rect 2489 28955 2496 29010
rect 2132 28927 2196 28936
rect 2132 28872 2139 28927
rect 2139 28872 2195 28927
rect 2195 28872 2196 28927
rect 2232 28927 2296 28936
rect 2232 28872 2237 28927
rect 2237 28872 2293 28927
rect 2293 28872 2296 28927
rect 2332 28927 2396 28936
rect 2332 28872 2335 28927
rect 2335 28872 2391 28927
rect 2391 28872 2396 28927
rect 2432 28927 2496 28936
rect 2432 28872 2433 28927
rect 2433 28872 2489 28927
rect 2489 28872 2496 28927
rect 4083 34617 4147 34681
rect 4165 34617 4229 34681
rect 4247 34617 4311 34681
rect 4329 34617 4393 34681
rect 4410 34617 4474 34681
rect 4491 34617 4555 34681
rect 4572 34617 4636 34681
rect 4653 34617 4717 34681
rect 4083 34529 4147 34593
rect 4165 34529 4229 34593
rect 4247 34529 4311 34593
rect 4329 34529 4393 34593
rect 4410 34529 4474 34593
rect 4491 34529 4555 34593
rect 4572 34529 4636 34593
rect 4653 34529 4717 34593
rect 4083 34441 4147 34505
rect 4165 34441 4229 34505
rect 4247 34441 4311 34505
rect 4329 34441 4393 34505
rect 4410 34441 4474 34505
rect 4491 34441 4555 34505
rect 4572 34441 4636 34505
rect 4653 34441 4717 34505
rect 4083 34353 4147 34417
rect 4165 34353 4229 34417
rect 4247 34353 4311 34417
rect 4329 34353 4393 34417
rect 4410 34353 4474 34417
rect 4491 34353 4555 34417
rect 4572 34353 4636 34417
rect 4653 34353 4717 34417
rect 4083 34265 4147 34329
rect 4165 34265 4229 34329
rect 4247 34265 4311 34329
rect 4329 34265 4393 34329
rect 4410 34265 4474 34329
rect 4491 34265 4555 34329
rect 4572 34265 4636 34329
rect 4653 34265 4717 34329
rect 4083 34177 4147 34241
rect 4165 34177 4229 34241
rect 4247 34177 4311 34241
rect 4329 34177 4393 34241
rect 4410 34177 4474 34241
rect 4491 34177 4555 34241
rect 4572 34177 4636 34241
rect 4653 34177 4717 34241
rect 5110 36385 5174 36449
rect 5190 36385 5254 36449
rect 5270 36385 5334 36449
rect 5350 36385 5414 36449
rect 5430 36385 5494 36449
rect 5510 36385 5574 36449
rect 5590 36385 5654 36449
rect 5670 36385 5734 36449
rect 5750 36385 5814 36449
rect 5830 36385 5894 36449
rect 5910 36385 5974 36449
rect 5990 36385 6054 36449
rect 6070 36385 6134 36449
rect 6150 36385 6214 36449
rect 6230 36385 6294 36449
rect 5110 36304 5174 36368
rect 5190 36304 5254 36368
rect 5270 36304 5334 36368
rect 5350 36304 5414 36368
rect 5430 36304 5494 36368
rect 5510 36304 5574 36368
rect 5590 36304 5654 36368
rect 5670 36304 5734 36368
rect 5750 36304 5814 36368
rect 5830 36304 5894 36368
rect 5910 36304 5974 36368
rect 5990 36304 6054 36368
rect 6070 36304 6134 36368
rect 6150 36304 6214 36368
rect 6230 36304 6294 36368
rect 5110 36223 5174 36287
rect 5190 36223 5254 36287
rect 5270 36223 5334 36287
rect 5350 36223 5414 36287
rect 5430 36223 5494 36287
rect 5510 36223 5574 36287
rect 5590 36223 5654 36287
rect 5670 36223 5734 36287
rect 5750 36223 5814 36287
rect 5830 36223 5894 36287
rect 5910 36223 5974 36287
rect 5990 36223 6054 36287
rect 6070 36223 6134 36287
rect 6150 36223 6214 36287
rect 6230 36223 6294 36287
rect 5110 36142 5174 36206
rect 5190 36142 5254 36206
rect 5270 36142 5334 36206
rect 5350 36142 5414 36206
rect 5430 36142 5494 36206
rect 5510 36142 5574 36206
rect 5590 36142 5654 36206
rect 5670 36142 5734 36206
rect 5750 36142 5814 36206
rect 5830 36142 5894 36206
rect 5910 36142 5974 36206
rect 5990 36142 6054 36206
rect 6070 36142 6134 36206
rect 6150 36142 6214 36206
rect 6230 36142 6294 36206
rect 5110 36060 5174 36124
rect 5190 36060 5254 36124
rect 5270 36060 5334 36124
rect 5350 36060 5414 36124
rect 5430 36060 5494 36124
rect 5510 36060 5574 36124
rect 5590 36060 5654 36124
rect 5670 36060 5734 36124
rect 5750 36060 5814 36124
rect 5830 36060 5894 36124
rect 5910 36060 5974 36124
rect 5990 36060 6054 36124
rect 6070 36060 6134 36124
rect 6150 36060 6214 36124
rect 6230 36060 6294 36124
rect 5110 35978 5174 36042
rect 5190 35978 5254 36042
rect 5270 35978 5334 36042
rect 5350 35978 5414 36042
rect 5430 35978 5494 36042
rect 5510 35978 5574 36042
rect 5590 35978 5654 36042
rect 5670 35978 5734 36042
rect 5750 35978 5814 36042
rect 5830 35978 5894 36042
rect 5910 35978 5974 36042
rect 5990 35978 6054 36042
rect 6070 35978 6134 36042
rect 6150 35978 6214 36042
rect 6230 35978 6294 36042
rect 5110 35896 5174 35960
rect 5190 35896 5254 35960
rect 5270 35896 5334 35960
rect 5350 35896 5414 35960
rect 5430 35896 5494 35960
rect 5510 35896 5574 35960
rect 5590 35896 5654 35960
rect 5670 35896 5734 35960
rect 5750 35896 5814 35960
rect 5830 35896 5894 35960
rect 5910 35896 5974 35960
rect 5990 35896 6054 35960
rect 6070 35896 6134 35960
rect 6150 35896 6214 35960
rect 6230 35896 6294 35960
rect 5110 35814 5174 35878
rect 5190 35814 5254 35878
rect 5270 35814 5334 35878
rect 5350 35814 5414 35878
rect 5430 35814 5494 35878
rect 5510 35814 5574 35878
rect 5590 35814 5654 35878
rect 5670 35814 5734 35878
rect 5750 35814 5814 35878
rect 5830 35814 5894 35878
rect 5910 35814 5974 35878
rect 5990 35814 6054 35878
rect 6070 35814 6134 35878
rect 6150 35814 6214 35878
rect 6230 35814 6294 35878
rect 5110 35732 5174 35796
rect 5190 35732 5254 35796
rect 5270 35732 5334 35796
rect 5350 35732 5414 35796
rect 5430 35732 5494 35796
rect 5510 35732 5574 35796
rect 5590 35732 5654 35796
rect 5670 35732 5734 35796
rect 5750 35732 5814 35796
rect 5830 35732 5894 35796
rect 5910 35732 5974 35796
rect 5990 35732 6054 35796
rect 6070 35732 6134 35796
rect 6150 35732 6214 35796
rect 6230 35732 6294 35796
rect 5110 35650 5174 35714
rect 5190 35650 5254 35714
rect 5270 35650 5334 35714
rect 5350 35650 5414 35714
rect 5430 35650 5494 35714
rect 5510 35650 5574 35714
rect 5590 35650 5654 35714
rect 5670 35650 5734 35714
rect 5750 35650 5814 35714
rect 5830 35650 5894 35714
rect 5910 35650 5974 35714
rect 5990 35650 6054 35714
rect 6070 35650 6134 35714
rect 6150 35650 6214 35714
rect 6230 35650 6294 35714
rect 5110 35568 5174 35632
rect 5190 35568 5254 35632
rect 5270 35568 5334 35632
rect 5350 35568 5414 35632
rect 5430 35568 5494 35632
rect 5510 35568 5574 35632
rect 5590 35568 5654 35632
rect 5670 35568 5734 35632
rect 5750 35568 5814 35632
rect 5830 35568 5894 35632
rect 5910 35568 5974 35632
rect 5990 35568 6054 35632
rect 6070 35568 6134 35632
rect 6150 35568 6214 35632
rect 6230 35568 6294 35632
rect 5110 35486 5174 35550
rect 5190 35486 5254 35550
rect 5270 35486 5334 35550
rect 5350 35486 5414 35550
rect 5430 35486 5494 35550
rect 5510 35486 5574 35550
rect 5590 35486 5654 35550
rect 5670 35486 5734 35550
rect 5750 35486 5814 35550
rect 5830 35486 5894 35550
rect 5910 35486 5974 35550
rect 5990 35486 6054 35550
rect 6070 35486 6134 35550
rect 6150 35486 6214 35550
rect 6230 35486 6294 35550
rect 5110 35404 5174 35468
rect 5190 35404 5254 35468
rect 5270 35404 5334 35468
rect 5350 35404 5414 35468
rect 5430 35404 5494 35468
rect 5510 35404 5574 35468
rect 5590 35404 5654 35468
rect 5670 35404 5734 35468
rect 5750 35404 5814 35468
rect 5830 35404 5894 35468
rect 5910 35404 5974 35468
rect 5990 35404 6054 35468
rect 6070 35404 6134 35468
rect 6150 35404 6214 35468
rect 6230 35404 6294 35468
rect 5110 35322 5174 35386
rect 5190 35322 5254 35386
rect 5270 35322 5334 35386
rect 5350 35322 5414 35386
rect 5430 35322 5494 35386
rect 5510 35322 5574 35386
rect 5590 35322 5654 35386
rect 5670 35322 5734 35386
rect 5750 35322 5814 35386
rect 5830 35322 5894 35386
rect 5910 35322 5974 35386
rect 5990 35322 6054 35386
rect 6070 35322 6134 35386
rect 6150 35322 6214 35386
rect 6230 35322 6294 35386
rect 5110 35240 5174 35304
rect 5190 35240 5254 35304
rect 5270 35240 5334 35304
rect 5350 35240 5414 35304
rect 5430 35240 5494 35304
rect 5510 35240 5574 35304
rect 5590 35240 5654 35304
rect 5670 35240 5734 35304
rect 5750 35240 5814 35304
rect 5830 35240 5894 35304
rect 5910 35240 5974 35304
rect 5990 35240 6054 35304
rect 6070 35240 6134 35304
rect 6150 35240 6214 35304
rect 6230 35240 6294 35304
rect 5110 35158 5174 35222
rect 5190 35158 5254 35222
rect 5270 35158 5334 35222
rect 5350 35158 5414 35222
rect 5430 35158 5494 35222
rect 5510 35158 5574 35222
rect 5590 35158 5654 35222
rect 5670 35158 5734 35222
rect 5750 35158 5814 35222
rect 5830 35158 5894 35222
rect 5910 35158 5974 35222
rect 5990 35158 6054 35222
rect 6070 35158 6134 35222
rect 6150 35158 6214 35222
rect 6230 35158 6294 35222
rect 6607 39301 6671 39365
rect 6687 39301 6751 39365
rect 6767 39301 6831 39365
rect 6847 39301 6911 39365
rect 6927 39301 6991 39365
rect 7007 39301 7071 39365
rect 7087 39301 7151 39365
rect 7167 39301 7231 39365
rect 7247 39301 7311 39365
rect 7327 39301 7391 39365
rect 7407 39301 7471 39365
rect 7487 39301 7551 39365
rect 7567 39301 7631 39365
rect 7647 39301 7711 39365
rect 7727 39301 7791 39365
rect 6607 39220 6671 39284
rect 6687 39220 6751 39284
rect 6767 39220 6831 39284
rect 6847 39220 6911 39284
rect 6927 39220 6991 39284
rect 7007 39220 7071 39284
rect 7087 39220 7151 39284
rect 7167 39220 7231 39284
rect 7247 39220 7311 39284
rect 7327 39220 7391 39284
rect 7407 39220 7471 39284
rect 7487 39220 7551 39284
rect 7567 39220 7631 39284
rect 7647 39220 7711 39284
rect 7727 39220 7791 39284
rect 6607 39139 6671 39203
rect 6687 39139 6751 39203
rect 6767 39139 6831 39203
rect 6847 39139 6911 39203
rect 6927 39139 6991 39203
rect 7007 39139 7071 39203
rect 7087 39139 7151 39203
rect 7167 39139 7231 39203
rect 7247 39139 7311 39203
rect 7327 39139 7391 39203
rect 7407 39139 7471 39203
rect 7487 39139 7551 39203
rect 7567 39139 7631 39203
rect 7647 39139 7711 39203
rect 7727 39139 7791 39203
rect 6607 39058 6671 39122
rect 6687 39058 6751 39122
rect 6767 39058 6831 39122
rect 6847 39058 6911 39122
rect 6927 39058 6991 39122
rect 7007 39058 7071 39122
rect 7087 39058 7151 39122
rect 7167 39058 7231 39122
rect 7247 39058 7311 39122
rect 7327 39058 7391 39122
rect 7407 39058 7471 39122
rect 7487 39058 7551 39122
rect 7567 39058 7631 39122
rect 7647 39058 7711 39122
rect 7727 39058 7791 39122
rect 6607 38977 6671 39041
rect 6687 38977 6751 39041
rect 6767 38977 6831 39041
rect 6847 38977 6911 39041
rect 6927 38977 6991 39041
rect 7007 38977 7071 39041
rect 7087 38977 7151 39041
rect 7167 38977 7231 39041
rect 7247 38977 7311 39041
rect 7327 38977 7391 39041
rect 7407 38977 7471 39041
rect 7487 38977 7551 39041
rect 7567 38977 7631 39041
rect 7647 38977 7711 39041
rect 7727 38977 7791 39041
rect 6607 38896 6671 38960
rect 6687 38896 6751 38960
rect 6767 38896 6831 38960
rect 6847 38896 6911 38960
rect 6927 38896 6991 38960
rect 7007 38896 7071 38960
rect 7087 38896 7151 38960
rect 7167 38896 7231 38960
rect 7247 38896 7311 38960
rect 7327 38896 7391 38960
rect 7407 38896 7471 38960
rect 7487 38896 7551 38960
rect 7567 38896 7631 38960
rect 7647 38896 7711 38960
rect 7727 38896 7791 38960
rect 6607 38815 6671 38879
rect 6687 38815 6751 38879
rect 6767 38815 6831 38879
rect 6847 38815 6911 38879
rect 6927 38815 6991 38879
rect 7007 38815 7071 38879
rect 7087 38815 7151 38879
rect 7167 38815 7231 38879
rect 7247 38815 7311 38879
rect 7327 38815 7391 38879
rect 7407 38815 7471 38879
rect 7487 38815 7551 38879
rect 7567 38815 7631 38879
rect 7647 38815 7711 38879
rect 7727 38815 7791 38879
rect 6607 38734 6671 38798
rect 6687 38734 6751 38798
rect 6767 38734 6831 38798
rect 6847 38734 6911 38798
rect 6927 38734 6991 38798
rect 7007 38734 7071 38798
rect 7087 38734 7151 38798
rect 7167 38734 7231 38798
rect 7247 38734 7311 38798
rect 7327 38734 7391 38798
rect 7407 38734 7471 38798
rect 7487 38734 7551 38798
rect 7567 38734 7631 38798
rect 7647 38734 7711 38798
rect 7727 38734 7791 38798
rect 6607 38653 6671 38717
rect 6687 38653 6751 38717
rect 6767 38653 6831 38717
rect 6847 38653 6911 38717
rect 6927 38653 6991 38717
rect 7007 38653 7071 38717
rect 7087 38653 7151 38717
rect 7167 38653 7231 38717
rect 7247 38653 7311 38717
rect 7327 38653 7391 38717
rect 7407 38653 7471 38717
rect 7487 38653 7551 38717
rect 7567 38653 7631 38717
rect 7647 38653 7711 38717
rect 7727 38653 7791 38717
rect 6607 38572 6671 38636
rect 6687 38572 6751 38636
rect 6767 38572 6831 38636
rect 6847 38572 6911 38636
rect 6927 38572 6991 38636
rect 7007 38572 7071 38636
rect 7087 38572 7151 38636
rect 7167 38572 7231 38636
rect 7247 38572 7311 38636
rect 7327 38572 7391 38636
rect 7407 38572 7471 38636
rect 7487 38572 7551 38636
rect 7567 38572 7631 38636
rect 7647 38572 7711 38636
rect 7727 38572 7791 38636
rect 6607 38491 6671 38555
rect 6687 38491 6751 38555
rect 6767 38491 6831 38555
rect 6847 38491 6911 38555
rect 6927 38491 6991 38555
rect 7007 38491 7071 38555
rect 7087 38491 7151 38555
rect 7167 38491 7231 38555
rect 7247 38491 7311 38555
rect 7327 38491 7391 38555
rect 7407 38491 7471 38555
rect 7487 38491 7551 38555
rect 7567 38491 7631 38555
rect 7647 38491 7711 38555
rect 7727 38491 7791 38555
rect 6607 38410 6671 38474
rect 6687 38410 6751 38474
rect 6767 38410 6831 38474
rect 6847 38410 6911 38474
rect 6927 38410 6991 38474
rect 7007 38410 7071 38474
rect 7087 38410 7151 38474
rect 7167 38410 7231 38474
rect 7247 38410 7311 38474
rect 7327 38410 7391 38474
rect 7407 38410 7471 38474
rect 7487 38410 7551 38474
rect 7567 38410 7631 38474
rect 7647 38410 7711 38474
rect 7727 38410 7791 38474
rect 6607 38329 6671 38393
rect 6687 38329 6751 38393
rect 6767 38329 6831 38393
rect 6847 38329 6911 38393
rect 6927 38329 6991 38393
rect 7007 38329 7071 38393
rect 7087 38329 7151 38393
rect 7167 38329 7231 38393
rect 7247 38329 7311 38393
rect 7327 38329 7391 38393
rect 7407 38329 7471 38393
rect 7487 38329 7551 38393
rect 7567 38329 7631 38393
rect 7647 38329 7711 38393
rect 7727 38329 7791 38393
rect 6607 38248 6671 38312
rect 6687 38248 6751 38312
rect 6767 38248 6831 38312
rect 6847 38248 6911 38312
rect 6927 38248 6991 38312
rect 7007 38248 7071 38312
rect 7087 38248 7151 38312
rect 7167 38248 7231 38312
rect 7247 38248 7311 38312
rect 7327 38248 7391 38312
rect 7407 38248 7471 38312
rect 7487 38248 7551 38312
rect 7567 38248 7631 38312
rect 7647 38248 7711 38312
rect 7727 38248 7791 38312
rect 6607 38167 6671 38231
rect 6687 38167 6751 38231
rect 6767 38167 6831 38231
rect 6847 38167 6911 38231
rect 6927 38167 6991 38231
rect 7007 38167 7071 38231
rect 7087 38167 7151 38231
rect 7167 38167 7231 38231
rect 7247 38167 7311 38231
rect 7327 38167 7391 38231
rect 7407 38167 7471 38231
rect 7487 38167 7551 38231
rect 7567 38167 7631 38231
rect 7647 38167 7711 38231
rect 7727 38167 7791 38231
rect 6607 38086 6671 38150
rect 6687 38086 6751 38150
rect 6767 38086 6831 38150
rect 6847 38086 6911 38150
rect 6927 38086 6991 38150
rect 7007 38086 7071 38150
rect 7087 38086 7151 38150
rect 7167 38086 7231 38150
rect 7247 38086 7311 38150
rect 7327 38086 7391 38150
rect 7407 38086 7471 38150
rect 7487 38086 7551 38150
rect 7567 38086 7631 38150
rect 7647 38086 7711 38150
rect 7727 38086 7791 38150
rect 6607 38005 6671 38069
rect 6687 38005 6751 38069
rect 6767 38005 6831 38069
rect 6847 38005 6911 38069
rect 6927 38005 6991 38069
rect 7007 38005 7071 38069
rect 7087 38005 7151 38069
rect 7167 38005 7231 38069
rect 7247 38005 7311 38069
rect 7327 38005 7391 38069
rect 7407 38005 7471 38069
rect 7487 38005 7551 38069
rect 7567 38005 7631 38069
rect 7647 38005 7711 38069
rect 7727 38005 7791 38069
rect 6607 37924 6671 37988
rect 6687 37924 6751 37988
rect 6767 37924 6831 37988
rect 6847 37924 6911 37988
rect 6927 37924 6991 37988
rect 7007 37924 7071 37988
rect 7087 37924 7151 37988
rect 7167 37924 7231 37988
rect 7247 37924 7311 37988
rect 7327 37924 7391 37988
rect 7407 37924 7471 37988
rect 7487 37924 7551 37988
rect 7567 37924 7631 37988
rect 7647 37924 7711 37988
rect 7727 37924 7791 37988
rect 6607 37843 6671 37907
rect 6687 37843 6751 37907
rect 6767 37843 6831 37907
rect 6847 37843 6911 37907
rect 6927 37843 6991 37907
rect 7007 37843 7071 37907
rect 7087 37843 7151 37907
rect 7167 37843 7231 37907
rect 7247 37843 7311 37907
rect 7327 37843 7391 37907
rect 7407 37843 7471 37907
rect 7487 37843 7551 37907
rect 7567 37843 7631 37907
rect 7647 37843 7711 37907
rect 7727 37843 7791 37907
rect 6607 37762 6671 37826
rect 6687 37762 6751 37826
rect 6767 37762 6831 37826
rect 6847 37762 6911 37826
rect 6927 37762 6991 37826
rect 7007 37762 7071 37826
rect 7087 37762 7151 37826
rect 7167 37762 7231 37826
rect 7247 37762 7311 37826
rect 7327 37762 7391 37826
rect 7407 37762 7471 37826
rect 7487 37762 7551 37826
rect 7567 37762 7631 37826
rect 7647 37762 7711 37826
rect 7727 37762 7791 37826
rect 6607 37681 6671 37745
rect 6687 37681 6751 37745
rect 6767 37681 6831 37745
rect 6847 37681 6911 37745
rect 6927 37681 6991 37745
rect 7007 37681 7071 37745
rect 7087 37681 7151 37745
rect 7167 37681 7231 37745
rect 7247 37681 7311 37745
rect 7327 37681 7391 37745
rect 7407 37681 7471 37745
rect 7487 37681 7551 37745
rect 7567 37681 7631 37745
rect 7647 37681 7711 37745
rect 7727 37681 7791 37745
rect 6607 37600 6671 37664
rect 6687 37600 6751 37664
rect 6767 37600 6831 37664
rect 6847 37600 6911 37664
rect 6927 37600 6991 37664
rect 7007 37600 7071 37664
rect 7087 37600 7151 37664
rect 7167 37600 7231 37664
rect 7247 37600 7311 37664
rect 7327 37600 7391 37664
rect 7407 37600 7471 37664
rect 7487 37600 7551 37664
rect 7567 37600 7631 37664
rect 7647 37600 7711 37664
rect 7727 37600 7791 37664
rect 6607 37519 6671 37583
rect 6687 37519 6751 37583
rect 6767 37519 6831 37583
rect 6847 37519 6911 37583
rect 6927 37519 6991 37583
rect 7007 37519 7071 37583
rect 7087 37519 7151 37583
rect 7167 37519 7231 37583
rect 7247 37519 7311 37583
rect 7327 37519 7391 37583
rect 7407 37519 7471 37583
rect 7487 37519 7551 37583
rect 7567 37519 7631 37583
rect 7647 37519 7711 37583
rect 7727 37519 7791 37583
rect 6607 37438 6671 37502
rect 6687 37438 6751 37502
rect 6767 37438 6831 37502
rect 6847 37438 6911 37502
rect 6927 37438 6991 37502
rect 7007 37438 7071 37502
rect 7087 37438 7151 37502
rect 7167 37438 7231 37502
rect 7247 37438 7311 37502
rect 7327 37438 7391 37502
rect 7407 37438 7471 37502
rect 7487 37438 7551 37502
rect 7567 37438 7631 37502
rect 7647 37438 7711 37502
rect 7727 37438 7791 37502
rect 6607 37357 6671 37421
rect 6687 37357 6751 37421
rect 6767 37357 6831 37421
rect 6847 37357 6911 37421
rect 6927 37357 6991 37421
rect 7007 37357 7071 37421
rect 7087 37357 7151 37421
rect 7167 37357 7231 37421
rect 7247 37357 7311 37421
rect 7327 37357 7391 37421
rect 7407 37357 7471 37421
rect 7487 37357 7551 37421
rect 7567 37357 7631 37421
rect 7647 37357 7711 37421
rect 7727 37357 7791 37421
rect 6607 37276 6671 37340
rect 6687 37276 6751 37340
rect 6767 37276 6831 37340
rect 6847 37276 6911 37340
rect 6927 37276 6991 37340
rect 7007 37276 7071 37340
rect 7087 37276 7151 37340
rect 7167 37276 7231 37340
rect 7247 37276 7311 37340
rect 7327 37276 7391 37340
rect 7407 37276 7471 37340
rect 7487 37276 7551 37340
rect 7567 37276 7631 37340
rect 7647 37276 7711 37340
rect 7727 37276 7791 37340
rect 6607 37195 6671 37259
rect 6687 37195 6751 37259
rect 6767 37195 6831 37259
rect 6847 37195 6911 37259
rect 6927 37195 6991 37259
rect 7007 37195 7071 37259
rect 7087 37195 7151 37259
rect 7167 37195 7231 37259
rect 7247 37195 7311 37259
rect 7327 37195 7391 37259
rect 7407 37195 7471 37259
rect 7487 37195 7551 37259
rect 7567 37195 7631 37259
rect 7647 37195 7711 37259
rect 7727 37195 7791 37259
rect 6607 37114 6671 37178
rect 6687 37114 6751 37178
rect 6767 37114 6831 37178
rect 6847 37114 6911 37178
rect 6927 37114 6991 37178
rect 7007 37114 7071 37178
rect 7087 37114 7151 37178
rect 7167 37114 7231 37178
rect 7247 37114 7311 37178
rect 7327 37114 7391 37178
rect 7407 37114 7471 37178
rect 7487 37114 7551 37178
rect 7567 37114 7631 37178
rect 7647 37114 7711 37178
rect 7727 37114 7791 37178
rect 6607 37033 6671 37097
rect 6687 37033 6751 37097
rect 6767 37033 6831 37097
rect 6847 37033 6911 37097
rect 6927 37033 6991 37097
rect 7007 37033 7071 37097
rect 7087 37033 7151 37097
rect 7167 37033 7231 37097
rect 7247 37033 7311 37097
rect 7327 37033 7391 37097
rect 7407 37033 7471 37097
rect 7487 37033 7551 37097
rect 7567 37033 7631 37097
rect 7647 37033 7711 37097
rect 7727 37033 7791 37097
rect 6607 36952 6671 37016
rect 6687 36952 6751 37016
rect 6767 36952 6831 37016
rect 6847 36952 6911 37016
rect 6927 36952 6991 37016
rect 7007 36952 7071 37016
rect 7087 36952 7151 37016
rect 7167 36952 7231 37016
rect 7247 36952 7311 37016
rect 7327 36952 7391 37016
rect 7407 36952 7471 37016
rect 7487 36952 7551 37016
rect 7567 36952 7631 37016
rect 7647 36952 7711 37016
rect 7727 36952 7791 37016
rect 6607 36871 6671 36935
rect 6687 36871 6751 36935
rect 6767 36871 6831 36935
rect 6847 36871 6911 36935
rect 6927 36871 6991 36935
rect 7007 36871 7071 36935
rect 7087 36871 7151 36935
rect 7167 36871 7231 36935
rect 7247 36871 7311 36935
rect 7327 36871 7391 36935
rect 7407 36871 7471 36935
rect 7487 36871 7551 36935
rect 7567 36871 7631 36935
rect 7647 36871 7711 36935
rect 7727 36871 7791 36935
rect 6607 36790 6671 36854
rect 6687 36790 6751 36854
rect 6767 36790 6831 36854
rect 6847 36790 6911 36854
rect 6927 36790 6991 36854
rect 7007 36790 7071 36854
rect 7087 36790 7151 36854
rect 7167 36790 7231 36854
rect 7247 36790 7311 36854
rect 7327 36790 7391 36854
rect 7407 36790 7471 36854
rect 7487 36790 7551 36854
rect 7567 36790 7631 36854
rect 7647 36790 7711 36854
rect 7727 36790 7791 36854
rect 6607 36709 6671 36773
rect 6687 36709 6751 36773
rect 6767 36709 6831 36773
rect 6847 36709 6911 36773
rect 6927 36709 6991 36773
rect 7007 36709 7071 36773
rect 7087 36709 7151 36773
rect 7167 36709 7231 36773
rect 7247 36709 7311 36773
rect 7327 36709 7391 36773
rect 7407 36709 7471 36773
rect 7487 36709 7551 36773
rect 7567 36709 7631 36773
rect 7647 36709 7711 36773
rect 7727 36709 7791 36773
rect 6607 36628 6671 36692
rect 6687 36628 6751 36692
rect 6767 36628 6831 36692
rect 6847 36628 6911 36692
rect 6927 36628 6991 36692
rect 7007 36628 7071 36692
rect 7087 36628 7151 36692
rect 7167 36628 7231 36692
rect 7247 36628 7311 36692
rect 7327 36628 7391 36692
rect 7407 36628 7471 36692
rect 7487 36628 7551 36692
rect 7567 36628 7631 36692
rect 7647 36628 7711 36692
rect 7727 36628 7791 36692
rect 6607 36547 6671 36611
rect 6687 36547 6751 36611
rect 6767 36547 6831 36611
rect 6847 36547 6911 36611
rect 6927 36547 6991 36611
rect 7007 36547 7071 36611
rect 7087 36547 7151 36611
rect 7167 36547 7231 36611
rect 7247 36547 7311 36611
rect 7327 36547 7391 36611
rect 7407 36547 7471 36611
rect 7487 36547 7551 36611
rect 7567 36547 7631 36611
rect 7647 36547 7711 36611
rect 7727 36547 7791 36611
rect 6607 36466 6671 36530
rect 6687 36466 6751 36530
rect 6767 36466 6831 36530
rect 6847 36466 6911 36530
rect 6927 36466 6991 36530
rect 7007 36466 7071 36530
rect 7087 36466 7151 36530
rect 7167 36466 7231 36530
rect 7247 36466 7311 36530
rect 7327 36466 7391 36530
rect 7407 36466 7471 36530
rect 7487 36466 7551 36530
rect 7567 36466 7631 36530
rect 7647 36466 7711 36530
rect 7727 36466 7791 36530
rect 6607 36385 6671 36449
rect 6687 36385 6751 36449
rect 6767 36385 6831 36449
rect 6847 36385 6911 36449
rect 6927 36385 6991 36449
rect 7007 36385 7071 36449
rect 7087 36385 7151 36449
rect 7167 36385 7231 36449
rect 7247 36385 7311 36449
rect 7327 36385 7391 36449
rect 7407 36385 7471 36449
rect 7487 36385 7551 36449
rect 7567 36385 7631 36449
rect 7647 36385 7711 36449
rect 7727 36385 7791 36449
rect 6607 36304 6671 36368
rect 6687 36304 6751 36368
rect 6767 36304 6831 36368
rect 6847 36304 6911 36368
rect 6927 36304 6991 36368
rect 7007 36304 7071 36368
rect 7087 36304 7151 36368
rect 7167 36304 7231 36368
rect 7247 36304 7311 36368
rect 7327 36304 7391 36368
rect 7407 36304 7471 36368
rect 7487 36304 7551 36368
rect 7567 36304 7631 36368
rect 7647 36304 7711 36368
rect 7727 36304 7791 36368
rect 6607 36223 6671 36287
rect 6687 36223 6751 36287
rect 6767 36223 6831 36287
rect 6847 36223 6911 36287
rect 6927 36223 6991 36287
rect 7007 36223 7071 36287
rect 7087 36223 7151 36287
rect 7167 36223 7231 36287
rect 7247 36223 7311 36287
rect 7327 36223 7391 36287
rect 7407 36223 7471 36287
rect 7487 36223 7551 36287
rect 7567 36223 7631 36287
rect 7647 36223 7711 36287
rect 7727 36223 7791 36287
rect 6607 36142 6671 36206
rect 6687 36142 6751 36206
rect 6767 36142 6831 36206
rect 6847 36142 6911 36206
rect 6927 36142 6991 36206
rect 7007 36142 7071 36206
rect 7087 36142 7151 36206
rect 7167 36142 7231 36206
rect 7247 36142 7311 36206
rect 7327 36142 7391 36206
rect 7407 36142 7471 36206
rect 7487 36142 7551 36206
rect 7567 36142 7631 36206
rect 7647 36142 7711 36206
rect 7727 36142 7791 36206
rect 6607 36060 6671 36124
rect 6687 36060 6751 36124
rect 6767 36060 6831 36124
rect 6847 36060 6911 36124
rect 6927 36060 6991 36124
rect 7007 36060 7071 36124
rect 7087 36060 7151 36124
rect 7167 36060 7231 36124
rect 7247 36060 7311 36124
rect 7327 36060 7391 36124
rect 7407 36060 7471 36124
rect 7487 36060 7551 36124
rect 7567 36060 7631 36124
rect 7647 36060 7711 36124
rect 7727 36060 7791 36124
rect 6607 35978 6671 36042
rect 6687 35978 6751 36042
rect 6767 35978 6831 36042
rect 6847 35978 6911 36042
rect 6927 35978 6991 36042
rect 7007 35978 7071 36042
rect 7087 35978 7151 36042
rect 7167 35978 7231 36042
rect 7247 35978 7311 36042
rect 7327 35978 7391 36042
rect 7407 35978 7471 36042
rect 7487 35978 7551 36042
rect 7567 35978 7631 36042
rect 7647 35978 7711 36042
rect 7727 35978 7791 36042
rect 6607 35896 6671 35960
rect 6687 35896 6751 35960
rect 6767 35896 6831 35960
rect 6847 35896 6911 35960
rect 6927 35896 6991 35960
rect 7007 35896 7071 35960
rect 7087 35896 7151 35960
rect 7167 35896 7231 35960
rect 7247 35896 7311 35960
rect 7327 35896 7391 35960
rect 7407 35896 7471 35960
rect 7487 35896 7551 35960
rect 7567 35896 7631 35960
rect 7647 35896 7711 35960
rect 7727 35896 7791 35960
rect 6607 35814 6671 35878
rect 6687 35814 6751 35878
rect 6767 35814 6831 35878
rect 6847 35814 6911 35878
rect 6927 35814 6991 35878
rect 7007 35814 7071 35878
rect 7087 35814 7151 35878
rect 7167 35814 7231 35878
rect 7247 35814 7311 35878
rect 7327 35814 7391 35878
rect 7407 35814 7471 35878
rect 7487 35814 7551 35878
rect 7567 35814 7631 35878
rect 7647 35814 7711 35878
rect 7727 35814 7791 35878
rect 6607 35732 6671 35796
rect 6687 35732 6751 35796
rect 6767 35732 6831 35796
rect 6847 35732 6911 35796
rect 6927 35732 6991 35796
rect 7007 35732 7071 35796
rect 7087 35732 7151 35796
rect 7167 35732 7231 35796
rect 7247 35732 7311 35796
rect 7327 35732 7391 35796
rect 7407 35732 7471 35796
rect 7487 35732 7551 35796
rect 7567 35732 7631 35796
rect 7647 35732 7711 35796
rect 7727 35732 7791 35796
rect 6607 35650 6671 35714
rect 6687 35650 6751 35714
rect 6767 35650 6831 35714
rect 6847 35650 6911 35714
rect 6927 35650 6991 35714
rect 7007 35650 7071 35714
rect 7087 35650 7151 35714
rect 7167 35650 7231 35714
rect 7247 35650 7311 35714
rect 7327 35650 7391 35714
rect 7407 35650 7471 35714
rect 7487 35650 7551 35714
rect 7567 35650 7631 35714
rect 7647 35650 7711 35714
rect 7727 35650 7791 35714
rect 6607 35568 6671 35632
rect 6687 35568 6751 35632
rect 6767 35568 6831 35632
rect 6847 35568 6911 35632
rect 6927 35568 6991 35632
rect 7007 35568 7071 35632
rect 7087 35568 7151 35632
rect 7167 35568 7231 35632
rect 7247 35568 7311 35632
rect 7327 35568 7391 35632
rect 7407 35568 7471 35632
rect 7487 35568 7551 35632
rect 7567 35568 7631 35632
rect 7647 35568 7711 35632
rect 7727 35568 7791 35632
rect 6607 35486 6671 35550
rect 6687 35486 6751 35550
rect 6767 35486 6831 35550
rect 6847 35486 6911 35550
rect 6927 35486 6991 35550
rect 7007 35486 7071 35550
rect 7087 35486 7151 35550
rect 7167 35486 7231 35550
rect 7247 35486 7311 35550
rect 7327 35486 7391 35550
rect 7407 35486 7471 35550
rect 7487 35486 7551 35550
rect 7567 35486 7631 35550
rect 7647 35486 7711 35550
rect 7727 35486 7791 35550
rect 6607 35404 6671 35468
rect 6687 35404 6751 35468
rect 6767 35404 6831 35468
rect 6847 35404 6911 35468
rect 6927 35404 6991 35468
rect 7007 35404 7071 35468
rect 7087 35404 7151 35468
rect 7167 35404 7231 35468
rect 7247 35404 7311 35468
rect 7327 35404 7391 35468
rect 7407 35404 7471 35468
rect 7487 35404 7551 35468
rect 7567 35404 7631 35468
rect 7647 35404 7711 35468
rect 7727 35404 7791 35468
rect 6607 35322 6671 35386
rect 6687 35322 6751 35386
rect 6767 35322 6831 35386
rect 6847 35322 6911 35386
rect 6927 35322 6991 35386
rect 7007 35322 7071 35386
rect 7087 35322 7151 35386
rect 7167 35322 7231 35386
rect 7247 35322 7311 35386
rect 7327 35322 7391 35386
rect 7407 35322 7471 35386
rect 7487 35322 7551 35386
rect 7567 35322 7631 35386
rect 7647 35322 7711 35386
rect 7727 35322 7791 35386
rect 6607 35240 6671 35304
rect 6687 35240 6751 35304
rect 6767 35240 6831 35304
rect 6847 35240 6911 35304
rect 6927 35240 6991 35304
rect 7007 35240 7071 35304
rect 7087 35240 7151 35304
rect 7167 35240 7231 35304
rect 7247 35240 7311 35304
rect 7327 35240 7391 35304
rect 7407 35240 7471 35304
rect 7487 35240 7551 35304
rect 7567 35240 7631 35304
rect 7647 35240 7711 35304
rect 7727 35240 7791 35304
rect 6607 35158 6671 35222
rect 6687 35158 6751 35222
rect 6767 35158 6831 35222
rect 6847 35158 6911 35222
rect 6927 35158 6991 35222
rect 7007 35158 7071 35222
rect 7087 35158 7151 35222
rect 7167 35158 7231 35222
rect 7247 35158 7311 35222
rect 7327 35158 7391 35222
rect 7407 35158 7471 35222
rect 7487 35158 7551 35222
rect 7567 35158 7631 35222
rect 7647 35158 7711 35222
rect 7727 35158 7791 35222
rect 8100 39301 8164 39365
rect 8180 39301 8244 39365
rect 8260 39301 8324 39365
rect 8340 39301 8404 39365
rect 8420 39301 8484 39365
rect 8500 39301 8564 39365
rect 8580 39301 8644 39365
rect 8660 39301 8724 39365
rect 8740 39301 8804 39365
rect 8820 39301 8884 39365
rect 8900 39301 8964 39365
rect 8980 39301 9044 39365
rect 9060 39301 9124 39365
rect 9140 39301 9204 39365
rect 9220 39301 9284 39365
rect 8100 39220 8164 39284
rect 8180 39220 8244 39284
rect 8260 39220 8324 39284
rect 8340 39220 8404 39284
rect 8420 39220 8484 39284
rect 8500 39220 8564 39284
rect 8580 39220 8644 39284
rect 8660 39220 8724 39284
rect 8740 39220 8804 39284
rect 8820 39220 8884 39284
rect 8900 39220 8964 39284
rect 8980 39220 9044 39284
rect 9060 39220 9124 39284
rect 9140 39220 9204 39284
rect 9220 39220 9284 39284
rect 8100 39139 8164 39203
rect 8180 39139 8244 39203
rect 8260 39139 8324 39203
rect 8340 39139 8404 39203
rect 8420 39139 8484 39203
rect 8500 39139 8564 39203
rect 8580 39139 8644 39203
rect 8660 39139 8724 39203
rect 8740 39139 8804 39203
rect 8820 39139 8884 39203
rect 8900 39139 8964 39203
rect 8980 39139 9044 39203
rect 9060 39139 9124 39203
rect 9140 39139 9204 39203
rect 9220 39139 9284 39203
rect 8100 39058 8164 39122
rect 8180 39058 8244 39122
rect 8260 39058 8324 39122
rect 8340 39058 8404 39122
rect 8420 39058 8484 39122
rect 8500 39058 8564 39122
rect 8580 39058 8644 39122
rect 8660 39058 8724 39122
rect 8740 39058 8804 39122
rect 8820 39058 8884 39122
rect 8900 39058 8964 39122
rect 8980 39058 9044 39122
rect 9060 39058 9124 39122
rect 9140 39058 9204 39122
rect 9220 39058 9284 39122
rect 8100 38977 8164 39041
rect 8180 38977 8244 39041
rect 8260 38977 8324 39041
rect 8340 38977 8404 39041
rect 8420 38977 8484 39041
rect 8500 38977 8564 39041
rect 8580 38977 8644 39041
rect 8660 38977 8724 39041
rect 8740 38977 8804 39041
rect 8820 38977 8884 39041
rect 8900 38977 8964 39041
rect 8980 38977 9044 39041
rect 9060 38977 9124 39041
rect 9140 38977 9204 39041
rect 9220 38977 9284 39041
rect 8100 38896 8164 38960
rect 8180 38896 8244 38960
rect 8260 38896 8324 38960
rect 8340 38896 8404 38960
rect 8420 38896 8484 38960
rect 8500 38896 8564 38960
rect 8580 38896 8644 38960
rect 8660 38896 8724 38960
rect 8740 38896 8804 38960
rect 8820 38896 8884 38960
rect 8900 38896 8964 38960
rect 8980 38896 9044 38960
rect 9060 38896 9124 38960
rect 9140 38896 9204 38960
rect 9220 38896 9284 38960
rect 8100 38815 8164 38879
rect 8180 38815 8244 38879
rect 8260 38815 8324 38879
rect 8340 38815 8404 38879
rect 8420 38815 8484 38879
rect 8500 38815 8564 38879
rect 8580 38815 8644 38879
rect 8660 38815 8724 38879
rect 8740 38815 8804 38879
rect 8820 38815 8884 38879
rect 8900 38815 8964 38879
rect 8980 38815 9044 38879
rect 9060 38815 9124 38879
rect 9140 38815 9204 38879
rect 9220 38815 9284 38879
rect 8100 38734 8164 38798
rect 8180 38734 8244 38798
rect 8260 38734 8324 38798
rect 8340 38734 8404 38798
rect 8420 38734 8484 38798
rect 8500 38734 8564 38798
rect 8580 38734 8644 38798
rect 8660 38734 8724 38798
rect 8740 38734 8804 38798
rect 8820 38734 8884 38798
rect 8900 38734 8964 38798
rect 8980 38734 9044 38798
rect 9060 38734 9124 38798
rect 9140 38734 9204 38798
rect 9220 38734 9284 38798
rect 8100 38653 8164 38717
rect 8180 38653 8244 38717
rect 8260 38653 8324 38717
rect 8340 38653 8404 38717
rect 8420 38653 8484 38717
rect 8500 38653 8564 38717
rect 8580 38653 8644 38717
rect 8660 38653 8724 38717
rect 8740 38653 8804 38717
rect 8820 38653 8884 38717
rect 8900 38653 8964 38717
rect 8980 38653 9044 38717
rect 9060 38653 9124 38717
rect 9140 38653 9204 38717
rect 9220 38653 9284 38717
rect 8100 38572 8164 38636
rect 8180 38572 8244 38636
rect 8260 38572 8324 38636
rect 8340 38572 8404 38636
rect 8420 38572 8484 38636
rect 8500 38572 8564 38636
rect 8580 38572 8644 38636
rect 8660 38572 8724 38636
rect 8740 38572 8804 38636
rect 8820 38572 8884 38636
rect 8900 38572 8964 38636
rect 8980 38572 9044 38636
rect 9060 38572 9124 38636
rect 9140 38572 9204 38636
rect 9220 38572 9284 38636
rect 8100 38491 8164 38555
rect 8180 38491 8244 38555
rect 8260 38491 8324 38555
rect 8340 38491 8404 38555
rect 8420 38491 8484 38555
rect 8500 38491 8564 38555
rect 8580 38491 8644 38555
rect 8660 38491 8724 38555
rect 8740 38491 8804 38555
rect 8820 38491 8884 38555
rect 8900 38491 8964 38555
rect 8980 38491 9044 38555
rect 9060 38491 9124 38555
rect 9140 38491 9204 38555
rect 9220 38491 9284 38555
rect 8100 38410 8164 38474
rect 8180 38410 8244 38474
rect 8260 38410 8324 38474
rect 8340 38410 8404 38474
rect 8420 38410 8484 38474
rect 8500 38410 8564 38474
rect 8580 38410 8644 38474
rect 8660 38410 8724 38474
rect 8740 38410 8804 38474
rect 8820 38410 8884 38474
rect 8900 38410 8964 38474
rect 8980 38410 9044 38474
rect 9060 38410 9124 38474
rect 9140 38410 9204 38474
rect 9220 38410 9284 38474
rect 8100 38329 8164 38393
rect 8180 38329 8244 38393
rect 8260 38329 8324 38393
rect 8340 38329 8404 38393
rect 8420 38329 8484 38393
rect 8500 38329 8564 38393
rect 8580 38329 8644 38393
rect 8660 38329 8724 38393
rect 8740 38329 8804 38393
rect 8820 38329 8884 38393
rect 8900 38329 8964 38393
rect 8980 38329 9044 38393
rect 9060 38329 9124 38393
rect 9140 38329 9204 38393
rect 9220 38329 9284 38393
rect 8100 38248 8164 38312
rect 8180 38248 8244 38312
rect 8260 38248 8324 38312
rect 8340 38248 8404 38312
rect 8420 38248 8484 38312
rect 8500 38248 8564 38312
rect 8580 38248 8644 38312
rect 8660 38248 8724 38312
rect 8740 38248 8804 38312
rect 8820 38248 8884 38312
rect 8900 38248 8964 38312
rect 8980 38248 9044 38312
rect 9060 38248 9124 38312
rect 9140 38248 9204 38312
rect 9220 38248 9284 38312
rect 8100 38167 8164 38231
rect 8180 38167 8244 38231
rect 8260 38167 8324 38231
rect 8340 38167 8404 38231
rect 8420 38167 8484 38231
rect 8500 38167 8564 38231
rect 8580 38167 8644 38231
rect 8660 38167 8724 38231
rect 8740 38167 8804 38231
rect 8820 38167 8884 38231
rect 8900 38167 8964 38231
rect 8980 38167 9044 38231
rect 9060 38167 9124 38231
rect 9140 38167 9204 38231
rect 9220 38167 9284 38231
rect 8100 38086 8164 38150
rect 8180 38086 8244 38150
rect 8260 38086 8324 38150
rect 8340 38086 8404 38150
rect 8420 38086 8484 38150
rect 8500 38086 8564 38150
rect 8580 38086 8644 38150
rect 8660 38086 8724 38150
rect 8740 38086 8804 38150
rect 8820 38086 8884 38150
rect 8900 38086 8964 38150
rect 8980 38086 9044 38150
rect 9060 38086 9124 38150
rect 9140 38086 9204 38150
rect 9220 38086 9284 38150
rect 8100 38005 8164 38069
rect 8180 38005 8244 38069
rect 8260 38005 8324 38069
rect 8340 38005 8404 38069
rect 8420 38005 8484 38069
rect 8500 38005 8564 38069
rect 8580 38005 8644 38069
rect 8660 38005 8724 38069
rect 8740 38005 8804 38069
rect 8820 38005 8884 38069
rect 8900 38005 8964 38069
rect 8980 38005 9044 38069
rect 9060 38005 9124 38069
rect 9140 38005 9204 38069
rect 9220 38005 9284 38069
rect 8100 37924 8164 37988
rect 8180 37924 8244 37988
rect 8260 37924 8324 37988
rect 8340 37924 8404 37988
rect 8420 37924 8484 37988
rect 8500 37924 8564 37988
rect 8580 37924 8644 37988
rect 8660 37924 8724 37988
rect 8740 37924 8804 37988
rect 8820 37924 8884 37988
rect 8900 37924 8964 37988
rect 8980 37924 9044 37988
rect 9060 37924 9124 37988
rect 9140 37924 9204 37988
rect 9220 37924 9284 37988
rect 8100 37843 8164 37907
rect 8180 37843 8244 37907
rect 8260 37843 8324 37907
rect 8340 37843 8404 37907
rect 8420 37843 8484 37907
rect 8500 37843 8564 37907
rect 8580 37843 8644 37907
rect 8660 37843 8724 37907
rect 8740 37843 8804 37907
rect 8820 37843 8884 37907
rect 8900 37843 8964 37907
rect 8980 37843 9044 37907
rect 9060 37843 9124 37907
rect 9140 37843 9204 37907
rect 9220 37843 9284 37907
rect 8100 37762 8164 37826
rect 8180 37762 8244 37826
rect 8260 37762 8324 37826
rect 8340 37762 8404 37826
rect 8420 37762 8484 37826
rect 8500 37762 8564 37826
rect 8580 37762 8644 37826
rect 8660 37762 8724 37826
rect 8740 37762 8804 37826
rect 8820 37762 8884 37826
rect 8900 37762 8964 37826
rect 8980 37762 9044 37826
rect 9060 37762 9124 37826
rect 9140 37762 9204 37826
rect 9220 37762 9284 37826
rect 8100 37681 8164 37745
rect 8180 37681 8244 37745
rect 8260 37681 8324 37745
rect 8340 37681 8404 37745
rect 8420 37681 8484 37745
rect 8500 37681 8564 37745
rect 8580 37681 8644 37745
rect 8660 37681 8724 37745
rect 8740 37681 8804 37745
rect 8820 37681 8884 37745
rect 8900 37681 8964 37745
rect 8980 37681 9044 37745
rect 9060 37681 9124 37745
rect 9140 37681 9204 37745
rect 9220 37681 9284 37745
rect 8100 37600 8164 37664
rect 8180 37600 8244 37664
rect 8260 37600 8324 37664
rect 8340 37600 8404 37664
rect 8420 37600 8484 37664
rect 8500 37600 8564 37664
rect 8580 37600 8644 37664
rect 8660 37600 8724 37664
rect 8740 37600 8804 37664
rect 8820 37600 8884 37664
rect 8900 37600 8964 37664
rect 8980 37600 9044 37664
rect 9060 37600 9124 37664
rect 9140 37600 9204 37664
rect 9220 37600 9284 37664
rect 8100 37519 8164 37583
rect 8180 37519 8244 37583
rect 8260 37519 8324 37583
rect 8340 37519 8404 37583
rect 8420 37519 8484 37583
rect 8500 37519 8564 37583
rect 8580 37519 8644 37583
rect 8660 37519 8724 37583
rect 8740 37519 8804 37583
rect 8820 37519 8884 37583
rect 8900 37519 8964 37583
rect 8980 37519 9044 37583
rect 9060 37519 9124 37583
rect 9140 37519 9204 37583
rect 9220 37519 9284 37583
rect 8100 37438 8164 37502
rect 8180 37438 8244 37502
rect 8260 37438 8324 37502
rect 8340 37438 8404 37502
rect 8420 37438 8484 37502
rect 8500 37438 8564 37502
rect 8580 37438 8644 37502
rect 8660 37438 8724 37502
rect 8740 37438 8804 37502
rect 8820 37438 8884 37502
rect 8900 37438 8964 37502
rect 8980 37438 9044 37502
rect 9060 37438 9124 37502
rect 9140 37438 9204 37502
rect 9220 37438 9284 37502
rect 8100 37357 8164 37421
rect 8180 37357 8244 37421
rect 8260 37357 8324 37421
rect 8340 37357 8404 37421
rect 8420 37357 8484 37421
rect 8500 37357 8564 37421
rect 8580 37357 8644 37421
rect 8660 37357 8724 37421
rect 8740 37357 8804 37421
rect 8820 37357 8884 37421
rect 8900 37357 8964 37421
rect 8980 37357 9044 37421
rect 9060 37357 9124 37421
rect 9140 37357 9204 37421
rect 9220 37357 9284 37421
rect 8100 37276 8164 37340
rect 8180 37276 8244 37340
rect 8260 37276 8324 37340
rect 8340 37276 8404 37340
rect 8420 37276 8484 37340
rect 8500 37276 8564 37340
rect 8580 37276 8644 37340
rect 8660 37276 8724 37340
rect 8740 37276 8804 37340
rect 8820 37276 8884 37340
rect 8900 37276 8964 37340
rect 8980 37276 9044 37340
rect 9060 37276 9124 37340
rect 9140 37276 9204 37340
rect 9220 37276 9284 37340
rect 8100 37195 8164 37259
rect 8180 37195 8244 37259
rect 8260 37195 8324 37259
rect 8340 37195 8404 37259
rect 8420 37195 8484 37259
rect 8500 37195 8564 37259
rect 8580 37195 8644 37259
rect 8660 37195 8724 37259
rect 8740 37195 8804 37259
rect 8820 37195 8884 37259
rect 8900 37195 8964 37259
rect 8980 37195 9044 37259
rect 9060 37195 9124 37259
rect 9140 37195 9204 37259
rect 9220 37195 9284 37259
rect 8100 37114 8164 37178
rect 8180 37114 8244 37178
rect 8260 37114 8324 37178
rect 8340 37114 8404 37178
rect 8420 37114 8484 37178
rect 8500 37114 8564 37178
rect 8580 37114 8644 37178
rect 8660 37114 8724 37178
rect 8740 37114 8804 37178
rect 8820 37114 8884 37178
rect 8900 37114 8964 37178
rect 8980 37114 9044 37178
rect 9060 37114 9124 37178
rect 9140 37114 9204 37178
rect 9220 37114 9284 37178
rect 8100 37033 8164 37097
rect 8180 37033 8244 37097
rect 8260 37033 8324 37097
rect 8340 37033 8404 37097
rect 8420 37033 8484 37097
rect 8500 37033 8564 37097
rect 8580 37033 8644 37097
rect 8660 37033 8724 37097
rect 8740 37033 8804 37097
rect 8820 37033 8884 37097
rect 8900 37033 8964 37097
rect 8980 37033 9044 37097
rect 9060 37033 9124 37097
rect 9140 37033 9204 37097
rect 9220 37033 9284 37097
rect 8100 36952 8164 37016
rect 8180 36952 8244 37016
rect 8260 36952 8324 37016
rect 8340 36952 8404 37016
rect 8420 36952 8484 37016
rect 8500 36952 8564 37016
rect 8580 36952 8644 37016
rect 8660 36952 8724 37016
rect 8740 36952 8804 37016
rect 8820 36952 8884 37016
rect 8900 36952 8964 37016
rect 8980 36952 9044 37016
rect 9060 36952 9124 37016
rect 9140 36952 9204 37016
rect 9220 36952 9284 37016
rect 8100 36871 8164 36935
rect 8180 36871 8244 36935
rect 8260 36871 8324 36935
rect 8340 36871 8404 36935
rect 8420 36871 8484 36935
rect 8500 36871 8564 36935
rect 8580 36871 8644 36935
rect 8660 36871 8724 36935
rect 8740 36871 8804 36935
rect 8820 36871 8884 36935
rect 8900 36871 8964 36935
rect 8980 36871 9044 36935
rect 9060 36871 9124 36935
rect 9140 36871 9204 36935
rect 9220 36871 9284 36935
rect 8100 36790 8164 36854
rect 8180 36790 8244 36854
rect 8260 36790 8324 36854
rect 8340 36790 8404 36854
rect 8420 36790 8484 36854
rect 8500 36790 8564 36854
rect 8580 36790 8644 36854
rect 8660 36790 8724 36854
rect 8740 36790 8804 36854
rect 8820 36790 8884 36854
rect 8900 36790 8964 36854
rect 8980 36790 9044 36854
rect 9060 36790 9124 36854
rect 9140 36790 9204 36854
rect 9220 36790 9284 36854
rect 8100 36709 8164 36773
rect 8180 36709 8244 36773
rect 8260 36709 8324 36773
rect 8340 36709 8404 36773
rect 8420 36709 8484 36773
rect 8500 36709 8564 36773
rect 8580 36709 8644 36773
rect 8660 36709 8724 36773
rect 8740 36709 8804 36773
rect 8820 36709 8884 36773
rect 8900 36709 8964 36773
rect 8980 36709 9044 36773
rect 9060 36709 9124 36773
rect 9140 36709 9204 36773
rect 9220 36709 9284 36773
rect 8100 36628 8164 36692
rect 8180 36628 8244 36692
rect 8260 36628 8324 36692
rect 8340 36628 8404 36692
rect 8420 36628 8484 36692
rect 8500 36628 8564 36692
rect 8580 36628 8644 36692
rect 8660 36628 8724 36692
rect 8740 36628 8804 36692
rect 8820 36628 8884 36692
rect 8900 36628 8964 36692
rect 8980 36628 9044 36692
rect 9060 36628 9124 36692
rect 9140 36628 9204 36692
rect 9220 36628 9284 36692
rect 8100 36547 8164 36611
rect 8180 36547 8244 36611
rect 8260 36547 8324 36611
rect 8340 36547 8404 36611
rect 8420 36547 8484 36611
rect 8500 36547 8564 36611
rect 8580 36547 8644 36611
rect 8660 36547 8724 36611
rect 8740 36547 8804 36611
rect 8820 36547 8884 36611
rect 8900 36547 8964 36611
rect 8980 36547 9044 36611
rect 9060 36547 9124 36611
rect 9140 36547 9204 36611
rect 9220 36547 9284 36611
rect 8100 36466 8164 36530
rect 8180 36466 8244 36530
rect 8260 36466 8324 36530
rect 8340 36466 8404 36530
rect 8420 36466 8484 36530
rect 8500 36466 8564 36530
rect 8580 36466 8644 36530
rect 8660 36466 8724 36530
rect 8740 36466 8804 36530
rect 8820 36466 8884 36530
rect 8900 36466 8964 36530
rect 8980 36466 9044 36530
rect 9060 36466 9124 36530
rect 9140 36466 9204 36530
rect 9220 36466 9284 36530
rect 8100 36385 8164 36449
rect 8180 36385 8244 36449
rect 8260 36385 8324 36449
rect 8340 36385 8404 36449
rect 8420 36385 8484 36449
rect 8500 36385 8564 36449
rect 8580 36385 8644 36449
rect 8660 36385 8724 36449
rect 8740 36385 8804 36449
rect 8820 36385 8884 36449
rect 8900 36385 8964 36449
rect 8980 36385 9044 36449
rect 9060 36385 9124 36449
rect 9140 36385 9204 36449
rect 9220 36385 9284 36449
rect 8100 36304 8164 36368
rect 8180 36304 8244 36368
rect 8260 36304 8324 36368
rect 8340 36304 8404 36368
rect 8420 36304 8484 36368
rect 8500 36304 8564 36368
rect 8580 36304 8644 36368
rect 8660 36304 8724 36368
rect 8740 36304 8804 36368
rect 8820 36304 8884 36368
rect 8900 36304 8964 36368
rect 8980 36304 9044 36368
rect 9060 36304 9124 36368
rect 9140 36304 9204 36368
rect 9220 36304 9284 36368
rect 8100 36223 8164 36287
rect 8180 36223 8244 36287
rect 8260 36223 8324 36287
rect 8340 36223 8404 36287
rect 8420 36223 8484 36287
rect 8500 36223 8564 36287
rect 8580 36223 8644 36287
rect 8660 36223 8724 36287
rect 8740 36223 8804 36287
rect 8820 36223 8884 36287
rect 8900 36223 8964 36287
rect 8980 36223 9044 36287
rect 9060 36223 9124 36287
rect 9140 36223 9204 36287
rect 9220 36223 9284 36287
rect 8100 36142 8164 36206
rect 8180 36142 8244 36206
rect 8260 36142 8324 36206
rect 8340 36142 8404 36206
rect 8420 36142 8484 36206
rect 8500 36142 8564 36206
rect 8580 36142 8644 36206
rect 8660 36142 8724 36206
rect 8740 36142 8804 36206
rect 8820 36142 8884 36206
rect 8900 36142 8964 36206
rect 8980 36142 9044 36206
rect 9060 36142 9124 36206
rect 9140 36142 9204 36206
rect 9220 36142 9284 36206
rect 8100 36060 8164 36124
rect 8180 36060 8244 36124
rect 8260 36060 8324 36124
rect 8340 36060 8404 36124
rect 8420 36060 8484 36124
rect 8500 36060 8564 36124
rect 8580 36060 8644 36124
rect 8660 36060 8724 36124
rect 8740 36060 8804 36124
rect 8820 36060 8884 36124
rect 8900 36060 8964 36124
rect 8980 36060 9044 36124
rect 9060 36060 9124 36124
rect 9140 36060 9204 36124
rect 9220 36060 9284 36124
rect 8100 35978 8164 36042
rect 8180 35978 8244 36042
rect 8260 35978 8324 36042
rect 8340 35978 8404 36042
rect 8420 35978 8484 36042
rect 8500 35978 8564 36042
rect 8580 35978 8644 36042
rect 8660 35978 8724 36042
rect 8740 35978 8804 36042
rect 8820 35978 8884 36042
rect 8900 35978 8964 36042
rect 8980 35978 9044 36042
rect 9060 35978 9124 36042
rect 9140 35978 9204 36042
rect 9220 35978 9284 36042
rect 8100 35896 8164 35960
rect 8180 35896 8244 35960
rect 8260 35896 8324 35960
rect 8340 35896 8404 35960
rect 8420 35896 8484 35960
rect 8500 35896 8564 35960
rect 8580 35896 8644 35960
rect 8660 35896 8724 35960
rect 8740 35896 8804 35960
rect 8820 35896 8884 35960
rect 8900 35896 8964 35960
rect 8980 35896 9044 35960
rect 9060 35896 9124 35960
rect 9140 35896 9204 35960
rect 9220 35896 9284 35960
rect 8100 35814 8164 35878
rect 8180 35814 8244 35878
rect 8260 35814 8324 35878
rect 8340 35814 8404 35878
rect 8420 35814 8484 35878
rect 8500 35814 8564 35878
rect 8580 35814 8644 35878
rect 8660 35814 8724 35878
rect 8740 35814 8804 35878
rect 8820 35814 8884 35878
rect 8900 35814 8964 35878
rect 8980 35814 9044 35878
rect 9060 35814 9124 35878
rect 9140 35814 9204 35878
rect 9220 35814 9284 35878
rect 8100 35732 8164 35796
rect 8180 35732 8244 35796
rect 8260 35732 8324 35796
rect 8340 35732 8404 35796
rect 8420 35732 8484 35796
rect 8500 35732 8564 35796
rect 8580 35732 8644 35796
rect 8660 35732 8724 35796
rect 8740 35732 8804 35796
rect 8820 35732 8884 35796
rect 8900 35732 8964 35796
rect 8980 35732 9044 35796
rect 9060 35732 9124 35796
rect 9140 35732 9204 35796
rect 9220 35732 9284 35796
rect 8100 35650 8164 35714
rect 8180 35650 8244 35714
rect 8260 35650 8324 35714
rect 8340 35650 8404 35714
rect 8420 35650 8484 35714
rect 8500 35650 8564 35714
rect 8580 35650 8644 35714
rect 8660 35650 8724 35714
rect 8740 35650 8804 35714
rect 8820 35650 8884 35714
rect 8900 35650 8964 35714
rect 8980 35650 9044 35714
rect 9060 35650 9124 35714
rect 9140 35650 9204 35714
rect 9220 35650 9284 35714
rect 8100 35568 8164 35632
rect 8180 35568 8244 35632
rect 8260 35568 8324 35632
rect 8340 35568 8404 35632
rect 8420 35568 8484 35632
rect 8500 35568 8564 35632
rect 8580 35568 8644 35632
rect 8660 35568 8724 35632
rect 8740 35568 8804 35632
rect 8820 35568 8884 35632
rect 8900 35568 8964 35632
rect 8980 35568 9044 35632
rect 9060 35568 9124 35632
rect 9140 35568 9204 35632
rect 9220 35568 9284 35632
rect 8100 35486 8164 35550
rect 8180 35486 8244 35550
rect 8260 35486 8324 35550
rect 8340 35486 8404 35550
rect 8420 35486 8484 35550
rect 8500 35486 8564 35550
rect 8580 35486 8644 35550
rect 8660 35486 8724 35550
rect 8740 35486 8804 35550
rect 8820 35486 8884 35550
rect 8900 35486 8964 35550
rect 8980 35486 9044 35550
rect 9060 35486 9124 35550
rect 9140 35486 9204 35550
rect 9220 35486 9284 35550
rect 8100 35404 8164 35468
rect 8180 35404 8244 35468
rect 8260 35404 8324 35468
rect 8340 35404 8404 35468
rect 8420 35404 8484 35468
rect 8500 35404 8564 35468
rect 8580 35404 8644 35468
rect 8660 35404 8724 35468
rect 8740 35404 8804 35468
rect 8820 35404 8884 35468
rect 8900 35404 8964 35468
rect 8980 35404 9044 35468
rect 9060 35404 9124 35468
rect 9140 35404 9204 35468
rect 9220 35404 9284 35468
rect 8100 35322 8164 35386
rect 8180 35322 8244 35386
rect 8260 35322 8324 35386
rect 8340 35322 8404 35386
rect 8420 35322 8484 35386
rect 8500 35322 8564 35386
rect 8580 35322 8644 35386
rect 8660 35322 8724 35386
rect 8740 35322 8804 35386
rect 8820 35322 8884 35386
rect 8900 35322 8964 35386
rect 8980 35322 9044 35386
rect 9060 35322 9124 35386
rect 9140 35322 9204 35386
rect 9220 35322 9284 35386
rect 8100 35240 8164 35304
rect 8180 35240 8244 35304
rect 8260 35240 8324 35304
rect 8340 35240 8404 35304
rect 8420 35240 8484 35304
rect 8500 35240 8564 35304
rect 8580 35240 8644 35304
rect 8660 35240 8724 35304
rect 8740 35240 8804 35304
rect 8820 35240 8884 35304
rect 8900 35240 8964 35304
rect 8980 35240 9044 35304
rect 9060 35240 9124 35304
rect 9140 35240 9204 35304
rect 9220 35240 9284 35304
rect 8100 35158 8164 35222
rect 8180 35158 8244 35222
rect 8260 35158 8324 35222
rect 8340 35158 8404 35222
rect 8420 35158 8484 35222
rect 8500 35158 8564 35222
rect 8580 35158 8644 35222
rect 8660 35158 8724 35222
rect 8740 35158 8804 35222
rect 8820 35158 8884 35222
rect 8900 35158 8964 35222
rect 8980 35158 9044 35222
rect 9060 35158 9124 35222
rect 9140 35158 9204 35222
rect 9220 35158 9284 35222
rect 9597 39301 9661 39365
rect 9677 39301 9741 39365
rect 9757 39301 9821 39365
rect 9837 39301 9901 39365
rect 9917 39301 9981 39365
rect 9997 39301 10061 39365
rect 10077 39301 10141 39365
rect 10157 39301 10221 39365
rect 10237 39301 10301 39365
rect 10317 39301 10381 39365
rect 10397 39301 10461 39365
rect 10477 39301 10541 39365
rect 10557 39301 10621 39365
rect 10637 39301 10701 39365
rect 10717 39301 10781 39365
rect 9597 39220 9661 39284
rect 9677 39220 9741 39284
rect 9757 39220 9821 39284
rect 9837 39220 9901 39284
rect 9917 39220 9981 39284
rect 9997 39220 10061 39284
rect 10077 39220 10141 39284
rect 10157 39220 10221 39284
rect 10237 39220 10301 39284
rect 10317 39220 10381 39284
rect 10397 39220 10461 39284
rect 10477 39220 10541 39284
rect 10557 39220 10621 39284
rect 10637 39220 10701 39284
rect 10717 39220 10781 39284
rect 9597 39139 9661 39203
rect 9677 39139 9741 39203
rect 9757 39139 9821 39203
rect 9837 39139 9901 39203
rect 9917 39139 9981 39203
rect 9997 39139 10061 39203
rect 10077 39139 10141 39203
rect 10157 39139 10221 39203
rect 10237 39139 10301 39203
rect 10317 39139 10381 39203
rect 10397 39139 10461 39203
rect 10477 39139 10541 39203
rect 10557 39139 10621 39203
rect 10637 39139 10701 39203
rect 10717 39139 10781 39203
rect 9597 39058 9661 39122
rect 9677 39058 9741 39122
rect 9757 39058 9821 39122
rect 9837 39058 9901 39122
rect 9917 39058 9981 39122
rect 9997 39058 10061 39122
rect 10077 39058 10141 39122
rect 10157 39058 10221 39122
rect 10237 39058 10301 39122
rect 10317 39058 10381 39122
rect 10397 39058 10461 39122
rect 10477 39058 10541 39122
rect 10557 39058 10621 39122
rect 10637 39058 10701 39122
rect 10717 39058 10781 39122
rect 9597 38977 9661 39041
rect 9677 38977 9741 39041
rect 9757 38977 9821 39041
rect 9837 38977 9901 39041
rect 9917 38977 9981 39041
rect 9997 38977 10061 39041
rect 10077 38977 10141 39041
rect 10157 38977 10221 39041
rect 10237 38977 10301 39041
rect 10317 38977 10381 39041
rect 10397 38977 10461 39041
rect 10477 38977 10541 39041
rect 10557 38977 10621 39041
rect 10637 38977 10701 39041
rect 10717 38977 10781 39041
rect 9597 38896 9661 38960
rect 9677 38896 9741 38960
rect 9757 38896 9821 38960
rect 9837 38896 9901 38960
rect 9917 38896 9981 38960
rect 9997 38896 10061 38960
rect 10077 38896 10141 38960
rect 10157 38896 10221 38960
rect 10237 38896 10301 38960
rect 10317 38896 10381 38960
rect 10397 38896 10461 38960
rect 10477 38896 10541 38960
rect 10557 38896 10621 38960
rect 10637 38896 10701 38960
rect 10717 38896 10781 38960
rect 9597 38815 9661 38879
rect 9677 38815 9741 38879
rect 9757 38815 9821 38879
rect 9837 38815 9901 38879
rect 9917 38815 9981 38879
rect 9997 38815 10061 38879
rect 10077 38815 10141 38879
rect 10157 38815 10221 38879
rect 10237 38815 10301 38879
rect 10317 38815 10381 38879
rect 10397 38815 10461 38879
rect 10477 38815 10541 38879
rect 10557 38815 10621 38879
rect 10637 38815 10701 38879
rect 10717 38815 10781 38879
rect 9597 38734 9661 38798
rect 9677 38734 9741 38798
rect 9757 38734 9821 38798
rect 9837 38734 9901 38798
rect 9917 38734 9981 38798
rect 9997 38734 10061 38798
rect 10077 38734 10141 38798
rect 10157 38734 10221 38798
rect 10237 38734 10301 38798
rect 10317 38734 10381 38798
rect 10397 38734 10461 38798
rect 10477 38734 10541 38798
rect 10557 38734 10621 38798
rect 10637 38734 10701 38798
rect 10717 38734 10781 38798
rect 9597 38653 9661 38717
rect 9677 38653 9741 38717
rect 9757 38653 9821 38717
rect 9837 38653 9901 38717
rect 9917 38653 9981 38717
rect 9997 38653 10061 38717
rect 10077 38653 10141 38717
rect 10157 38653 10221 38717
rect 10237 38653 10301 38717
rect 10317 38653 10381 38717
rect 10397 38653 10461 38717
rect 10477 38653 10541 38717
rect 10557 38653 10621 38717
rect 10637 38653 10701 38717
rect 10717 38653 10781 38717
rect 9597 38572 9661 38636
rect 9677 38572 9741 38636
rect 9757 38572 9821 38636
rect 9837 38572 9901 38636
rect 9917 38572 9981 38636
rect 9997 38572 10061 38636
rect 10077 38572 10141 38636
rect 10157 38572 10221 38636
rect 10237 38572 10301 38636
rect 10317 38572 10381 38636
rect 10397 38572 10461 38636
rect 10477 38572 10541 38636
rect 10557 38572 10621 38636
rect 10637 38572 10701 38636
rect 10717 38572 10781 38636
rect 9597 38491 9661 38555
rect 9677 38491 9741 38555
rect 9757 38491 9821 38555
rect 9837 38491 9901 38555
rect 9917 38491 9981 38555
rect 9997 38491 10061 38555
rect 10077 38491 10141 38555
rect 10157 38491 10221 38555
rect 10237 38491 10301 38555
rect 10317 38491 10381 38555
rect 10397 38491 10461 38555
rect 10477 38491 10541 38555
rect 10557 38491 10621 38555
rect 10637 38491 10701 38555
rect 10717 38491 10781 38555
rect 9597 38410 9661 38474
rect 9677 38410 9741 38474
rect 9757 38410 9821 38474
rect 9837 38410 9901 38474
rect 9917 38410 9981 38474
rect 9997 38410 10061 38474
rect 10077 38410 10141 38474
rect 10157 38410 10221 38474
rect 10237 38410 10301 38474
rect 10317 38410 10381 38474
rect 10397 38410 10461 38474
rect 10477 38410 10541 38474
rect 10557 38410 10621 38474
rect 10637 38410 10701 38474
rect 10717 38410 10781 38474
rect 9597 38329 9661 38393
rect 9677 38329 9741 38393
rect 9757 38329 9821 38393
rect 9837 38329 9901 38393
rect 9917 38329 9981 38393
rect 9997 38329 10061 38393
rect 10077 38329 10141 38393
rect 10157 38329 10221 38393
rect 10237 38329 10301 38393
rect 10317 38329 10381 38393
rect 10397 38329 10461 38393
rect 10477 38329 10541 38393
rect 10557 38329 10621 38393
rect 10637 38329 10701 38393
rect 10717 38329 10781 38393
rect 9597 38248 9661 38312
rect 9677 38248 9741 38312
rect 9757 38248 9821 38312
rect 9837 38248 9901 38312
rect 9917 38248 9981 38312
rect 9997 38248 10061 38312
rect 10077 38248 10141 38312
rect 10157 38248 10221 38312
rect 10237 38248 10301 38312
rect 10317 38248 10381 38312
rect 10397 38248 10461 38312
rect 10477 38248 10541 38312
rect 10557 38248 10621 38312
rect 10637 38248 10701 38312
rect 10717 38248 10781 38312
rect 9597 38167 9661 38231
rect 9677 38167 9741 38231
rect 9757 38167 9821 38231
rect 9837 38167 9901 38231
rect 9917 38167 9981 38231
rect 9997 38167 10061 38231
rect 10077 38167 10141 38231
rect 10157 38167 10221 38231
rect 10237 38167 10301 38231
rect 10317 38167 10381 38231
rect 10397 38167 10461 38231
rect 10477 38167 10541 38231
rect 10557 38167 10621 38231
rect 10637 38167 10701 38231
rect 10717 38167 10781 38231
rect 9597 38086 9661 38150
rect 9677 38086 9741 38150
rect 9757 38086 9821 38150
rect 9837 38086 9901 38150
rect 9917 38086 9981 38150
rect 9997 38086 10061 38150
rect 10077 38086 10141 38150
rect 10157 38086 10221 38150
rect 10237 38086 10301 38150
rect 10317 38086 10381 38150
rect 10397 38086 10461 38150
rect 10477 38086 10541 38150
rect 10557 38086 10621 38150
rect 10637 38086 10701 38150
rect 10717 38086 10781 38150
rect 9597 38005 9661 38069
rect 9677 38005 9741 38069
rect 9757 38005 9821 38069
rect 9837 38005 9901 38069
rect 9917 38005 9981 38069
rect 9997 38005 10061 38069
rect 10077 38005 10141 38069
rect 10157 38005 10221 38069
rect 10237 38005 10301 38069
rect 10317 38005 10381 38069
rect 10397 38005 10461 38069
rect 10477 38005 10541 38069
rect 10557 38005 10621 38069
rect 10637 38005 10701 38069
rect 10717 38005 10781 38069
rect 9597 37924 9661 37988
rect 9677 37924 9741 37988
rect 9757 37924 9821 37988
rect 9837 37924 9901 37988
rect 9917 37924 9981 37988
rect 9997 37924 10061 37988
rect 10077 37924 10141 37988
rect 10157 37924 10221 37988
rect 10237 37924 10301 37988
rect 10317 37924 10381 37988
rect 10397 37924 10461 37988
rect 10477 37924 10541 37988
rect 10557 37924 10621 37988
rect 10637 37924 10701 37988
rect 10717 37924 10781 37988
rect 9597 37843 9661 37907
rect 9677 37843 9741 37907
rect 9757 37843 9821 37907
rect 9837 37843 9901 37907
rect 9917 37843 9981 37907
rect 9997 37843 10061 37907
rect 10077 37843 10141 37907
rect 10157 37843 10221 37907
rect 10237 37843 10301 37907
rect 10317 37843 10381 37907
rect 10397 37843 10461 37907
rect 10477 37843 10541 37907
rect 10557 37843 10621 37907
rect 10637 37843 10701 37907
rect 10717 37843 10781 37907
rect 9597 37762 9661 37826
rect 9677 37762 9741 37826
rect 9757 37762 9821 37826
rect 9837 37762 9901 37826
rect 9917 37762 9981 37826
rect 9997 37762 10061 37826
rect 10077 37762 10141 37826
rect 10157 37762 10221 37826
rect 10237 37762 10301 37826
rect 10317 37762 10381 37826
rect 10397 37762 10461 37826
rect 10477 37762 10541 37826
rect 10557 37762 10621 37826
rect 10637 37762 10701 37826
rect 10717 37762 10781 37826
rect 9597 37681 9661 37745
rect 9677 37681 9741 37745
rect 9757 37681 9821 37745
rect 9837 37681 9901 37745
rect 9917 37681 9981 37745
rect 9997 37681 10061 37745
rect 10077 37681 10141 37745
rect 10157 37681 10221 37745
rect 10237 37681 10301 37745
rect 10317 37681 10381 37745
rect 10397 37681 10461 37745
rect 10477 37681 10541 37745
rect 10557 37681 10621 37745
rect 10637 37681 10701 37745
rect 10717 37681 10781 37745
rect 9597 37600 9661 37664
rect 9677 37600 9741 37664
rect 9757 37600 9821 37664
rect 9837 37600 9901 37664
rect 9917 37600 9981 37664
rect 9997 37600 10061 37664
rect 10077 37600 10141 37664
rect 10157 37600 10221 37664
rect 10237 37600 10301 37664
rect 10317 37600 10381 37664
rect 10397 37600 10461 37664
rect 10477 37600 10541 37664
rect 10557 37600 10621 37664
rect 10637 37600 10701 37664
rect 10717 37600 10781 37664
rect 9597 37519 9661 37583
rect 9677 37519 9741 37583
rect 9757 37519 9821 37583
rect 9837 37519 9901 37583
rect 9917 37519 9981 37583
rect 9997 37519 10061 37583
rect 10077 37519 10141 37583
rect 10157 37519 10221 37583
rect 10237 37519 10301 37583
rect 10317 37519 10381 37583
rect 10397 37519 10461 37583
rect 10477 37519 10541 37583
rect 10557 37519 10621 37583
rect 10637 37519 10701 37583
rect 10717 37519 10781 37583
rect 9597 37438 9661 37502
rect 9677 37438 9741 37502
rect 9757 37438 9821 37502
rect 9837 37438 9901 37502
rect 9917 37438 9981 37502
rect 9997 37438 10061 37502
rect 10077 37438 10141 37502
rect 10157 37438 10221 37502
rect 10237 37438 10301 37502
rect 10317 37438 10381 37502
rect 10397 37438 10461 37502
rect 10477 37438 10541 37502
rect 10557 37438 10621 37502
rect 10637 37438 10701 37502
rect 10717 37438 10781 37502
rect 9597 37357 9661 37421
rect 9677 37357 9741 37421
rect 9757 37357 9821 37421
rect 9837 37357 9901 37421
rect 9917 37357 9981 37421
rect 9997 37357 10061 37421
rect 10077 37357 10141 37421
rect 10157 37357 10221 37421
rect 10237 37357 10301 37421
rect 10317 37357 10381 37421
rect 10397 37357 10461 37421
rect 10477 37357 10541 37421
rect 10557 37357 10621 37421
rect 10637 37357 10701 37421
rect 10717 37357 10781 37421
rect 9597 37276 9661 37340
rect 9677 37276 9741 37340
rect 9757 37276 9821 37340
rect 9837 37276 9901 37340
rect 9917 37276 9981 37340
rect 9997 37276 10061 37340
rect 10077 37276 10141 37340
rect 10157 37276 10221 37340
rect 10237 37276 10301 37340
rect 10317 37276 10381 37340
rect 10397 37276 10461 37340
rect 10477 37276 10541 37340
rect 10557 37276 10621 37340
rect 10637 37276 10701 37340
rect 10717 37276 10781 37340
rect 9597 37195 9661 37259
rect 9677 37195 9741 37259
rect 9757 37195 9821 37259
rect 9837 37195 9901 37259
rect 9917 37195 9981 37259
rect 9997 37195 10061 37259
rect 10077 37195 10141 37259
rect 10157 37195 10221 37259
rect 10237 37195 10301 37259
rect 10317 37195 10381 37259
rect 10397 37195 10461 37259
rect 10477 37195 10541 37259
rect 10557 37195 10621 37259
rect 10637 37195 10701 37259
rect 10717 37195 10781 37259
rect 9597 37114 9661 37178
rect 9677 37114 9741 37178
rect 9757 37114 9821 37178
rect 9837 37114 9901 37178
rect 9917 37114 9981 37178
rect 9997 37114 10061 37178
rect 10077 37114 10141 37178
rect 10157 37114 10221 37178
rect 10237 37114 10301 37178
rect 10317 37114 10381 37178
rect 10397 37114 10461 37178
rect 10477 37114 10541 37178
rect 10557 37114 10621 37178
rect 10637 37114 10701 37178
rect 10717 37114 10781 37178
rect 9597 37033 9661 37097
rect 9677 37033 9741 37097
rect 9757 37033 9821 37097
rect 9837 37033 9901 37097
rect 9917 37033 9981 37097
rect 9997 37033 10061 37097
rect 10077 37033 10141 37097
rect 10157 37033 10221 37097
rect 10237 37033 10301 37097
rect 10317 37033 10381 37097
rect 10397 37033 10461 37097
rect 10477 37033 10541 37097
rect 10557 37033 10621 37097
rect 10637 37033 10701 37097
rect 10717 37033 10781 37097
rect 9597 36952 9661 37016
rect 9677 36952 9741 37016
rect 9757 36952 9821 37016
rect 9837 36952 9901 37016
rect 9917 36952 9981 37016
rect 9997 36952 10061 37016
rect 10077 36952 10141 37016
rect 10157 36952 10221 37016
rect 10237 36952 10301 37016
rect 10317 36952 10381 37016
rect 10397 36952 10461 37016
rect 10477 36952 10541 37016
rect 10557 36952 10621 37016
rect 10637 36952 10701 37016
rect 10717 36952 10781 37016
rect 9597 36871 9661 36935
rect 9677 36871 9741 36935
rect 9757 36871 9821 36935
rect 9837 36871 9901 36935
rect 9917 36871 9981 36935
rect 9997 36871 10061 36935
rect 10077 36871 10141 36935
rect 10157 36871 10221 36935
rect 10237 36871 10301 36935
rect 10317 36871 10381 36935
rect 10397 36871 10461 36935
rect 10477 36871 10541 36935
rect 10557 36871 10621 36935
rect 10637 36871 10701 36935
rect 10717 36871 10781 36935
rect 9597 36790 9661 36854
rect 9677 36790 9741 36854
rect 9757 36790 9821 36854
rect 9837 36790 9901 36854
rect 9917 36790 9981 36854
rect 9997 36790 10061 36854
rect 10077 36790 10141 36854
rect 10157 36790 10221 36854
rect 10237 36790 10301 36854
rect 10317 36790 10381 36854
rect 10397 36790 10461 36854
rect 10477 36790 10541 36854
rect 10557 36790 10621 36854
rect 10637 36790 10701 36854
rect 10717 36790 10781 36854
rect 9597 36709 9661 36773
rect 9677 36709 9741 36773
rect 9757 36709 9821 36773
rect 9837 36709 9901 36773
rect 9917 36709 9981 36773
rect 9997 36709 10061 36773
rect 10077 36709 10141 36773
rect 10157 36709 10221 36773
rect 10237 36709 10301 36773
rect 10317 36709 10381 36773
rect 10397 36709 10461 36773
rect 10477 36709 10541 36773
rect 10557 36709 10621 36773
rect 10637 36709 10701 36773
rect 10717 36709 10781 36773
rect 9597 36628 9661 36692
rect 9677 36628 9741 36692
rect 9757 36628 9821 36692
rect 9837 36628 9901 36692
rect 9917 36628 9981 36692
rect 9997 36628 10061 36692
rect 10077 36628 10141 36692
rect 10157 36628 10221 36692
rect 10237 36628 10301 36692
rect 10317 36628 10381 36692
rect 10397 36628 10461 36692
rect 10477 36628 10541 36692
rect 10557 36628 10621 36692
rect 10637 36628 10701 36692
rect 10717 36628 10781 36692
rect 9597 36547 9661 36611
rect 9677 36547 9741 36611
rect 9757 36547 9821 36611
rect 9837 36547 9901 36611
rect 9917 36547 9981 36611
rect 9997 36547 10061 36611
rect 10077 36547 10141 36611
rect 10157 36547 10221 36611
rect 10237 36547 10301 36611
rect 10317 36547 10381 36611
rect 10397 36547 10461 36611
rect 10477 36547 10541 36611
rect 10557 36547 10621 36611
rect 10637 36547 10701 36611
rect 10717 36547 10781 36611
rect 9597 36466 9661 36530
rect 9677 36466 9741 36530
rect 9757 36466 9821 36530
rect 9837 36466 9901 36530
rect 9917 36466 9981 36530
rect 9997 36466 10061 36530
rect 10077 36466 10141 36530
rect 10157 36466 10221 36530
rect 10237 36466 10301 36530
rect 10317 36466 10381 36530
rect 10397 36466 10461 36530
rect 10477 36466 10541 36530
rect 10557 36466 10621 36530
rect 10637 36466 10701 36530
rect 10717 36466 10781 36530
rect 9597 36385 9661 36449
rect 9677 36385 9741 36449
rect 9757 36385 9821 36449
rect 9837 36385 9901 36449
rect 9917 36385 9981 36449
rect 9997 36385 10061 36449
rect 10077 36385 10141 36449
rect 10157 36385 10221 36449
rect 10237 36385 10301 36449
rect 10317 36385 10381 36449
rect 10397 36385 10461 36449
rect 10477 36385 10541 36449
rect 10557 36385 10621 36449
rect 10637 36385 10701 36449
rect 10717 36385 10781 36449
rect 9597 36304 9661 36368
rect 9677 36304 9741 36368
rect 9757 36304 9821 36368
rect 9837 36304 9901 36368
rect 9917 36304 9981 36368
rect 9997 36304 10061 36368
rect 10077 36304 10141 36368
rect 10157 36304 10221 36368
rect 10237 36304 10301 36368
rect 10317 36304 10381 36368
rect 10397 36304 10461 36368
rect 10477 36304 10541 36368
rect 10557 36304 10621 36368
rect 10637 36304 10701 36368
rect 10717 36304 10781 36368
rect 9597 36223 9661 36287
rect 9677 36223 9741 36287
rect 9757 36223 9821 36287
rect 9837 36223 9901 36287
rect 9917 36223 9981 36287
rect 9997 36223 10061 36287
rect 10077 36223 10141 36287
rect 10157 36223 10221 36287
rect 10237 36223 10301 36287
rect 10317 36223 10381 36287
rect 10397 36223 10461 36287
rect 10477 36223 10541 36287
rect 10557 36223 10621 36287
rect 10637 36223 10701 36287
rect 10717 36223 10781 36287
rect 9597 36142 9661 36206
rect 9677 36142 9741 36206
rect 9757 36142 9821 36206
rect 9837 36142 9901 36206
rect 9917 36142 9981 36206
rect 9997 36142 10061 36206
rect 10077 36142 10141 36206
rect 10157 36142 10221 36206
rect 10237 36142 10301 36206
rect 10317 36142 10381 36206
rect 10397 36142 10461 36206
rect 10477 36142 10541 36206
rect 10557 36142 10621 36206
rect 10637 36142 10701 36206
rect 10717 36142 10781 36206
rect 9597 36060 9661 36124
rect 9677 36060 9741 36124
rect 9757 36060 9821 36124
rect 9837 36060 9901 36124
rect 9917 36060 9981 36124
rect 9997 36060 10061 36124
rect 10077 36060 10141 36124
rect 10157 36060 10221 36124
rect 10237 36060 10301 36124
rect 10317 36060 10381 36124
rect 10397 36060 10461 36124
rect 10477 36060 10541 36124
rect 10557 36060 10621 36124
rect 10637 36060 10701 36124
rect 10717 36060 10781 36124
rect 9597 35978 9661 36042
rect 9677 35978 9741 36042
rect 9757 35978 9821 36042
rect 9837 35978 9901 36042
rect 9917 35978 9981 36042
rect 9997 35978 10061 36042
rect 10077 35978 10141 36042
rect 10157 35978 10221 36042
rect 10237 35978 10301 36042
rect 10317 35978 10381 36042
rect 10397 35978 10461 36042
rect 10477 35978 10541 36042
rect 10557 35978 10621 36042
rect 10637 35978 10701 36042
rect 10717 35978 10781 36042
rect 9597 35896 9661 35960
rect 9677 35896 9741 35960
rect 9757 35896 9821 35960
rect 9837 35896 9901 35960
rect 9917 35896 9981 35960
rect 9997 35896 10061 35960
rect 10077 35896 10141 35960
rect 10157 35896 10221 35960
rect 10237 35896 10301 35960
rect 10317 35896 10381 35960
rect 10397 35896 10461 35960
rect 10477 35896 10541 35960
rect 10557 35896 10621 35960
rect 10637 35896 10701 35960
rect 10717 35896 10781 35960
rect 9597 35814 9661 35878
rect 9677 35814 9741 35878
rect 9757 35814 9821 35878
rect 9837 35814 9901 35878
rect 9917 35814 9981 35878
rect 9997 35814 10061 35878
rect 10077 35814 10141 35878
rect 10157 35814 10221 35878
rect 10237 35814 10301 35878
rect 10317 35814 10381 35878
rect 10397 35814 10461 35878
rect 10477 35814 10541 35878
rect 10557 35814 10621 35878
rect 10637 35814 10701 35878
rect 10717 35814 10781 35878
rect 9597 35732 9661 35796
rect 9677 35732 9741 35796
rect 9757 35732 9821 35796
rect 9837 35732 9901 35796
rect 9917 35732 9981 35796
rect 9997 35732 10061 35796
rect 10077 35732 10141 35796
rect 10157 35732 10221 35796
rect 10237 35732 10301 35796
rect 10317 35732 10381 35796
rect 10397 35732 10461 35796
rect 10477 35732 10541 35796
rect 10557 35732 10621 35796
rect 10637 35732 10701 35796
rect 10717 35732 10781 35796
rect 9597 35650 9661 35714
rect 9677 35650 9741 35714
rect 9757 35650 9821 35714
rect 9837 35650 9901 35714
rect 9917 35650 9981 35714
rect 9997 35650 10061 35714
rect 10077 35650 10141 35714
rect 10157 35650 10221 35714
rect 10237 35650 10301 35714
rect 10317 35650 10381 35714
rect 10397 35650 10461 35714
rect 10477 35650 10541 35714
rect 10557 35650 10621 35714
rect 10637 35650 10701 35714
rect 10717 35650 10781 35714
rect 9597 35568 9661 35632
rect 9677 35568 9741 35632
rect 9757 35568 9821 35632
rect 9837 35568 9901 35632
rect 9917 35568 9981 35632
rect 9997 35568 10061 35632
rect 10077 35568 10141 35632
rect 10157 35568 10221 35632
rect 10237 35568 10301 35632
rect 10317 35568 10381 35632
rect 10397 35568 10461 35632
rect 10477 35568 10541 35632
rect 10557 35568 10621 35632
rect 10637 35568 10701 35632
rect 10717 35568 10781 35632
rect 9597 35486 9661 35550
rect 9677 35486 9741 35550
rect 9757 35486 9821 35550
rect 9837 35486 9901 35550
rect 9917 35486 9981 35550
rect 9997 35486 10061 35550
rect 10077 35486 10141 35550
rect 10157 35486 10221 35550
rect 10237 35486 10301 35550
rect 10317 35486 10381 35550
rect 10397 35486 10461 35550
rect 10477 35486 10541 35550
rect 10557 35486 10621 35550
rect 10637 35486 10701 35550
rect 10717 35486 10781 35550
rect 9597 35404 9661 35468
rect 9677 35404 9741 35468
rect 9757 35404 9821 35468
rect 9837 35404 9901 35468
rect 9917 35404 9981 35468
rect 9997 35404 10061 35468
rect 10077 35404 10141 35468
rect 10157 35404 10221 35468
rect 10237 35404 10301 35468
rect 10317 35404 10381 35468
rect 10397 35404 10461 35468
rect 10477 35404 10541 35468
rect 10557 35404 10621 35468
rect 10637 35404 10701 35468
rect 10717 35404 10781 35468
rect 9597 35322 9661 35386
rect 9677 35322 9741 35386
rect 9757 35322 9821 35386
rect 9837 35322 9901 35386
rect 9917 35322 9981 35386
rect 9997 35322 10061 35386
rect 10077 35322 10141 35386
rect 10157 35322 10221 35386
rect 10237 35322 10301 35386
rect 10317 35322 10381 35386
rect 10397 35322 10461 35386
rect 10477 35322 10541 35386
rect 10557 35322 10621 35386
rect 10637 35322 10701 35386
rect 10717 35322 10781 35386
rect 9597 35240 9661 35304
rect 9677 35240 9741 35304
rect 9757 35240 9821 35304
rect 9837 35240 9901 35304
rect 9917 35240 9981 35304
rect 9997 35240 10061 35304
rect 10077 35240 10141 35304
rect 10157 35240 10221 35304
rect 10237 35240 10301 35304
rect 10317 35240 10381 35304
rect 10397 35240 10461 35304
rect 10477 35240 10541 35304
rect 10557 35240 10621 35304
rect 10637 35240 10701 35304
rect 10717 35240 10781 35304
rect 9597 35158 9661 35222
rect 9677 35158 9741 35222
rect 9757 35158 9821 35222
rect 9837 35158 9901 35222
rect 9917 35158 9981 35222
rect 9997 35158 10061 35222
rect 10077 35158 10141 35222
rect 10157 35158 10221 35222
rect 10237 35158 10301 35222
rect 10317 35158 10381 35222
rect 10397 35158 10461 35222
rect 10477 35158 10541 35222
rect 10557 35158 10621 35222
rect 10637 35158 10701 35222
rect 10717 35158 10781 35222
rect 11098 39301 11162 39365
rect 11178 39301 11242 39365
rect 11258 39301 11322 39365
rect 11338 39301 11402 39365
rect 11418 39301 11482 39365
rect 11498 39301 11562 39365
rect 11578 39301 11642 39365
rect 11658 39301 11722 39365
rect 11738 39301 11802 39365
rect 11818 39301 11882 39365
rect 11898 39301 11962 39365
rect 11978 39301 12042 39365
rect 12058 39301 12122 39365
rect 12138 39301 12202 39365
rect 12218 39301 12282 39365
rect 11098 39220 11162 39284
rect 11178 39220 11242 39284
rect 11258 39220 11322 39284
rect 11338 39220 11402 39284
rect 11418 39220 11482 39284
rect 11498 39220 11562 39284
rect 11578 39220 11642 39284
rect 11658 39220 11722 39284
rect 11738 39220 11802 39284
rect 11818 39220 11882 39284
rect 11898 39220 11962 39284
rect 11978 39220 12042 39284
rect 12058 39220 12122 39284
rect 12138 39220 12202 39284
rect 12218 39220 12282 39284
rect 11098 39139 11162 39203
rect 11178 39139 11242 39203
rect 11258 39139 11322 39203
rect 11338 39139 11402 39203
rect 11418 39139 11482 39203
rect 11498 39139 11562 39203
rect 11578 39139 11642 39203
rect 11658 39139 11722 39203
rect 11738 39139 11802 39203
rect 11818 39139 11882 39203
rect 11898 39139 11962 39203
rect 11978 39139 12042 39203
rect 12058 39139 12122 39203
rect 12138 39139 12202 39203
rect 12218 39139 12282 39203
rect 11098 39058 11162 39122
rect 11178 39058 11242 39122
rect 11258 39058 11322 39122
rect 11338 39058 11402 39122
rect 11418 39058 11482 39122
rect 11498 39058 11562 39122
rect 11578 39058 11642 39122
rect 11658 39058 11722 39122
rect 11738 39058 11802 39122
rect 11818 39058 11882 39122
rect 11898 39058 11962 39122
rect 11978 39058 12042 39122
rect 12058 39058 12122 39122
rect 12138 39058 12202 39122
rect 12218 39058 12282 39122
rect 11098 38977 11162 39041
rect 11178 38977 11242 39041
rect 11258 38977 11322 39041
rect 11338 38977 11402 39041
rect 11418 38977 11482 39041
rect 11498 38977 11562 39041
rect 11578 38977 11642 39041
rect 11658 38977 11722 39041
rect 11738 38977 11802 39041
rect 11818 38977 11882 39041
rect 11898 38977 11962 39041
rect 11978 38977 12042 39041
rect 12058 38977 12122 39041
rect 12138 38977 12202 39041
rect 12218 38977 12282 39041
rect 11098 38896 11162 38960
rect 11178 38896 11242 38960
rect 11258 38896 11322 38960
rect 11338 38896 11402 38960
rect 11418 38896 11482 38960
rect 11498 38896 11562 38960
rect 11578 38896 11642 38960
rect 11658 38896 11722 38960
rect 11738 38896 11802 38960
rect 11818 38896 11882 38960
rect 11898 38896 11962 38960
rect 11978 38896 12042 38960
rect 12058 38896 12122 38960
rect 12138 38896 12202 38960
rect 12218 38896 12282 38960
rect 11098 38815 11162 38879
rect 11178 38815 11242 38879
rect 11258 38815 11322 38879
rect 11338 38815 11402 38879
rect 11418 38815 11482 38879
rect 11498 38815 11562 38879
rect 11578 38815 11642 38879
rect 11658 38815 11722 38879
rect 11738 38815 11802 38879
rect 11818 38815 11882 38879
rect 11898 38815 11962 38879
rect 11978 38815 12042 38879
rect 12058 38815 12122 38879
rect 12138 38815 12202 38879
rect 12218 38815 12282 38879
rect 11098 38734 11162 38798
rect 11178 38734 11242 38798
rect 11258 38734 11322 38798
rect 11338 38734 11402 38798
rect 11418 38734 11482 38798
rect 11498 38734 11562 38798
rect 11578 38734 11642 38798
rect 11658 38734 11722 38798
rect 11738 38734 11802 38798
rect 11818 38734 11882 38798
rect 11898 38734 11962 38798
rect 11978 38734 12042 38798
rect 12058 38734 12122 38798
rect 12138 38734 12202 38798
rect 12218 38734 12282 38798
rect 11098 38653 11162 38717
rect 11178 38653 11242 38717
rect 11258 38653 11322 38717
rect 11338 38653 11402 38717
rect 11418 38653 11482 38717
rect 11498 38653 11562 38717
rect 11578 38653 11642 38717
rect 11658 38653 11722 38717
rect 11738 38653 11802 38717
rect 11818 38653 11882 38717
rect 11898 38653 11962 38717
rect 11978 38653 12042 38717
rect 12058 38653 12122 38717
rect 12138 38653 12202 38717
rect 12218 38653 12282 38717
rect 11098 38572 11162 38636
rect 11178 38572 11242 38636
rect 11258 38572 11322 38636
rect 11338 38572 11402 38636
rect 11418 38572 11482 38636
rect 11498 38572 11562 38636
rect 11578 38572 11642 38636
rect 11658 38572 11722 38636
rect 11738 38572 11802 38636
rect 11818 38572 11882 38636
rect 11898 38572 11962 38636
rect 11978 38572 12042 38636
rect 12058 38572 12122 38636
rect 12138 38572 12202 38636
rect 12218 38572 12282 38636
rect 11098 38491 11162 38555
rect 11178 38491 11242 38555
rect 11258 38491 11322 38555
rect 11338 38491 11402 38555
rect 11418 38491 11482 38555
rect 11498 38491 11562 38555
rect 11578 38491 11642 38555
rect 11658 38491 11722 38555
rect 11738 38491 11802 38555
rect 11818 38491 11882 38555
rect 11898 38491 11962 38555
rect 11978 38491 12042 38555
rect 12058 38491 12122 38555
rect 12138 38491 12202 38555
rect 12218 38491 12282 38555
rect 11098 38410 11162 38474
rect 11178 38410 11242 38474
rect 11258 38410 11322 38474
rect 11338 38410 11402 38474
rect 11418 38410 11482 38474
rect 11498 38410 11562 38474
rect 11578 38410 11642 38474
rect 11658 38410 11722 38474
rect 11738 38410 11802 38474
rect 11818 38410 11882 38474
rect 11898 38410 11962 38474
rect 11978 38410 12042 38474
rect 12058 38410 12122 38474
rect 12138 38410 12202 38474
rect 12218 38410 12282 38474
rect 11098 38329 11162 38393
rect 11178 38329 11242 38393
rect 11258 38329 11322 38393
rect 11338 38329 11402 38393
rect 11418 38329 11482 38393
rect 11498 38329 11562 38393
rect 11578 38329 11642 38393
rect 11658 38329 11722 38393
rect 11738 38329 11802 38393
rect 11818 38329 11882 38393
rect 11898 38329 11962 38393
rect 11978 38329 12042 38393
rect 12058 38329 12122 38393
rect 12138 38329 12202 38393
rect 12218 38329 12282 38393
rect 11098 38248 11162 38312
rect 11178 38248 11242 38312
rect 11258 38248 11322 38312
rect 11338 38248 11402 38312
rect 11418 38248 11482 38312
rect 11498 38248 11562 38312
rect 11578 38248 11642 38312
rect 11658 38248 11722 38312
rect 11738 38248 11802 38312
rect 11818 38248 11882 38312
rect 11898 38248 11962 38312
rect 11978 38248 12042 38312
rect 12058 38248 12122 38312
rect 12138 38248 12202 38312
rect 12218 38248 12282 38312
rect 11098 38167 11162 38231
rect 11178 38167 11242 38231
rect 11258 38167 11322 38231
rect 11338 38167 11402 38231
rect 11418 38167 11482 38231
rect 11498 38167 11562 38231
rect 11578 38167 11642 38231
rect 11658 38167 11722 38231
rect 11738 38167 11802 38231
rect 11818 38167 11882 38231
rect 11898 38167 11962 38231
rect 11978 38167 12042 38231
rect 12058 38167 12122 38231
rect 12138 38167 12202 38231
rect 12218 38167 12282 38231
rect 11098 38086 11162 38150
rect 11178 38086 11242 38150
rect 11258 38086 11322 38150
rect 11338 38086 11402 38150
rect 11418 38086 11482 38150
rect 11498 38086 11562 38150
rect 11578 38086 11642 38150
rect 11658 38086 11722 38150
rect 11738 38086 11802 38150
rect 11818 38086 11882 38150
rect 11898 38086 11962 38150
rect 11978 38086 12042 38150
rect 12058 38086 12122 38150
rect 12138 38086 12202 38150
rect 12218 38086 12282 38150
rect 11098 38005 11162 38069
rect 11178 38005 11242 38069
rect 11258 38005 11322 38069
rect 11338 38005 11402 38069
rect 11418 38005 11482 38069
rect 11498 38005 11562 38069
rect 11578 38005 11642 38069
rect 11658 38005 11722 38069
rect 11738 38005 11802 38069
rect 11818 38005 11882 38069
rect 11898 38005 11962 38069
rect 11978 38005 12042 38069
rect 12058 38005 12122 38069
rect 12138 38005 12202 38069
rect 12218 38005 12282 38069
rect 11098 37924 11162 37988
rect 11178 37924 11242 37988
rect 11258 37924 11322 37988
rect 11338 37924 11402 37988
rect 11418 37924 11482 37988
rect 11498 37924 11562 37988
rect 11578 37924 11642 37988
rect 11658 37924 11722 37988
rect 11738 37924 11802 37988
rect 11818 37924 11882 37988
rect 11898 37924 11962 37988
rect 11978 37924 12042 37988
rect 12058 37924 12122 37988
rect 12138 37924 12202 37988
rect 12218 37924 12282 37988
rect 11098 37843 11162 37907
rect 11178 37843 11242 37907
rect 11258 37843 11322 37907
rect 11338 37843 11402 37907
rect 11418 37843 11482 37907
rect 11498 37843 11562 37907
rect 11578 37843 11642 37907
rect 11658 37843 11722 37907
rect 11738 37843 11802 37907
rect 11818 37843 11882 37907
rect 11898 37843 11962 37907
rect 11978 37843 12042 37907
rect 12058 37843 12122 37907
rect 12138 37843 12202 37907
rect 12218 37843 12282 37907
rect 11098 37762 11162 37826
rect 11178 37762 11242 37826
rect 11258 37762 11322 37826
rect 11338 37762 11402 37826
rect 11418 37762 11482 37826
rect 11498 37762 11562 37826
rect 11578 37762 11642 37826
rect 11658 37762 11722 37826
rect 11738 37762 11802 37826
rect 11818 37762 11882 37826
rect 11898 37762 11962 37826
rect 11978 37762 12042 37826
rect 12058 37762 12122 37826
rect 12138 37762 12202 37826
rect 12218 37762 12282 37826
rect 11098 37681 11162 37745
rect 11178 37681 11242 37745
rect 11258 37681 11322 37745
rect 11338 37681 11402 37745
rect 11418 37681 11482 37745
rect 11498 37681 11562 37745
rect 11578 37681 11642 37745
rect 11658 37681 11722 37745
rect 11738 37681 11802 37745
rect 11818 37681 11882 37745
rect 11898 37681 11962 37745
rect 11978 37681 12042 37745
rect 12058 37681 12122 37745
rect 12138 37681 12202 37745
rect 12218 37681 12282 37745
rect 11098 37600 11162 37664
rect 11178 37600 11242 37664
rect 11258 37600 11322 37664
rect 11338 37600 11402 37664
rect 11418 37600 11482 37664
rect 11498 37600 11562 37664
rect 11578 37600 11642 37664
rect 11658 37600 11722 37664
rect 11738 37600 11802 37664
rect 11818 37600 11882 37664
rect 11898 37600 11962 37664
rect 11978 37600 12042 37664
rect 12058 37600 12122 37664
rect 12138 37600 12202 37664
rect 12218 37600 12282 37664
rect 11098 37519 11162 37583
rect 11178 37519 11242 37583
rect 11258 37519 11322 37583
rect 11338 37519 11402 37583
rect 11418 37519 11482 37583
rect 11498 37519 11562 37583
rect 11578 37519 11642 37583
rect 11658 37519 11722 37583
rect 11738 37519 11802 37583
rect 11818 37519 11882 37583
rect 11898 37519 11962 37583
rect 11978 37519 12042 37583
rect 12058 37519 12122 37583
rect 12138 37519 12202 37583
rect 12218 37519 12282 37583
rect 11098 37438 11162 37502
rect 11178 37438 11242 37502
rect 11258 37438 11322 37502
rect 11338 37438 11402 37502
rect 11418 37438 11482 37502
rect 11498 37438 11562 37502
rect 11578 37438 11642 37502
rect 11658 37438 11722 37502
rect 11738 37438 11802 37502
rect 11818 37438 11882 37502
rect 11898 37438 11962 37502
rect 11978 37438 12042 37502
rect 12058 37438 12122 37502
rect 12138 37438 12202 37502
rect 12218 37438 12282 37502
rect 11098 37357 11162 37421
rect 11178 37357 11242 37421
rect 11258 37357 11322 37421
rect 11338 37357 11402 37421
rect 11418 37357 11482 37421
rect 11498 37357 11562 37421
rect 11578 37357 11642 37421
rect 11658 37357 11722 37421
rect 11738 37357 11802 37421
rect 11818 37357 11882 37421
rect 11898 37357 11962 37421
rect 11978 37357 12042 37421
rect 12058 37357 12122 37421
rect 12138 37357 12202 37421
rect 12218 37357 12282 37421
rect 11098 37276 11162 37340
rect 11178 37276 11242 37340
rect 11258 37276 11322 37340
rect 11338 37276 11402 37340
rect 11418 37276 11482 37340
rect 11498 37276 11562 37340
rect 11578 37276 11642 37340
rect 11658 37276 11722 37340
rect 11738 37276 11802 37340
rect 11818 37276 11882 37340
rect 11898 37276 11962 37340
rect 11978 37276 12042 37340
rect 12058 37276 12122 37340
rect 12138 37276 12202 37340
rect 12218 37276 12282 37340
rect 11098 37195 11162 37259
rect 11178 37195 11242 37259
rect 11258 37195 11322 37259
rect 11338 37195 11402 37259
rect 11418 37195 11482 37259
rect 11498 37195 11562 37259
rect 11578 37195 11642 37259
rect 11658 37195 11722 37259
rect 11738 37195 11802 37259
rect 11818 37195 11882 37259
rect 11898 37195 11962 37259
rect 11978 37195 12042 37259
rect 12058 37195 12122 37259
rect 12138 37195 12202 37259
rect 12218 37195 12282 37259
rect 11098 37114 11162 37178
rect 11178 37114 11242 37178
rect 11258 37114 11322 37178
rect 11338 37114 11402 37178
rect 11418 37114 11482 37178
rect 11498 37114 11562 37178
rect 11578 37114 11642 37178
rect 11658 37114 11722 37178
rect 11738 37114 11802 37178
rect 11818 37114 11882 37178
rect 11898 37114 11962 37178
rect 11978 37114 12042 37178
rect 12058 37114 12122 37178
rect 12138 37114 12202 37178
rect 12218 37114 12282 37178
rect 11098 37033 11162 37097
rect 11178 37033 11242 37097
rect 11258 37033 11322 37097
rect 11338 37033 11402 37097
rect 11418 37033 11482 37097
rect 11498 37033 11562 37097
rect 11578 37033 11642 37097
rect 11658 37033 11722 37097
rect 11738 37033 11802 37097
rect 11818 37033 11882 37097
rect 11898 37033 11962 37097
rect 11978 37033 12042 37097
rect 12058 37033 12122 37097
rect 12138 37033 12202 37097
rect 12218 37033 12282 37097
rect 11098 36952 11162 37016
rect 11178 36952 11242 37016
rect 11258 36952 11322 37016
rect 11338 36952 11402 37016
rect 11418 36952 11482 37016
rect 11498 36952 11562 37016
rect 11578 36952 11642 37016
rect 11658 36952 11722 37016
rect 11738 36952 11802 37016
rect 11818 36952 11882 37016
rect 11898 36952 11962 37016
rect 11978 36952 12042 37016
rect 12058 36952 12122 37016
rect 12138 36952 12202 37016
rect 12218 36952 12282 37016
rect 11098 36871 11162 36935
rect 11178 36871 11242 36935
rect 11258 36871 11322 36935
rect 11338 36871 11402 36935
rect 11418 36871 11482 36935
rect 11498 36871 11562 36935
rect 11578 36871 11642 36935
rect 11658 36871 11722 36935
rect 11738 36871 11802 36935
rect 11818 36871 11882 36935
rect 11898 36871 11962 36935
rect 11978 36871 12042 36935
rect 12058 36871 12122 36935
rect 12138 36871 12202 36935
rect 12218 36871 12282 36935
rect 11098 36790 11162 36854
rect 11178 36790 11242 36854
rect 11258 36790 11322 36854
rect 11338 36790 11402 36854
rect 11418 36790 11482 36854
rect 11498 36790 11562 36854
rect 11578 36790 11642 36854
rect 11658 36790 11722 36854
rect 11738 36790 11802 36854
rect 11818 36790 11882 36854
rect 11898 36790 11962 36854
rect 11978 36790 12042 36854
rect 12058 36790 12122 36854
rect 12138 36790 12202 36854
rect 12218 36790 12282 36854
rect 11098 36709 11162 36773
rect 11178 36709 11242 36773
rect 11258 36709 11322 36773
rect 11338 36709 11402 36773
rect 11418 36709 11482 36773
rect 11498 36709 11562 36773
rect 11578 36709 11642 36773
rect 11658 36709 11722 36773
rect 11738 36709 11802 36773
rect 11818 36709 11882 36773
rect 11898 36709 11962 36773
rect 11978 36709 12042 36773
rect 12058 36709 12122 36773
rect 12138 36709 12202 36773
rect 12218 36709 12282 36773
rect 11098 36628 11162 36692
rect 11178 36628 11242 36692
rect 11258 36628 11322 36692
rect 11338 36628 11402 36692
rect 11418 36628 11482 36692
rect 11498 36628 11562 36692
rect 11578 36628 11642 36692
rect 11658 36628 11722 36692
rect 11738 36628 11802 36692
rect 11818 36628 11882 36692
rect 11898 36628 11962 36692
rect 11978 36628 12042 36692
rect 12058 36628 12122 36692
rect 12138 36628 12202 36692
rect 12218 36628 12282 36692
rect 11098 36547 11162 36611
rect 11178 36547 11242 36611
rect 11258 36547 11322 36611
rect 11338 36547 11402 36611
rect 11418 36547 11482 36611
rect 11498 36547 11562 36611
rect 11578 36547 11642 36611
rect 11658 36547 11722 36611
rect 11738 36547 11802 36611
rect 11818 36547 11882 36611
rect 11898 36547 11962 36611
rect 11978 36547 12042 36611
rect 12058 36547 12122 36611
rect 12138 36547 12202 36611
rect 12218 36547 12282 36611
rect 11098 36466 11162 36530
rect 11178 36466 11242 36530
rect 11258 36466 11322 36530
rect 11338 36466 11402 36530
rect 11418 36466 11482 36530
rect 11498 36466 11562 36530
rect 11578 36466 11642 36530
rect 11658 36466 11722 36530
rect 11738 36466 11802 36530
rect 11818 36466 11882 36530
rect 11898 36466 11962 36530
rect 11978 36466 12042 36530
rect 12058 36466 12122 36530
rect 12138 36466 12202 36530
rect 12218 36466 12282 36530
rect 11098 36385 11162 36449
rect 11178 36385 11242 36449
rect 11258 36385 11322 36449
rect 11338 36385 11402 36449
rect 11418 36385 11482 36449
rect 11498 36385 11562 36449
rect 11578 36385 11642 36449
rect 11658 36385 11722 36449
rect 11738 36385 11802 36449
rect 11818 36385 11882 36449
rect 11898 36385 11962 36449
rect 11978 36385 12042 36449
rect 12058 36385 12122 36449
rect 12138 36385 12202 36449
rect 12218 36385 12282 36449
rect 11098 36304 11162 36368
rect 11178 36304 11242 36368
rect 11258 36304 11322 36368
rect 11338 36304 11402 36368
rect 11418 36304 11482 36368
rect 11498 36304 11562 36368
rect 11578 36304 11642 36368
rect 11658 36304 11722 36368
rect 11738 36304 11802 36368
rect 11818 36304 11882 36368
rect 11898 36304 11962 36368
rect 11978 36304 12042 36368
rect 12058 36304 12122 36368
rect 12138 36304 12202 36368
rect 12218 36304 12282 36368
rect 11098 36223 11162 36287
rect 11178 36223 11242 36287
rect 11258 36223 11322 36287
rect 11338 36223 11402 36287
rect 11418 36223 11482 36287
rect 11498 36223 11562 36287
rect 11578 36223 11642 36287
rect 11658 36223 11722 36287
rect 11738 36223 11802 36287
rect 11818 36223 11882 36287
rect 11898 36223 11962 36287
rect 11978 36223 12042 36287
rect 12058 36223 12122 36287
rect 12138 36223 12202 36287
rect 12218 36223 12282 36287
rect 11098 36142 11162 36206
rect 11178 36142 11242 36206
rect 11258 36142 11322 36206
rect 11338 36142 11402 36206
rect 11418 36142 11482 36206
rect 11498 36142 11562 36206
rect 11578 36142 11642 36206
rect 11658 36142 11722 36206
rect 11738 36142 11802 36206
rect 11818 36142 11882 36206
rect 11898 36142 11962 36206
rect 11978 36142 12042 36206
rect 12058 36142 12122 36206
rect 12138 36142 12202 36206
rect 12218 36142 12282 36206
rect 11098 36060 11162 36124
rect 11178 36060 11242 36124
rect 11258 36060 11322 36124
rect 11338 36060 11402 36124
rect 11418 36060 11482 36124
rect 11498 36060 11562 36124
rect 11578 36060 11642 36124
rect 11658 36060 11722 36124
rect 11738 36060 11802 36124
rect 11818 36060 11882 36124
rect 11898 36060 11962 36124
rect 11978 36060 12042 36124
rect 12058 36060 12122 36124
rect 12138 36060 12202 36124
rect 12218 36060 12282 36124
rect 11098 35978 11162 36042
rect 11178 35978 11242 36042
rect 11258 35978 11322 36042
rect 11338 35978 11402 36042
rect 11418 35978 11482 36042
rect 11498 35978 11562 36042
rect 11578 35978 11642 36042
rect 11658 35978 11722 36042
rect 11738 35978 11802 36042
rect 11818 35978 11882 36042
rect 11898 35978 11962 36042
rect 11978 35978 12042 36042
rect 12058 35978 12122 36042
rect 12138 35978 12202 36042
rect 12218 35978 12282 36042
rect 11098 35896 11162 35960
rect 11178 35896 11242 35960
rect 11258 35896 11322 35960
rect 11338 35896 11402 35960
rect 11418 35896 11482 35960
rect 11498 35896 11562 35960
rect 11578 35896 11642 35960
rect 11658 35896 11722 35960
rect 11738 35896 11802 35960
rect 11818 35896 11882 35960
rect 11898 35896 11962 35960
rect 11978 35896 12042 35960
rect 12058 35896 12122 35960
rect 12138 35896 12202 35960
rect 12218 35896 12282 35960
rect 11098 35814 11162 35878
rect 11178 35814 11242 35878
rect 11258 35814 11322 35878
rect 11338 35814 11402 35878
rect 11418 35814 11482 35878
rect 11498 35814 11562 35878
rect 11578 35814 11642 35878
rect 11658 35814 11722 35878
rect 11738 35814 11802 35878
rect 11818 35814 11882 35878
rect 11898 35814 11962 35878
rect 11978 35814 12042 35878
rect 12058 35814 12122 35878
rect 12138 35814 12202 35878
rect 12218 35814 12282 35878
rect 11098 35732 11162 35796
rect 11178 35732 11242 35796
rect 11258 35732 11322 35796
rect 11338 35732 11402 35796
rect 11418 35732 11482 35796
rect 11498 35732 11562 35796
rect 11578 35732 11642 35796
rect 11658 35732 11722 35796
rect 11738 35732 11802 35796
rect 11818 35732 11882 35796
rect 11898 35732 11962 35796
rect 11978 35732 12042 35796
rect 12058 35732 12122 35796
rect 12138 35732 12202 35796
rect 12218 35732 12282 35796
rect 11098 35650 11162 35714
rect 11178 35650 11242 35714
rect 11258 35650 11322 35714
rect 11338 35650 11402 35714
rect 11418 35650 11482 35714
rect 11498 35650 11562 35714
rect 11578 35650 11642 35714
rect 11658 35650 11722 35714
rect 11738 35650 11802 35714
rect 11818 35650 11882 35714
rect 11898 35650 11962 35714
rect 11978 35650 12042 35714
rect 12058 35650 12122 35714
rect 12138 35650 12202 35714
rect 12218 35650 12282 35714
rect 11098 35568 11162 35632
rect 11178 35568 11242 35632
rect 11258 35568 11322 35632
rect 11338 35568 11402 35632
rect 11418 35568 11482 35632
rect 11498 35568 11562 35632
rect 11578 35568 11642 35632
rect 11658 35568 11722 35632
rect 11738 35568 11802 35632
rect 11818 35568 11882 35632
rect 11898 35568 11962 35632
rect 11978 35568 12042 35632
rect 12058 35568 12122 35632
rect 12138 35568 12202 35632
rect 12218 35568 12282 35632
rect 11098 35486 11162 35550
rect 11178 35486 11242 35550
rect 11258 35486 11322 35550
rect 11338 35486 11402 35550
rect 11418 35486 11482 35550
rect 11498 35486 11562 35550
rect 11578 35486 11642 35550
rect 11658 35486 11722 35550
rect 11738 35486 11802 35550
rect 11818 35486 11882 35550
rect 11898 35486 11962 35550
rect 11978 35486 12042 35550
rect 12058 35486 12122 35550
rect 12138 35486 12202 35550
rect 12218 35486 12282 35550
rect 11098 35404 11162 35468
rect 11178 35404 11242 35468
rect 11258 35404 11322 35468
rect 11338 35404 11402 35468
rect 11418 35404 11482 35468
rect 11498 35404 11562 35468
rect 11578 35404 11642 35468
rect 11658 35404 11722 35468
rect 11738 35404 11802 35468
rect 11818 35404 11882 35468
rect 11898 35404 11962 35468
rect 11978 35404 12042 35468
rect 12058 35404 12122 35468
rect 12138 35404 12202 35468
rect 12218 35404 12282 35468
rect 11098 35322 11162 35386
rect 11178 35322 11242 35386
rect 11258 35322 11322 35386
rect 11338 35322 11402 35386
rect 11418 35322 11482 35386
rect 11498 35322 11562 35386
rect 11578 35322 11642 35386
rect 11658 35322 11722 35386
rect 11738 35322 11802 35386
rect 11818 35322 11882 35386
rect 11898 35322 11962 35386
rect 11978 35322 12042 35386
rect 12058 35322 12122 35386
rect 12138 35322 12202 35386
rect 12218 35322 12282 35386
rect 11098 35240 11162 35304
rect 11178 35240 11242 35304
rect 11258 35240 11322 35304
rect 11338 35240 11402 35304
rect 11418 35240 11482 35304
rect 11498 35240 11562 35304
rect 11578 35240 11642 35304
rect 11658 35240 11722 35304
rect 11738 35240 11802 35304
rect 11818 35240 11882 35304
rect 11898 35240 11962 35304
rect 11978 35240 12042 35304
rect 12058 35240 12122 35304
rect 12138 35240 12202 35304
rect 12218 35240 12282 35304
rect 11098 35158 11162 35222
rect 11178 35158 11242 35222
rect 11258 35158 11322 35222
rect 11338 35158 11402 35222
rect 11418 35158 11482 35222
rect 11498 35158 11562 35222
rect 11578 35158 11642 35222
rect 11658 35158 11722 35222
rect 11738 35158 11802 35222
rect 11818 35158 11882 35222
rect 11898 35158 11962 35222
rect 11978 35158 12042 35222
rect 12058 35158 12122 35222
rect 12138 35158 12202 35222
rect 12218 35158 12282 35222
rect 12588 39308 12652 39372
rect 12676 39308 12740 39372
rect 12764 39308 12828 39372
rect 12852 39308 12916 39372
rect 12940 39308 13004 39372
rect 12588 39228 12652 39292
rect 12676 39228 12740 39292
rect 12764 39228 12828 39292
rect 12852 39228 12916 39292
rect 12940 39228 13004 39292
rect 12588 39148 12652 39212
rect 12676 39148 12740 39212
rect 12764 39148 12828 39212
rect 12852 39148 12916 39212
rect 12940 39148 13004 39212
rect 12588 39068 12652 39132
rect 12676 39068 12740 39132
rect 12764 39068 12828 39132
rect 12852 39068 12916 39132
rect 12940 39068 13004 39132
rect 12588 38988 12652 39052
rect 12676 38988 12740 39052
rect 12764 38988 12828 39052
rect 12852 38988 12916 39052
rect 12940 38988 13004 39052
rect 12588 38908 12652 38972
rect 12676 38908 12740 38972
rect 12764 38908 12828 38972
rect 12852 38908 12916 38972
rect 12940 38908 13004 38972
rect 12588 38828 12652 38892
rect 12676 38828 12740 38892
rect 12764 38828 12828 38892
rect 12852 38828 12916 38892
rect 12940 38828 13004 38892
rect 12588 38748 12652 38812
rect 12676 38748 12740 38812
rect 12764 38748 12828 38812
rect 12852 38748 12916 38812
rect 12940 38748 13004 38812
rect 12588 38667 12652 38731
rect 12676 38667 12740 38731
rect 12764 38667 12828 38731
rect 12852 38667 12916 38731
rect 12940 38667 13004 38731
rect 12588 38586 12652 38650
rect 12676 38586 12740 38650
rect 12764 38586 12828 38650
rect 12852 38586 12916 38650
rect 12940 38586 13004 38650
rect 12588 38505 12652 38569
rect 12676 38505 12740 38569
rect 12764 38505 12828 38569
rect 12852 38505 12916 38569
rect 12940 38505 13004 38569
rect 12588 38424 12652 38488
rect 12676 38424 12740 38488
rect 12764 38424 12828 38488
rect 12852 38424 12916 38488
rect 12940 38424 13004 38488
rect 12588 38343 12652 38407
rect 12676 38343 12740 38407
rect 12764 38343 12828 38407
rect 12852 38343 12916 38407
rect 12940 38343 13004 38407
rect 12588 38262 12652 38326
rect 12676 38262 12740 38326
rect 12764 38262 12828 38326
rect 12852 38262 12916 38326
rect 12940 38262 13004 38326
rect 12588 38181 12652 38245
rect 12676 38181 12740 38245
rect 12764 38181 12828 38245
rect 12852 38181 12916 38245
rect 12940 38181 13004 38245
rect 12588 38100 12652 38164
rect 12676 38100 12740 38164
rect 12764 38100 12828 38164
rect 12852 38100 12916 38164
rect 12940 38100 13004 38164
rect 12588 38019 12652 38083
rect 12676 38019 12740 38083
rect 12764 38019 12828 38083
rect 12852 38019 12916 38083
rect 12940 38019 13004 38083
rect 12588 37938 12652 38002
rect 12676 37938 12740 38002
rect 12764 37938 12828 38002
rect 12852 37938 12916 38002
rect 12940 37938 13004 38002
rect 12588 37857 12652 37921
rect 12676 37857 12740 37921
rect 12764 37857 12828 37921
rect 12852 37857 12916 37921
rect 12940 37857 13004 37921
rect 12588 37776 12652 37840
rect 12676 37776 12740 37840
rect 12764 37776 12828 37840
rect 12852 37776 12916 37840
rect 12940 37776 13004 37840
rect 12588 37695 12652 37759
rect 12676 37695 12740 37759
rect 12764 37695 12828 37759
rect 12852 37695 12916 37759
rect 12940 37695 13004 37759
rect 12588 37614 12652 37678
rect 12676 37614 12740 37678
rect 12764 37614 12828 37678
rect 12852 37614 12916 37678
rect 12940 37614 13004 37678
rect 12588 37533 12652 37597
rect 12676 37533 12740 37597
rect 12764 37533 12828 37597
rect 12852 37533 12916 37597
rect 12940 37533 13004 37597
rect 12588 37452 12652 37516
rect 12676 37452 12740 37516
rect 12764 37452 12828 37516
rect 12852 37452 12916 37516
rect 12940 37452 13004 37516
rect 12588 37371 12652 37435
rect 12676 37371 12740 37435
rect 12764 37371 12828 37435
rect 12852 37371 12916 37435
rect 12940 37371 13004 37435
rect 12588 37290 12652 37354
rect 12676 37290 12740 37354
rect 12764 37290 12828 37354
rect 12852 37290 12916 37354
rect 12940 37290 13004 37354
rect 12588 37209 12652 37273
rect 12676 37209 12740 37273
rect 12764 37209 12828 37273
rect 12852 37209 12916 37273
rect 12940 37209 13004 37273
rect 12588 37128 12652 37192
rect 12676 37128 12740 37192
rect 12764 37128 12828 37192
rect 12852 37128 12916 37192
rect 12940 37128 13004 37192
rect 12588 37047 12652 37111
rect 12676 37047 12740 37111
rect 12764 37047 12828 37111
rect 12852 37047 12916 37111
rect 12940 37047 13004 37111
rect 12588 36966 12652 37030
rect 12676 36966 12740 37030
rect 12764 36966 12828 37030
rect 12852 36966 12916 37030
rect 12940 36966 13004 37030
rect 12588 36885 12652 36949
rect 12676 36885 12740 36949
rect 12764 36885 12828 36949
rect 12852 36885 12916 36949
rect 12940 36885 13004 36949
rect 12588 36804 12652 36868
rect 12676 36804 12740 36868
rect 12764 36804 12828 36868
rect 12852 36804 12916 36868
rect 12940 36804 13004 36868
rect 12588 36723 12652 36787
rect 12676 36723 12740 36787
rect 12764 36723 12828 36787
rect 12852 36723 12916 36787
rect 12940 36723 13004 36787
rect 12588 36642 12652 36706
rect 12676 36642 12740 36706
rect 12764 36642 12828 36706
rect 12852 36642 12916 36706
rect 12940 36642 13004 36706
rect 12588 36561 12652 36625
rect 12676 36561 12740 36625
rect 12764 36561 12828 36625
rect 12852 36561 12916 36625
rect 12940 36561 13004 36625
rect 12588 36480 12652 36544
rect 12676 36480 12740 36544
rect 12764 36480 12828 36544
rect 12852 36480 12916 36544
rect 12940 36480 13004 36544
rect 12588 36399 12652 36463
rect 12676 36399 12740 36463
rect 12764 36399 12828 36463
rect 12852 36399 12916 36463
rect 12940 36399 13004 36463
rect 12588 36318 12652 36382
rect 12676 36318 12740 36382
rect 12764 36318 12828 36382
rect 12852 36318 12916 36382
rect 12940 36318 13004 36382
rect 12588 36237 12652 36301
rect 12676 36237 12740 36301
rect 12764 36237 12828 36301
rect 12852 36237 12916 36301
rect 12940 36237 13004 36301
rect 12588 36156 12652 36220
rect 12676 36156 12740 36220
rect 12764 36156 12828 36220
rect 12852 36156 12916 36220
rect 12940 36156 13004 36220
rect 12588 36075 12652 36139
rect 12676 36075 12740 36139
rect 12764 36075 12828 36139
rect 12852 36075 12916 36139
rect 12940 36075 13004 36139
rect 12588 35994 12652 36058
rect 12676 35994 12740 36058
rect 12764 35994 12828 36058
rect 12852 35994 12916 36058
rect 12940 35994 13004 36058
rect 12588 35913 12652 35977
rect 12676 35913 12740 35977
rect 12764 35913 12828 35977
rect 12852 35913 12916 35977
rect 12940 35913 13004 35977
rect 12598 35787 12662 35851
rect 12682 35787 12746 35851
rect 12766 35787 12830 35851
rect 12850 35787 12914 35851
rect 12933 35787 12997 35851
rect 13016 35787 13080 35851
rect 13099 35787 13163 35851
rect 13182 35787 13246 35851
rect 12598 35703 12662 35767
rect 12682 35703 12746 35767
rect 12766 35703 12830 35767
rect 12850 35703 12914 35767
rect 12933 35703 12997 35767
rect 13016 35703 13080 35767
rect 13099 35703 13163 35767
rect 13182 35703 13246 35767
rect 12598 35619 12662 35683
rect 12682 35619 12746 35683
rect 12766 35619 12830 35683
rect 12850 35619 12914 35683
rect 12933 35619 12997 35683
rect 13016 35619 13080 35683
rect 13099 35619 13163 35683
rect 13182 35619 13246 35683
rect 12598 35535 12662 35599
rect 12682 35535 12746 35599
rect 12766 35535 12830 35599
rect 12850 35535 12914 35599
rect 12933 35535 12997 35599
rect 13016 35535 13080 35599
rect 13099 35535 13163 35599
rect 13182 35535 13246 35599
rect 12598 35451 12662 35515
rect 12682 35451 12746 35515
rect 12766 35451 12830 35515
rect 12850 35451 12914 35515
rect 12933 35451 12997 35515
rect 13016 35451 13080 35515
rect 13099 35451 13163 35515
rect 13182 35451 13246 35515
rect 12598 35367 12662 35431
rect 12682 35367 12746 35431
rect 12766 35367 12830 35431
rect 12850 35367 12914 35431
rect 12933 35367 12997 35431
rect 13016 35367 13080 35431
rect 13099 35367 13163 35431
rect 13182 35367 13246 35431
rect 1977 25789 2041 25853
rect 2067 25789 2131 25853
rect 2157 25820 2221 25853
rect 2247 25820 2311 25853
rect 2337 25820 2401 25853
rect 2427 25820 2491 25853
rect 2157 25789 2170 25820
rect 2170 25789 2221 25820
rect 2247 25789 2252 25820
rect 2252 25789 2308 25820
rect 2308 25789 2311 25820
rect 2337 25789 2390 25820
rect 2390 25789 2401 25820
rect 2427 25789 2472 25820
rect 2472 25789 2491 25820
rect 1977 25706 2041 25770
rect 2067 25706 2131 25770
rect 2157 25764 2170 25770
rect 2170 25764 2221 25770
rect 2247 25764 2252 25770
rect 2252 25764 2308 25770
rect 2308 25764 2311 25770
rect 2337 25764 2390 25770
rect 2390 25764 2401 25770
rect 2427 25764 2472 25770
rect 2472 25764 2491 25770
rect 2157 25739 2221 25764
rect 2247 25739 2311 25764
rect 2337 25739 2401 25764
rect 2427 25739 2491 25764
rect 2157 25706 2170 25739
rect 2170 25706 2221 25739
rect 2247 25706 2252 25739
rect 2252 25706 2308 25739
rect 2308 25706 2311 25739
rect 2337 25706 2390 25739
rect 2390 25706 2401 25739
rect 2427 25706 2472 25739
rect 2472 25706 2491 25739
rect 1977 25623 2041 25687
rect 2067 25623 2131 25687
rect 2157 25683 2170 25687
rect 2170 25683 2221 25687
rect 2247 25683 2252 25687
rect 2252 25683 2308 25687
rect 2308 25683 2311 25687
rect 2337 25683 2390 25687
rect 2390 25683 2401 25687
rect 2427 25683 2472 25687
rect 2472 25683 2491 25687
rect 2157 25658 2221 25683
rect 2247 25658 2311 25683
rect 2337 25658 2401 25683
rect 2427 25658 2491 25683
rect 2157 25623 2170 25658
rect 2170 25623 2221 25658
rect 2247 25623 2252 25658
rect 2252 25623 2308 25658
rect 2308 25623 2311 25658
rect 2337 25623 2390 25658
rect 2390 25623 2401 25658
rect 2427 25623 2472 25658
rect 2472 25623 2491 25658
rect 1977 25540 2041 25604
rect 2067 25540 2131 25604
rect 2157 25602 2170 25604
rect 2170 25602 2221 25604
rect 2247 25602 2252 25604
rect 2252 25602 2308 25604
rect 2308 25602 2311 25604
rect 2337 25602 2390 25604
rect 2390 25602 2401 25604
rect 2427 25602 2472 25604
rect 2472 25602 2491 25604
rect 2157 25577 2221 25602
rect 2247 25577 2311 25602
rect 2337 25577 2401 25602
rect 2427 25577 2491 25602
rect 2157 25540 2170 25577
rect 2170 25540 2221 25577
rect 2247 25540 2252 25577
rect 2252 25540 2308 25577
rect 2308 25540 2311 25577
rect 2337 25540 2390 25577
rect 2390 25540 2401 25577
rect 2427 25540 2472 25577
rect 2472 25540 2491 25577
rect 1977 25457 2041 25521
rect 2067 25457 2131 25521
rect 2157 25496 2221 25521
rect 2247 25496 2311 25521
rect 2337 25496 2401 25521
rect 2427 25496 2491 25521
rect 2157 25457 2170 25496
rect 2170 25457 2221 25496
rect 2247 25457 2252 25496
rect 2252 25457 2308 25496
rect 2308 25457 2311 25496
rect 2337 25457 2390 25496
rect 2390 25457 2401 25496
rect 2427 25457 2472 25496
rect 2472 25457 2491 25496
rect 1977 25373 2041 25437
rect 2067 25373 2131 25437
rect 2157 25415 2221 25437
rect 2247 25415 2311 25437
rect 2337 25415 2401 25437
rect 2427 25415 2491 25437
rect 2157 25373 2170 25415
rect 2170 25373 2221 25415
rect 2247 25373 2252 25415
rect 2252 25373 2308 25415
rect 2308 25373 2311 25415
rect 2337 25373 2390 25415
rect 2390 25373 2401 25415
rect 2427 25373 2472 25415
rect 2472 25373 2491 25415
rect 1977 25289 2041 25353
rect 2067 25289 2131 25353
rect 2157 25334 2221 25353
rect 2247 25334 2311 25353
rect 2337 25334 2401 25353
rect 2427 25334 2491 25353
rect 2157 25289 2170 25334
rect 2170 25289 2221 25334
rect 2247 25289 2252 25334
rect 2252 25289 2308 25334
rect 2308 25289 2311 25334
rect 2337 25289 2390 25334
rect 2390 25289 2401 25334
rect 2427 25289 2472 25334
rect 2472 25289 2491 25334
rect 1977 25205 2041 25269
rect 2067 25205 2131 25269
rect 2157 25253 2221 25269
rect 2247 25253 2311 25269
rect 2337 25253 2401 25269
rect 2427 25253 2491 25269
rect 2157 25205 2170 25253
rect 2170 25205 2221 25253
rect 2247 25205 2252 25253
rect 2252 25205 2308 25253
rect 2308 25205 2311 25253
rect 2337 25205 2390 25253
rect 2390 25205 2401 25253
rect 2427 25205 2472 25253
rect 2472 25205 2491 25253
rect 1977 25121 2041 25185
rect 2067 25121 2131 25185
rect 2157 25172 2221 25185
rect 2247 25172 2311 25185
rect 2337 25172 2401 25185
rect 2427 25172 2491 25185
rect 2157 25121 2170 25172
rect 2170 25121 2221 25172
rect 2247 25121 2252 25172
rect 2252 25121 2308 25172
rect 2308 25121 2311 25172
rect 2337 25121 2390 25172
rect 2390 25121 2401 25172
rect 2427 25121 2472 25172
rect 2472 25121 2491 25172
rect 1977 25037 2041 25101
rect 2067 25037 2131 25101
rect 2157 25091 2221 25101
rect 2247 25091 2311 25101
rect 2337 25091 2401 25101
rect 2427 25091 2491 25101
rect 2157 25037 2170 25091
rect 2170 25037 2221 25091
rect 2247 25037 2252 25091
rect 2252 25037 2308 25091
rect 2308 25037 2311 25091
rect 2337 25037 2390 25091
rect 2390 25037 2401 25091
rect 2427 25037 2472 25091
rect 2472 25037 2491 25091
rect 1977 24953 2041 25017
rect 2067 24953 2131 25017
rect 2157 25010 2221 25017
rect 2247 25010 2311 25017
rect 2337 25010 2401 25017
rect 2427 25010 2491 25017
rect 2157 24954 2170 25010
rect 2170 24954 2221 25010
rect 2247 24954 2252 25010
rect 2252 24954 2308 25010
rect 2308 24954 2311 25010
rect 2337 24954 2390 25010
rect 2390 24954 2401 25010
rect 2427 24954 2472 25010
rect 2472 24954 2491 25010
rect 2157 24953 2221 24954
rect 2247 24953 2311 24954
rect 2337 24953 2401 24954
rect 2427 24953 2491 24954
rect 1977 24869 2041 24933
rect 2067 24869 2131 24933
rect 2157 24929 2221 24933
rect 2247 24929 2311 24933
rect 2337 24929 2401 24933
rect 2427 24929 2491 24933
rect 2157 24873 2170 24929
rect 2170 24873 2221 24929
rect 2247 24873 2252 24929
rect 2252 24873 2308 24929
rect 2308 24873 2311 24929
rect 2337 24873 2390 24929
rect 2390 24873 2401 24929
rect 2427 24873 2472 24929
rect 2472 24873 2491 24929
rect 2157 24869 2221 24873
rect 2247 24869 2311 24873
rect 2337 24869 2401 24873
rect 2427 24869 2491 24873
rect 1977 24785 2041 24849
rect 2067 24785 2131 24849
rect 2157 24848 2221 24849
rect 2247 24848 2311 24849
rect 2337 24848 2401 24849
rect 2427 24848 2491 24849
rect 2157 24792 2170 24848
rect 2170 24792 2221 24848
rect 2247 24792 2252 24848
rect 2252 24792 2308 24848
rect 2308 24792 2311 24848
rect 2337 24792 2390 24848
rect 2390 24792 2401 24848
rect 2427 24792 2472 24848
rect 2472 24792 2491 24848
rect 2157 24785 2221 24792
rect 2247 24785 2311 24792
rect 2337 24785 2401 24792
rect 2427 24785 2491 24792
rect 1977 24701 2041 24765
rect 2067 24701 2131 24765
rect 2157 24711 2170 24765
rect 2170 24711 2221 24765
rect 2247 24711 2252 24765
rect 2252 24711 2308 24765
rect 2308 24711 2311 24765
rect 2337 24711 2390 24765
rect 2390 24711 2401 24765
rect 2427 24711 2472 24765
rect 2472 24711 2491 24765
rect 2157 24701 2221 24711
rect 2247 24701 2311 24711
rect 2337 24701 2401 24711
rect 2427 24701 2491 24711
rect 1977 24617 2041 24681
rect 2067 24617 2131 24681
rect 2157 24630 2170 24681
rect 2170 24630 2221 24681
rect 2247 24630 2252 24681
rect 2252 24630 2308 24681
rect 2308 24630 2311 24681
rect 2337 24630 2390 24681
rect 2390 24630 2401 24681
rect 2427 24630 2472 24681
rect 2472 24630 2491 24681
rect 2157 24617 2221 24630
rect 2247 24617 2311 24630
rect 2337 24617 2401 24630
rect 2427 24617 2491 24630
rect 1977 24533 2041 24597
rect 2067 24533 2131 24597
rect 2157 24548 2170 24597
rect 2170 24548 2221 24597
rect 2247 24548 2252 24597
rect 2252 24548 2308 24597
rect 2308 24548 2311 24597
rect 2337 24548 2390 24597
rect 2390 24548 2401 24597
rect 2427 24548 2472 24597
rect 2472 24548 2491 24597
rect 2157 24533 2221 24548
rect 2247 24533 2311 24548
rect 2337 24533 2401 24548
rect 2427 24533 2491 24548
rect 1977 24449 2041 24513
rect 2067 24449 2131 24513
rect 2157 24466 2170 24513
rect 2170 24466 2221 24513
rect 2247 24466 2252 24513
rect 2252 24466 2308 24513
rect 2308 24466 2311 24513
rect 2337 24466 2390 24513
rect 2390 24466 2401 24513
rect 2427 24466 2472 24513
rect 2472 24466 2491 24513
rect 2157 24449 2221 24466
rect 2247 24449 2311 24466
rect 2337 24449 2401 24466
rect 2427 24449 2491 24466
rect 1977 24365 2041 24429
rect 2067 24365 2131 24429
rect 2157 24384 2170 24429
rect 2170 24384 2221 24429
rect 2247 24384 2252 24429
rect 2252 24384 2308 24429
rect 2308 24384 2311 24429
rect 2337 24384 2390 24429
rect 2390 24384 2401 24429
rect 2427 24384 2472 24429
rect 2472 24384 2491 24429
rect 2157 24365 2221 24384
rect 2247 24365 2311 24384
rect 2337 24365 2401 24384
rect 2427 24365 2491 24384
rect 1977 24281 2041 24345
rect 2067 24281 2131 24345
rect 2157 24302 2170 24345
rect 2170 24302 2221 24345
rect 2247 24302 2252 24345
rect 2252 24302 2308 24345
rect 2308 24302 2311 24345
rect 2337 24302 2390 24345
rect 2390 24302 2401 24345
rect 2427 24302 2472 24345
rect 2472 24302 2491 24345
rect 2157 24281 2221 24302
rect 2247 24281 2311 24302
rect 2337 24281 2401 24302
rect 2427 24281 2491 24302
rect 1977 24176 2041 24240
rect 2065 24176 2129 24240
rect 2153 24220 2170 24240
rect 2170 24220 2217 24240
rect 2241 24220 2252 24240
rect 2252 24220 2305 24240
rect 2328 24220 2334 24240
rect 2334 24220 2390 24240
rect 2390 24220 2392 24240
rect 2153 24194 2217 24220
rect 2241 24194 2305 24220
rect 2328 24194 2392 24220
rect 2153 24176 2170 24194
rect 2170 24176 2217 24194
rect 2241 24176 2252 24194
rect 2252 24176 2305 24194
rect 2328 24176 2334 24194
rect 2334 24176 2390 24194
rect 2390 24176 2392 24194
rect 2415 24220 2416 24240
rect 2416 24220 2472 24240
rect 2472 24220 2479 24240
rect 2415 24194 2479 24220
rect 2415 24176 2416 24194
rect 2416 24176 2472 24194
rect 2472 24176 2479 24194
rect 1977 24080 2041 24144
rect 2065 24080 2129 24144
rect 2153 24138 2170 24144
rect 2170 24138 2217 24144
rect 2241 24138 2252 24144
rect 2252 24138 2305 24144
rect 2328 24138 2334 24144
rect 2334 24138 2390 24144
rect 2390 24138 2392 24144
rect 2153 24112 2217 24138
rect 2241 24112 2305 24138
rect 2328 24112 2392 24138
rect 2153 24080 2170 24112
rect 2170 24080 2217 24112
rect 2241 24080 2252 24112
rect 2252 24080 2305 24112
rect 2328 24080 2334 24112
rect 2334 24080 2390 24112
rect 2390 24080 2392 24112
rect 2415 24138 2416 24144
rect 2416 24138 2472 24144
rect 2472 24138 2479 24144
rect 2415 24112 2479 24138
rect 2415 24080 2416 24112
rect 2416 24080 2472 24112
rect 2472 24080 2479 24112
rect 1739 23937 1803 24001
rect 1875 23937 1939 24001
rect 1977 23984 2041 24048
rect 2065 23984 2129 24048
rect 2153 24030 2217 24048
rect 2241 24030 2305 24048
rect 2328 24030 2392 24048
rect 2153 23984 2170 24030
rect 2170 23984 2217 24030
rect 2241 23984 2252 24030
rect 2252 23984 2305 24030
rect 2328 23984 2334 24030
rect 2334 23984 2390 24030
rect 2390 23984 2392 24030
rect 2415 24030 2479 24048
rect 2415 23984 2416 24030
rect 2416 23984 2472 24030
rect 2472 23984 2479 24030
rect 1977 23888 2041 23952
rect 2065 23888 2129 23952
rect 2153 23948 2217 23952
rect 2241 23948 2305 23952
rect 2328 23948 2392 23952
rect 2153 23892 2170 23948
rect 2170 23892 2217 23948
rect 2241 23892 2252 23948
rect 2252 23892 2305 23948
rect 2328 23892 2334 23948
rect 2334 23892 2390 23948
rect 2390 23892 2392 23948
rect 2153 23888 2217 23892
rect 2241 23888 2305 23892
rect 2328 23888 2392 23892
rect 2415 23948 2479 23952
rect 2415 23892 2416 23948
rect 2416 23892 2472 23948
rect 2472 23892 2479 23948
rect 2415 23888 2479 23892
rect 1739 23801 1803 23865
rect 1875 23801 1939 23865
rect 1977 23792 2041 23856
rect 2065 23792 2129 23856
rect 2153 23810 2170 23856
rect 2170 23810 2217 23856
rect 2241 23810 2252 23856
rect 2252 23810 2305 23856
rect 2328 23810 2334 23856
rect 2334 23810 2390 23856
rect 2390 23810 2392 23856
rect 2153 23792 2217 23810
rect 2241 23792 2305 23810
rect 2328 23792 2392 23810
rect 2415 23810 2416 23856
rect 2416 23810 2472 23856
rect 2472 23810 2479 23856
rect 2415 23792 2479 23810
rect 1094 23721 1158 23785
rect 1188 23721 1252 23785
rect 1282 23721 1346 23785
rect 1376 23721 1440 23785
rect 1094 23639 1158 23703
rect 1188 23639 1252 23703
rect 1282 23639 1346 23703
rect 1376 23639 1440 23703
rect 1094 23557 1158 23621
rect 1188 23557 1252 23621
rect 1282 23557 1346 23621
rect 1376 23557 1440 23621
rect 1094 23475 1158 23539
rect 1188 23475 1252 23539
rect 1282 23475 1346 23539
rect 1376 23475 1440 23539
rect 1094 23393 1158 23457
rect 1188 23393 1252 23457
rect 1282 23393 1346 23457
rect 1376 23393 1440 23457
rect 1094 23311 1158 23375
rect 1188 23311 1252 23375
rect 1282 23311 1346 23375
rect 1376 23311 1440 23375
rect 1094 23229 1158 23293
rect 1188 23229 1252 23293
rect 1282 23229 1346 23293
rect 1376 23229 1440 23293
rect 1094 23147 1158 23211
rect 1188 23147 1252 23211
rect 1282 23147 1346 23211
rect 1376 23147 1440 23211
rect 1094 23065 1158 23129
rect 1188 23065 1252 23129
rect 1282 23065 1346 23129
rect 1376 23065 1440 23129
rect 1094 22983 1158 23047
rect 1188 22983 1252 23047
rect 1282 22983 1346 23047
rect 1376 22983 1440 23047
rect 1094 22900 1158 22964
rect 1188 22900 1252 22964
rect 1282 22900 1346 22964
rect 1376 22900 1440 22964
rect 1094 22817 1158 22881
rect 1188 22817 1252 22881
rect 1282 22817 1346 22881
rect 1376 22817 1440 22881
rect 1094 22734 1158 22798
rect 1188 22734 1252 22798
rect 1282 22734 1346 22798
rect 1376 22734 1440 22798
rect 1094 22651 1158 22715
rect 1188 22651 1252 22715
rect 1282 22651 1346 22715
rect 1376 22651 1440 22715
rect 1094 22568 1158 22632
rect 1188 22568 1252 22632
rect 1282 22568 1346 22632
rect 1376 22568 1440 22632
rect 1094 22485 1158 22549
rect 1188 22485 1252 22549
rect 1282 22485 1346 22549
rect 1376 22485 1440 22549
rect 1094 22402 1158 22466
rect 1188 22402 1252 22466
rect 1282 22402 1346 22466
rect 1376 22402 1440 22466
rect 1094 22319 1158 22383
rect 1188 22319 1252 22383
rect 1282 22319 1346 22383
rect 1376 22319 1440 22383
rect 1094 22236 1158 22300
rect 1188 22236 1252 22300
rect 1282 22236 1346 22300
rect 1376 22236 1440 22300
rect 1094 22153 1158 22217
rect 1188 22153 1252 22217
rect 1282 22153 1346 22217
rect 1376 22153 1440 22217
rect 1094 22070 1158 22134
rect 1188 22070 1252 22134
rect 1282 22070 1346 22134
rect 1376 22070 1440 22134
rect 1094 21987 1158 22051
rect 1188 21987 1252 22051
rect 1282 21987 1346 22051
rect 1376 21987 1440 22051
rect 1094 21904 1158 21968
rect 1188 21904 1252 21968
rect 1282 21904 1346 21968
rect 1376 21904 1440 21968
rect 1094 21821 1158 21885
rect 1188 21821 1252 21885
rect 1282 21821 1346 21885
rect 1376 21821 1440 21885
rect 1094 21738 1158 21802
rect 1188 21738 1252 21802
rect 1282 21738 1346 21802
rect 1376 21738 1440 21802
rect 1094 21655 1158 21719
rect 1188 21655 1252 21719
rect 1282 21655 1346 21719
rect 1376 21655 1440 21719
rect 1094 21572 1158 21636
rect 1188 21572 1252 21636
rect 1282 21572 1346 21636
rect 1376 21572 1440 21636
rect 1094 21489 1158 21553
rect 1188 21489 1252 21553
rect 1282 21489 1346 21553
rect 1376 21489 1440 21553
rect 1094 21406 1158 21470
rect 1188 21406 1252 21470
rect 1282 21406 1346 21470
rect 1376 21406 1440 21470
rect 1094 21323 1158 21387
rect 1188 21323 1252 21387
rect 1282 21323 1346 21387
rect 1376 21323 1440 21387
rect 1474 23709 1538 23773
rect 1554 23709 1618 23773
rect 1634 23709 1698 23773
rect 1714 23709 1778 23773
rect 1794 23709 1858 23773
rect 1874 23709 1938 23773
rect 1954 23709 2018 23773
rect 2034 23709 2098 23773
rect 2114 23728 2170 23773
rect 2170 23728 2178 23773
rect 2194 23728 2226 23773
rect 2226 23728 2252 23773
rect 2252 23728 2258 23773
rect 2274 23728 2308 23773
rect 2308 23728 2334 23773
rect 2334 23728 2338 23773
rect 2354 23728 2390 23773
rect 2390 23728 2416 23773
rect 2416 23728 2418 23773
rect 2434 23728 2472 23773
rect 2472 23728 2498 23773
rect 2114 23709 2178 23728
rect 2194 23709 2258 23728
rect 2274 23709 2338 23728
rect 2354 23709 2418 23728
rect 2434 23709 2498 23728
rect 1474 23627 1538 23691
rect 1554 23627 1618 23691
rect 1634 23627 1698 23691
rect 1714 23627 1778 23691
rect 1794 23627 1858 23691
rect 1874 23627 1938 23691
rect 1954 23627 2018 23691
rect 2034 23627 2098 23691
rect 2114 23646 2170 23691
rect 2170 23646 2178 23691
rect 2194 23646 2226 23691
rect 2226 23646 2252 23691
rect 2252 23646 2258 23691
rect 2274 23646 2308 23691
rect 2308 23646 2334 23691
rect 2334 23646 2338 23691
rect 2354 23646 2390 23691
rect 2390 23646 2416 23691
rect 2416 23646 2418 23691
rect 2434 23646 2472 23691
rect 2472 23646 2498 23691
rect 2114 23627 2178 23646
rect 2194 23627 2258 23646
rect 2274 23627 2338 23646
rect 2354 23627 2418 23646
rect 2434 23627 2498 23646
rect 1474 23545 1538 23609
rect 1554 23545 1618 23609
rect 1634 23545 1698 23609
rect 1714 23545 1778 23609
rect 1794 23545 1858 23609
rect 1874 23545 1938 23609
rect 1954 23545 2018 23609
rect 2034 23545 2098 23609
rect 2114 23564 2170 23609
rect 2170 23564 2178 23609
rect 2194 23564 2226 23609
rect 2226 23564 2252 23609
rect 2252 23564 2258 23609
rect 2274 23564 2308 23609
rect 2308 23564 2334 23609
rect 2334 23564 2338 23609
rect 2354 23564 2390 23609
rect 2390 23564 2416 23609
rect 2416 23564 2418 23609
rect 2434 23564 2472 23609
rect 2472 23564 2498 23609
rect 2114 23545 2178 23564
rect 2194 23545 2258 23564
rect 2274 23545 2338 23564
rect 2354 23545 2418 23564
rect 2434 23545 2498 23564
rect 1474 23463 1538 23527
rect 1554 23463 1618 23527
rect 1634 23463 1698 23527
rect 1714 23463 1778 23527
rect 1794 23463 1858 23527
rect 1874 23463 1938 23527
rect 1954 23463 2018 23527
rect 2034 23463 2098 23527
rect 2114 23482 2170 23527
rect 2170 23482 2178 23527
rect 2194 23482 2226 23527
rect 2226 23482 2252 23527
rect 2252 23482 2258 23527
rect 2274 23482 2308 23527
rect 2308 23482 2334 23527
rect 2334 23482 2338 23527
rect 2354 23482 2390 23527
rect 2390 23482 2416 23527
rect 2416 23482 2418 23527
rect 2434 23482 2472 23527
rect 2472 23482 2498 23527
rect 2114 23463 2178 23482
rect 2194 23463 2258 23482
rect 2274 23463 2338 23482
rect 2354 23463 2418 23482
rect 2434 23463 2498 23482
rect 1474 23381 1538 23445
rect 1554 23381 1618 23445
rect 1634 23381 1698 23445
rect 1714 23381 1778 23445
rect 1794 23381 1858 23445
rect 1874 23381 1938 23445
rect 1954 23381 2018 23445
rect 2034 23381 2098 23445
rect 2114 23400 2170 23445
rect 2170 23400 2178 23445
rect 2194 23400 2226 23445
rect 2226 23400 2252 23445
rect 2252 23400 2258 23445
rect 2274 23400 2308 23445
rect 2308 23400 2334 23445
rect 2334 23400 2338 23445
rect 2354 23400 2390 23445
rect 2390 23400 2416 23445
rect 2416 23400 2418 23445
rect 2434 23400 2472 23445
rect 2472 23400 2498 23445
rect 2114 23381 2178 23400
rect 2194 23381 2258 23400
rect 2274 23381 2338 23400
rect 2354 23381 2418 23400
rect 2434 23381 2498 23400
rect 1474 23299 1538 23363
rect 1554 23299 1618 23363
rect 1634 23299 1698 23363
rect 1714 23299 1778 23363
rect 1794 23299 1858 23363
rect 1874 23299 1938 23363
rect 1954 23299 2018 23363
rect 2034 23299 2098 23363
rect 2114 23318 2170 23363
rect 2170 23318 2178 23363
rect 2194 23318 2226 23363
rect 2226 23318 2252 23363
rect 2252 23318 2258 23363
rect 2274 23318 2308 23363
rect 2308 23318 2334 23363
rect 2334 23318 2338 23363
rect 2354 23318 2390 23363
rect 2390 23318 2416 23363
rect 2416 23318 2418 23363
rect 2434 23318 2472 23363
rect 2472 23318 2498 23363
rect 2114 23299 2178 23318
rect 2194 23299 2258 23318
rect 2274 23299 2338 23318
rect 2354 23299 2418 23318
rect 2434 23299 2498 23318
rect 1474 23217 1538 23281
rect 1554 23217 1618 23281
rect 1634 23217 1698 23281
rect 1714 23217 1778 23281
rect 1794 23217 1858 23281
rect 1874 23217 1938 23281
rect 1954 23217 2018 23281
rect 2034 23217 2098 23281
rect 2114 23236 2170 23281
rect 2170 23236 2178 23281
rect 2194 23236 2226 23281
rect 2226 23236 2252 23281
rect 2252 23236 2258 23281
rect 2274 23236 2308 23281
rect 2308 23236 2334 23281
rect 2334 23236 2338 23281
rect 2354 23236 2390 23281
rect 2390 23236 2416 23281
rect 2416 23236 2418 23281
rect 2434 23236 2472 23281
rect 2472 23236 2498 23281
rect 2114 23217 2178 23236
rect 2194 23217 2258 23236
rect 2274 23217 2338 23236
rect 2354 23217 2418 23236
rect 2434 23217 2498 23236
rect 1474 23135 1538 23199
rect 1554 23135 1618 23199
rect 1634 23135 1698 23199
rect 1714 23135 1778 23199
rect 1794 23135 1858 23199
rect 1874 23135 1938 23199
rect 1954 23135 2018 23199
rect 2034 23135 2098 23199
rect 2114 23154 2170 23199
rect 2170 23154 2178 23199
rect 2194 23154 2226 23199
rect 2226 23154 2252 23199
rect 2252 23154 2258 23199
rect 2274 23154 2308 23199
rect 2308 23154 2334 23199
rect 2334 23154 2338 23199
rect 2354 23154 2390 23199
rect 2390 23154 2416 23199
rect 2416 23154 2418 23199
rect 2434 23154 2472 23199
rect 2472 23154 2498 23199
rect 2114 23135 2178 23154
rect 2194 23135 2258 23154
rect 2274 23135 2338 23154
rect 2354 23135 2418 23154
rect 2434 23135 2498 23154
rect 1474 23053 1538 23117
rect 1554 23053 1618 23117
rect 1634 23053 1698 23117
rect 1714 23053 1778 23117
rect 1794 23053 1858 23117
rect 1874 23053 1938 23117
rect 1954 23053 2018 23117
rect 2034 23053 2098 23117
rect 2114 23053 2178 23117
rect 2194 23053 2258 23117
rect 2274 23053 2338 23117
rect 2354 23053 2418 23117
rect 2434 23053 2498 23117
rect 1474 22971 1538 23035
rect 1554 22971 1618 23035
rect 1634 22971 1698 23035
rect 1714 22971 1778 23035
rect 1794 22971 1858 23035
rect 1874 22971 1938 23035
rect 1954 22971 2018 23035
rect 2034 22971 2098 23035
rect 2114 22971 2178 23035
rect 2194 22971 2258 23035
rect 2274 22971 2338 23035
rect 2354 22971 2418 23035
rect 2434 22971 2498 23035
rect 1474 22889 1538 22953
rect 1554 22889 1618 22953
rect 1634 22889 1698 22953
rect 1714 22889 1778 22953
rect 1794 22889 1858 22953
rect 1874 22889 1938 22953
rect 1954 22889 2018 22953
rect 2034 22889 2098 22953
rect 2114 22889 2178 22953
rect 2194 22889 2258 22953
rect 2274 22889 2338 22953
rect 2354 22889 2418 22953
rect 2434 22889 2498 22953
rect 1474 22807 1538 22871
rect 1554 22807 1618 22871
rect 1634 22807 1698 22871
rect 1714 22807 1778 22871
rect 1794 22807 1858 22871
rect 1874 22807 1938 22871
rect 1954 22807 2018 22871
rect 2034 22807 2098 22871
rect 2114 22807 2178 22871
rect 2194 22807 2258 22871
rect 2274 22807 2338 22871
rect 2354 22807 2418 22871
rect 2434 22807 2498 22871
rect 1474 22725 1538 22789
rect 1554 22725 1618 22789
rect 1634 22725 1698 22789
rect 1714 22725 1778 22789
rect 1794 22725 1858 22789
rect 1874 22725 1938 22789
rect 1954 22725 2018 22789
rect 2034 22725 2098 22789
rect 2114 22725 2178 22789
rect 2194 22725 2258 22789
rect 2274 22725 2338 22789
rect 2354 22725 2418 22789
rect 2434 22725 2498 22789
rect 1474 22643 1538 22707
rect 1554 22643 1618 22707
rect 1634 22643 1698 22707
rect 1714 22643 1778 22707
rect 1794 22643 1858 22707
rect 1874 22643 1938 22707
rect 1954 22643 2018 22707
rect 2034 22643 2098 22707
rect 2114 22643 2178 22707
rect 2194 22643 2258 22707
rect 2274 22643 2338 22707
rect 2354 22643 2418 22707
rect 2434 22643 2498 22707
rect 1474 22561 1538 22625
rect 1554 22561 1618 22625
rect 1634 22561 1698 22625
rect 1714 22561 1778 22625
rect 1794 22561 1858 22625
rect 1874 22561 1938 22625
rect 1954 22561 2018 22625
rect 2034 22561 2098 22625
rect 2114 22561 2178 22625
rect 2194 22561 2258 22625
rect 2274 22561 2338 22625
rect 2354 22561 2418 22625
rect 2434 22561 2498 22625
rect 1474 22479 1538 22543
rect 1554 22479 1618 22543
rect 1634 22479 1698 22543
rect 1714 22479 1778 22543
rect 1794 22479 1858 22543
rect 1874 22479 1938 22543
rect 1954 22479 2018 22543
rect 2034 22479 2098 22543
rect 2114 22479 2178 22543
rect 2194 22479 2258 22543
rect 2274 22479 2338 22543
rect 2354 22479 2418 22543
rect 2434 22479 2498 22543
rect 1474 22397 1538 22461
rect 1554 22397 1618 22461
rect 1634 22397 1698 22461
rect 1714 22397 1778 22461
rect 1794 22397 1858 22461
rect 1874 22397 1938 22461
rect 1954 22397 2018 22461
rect 2034 22397 2098 22461
rect 2114 22397 2178 22461
rect 2194 22397 2258 22461
rect 2274 22397 2338 22461
rect 2354 22397 2418 22461
rect 2434 22397 2498 22461
rect 1474 22315 1538 22379
rect 1554 22315 1618 22379
rect 1634 22315 1698 22379
rect 1714 22315 1778 22379
rect 1794 22315 1858 22379
rect 1874 22315 1938 22379
rect 1954 22315 2018 22379
rect 2034 22315 2098 22379
rect 2114 22315 2178 22379
rect 2194 22315 2258 22379
rect 2274 22315 2338 22379
rect 2354 22315 2418 22379
rect 2434 22315 2498 22379
rect 1474 22233 1538 22297
rect 1554 22233 1618 22297
rect 1634 22233 1698 22297
rect 1714 22233 1778 22297
rect 1794 22233 1858 22297
rect 1874 22233 1938 22297
rect 1954 22233 2018 22297
rect 2034 22233 2098 22297
rect 2114 22233 2178 22297
rect 2194 22233 2258 22297
rect 2274 22233 2338 22297
rect 2354 22233 2418 22297
rect 2434 22233 2498 22297
rect 1474 22151 1538 22215
rect 1554 22151 1618 22215
rect 1634 22151 1698 22215
rect 1714 22151 1778 22215
rect 1794 22151 1858 22215
rect 1874 22151 1938 22215
rect 1954 22151 2018 22215
rect 2034 22151 2098 22215
rect 2114 22151 2178 22215
rect 2194 22151 2258 22215
rect 2274 22151 2338 22215
rect 2354 22151 2418 22215
rect 2434 22151 2498 22215
rect 1474 22069 1538 22133
rect 1554 22069 1618 22133
rect 1634 22069 1698 22133
rect 1714 22069 1778 22133
rect 1794 22069 1858 22133
rect 1874 22069 1938 22133
rect 1954 22069 2018 22133
rect 2034 22069 2098 22133
rect 2114 22069 2178 22133
rect 2194 22069 2258 22133
rect 2274 22069 2338 22133
rect 2354 22069 2418 22133
rect 2434 22069 2498 22133
rect 1474 21987 1538 22051
rect 1554 21987 1618 22051
rect 1634 21987 1698 22051
rect 1714 21987 1778 22051
rect 1794 21987 1858 22051
rect 1874 21987 1938 22051
rect 1954 21987 2018 22051
rect 2034 21987 2098 22051
rect 2114 21987 2178 22051
rect 2194 21987 2258 22051
rect 2274 21987 2338 22051
rect 2354 21987 2418 22051
rect 2434 21987 2498 22051
rect 1474 21904 1538 21968
rect 1554 21904 1618 21968
rect 1634 21904 1698 21968
rect 1714 21904 1778 21968
rect 1794 21904 1858 21968
rect 1874 21904 1938 21968
rect 1954 21904 2018 21968
rect 2034 21904 2098 21968
rect 2114 21904 2178 21968
rect 2194 21904 2258 21968
rect 2274 21904 2338 21968
rect 2354 21904 2418 21968
rect 2434 21904 2498 21968
rect 1474 21821 1538 21885
rect 1554 21821 1618 21885
rect 1634 21821 1698 21885
rect 1714 21821 1778 21885
rect 1794 21821 1858 21885
rect 1874 21821 1938 21885
rect 1954 21821 2018 21885
rect 2034 21821 2098 21885
rect 2114 21821 2178 21885
rect 2194 21821 2258 21885
rect 2274 21821 2338 21885
rect 2354 21821 2418 21885
rect 2434 21821 2498 21885
rect 1474 21738 1538 21802
rect 1554 21738 1618 21802
rect 1634 21738 1698 21802
rect 1714 21738 1778 21802
rect 1794 21738 1858 21802
rect 1874 21738 1938 21802
rect 1954 21738 2018 21802
rect 2034 21738 2098 21802
rect 2114 21738 2178 21802
rect 2194 21738 2258 21802
rect 2274 21738 2338 21802
rect 2354 21738 2418 21802
rect 2434 21738 2498 21802
rect 1474 21655 1538 21719
rect 1554 21655 1618 21719
rect 1634 21655 1698 21719
rect 1714 21655 1778 21719
rect 1794 21655 1858 21719
rect 1874 21655 1938 21719
rect 1954 21655 2018 21719
rect 2034 21655 2098 21719
rect 2114 21655 2178 21719
rect 2194 21655 2258 21719
rect 2274 21655 2338 21719
rect 2354 21655 2418 21719
rect 2434 21655 2498 21719
rect 1474 21572 1538 21636
rect 1554 21572 1618 21636
rect 1634 21572 1698 21636
rect 1714 21572 1778 21636
rect 1794 21572 1858 21636
rect 1874 21572 1938 21636
rect 1954 21572 2018 21636
rect 2034 21572 2098 21636
rect 2114 21572 2178 21636
rect 2194 21572 2258 21636
rect 2274 21572 2338 21636
rect 2354 21572 2418 21636
rect 2434 21572 2498 21636
rect 1474 21489 1538 21553
rect 1554 21489 1618 21553
rect 1634 21489 1698 21553
rect 1714 21489 1778 21553
rect 1794 21489 1858 21553
rect 1874 21489 1938 21553
rect 1954 21489 2018 21553
rect 2034 21489 2098 21553
rect 2114 21489 2178 21553
rect 2194 21489 2258 21553
rect 2274 21489 2338 21553
rect 2354 21489 2418 21553
rect 2434 21489 2498 21553
rect 1474 21406 1538 21470
rect 1554 21406 1618 21470
rect 1634 21406 1698 21470
rect 1714 21406 1778 21470
rect 1794 21406 1858 21470
rect 1874 21406 1938 21470
rect 1954 21406 2018 21470
rect 2034 21406 2098 21470
rect 2114 21406 2178 21470
rect 2194 21406 2258 21470
rect 2274 21406 2338 21470
rect 2354 21406 2418 21470
rect 2434 21406 2498 21470
rect 1474 21323 1538 21387
rect 1554 21323 1618 21387
rect 1634 21323 1698 21387
rect 1714 21323 1778 21387
rect 1794 21323 1858 21387
rect 1874 21323 1938 21387
rect 1954 21323 2018 21387
rect 2034 21323 2098 21387
rect 2114 21323 2178 21387
rect 2194 21323 2258 21387
rect 2274 21323 2338 21387
rect 2354 21323 2418 21387
rect 2434 21323 2498 21387
rect 14508 31164 15292 31178
rect 14508 31108 14514 31164
rect 14514 31108 14570 31164
rect 14570 31108 14594 31164
rect 14594 31108 14650 31164
rect 14650 31108 14674 31164
rect 14674 31108 14730 31164
rect 14730 31108 14754 31164
rect 14754 31108 14810 31164
rect 14810 31108 14834 31164
rect 14834 31108 14890 31164
rect 14890 31108 14914 31164
rect 14914 31108 14970 31164
rect 14970 31108 14994 31164
rect 14994 31108 15050 31164
rect 15050 31108 15074 31164
rect 15074 31108 15130 31164
rect 15130 31108 15154 31164
rect 15154 31108 15210 31164
rect 15210 31108 15234 31164
rect 15234 31108 15290 31164
rect 15290 31108 15292 31164
rect 14508 31082 15292 31108
rect 14508 31026 14514 31082
rect 14514 31026 14570 31082
rect 14570 31026 14594 31082
rect 14594 31026 14650 31082
rect 14650 31026 14674 31082
rect 14674 31026 14730 31082
rect 14730 31026 14754 31082
rect 14754 31026 14810 31082
rect 14810 31026 14834 31082
rect 14834 31026 14890 31082
rect 14890 31026 14914 31082
rect 14914 31026 14970 31082
rect 14970 31026 14994 31082
rect 14994 31026 15050 31082
rect 15050 31026 15074 31082
rect 15074 31026 15130 31082
rect 15130 31026 15154 31082
rect 15154 31026 15210 31082
rect 15210 31026 15234 31082
rect 15234 31026 15290 31082
rect 15290 31026 15292 31082
rect 14508 31000 15292 31026
rect 14508 30944 14514 31000
rect 14514 30944 14570 31000
rect 14570 30944 14594 31000
rect 14594 30944 14650 31000
rect 14650 30944 14674 31000
rect 14674 30944 14730 31000
rect 14730 30944 14754 31000
rect 14754 30944 14810 31000
rect 14810 30944 14834 31000
rect 14834 30944 14890 31000
rect 14890 30944 14914 31000
rect 14914 30944 14970 31000
rect 14970 30944 14994 31000
rect 14994 30944 15050 31000
rect 15050 30944 15074 31000
rect 15074 30944 15130 31000
rect 15130 30944 15154 31000
rect 15154 30944 15210 31000
rect 15210 30944 15234 31000
rect 15234 30944 15290 31000
rect 15290 30944 15292 31000
rect 14508 30918 15292 30944
rect 14508 30862 14514 30918
rect 14514 30862 14570 30918
rect 14570 30862 14594 30918
rect 14594 30862 14650 30918
rect 14650 30862 14674 30918
rect 14674 30862 14730 30918
rect 14730 30862 14754 30918
rect 14754 30862 14810 30918
rect 14810 30862 14834 30918
rect 14834 30862 14890 30918
rect 14890 30862 14914 30918
rect 14914 30862 14970 30918
rect 14970 30862 14994 30918
rect 14994 30862 15050 30918
rect 15050 30862 15074 30918
rect 15074 30862 15130 30918
rect 15130 30862 15154 30918
rect 15154 30862 15210 30918
rect 15210 30862 15234 30918
rect 15234 30862 15290 30918
rect 15290 30862 15292 30918
rect 14508 30836 15292 30862
rect 14508 30780 14514 30836
rect 14514 30780 14570 30836
rect 14570 30780 14594 30836
rect 14594 30780 14650 30836
rect 14650 30780 14674 30836
rect 14674 30780 14730 30836
rect 14730 30780 14754 30836
rect 14754 30780 14810 30836
rect 14810 30780 14834 30836
rect 14834 30780 14890 30836
rect 14890 30780 14914 30836
rect 14914 30780 14970 30836
rect 14970 30780 14994 30836
rect 14994 30780 15050 30836
rect 15050 30780 15074 30836
rect 15074 30780 15130 30836
rect 15130 30780 15154 30836
rect 15154 30780 15210 30836
rect 15210 30780 15234 30836
rect 15234 30780 15290 30836
rect 15290 30780 15292 30836
rect 14508 30753 15292 30780
rect 14508 30697 14514 30753
rect 14514 30697 14570 30753
rect 14570 30697 14594 30753
rect 14594 30697 14650 30753
rect 14650 30697 14674 30753
rect 14674 30697 14730 30753
rect 14730 30697 14754 30753
rect 14754 30697 14810 30753
rect 14810 30697 14834 30753
rect 14834 30697 14890 30753
rect 14890 30697 14914 30753
rect 14914 30697 14970 30753
rect 14970 30697 14994 30753
rect 14994 30697 15050 30753
rect 15050 30697 15074 30753
rect 15074 30697 15130 30753
rect 15130 30697 15154 30753
rect 15154 30697 15210 30753
rect 15210 30697 15234 30753
rect 15234 30697 15290 30753
rect 15290 30697 15292 30753
rect 14508 30670 15292 30697
rect 14508 30614 14514 30670
rect 14514 30614 14570 30670
rect 14570 30614 14594 30670
rect 14594 30614 14650 30670
rect 14650 30614 14674 30670
rect 14674 30614 14730 30670
rect 14730 30614 14754 30670
rect 14754 30614 14810 30670
rect 14810 30614 14834 30670
rect 14834 30614 14890 30670
rect 14890 30614 14914 30670
rect 14914 30614 14970 30670
rect 14970 30614 14994 30670
rect 14994 30614 15050 30670
rect 15050 30614 15074 30670
rect 15074 30614 15130 30670
rect 15130 30614 15154 30670
rect 15154 30614 15210 30670
rect 15210 30614 15234 30670
rect 15234 30614 15290 30670
rect 15290 30614 15292 30670
rect 14508 30587 15292 30614
rect 14508 30531 14514 30587
rect 14514 30531 14570 30587
rect 14570 30531 14594 30587
rect 14594 30531 14650 30587
rect 14650 30531 14674 30587
rect 14674 30531 14730 30587
rect 14730 30531 14754 30587
rect 14754 30531 14810 30587
rect 14810 30531 14834 30587
rect 14834 30531 14890 30587
rect 14890 30531 14914 30587
rect 14914 30531 14970 30587
rect 14970 30531 14994 30587
rect 14994 30531 15050 30587
rect 15050 30531 15074 30587
rect 15074 30531 15130 30587
rect 15130 30531 15154 30587
rect 15154 30531 15210 30587
rect 15210 30531 15234 30587
rect 15234 30531 15290 30587
rect 15290 30531 15292 30587
rect 14508 30504 15292 30531
rect 14508 30448 14514 30504
rect 14514 30448 14570 30504
rect 14570 30448 14594 30504
rect 14594 30448 14650 30504
rect 14650 30448 14674 30504
rect 14674 30448 14730 30504
rect 14730 30448 14754 30504
rect 14754 30448 14810 30504
rect 14810 30448 14834 30504
rect 14834 30448 14890 30504
rect 14890 30448 14914 30504
rect 14914 30448 14970 30504
rect 14970 30448 14994 30504
rect 14994 30448 15050 30504
rect 15050 30448 15074 30504
rect 15074 30448 15130 30504
rect 15130 30448 15154 30504
rect 15154 30448 15210 30504
rect 15210 30448 15234 30504
rect 15234 30448 15290 30504
rect 15290 30448 15292 30504
rect 14508 30421 15292 30448
rect 14508 30365 14514 30421
rect 14514 30365 14570 30421
rect 14570 30365 14594 30421
rect 14594 30365 14650 30421
rect 14650 30365 14674 30421
rect 14674 30365 14730 30421
rect 14730 30365 14754 30421
rect 14754 30365 14810 30421
rect 14810 30365 14834 30421
rect 14834 30365 14890 30421
rect 14890 30365 14914 30421
rect 14914 30365 14970 30421
rect 14970 30365 14994 30421
rect 14994 30365 15050 30421
rect 15050 30365 15074 30421
rect 15074 30365 15130 30421
rect 15130 30365 15154 30421
rect 15154 30365 15210 30421
rect 15210 30365 15234 30421
rect 15234 30365 15290 30421
rect 15290 30365 15292 30421
rect 14508 30338 15292 30365
rect 14508 30282 14514 30338
rect 14514 30282 14570 30338
rect 14570 30282 14594 30338
rect 14594 30282 14650 30338
rect 14650 30282 14674 30338
rect 14674 30282 14730 30338
rect 14730 30282 14754 30338
rect 14754 30282 14810 30338
rect 14810 30282 14834 30338
rect 14834 30282 14890 30338
rect 14890 30282 14914 30338
rect 14914 30282 14970 30338
rect 14970 30282 14994 30338
rect 14994 30282 15050 30338
rect 15050 30282 15074 30338
rect 15074 30282 15130 30338
rect 15130 30282 15154 30338
rect 15154 30282 15210 30338
rect 15210 30282 15234 30338
rect 15234 30282 15290 30338
rect 15290 30282 15292 30338
rect 14508 30255 15292 30282
rect 14508 30199 14514 30255
rect 14514 30199 14570 30255
rect 14570 30199 14594 30255
rect 14594 30199 14650 30255
rect 14650 30199 14674 30255
rect 14674 30199 14730 30255
rect 14730 30199 14754 30255
rect 14754 30199 14810 30255
rect 14810 30199 14834 30255
rect 14834 30199 14890 30255
rect 14890 30199 14914 30255
rect 14914 30199 14970 30255
rect 14970 30199 14994 30255
rect 14994 30199 15050 30255
rect 15050 30199 15074 30255
rect 15074 30199 15130 30255
rect 15130 30199 15154 30255
rect 15154 30199 15210 30255
rect 15210 30199 15234 30255
rect 15234 30199 15290 30255
rect 15290 30199 15292 30255
rect 14508 30172 15292 30199
rect 14508 30116 14514 30172
rect 14514 30116 14570 30172
rect 14570 30116 14594 30172
rect 14594 30116 14650 30172
rect 14650 30116 14674 30172
rect 14674 30116 14730 30172
rect 14730 30116 14754 30172
rect 14754 30116 14810 30172
rect 14810 30116 14834 30172
rect 14834 30116 14890 30172
rect 14890 30116 14914 30172
rect 14914 30116 14970 30172
rect 14970 30116 14994 30172
rect 14994 30116 15050 30172
rect 15050 30116 15074 30172
rect 15074 30116 15130 30172
rect 15130 30116 15154 30172
rect 15154 30116 15210 30172
rect 15210 30116 15234 30172
rect 15234 30116 15290 30172
rect 15290 30116 15292 30172
rect 14508 30089 15292 30116
rect 14508 30033 14514 30089
rect 14514 30033 14570 30089
rect 14570 30033 14594 30089
rect 14594 30033 14650 30089
rect 14650 30033 14674 30089
rect 14674 30033 14730 30089
rect 14730 30033 14754 30089
rect 14754 30033 14810 30089
rect 14810 30033 14834 30089
rect 14834 30033 14890 30089
rect 14890 30033 14914 30089
rect 14914 30033 14970 30089
rect 14970 30033 14994 30089
rect 14994 30033 15050 30089
rect 15050 30033 15074 30089
rect 15074 30033 15130 30089
rect 15130 30033 15154 30089
rect 15154 30033 15210 30089
rect 15210 30033 15234 30089
rect 15234 30033 15290 30089
rect 15290 30033 15292 30089
rect 14508 30006 15292 30033
rect 14508 29950 14514 30006
rect 14514 29950 14570 30006
rect 14570 29950 14594 30006
rect 14594 29950 14650 30006
rect 14650 29950 14674 30006
rect 14674 29950 14730 30006
rect 14730 29950 14754 30006
rect 14754 29950 14810 30006
rect 14810 29950 14834 30006
rect 14834 29950 14890 30006
rect 14890 29950 14914 30006
rect 14914 29950 14970 30006
rect 14970 29950 14994 30006
rect 14994 29950 15050 30006
rect 15050 29950 15074 30006
rect 15074 29950 15130 30006
rect 15130 29950 15154 30006
rect 15154 29950 15210 30006
rect 15210 29950 15234 30006
rect 15234 29950 15290 30006
rect 15290 29950 15292 30006
rect 14508 29923 15292 29950
rect 14508 29867 14514 29923
rect 14514 29867 14570 29923
rect 14570 29867 14594 29923
rect 14594 29867 14650 29923
rect 14650 29867 14674 29923
rect 14674 29867 14730 29923
rect 14730 29867 14754 29923
rect 14754 29867 14810 29923
rect 14810 29867 14834 29923
rect 14834 29867 14890 29923
rect 14890 29867 14914 29923
rect 14914 29867 14970 29923
rect 14970 29867 14994 29923
rect 14994 29867 15050 29923
rect 15050 29867 15074 29923
rect 15074 29867 15130 29923
rect 15130 29867 15154 29923
rect 15154 29867 15210 29923
rect 15210 29867 15234 29923
rect 15234 29867 15290 29923
rect 15290 29867 15292 29923
rect 14508 29840 15292 29867
rect 14508 29784 14514 29840
rect 14514 29784 14570 29840
rect 14570 29784 14594 29840
rect 14594 29784 14650 29840
rect 14650 29784 14674 29840
rect 14674 29784 14730 29840
rect 14730 29784 14754 29840
rect 14754 29784 14810 29840
rect 14810 29784 14834 29840
rect 14834 29784 14890 29840
rect 14890 29784 14914 29840
rect 14914 29784 14970 29840
rect 14970 29784 14994 29840
rect 14994 29784 15050 29840
rect 15050 29784 15074 29840
rect 15074 29784 15130 29840
rect 15130 29784 15154 29840
rect 15154 29784 15210 29840
rect 15210 29784 15234 29840
rect 15234 29784 15290 29840
rect 15290 29784 15292 29840
rect 14508 29757 15292 29784
rect 14508 29701 14514 29757
rect 14514 29701 14570 29757
rect 14570 29701 14594 29757
rect 14594 29701 14650 29757
rect 14650 29701 14674 29757
rect 14674 29701 14730 29757
rect 14730 29701 14754 29757
rect 14754 29701 14810 29757
rect 14810 29701 14834 29757
rect 14834 29701 14890 29757
rect 14890 29701 14914 29757
rect 14914 29701 14970 29757
rect 14970 29701 14994 29757
rect 14994 29701 15050 29757
rect 15050 29701 15074 29757
rect 15074 29701 15130 29757
rect 15130 29701 15154 29757
rect 15154 29701 15210 29757
rect 15210 29701 15234 29757
rect 15234 29701 15290 29757
rect 15290 29701 15292 29757
rect 14508 29674 15292 29701
rect 14508 29618 14514 29674
rect 14514 29618 14570 29674
rect 14570 29618 14594 29674
rect 14594 29618 14650 29674
rect 14650 29618 14674 29674
rect 14674 29618 14730 29674
rect 14730 29618 14754 29674
rect 14754 29618 14810 29674
rect 14810 29618 14834 29674
rect 14834 29618 14890 29674
rect 14890 29618 14914 29674
rect 14914 29618 14970 29674
rect 14970 29618 14994 29674
rect 14994 29618 15050 29674
rect 15050 29618 15074 29674
rect 15074 29618 15130 29674
rect 15130 29618 15154 29674
rect 15154 29618 15210 29674
rect 15210 29618 15234 29674
rect 15234 29618 15290 29674
rect 15290 29618 15292 29674
rect 14508 29591 15292 29618
rect 14508 29535 14514 29591
rect 14514 29535 14570 29591
rect 14570 29535 14594 29591
rect 14594 29535 14650 29591
rect 14650 29535 14674 29591
rect 14674 29535 14730 29591
rect 14730 29535 14754 29591
rect 14754 29535 14810 29591
rect 14810 29535 14834 29591
rect 14834 29535 14890 29591
rect 14890 29535 14914 29591
rect 14914 29535 14970 29591
rect 14970 29535 14994 29591
rect 14994 29535 15050 29591
rect 15050 29535 15074 29591
rect 15074 29535 15130 29591
rect 15130 29535 15154 29591
rect 15154 29535 15210 29591
rect 15210 29535 15234 29591
rect 15234 29535 15290 29591
rect 15290 29535 15292 29591
rect 14508 29508 15292 29535
rect 14508 29452 14514 29508
rect 14514 29452 14570 29508
rect 14570 29452 14594 29508
rect 14594 29452 14650 29508
rect 14650 29452 14674 29508
rect 14674 29452 14730 29508
rect 14730 29452 14754 29508
rect 14754 29452 14810 29508
rect 14810 29452 14834 29508
rect 14834 29452 14890 29508
rect 14890 29452 14914 29508
rect 14914 29452 14970 29508
rect 14970 29452 14994 29508
rect 14994 29452 15050 29508
rect 15050 29452 15074 29508
rect 15074 29452 15130 29508
rect 15130 29452 15154 29508
rect 15154 29452 15210 29508
rect 15210 29452 15234 29508
rect 15234 29452 15290 29508
rect 15290 29452 15292 29508
rect 14508 29425 15292 29452
rect 14508 29369 14514 29425
rect 14514 29369 14570 29425
rect 14570 29369 14594 29425
rect 14594 29369 14650 29425
rect 14650 29369 14674 29425
rect 14674 29369 14730 29425
rect 14730 29369 14754 29425
rect 14754 29369 14810 29425
rect 14810 29369 14834 29425
rect 14834 29369 14890 29425
rect 14890 29369 14914 29425
rect 14914 29369 14970 29425
rect 14970 29369 14994 29425
rect 14994 29369 15050 29425
rect 15050 29369 15074 29425
rect 15074 29369 15130 29425
rect 15130 29369 15154 29425
rect 15154 29369 15210 29425
rect 15210 29369 15234 29425
rect 15234 29369 15290 29425
rect 15290 29369 15292 29425
rect 14508 29342 15292 29369
rect 14508 29286 14514 29342
rect 14514 29286 14570 29342
rect 14570 29286 14594 29342
rect 14594 29286 14650 29342
rect 14650 29286 14674 29342
rect 14674 29286 14730 29342
rect 14730 29286 14754 29342
rect 14754 29286 14810 29342
rect 14810 29286 14834 29342
rect 14834 29286 14890 29342
rect 14890 29286 14914 29342
rect 14914 29286 14970 29342
rect 14970 29286 14994 29342
rect 14994 29286 15050 29342
rect 15050 29286 15074 29342
rect 15074 29286 15130 29342
rect 15130 29286 15154 29342
rect 15154 29286 15210 29342
rect 15210 29286 15234 29342
rect 15234 29286 15290 29342
rect 15290 29286 15292 29342
rect 14508 29259 15292 29286
rect 14508 29203 14514 29259
rect 14514 29203 14570 29259
rect 14570 29203 14594 29259
rect 14594 29203 14650 29259
rect 14650 29203 14674 29259
rect 14674 29203 14730 29259
rect 14730 29203 14754 29259
rect 14754 29203 14810 29259
rect 14810 29203 14834 29259
rect 14834 29203 14890 29259
rect 14890 29203 14914 29259
rect 14914 29203 14970 29259
rect 14970 29203 14994 29259
rect 14994 29203 15050 29259
rect 15050 29203 15074 29259
rect 15074 29203 15130 29259
rect 15130 29203 15154 29259
rect 15154 29203 15210 29259
rect 15210 29203 15234 29259
rect 15234 29203 15290 29259
rect 15290 29203 15292 29259
rect 14508 29176 15292 29203
rect 14508 29120 14514 29176
rect 14514 29120 14570 29176
rect 14570 29120 14594 29176
rect 14594 29120 14650 29176
rect 14650 29120 14674 29176
rect 14674 29120 14730 29176
rect 14730 29120 14754 29176
rect 14754 29120 14810 29176
rect 14810 29120 14834 29176
rect 14834 29120 14890 29176
rect 14890 29120 14914 29176
rect 14914 29120 14970 29176
rect 14970 29120 14994 29176
rect 14994 29120 15050 29176
rect 15050 29120 15074 29176
rect 15074 29120 15130 29176
rect 15130 29120 15154 29176
rect 15154 29120 15210 29176
rect 15210 29120 15234 29176
rect 15234 29120 15290 29176
rect 15290 29120 15292 29176
rect 14508 29093 15292 29120
rect 14508 29037 14514 29093
rect 14514 29037 14570 29093
rect 14570 29037 14594 29093
rect 14594 29037 14650 29093
rect 14650 29037 14674 29093
rect 14674 29037 14730 29093
rect 14730 29037 14754 29093
rect 14754 29037 14810 29093
rect 14810 29037 14834 29093
rect 14834 29037 14890 29093
rect 14890 29037 14914 29093
rect 14914 29037 14970 29093
rect 14970 29037 14994 29093
rect 14994 29037 15050 29093
rect 15050 29037 15074 29093
rect 15074 29037 15130 29093
rect 15130 29037 15154 29093
rect 15154 29037 15210 29093
rect 15210 29037 15234 29093
rect 15234 29037 15290 29093
rect 15290 29037 15292 29093
rect 14508 29034 15292 29037
rect 14508 29010 14572 29017
rect 14508 28954 14514 29010
rect 14514 28954 14570 29010
rect 14570 28954 14572 29010
rect 14508 28953 14572 28954
rect 14588 29010 14652 29017
rect 14588 28954 14594 29010
rect 14594 28954 14650 29010
rect 14650 28954 14652 29010
rect 14588 28953 14652 28954
rect 14668 29010 14732 29017
rect 14668 28954 14674 29010
rect 14674 28954 14730 29010
rect 14730 28954 14732 29010
rect 14668 28953 14732 28954
rect 14748 29010 14812 29017
rect 14748 28954 14754 29010
rect 14754 28954 14810 29010
rect 14810 28954 14812 29010
rect 14748 28953 14812 28954
rect 14828 29010 14892 29017
rect 14828 28954 14834 29010
rect 14834 28954 14890 29010
rect 14890 28954 14892 29010
rect 14828 28953 14892 28954
rect 14908 29010 14972 29017
rect 14908 28954 14914 29010
rect 14914 28954 14970 29010
rect 14970 28954 14972 29010
rect 14908 28953 14972 28954
rect 14988 29010 15052 29017
rect 14988 28954 14994 29010
rect 14994 28954 15050 29010
rect 15050 28954 15052 29010
rect 14988 28953 15052 28954
rect 15068 29010 15132 29017
rect 15068 28954 15074 29010
rect 15074 28954 15130 29010
rect 15130 28954 15132 29010
rect 15068 28953 15132 28954
rect 15148 29010 15212 29017
rect 15148 28954 15154 29010
rect 15154 28954 15210 29010
rect 15210 28954 15212 29010
rect 15148 28953 15212 28954
rect 15228 29010 15292 29017
rect 15228 28954 15234 29010
rect 15234 28954 15290 29010
rect 15290 28954 15292 29010
rect 15228 28953 15292 28954
rect 14508 28927 14572 28936
rect 14508 28872 14514 28927
rect 14514 28872 14570 28927
rect 14570 28872 14572 28927
rect 14588 28927 14652 28936
rect 14588 28872 14594 28927
rect 14594 28872 14650 28927
rect 14650 28872 14652 28927
rect 14668 28927 14732 28936
rect 14668 28872 14674 28927
rect 14674 28872 14730 28927
rect 14730 28872 14732 28927
rect 14748 28927 14812 28936
rect 14748 28872 14754 28927
rect 14754 28872 14810 28927
rect 14810 28872 14812 28927
rect 14828 28927 14892 28936
rect 14828 28872 14834 28927
rect 14834 28872 14890 28927
rect 14890 28872 14892 28927
rect 14908 28927 14972 28936
rect 14908 28872 14914 28927
rect 14914 28872 14970 28927
rect 14970 28872 14972 28927
rect 14988 28927 15052 28936
rect 14988 28872 14994 28927
rect 14994 28872 15050 28927
rect 15050 28872 15052 28927
rect 15068 28927 15132 28936
rect 15068 28872 15074 28927
rect 15074 28872 15130 28927
rect 15130 28872 15132 28927
rect 15148 28927 15212 28936
rect 15148 28872 15154 28927
rect 15154 28872 15210 28927
rect 15210 28872 15212 28927
rect 15228 28927 15292 28936
rect 15228 28872 15234 28927
rect 15234 28872 15290 28927
rect 15290 28872 15292 28927
rect 14521 27574 14585 27593
rect 14521 27529 14522 27574
rect 14522 27529 14578 27574
rect 14578 27529 14585 27574
rect 14611 27574 14675 27593
rect 14611 27529 14612 27574
rect 14612 27529 14668 27574
rect 14668 27529 14675 27574
rect 14701 27574 14765 27593
rect 14701 27529 14702 27574
rect 14702 27529 14758 27574
rect 14758 27529 14765 27574
rect 14791 27574 14855 27593
rect 14881 27574 14945 27593
rect 14971 27574 15035 27593
rect 14791 27529 14847 27574
rect 14847 27529 14855 27574
rect 14881 27529 14936 27574
rect 14936 27529 14945 27574
rect 14971 27529 15025 27574
rect 15025 27529 15035 27574
rect 14521 27488 14585 27512
rect 14521 27448 14522 27488
rect 14522 27448 14578 27488
rect 14578 27448 14585 27488
rect 14611 27488 14675 27512
rect 14611 27448 14612 27488
rect 14612 27448 14668 27488
rect 14668 27448 14675 27488
rect 14701 27488 14765 27512
rect 14701 27448 14702 27488
rect 14702 27448 14758 27488
rect 14758 27448 14765 27488
rect 14791 27488 14855 27512
rect 14881 27488 14945 27512
rect 14971 27488 15035 27512
rect 14791 27448 14847 27488
rect 14847 27448 14855 27488
rect 14881 27448 14936 27488
rect 14936 27448 14945 27488
rect 14971 27448 15025 27488
rect 15025 27448 15035 27488
rect 14521 27402 14585 27431
rect 14521 27367 14522 27402
rect 14522 27367 14578 27402
rect 14578 27367 14585 27402
rect 14611 27402 14675 27431
rect 14611 27367 14612 27402
rect 14612 27367 14668 27402
rect 14668 27367 14675 27402
rect 14701 27402 14765 27431
rect 14701 27367 14702 27402
rect 14702 27367 14758 27402
rect 14758 27367 14765 27402
rect 14791 27402 14855 27431
rect 14881 27402 14945 27431
rect 14971 27402 15035 27431
rect 14791 27367 14847 27402
rect 14847 27367 14855 27402
rect 14881 27367 14936 27402
rect 14936 27367 14945 27402
rect 14971 27367 15025 27402
rect 15025 27367 15035 27402
rect 14521 27346 14522 27350
rect 14522 27346 14578 27350
rect 14578 27346 14585 27350
rect 14521 27316 14585 27346
rect 14521 27286 14522 27316
rect 14522 27286 14578 27316
rect 14578 27286 14585 27316
rect 14611 27346 14612 27350
rect 14612 27346 14668 27350
rect 14668 27346 14675 27350
rect 14611 27316 14675 27346
rect 14611 27286 14612 27316
rect 14612 27286 14668 27316
rect 14668 27286 14675 27316
rect 14701 27346 14702 27350
rect 14702 27346 14758 27350
rect 14758 27346 14765 27350
rect 14701 27316 14765 27346
rect 14701 27286 14702 27316
rect 14702 27286 14758 27316
rect 14758 27286 14765 27316
rect 14791 27346 14847 27350
rect 14847 27346 14855 27350
rect 14881 27346 14936 27350
rect 14936 27346 14945 27350
rect 14971 27346 15025 27350
rect 15025 27346 15035 27350
rect 14791 27316 14855 27346
rect 14881 27316 14945 27346
rect 14971 27316 15035 27346
rect 14791 27286 14847 27316
rect 14847 27286 14855 27316
rect 14881 27286 14936 27316
rect 14936 27286 14945 27316
rect 14971 27286 15025 27316
rect 15025 27286 15035 27316
rect 14521 27260 14522 27268
rect 14522 27260 14578 27268
rect 14578 27260 14585 27268
rect 14521 27230 14585 27260
rect 14521 27204 14522 27230
rect 14522 27204 14578 27230
rect 14578 27204 14585 27230
rect 14611 27260 14612 27268
rect 14612 27260 14668 27268
rect 14668 27260 14675 27268
rect 14611 27230 14675 27260
rect 14611 27204 14612 27230
rect 14612 27204 14668 27230
rect 14668 27204 14675 27230
rect 14701 27260 14702 27268
rect 14702 27260 14758 27268
rect 14758 27260 14765 27268
rect 14701 27230 14765 27260
rect 14701 27204 14702 27230
rect 14702 27204 14758 27230
rect 14758 27204 14765 27230
rect 14791 27260 14847 27268
rect 14847 27260 14855 27268
rect 14881 27260 14936 27268
rect 14936 27260 14945 27268
rect 14971 27260 15025 27268
rect 15025 27260 15035 27268
rect 14791 27230 14855 27260
rect 14881 27230 14945 27260
rect 14971 27230 15035 27260
rect 14791 27204 14847 27230
rect 14847 27204 14855 27230
rect 14881 27204 14936 27230
rect 14936 27204 14945 27230
rect 14971 27204 15025 27230
rect 15025 27204 15035 27230
rect 14521 27174 14522 27186
rect 14522 27174 14578 27186
rect 14578 27174 14585 27186
rect 14521 27144 14585 27174
rect 14521 27122 14522 27144
rect 14522 27122 14578 27144
rect 14578 27122 14585 27144
rect 14611 27174 14612 27186
rect 14612 27174 14668 27186
rect 14668 27174 14675 27186
rect 14611 27144 14675 27174
rect 14611 27122 14612 27144
rect 14612 27122 14668 27144
rect 14668 27122 14675 27144
rect 14701 27174 14702 27186
rect 14702 27174 14758 27186
rect 14758 27174 14765 27186
rect 14701 27144 14765 27174
rect 14701 27122 14702 27144
rect 14702 27122 14758 27144
rect 14758 27122 14765 27144
rect 14791 27174 14847 27186
rect 14847 27174 14855 27186
rect 14881 27174 14936 27186
rect 14936 27174 14945 27186
rect 14971 27174 15025 27186
rect 15025 27174 15035 27186
rect 14791 27144 14855 27174
rect 14881 27144 14945 27174
rect 14971 27144 15035 27174
rect 14791 27122 14847 27144
rect 14847 27122 14855 27144
rect 14881 27122 14936 27144
rect 14936 27122 14945 27144
rect 14971 27122 15025 27144
rect 15025 27122 15035 27144
rect 14521 27088 14522 27104
rect 14522 27088 14578 27104
rect 14578 27088 14585 27104
rect 14521 27040 14585 27088
rect 14611 27088 14612 27104
rect 14612 27088 14668 27104
rect 14668 27088 14675 27104
rect 14611 27040 14675 27088
rect 14701 27088 14702 27104
rect 14702 27088 14758 27104
rect 14758 27088 14765 27104
rect 14701 27040 14765 27088
rect 14791 27088 14847 27104
rect 14847 27088 14855 27104
rect 14881 27088 14936 27104
rect 14936 27088 14945 27104
rect 14971 27088 15025 27104
rect 15025 27088 15035 27104
rect 14791 27040 14855 27088
rect 14881 27040 14945 27088
rect 14971 27040 15035 27088
rect 14510 25766 14565 25809
rect 14565 25766 14574 25809
rect 14510 25745 14574 25766
rect 14602 25766 14603 25809
rect 14603 25766 14659 25809
rect 14659 25766 14666 25809
rect 14602 25745 14666 25766
rect 14694 25766 14697 25809
rect 14697 25766 14753 25809
rect 14753 25766 14758 25809
rect 14694 25745 14758 25766
rect 14786 25766 14791 25809
rect 14791 25766 14847 25809
rect 14847 25766 14850 25809
rect 14786 25745 14850 25766
rect 14878 25766 14885 25809
rect 14885 25766 14941 25809
rect 14941 25766 14942 25809
rect 14878 25745 14942 25766
rect 14970 25766 14979 25809
rect 14979 25766 15034 25809
rect 14970 25745 15034 25766
rect 14510 25685 14565 25729
rect 14565 25685 14574 25729
rect 14510 25665 14574 25685
rect 14602 25685 14603 25729
rect 14603 25685 14659 25729
rect 14659 25685 14666 25729
rect 14602 25665 14666 25685
rect 14694 25685 14697 25729
rect 14697 25685 14753 25729
rect 14753 25685 14758 25729
rect 14694 25665 14758 25685
rect 14786 25685 14791 25729
rect 14791 25685 14847 25729
rect 14847 25685 14850 25729
rect 14786 25665 14850 25685
rect 14878 25685 14885 25729
rect 14885 25685 14941 25729
rect 14941 25685 14942 25729
rect 14878 25665 14942 25685
rect 14970 25685 14979 25729
rect 14979 25685 15034 25729
rect 14970 25665 15034 25685
rect 14510 25604 14565 25648
rect 14565 25604 14574 25648
rect 14510 25584 14574 25604
rect 14602 25604 14603 25648
rect 14603 25604 14659 25648
rect 14659 25604 14666 25648
rect 14602 25584 14666 25604
rect 14694 25604 14697 25648
rect 14697 25604 14753 25648
rect 14753 25604 14758 25648
rect 14694 25584 14758 25604
rect 14786 25604 14791 25648
rect 14791 25604 14847 25648
rect 14847 25604 14850 25648
rect 14786 25584 14850 25604
rect 14878 25604 14885 25648
rect 14885 25604 14941 25648
rect 14941 25604 14942 25648
rect 14878 25584 14942 25604
rect 14970 25604 14979 25648
rect 14979 25604 15034 25648
rect 14970 25584 15034 25604
rect 14510 25523 14565 25567
rect 14565 25523 14574 25567
rect 14510 25503 14574 25523
rect 14602 25523 14603 25567
rect 14603 25523 14659 25567
rect 14659 25523 14666 25567
rect 14602 25503 14666 25523
rect 14694 25523 14697 25567
rect 14697 25523 14753 25567
rect 14753 25523 14758 25567
rect 14694 25503 14758 25523
rect 14786 25523 14791 25567
rect 14791 25523 14847 25567
rect 14847 25523 14850 25567
rect 14786 25503 14850 25523
rect 14878 25523 14885 25567
rect 14885 25523 14941 25567
rect 14941 25523 14942 25567
rect 14878 25503 14942 25523
rect 14970 25523 14979 25567
rect 14979 25523 15034 25567
rect 14970 25503 15034 25523
rect 14510 25442 14565 25486
rect 14565 25442 14574 25486
rect 14510 25422 14574 25442
rect 14602 25442 14603 25486
rect 14603 25442 14659 25486
rect 14659 25442 14666 25486
rect 14602 25422 14666 25442
rect 14694 25442 14697 25486
rect 14697 25442 14753 25486
rect 14753 25442 14758 25486
rect 14694 25422 14758 25442
rect 14786 25442 14791 25486
rect 14791 25442 14847 25486
rect 14847 25442 14850 25486
rect 14786 25422 14850 25442
rect 14878 25442 14885 25486
rect 14885 25442 14941 25486
rect 14941 25442 14942 25486
rect 14878 25422 14942 25442
rect 14970 25442 14979 25486
rect 14979 25442 15034 25486
rect 14970 25422 15034 25442
rect 14510 25361 14565 25405
rect 14565 25361 14574 25405
rect 14510 25341 14574 25361
rect 14602 25361 14603 25405
rect 14603 25361 14659 25405
rect 14659 25361 14666 25405
rect 14602 25341 14666 25361
rect 14694 25361 14697 25405
rect 14697 25361 14753 25405
rect 14753 25361 14758 25405
rect 14694 25341 14758 25361
rect 14786 25361 14791 25405
rect 14791 25361 14847 25405
rect 14847 25361 14850 25405
rect 14786 25341 14850 25361
rect 14878 25361 14885 25405
rect 14885 25361 14941 25405
rect 14941 25361 14942 25405
rect 14878 25341 14942 25361
rect 14970 25361 14979 25405
rect 14979 25361 15034 25405
rect 14970 25341 15034 25361
rect 14510 25280 14565 25324
rect 14565 25280 14574 25324
rect 14510 25260 14574 25280
rect 14602 25280 14603 25324
rect 14603 25280 14659 25324
rect 14659 25280 14666 25324
rect 14602 25260 14666 25280
rect 14694 25280 14697 25324
rect 14697 25280 14753 25324
rect 14753 25280 14758 25324
rect 14694 25260 14758 25280
rect 14786 25280 14791 25324
rect 14791 25280 14847 25324
rect 14847 25280 14850 25324
rect 14786 25260 14850 25280
rect 14878 25280 14885 25324
rect 14885 25280 14941 25324
rect 14941 25280 14942 25324
rect 14878 25260 14942 25280
rect 14970 25280 14979 25324
rect 14979 25280 15034 25324
rect 14970 25260 15034 25280
rect 14510 25199 14565 25243
rect 14565 25199 14574 25243
rect 14510 25179 14574 25199
rect 14602 25199 14603 25243
rect 14603 25199 14659 25243
rect 14659 25199 14666 25243
rect 14602 25179 14666 25199
rect 14694 25199 14697 25243
rect 14697 25199 14753 25243
rect 14753 25199 14758 25243
rect 14694 25179 14758 25199
rect 14786 25199 14791 25243
rect 14791 25199 14847 25243
rect 14847 25199 14850 25243
rect 14786 25179 14850 25199
rect 14878 25199 14885 25243
rect 14885 25199 14941 25243
rect 14941 25199 14942 25243
rect 14878 25179 14942 25199
rect 14970 25199 14979 25243
rect 14979 25199 15034 25243
rect 14970 25179 15034 25199
rect 14510 25118 14565 25162
rect 14565 25118 14574 25162
rect 14510 25098 14574 25118
rect 14602 25118 14603 25162
rect 14603 25118 14659 25162
rect 14659 25118 14666 25162
rect 14602 25098 14666 25118
rect 14694 25118 14697 25162
rect 14697 25118 14753 25162
rect 14753 25118 14758 25162
rect 14694 25098 14758 25118
rect 14786 25118 14791 25162
rect 14791 25118 14847 25162
rect 14847 25118 14850 25162
rect 14786 25098 14850 25118
rect 14878 25118 14885 25162
rect 14885 25118 14941 25162
rect 14941 25118 14942 25162
rect 14878 25098 14942 25118
rect 14970 25118 14979 25162
rect 14979 25118 15034 25162
rect 14970 25098 15034 25118
rect 14510 25037 14565 25081
rect 14565 25037 14574 25081
rect 14510 25017 14574 25037
rect 14602 25037 14603 25081
rect 14603 25037 14659 25081
rect 14659 25037 14666 25081
rect 14602 25017 14666 25037
rect 14694 25037 14697 25081
rect 14697 25037 14753 25081
rect 14753 25037 14758 25081
rect 14694 25017 14758 25037
rect 14786 25037 14791 25081
rect 14791 25037 14847 25081
rect 14847 25037 14850 25081
rect 14786 25017 14850 25037
rect 14878 25037 14885 25081
rect 14885 25037 14941 25081
rect 14941 25037 14942 25081
rect 14878 25017 14942 25037
rect 14970 25037 14979 25081
rect 14979 25037 15034 25081
rect 14970 25017 15034 25037
rect 14510 24955 14565 25000
rect 14565 24955 14574 25000
rect 14510 24936 14574 24955
rect 14602 24955 14603 25000
rect 14603 24955 14659 25000
rect 14659 24955 14666 25000
rect 14602 24936 14666 24955
rect 14694 24955 14697 25000
rect 14697 24955 14753 25000
rect 14753 24955 14758 25000
rect 14694 24936 14758 24955
rect 14786 24955 14791 25000
rect 14791 24955 14847 25000
rect 14847 24955 14850 25000
rect 14786 24936 14850 24955
rect 14878 24955 14885 25000
rect 14885 24955 14941 25000
rect 14941 24955 14942 25000
rect 14878 24936 14942 24955
rect 14970 24955 14979 25000
rect 14979 24955 15034 25000
rect 14970 24936 15034 24955
rect 14510 24873 14565 24919
rect 14565 24873 14574 24919
rect 14510 24855 14574 24873
rect 14602 24873 14603 24919
rect 14603 24873 14659 24919
rect 14659 24873 14666 24919
rect 14602 24855 14666 24873
rect 14694 24873 14697 24919
rect 14697 24873 14753 24919
rect 14753 24873 14758 24919
rect 14694 24855 14758 24873
rect 14786 24873 14791 24919
rect 14791 24873 14847 24919
rect 14847 24873 14850 24919
rect 14786 24855 14850 24873
rect 14878 24873 14885 24919
rect 14885 24873 14941 24919
rect 14941 24873 14942 24919
rect 14878 24855 14942 24873
rect 14970 24873 14979 24919
rect 14979 24873 15034 24919
rect 14970 24855 15034 24873
rect 14510 24791 14565 24838
rect 14565 24791 14574 24838
rect 14510 24774 14574 24791
rect 14602 24791 14603 24838
rect 14603 24791 14659 24838
rect 14659 24791 14666 24838
rect 14602 24774 14666 24791
rect 14694 24791 14697 24838
rect 14697 24791 14753 24838
rect 14753 24791 14758 24838
rect 14694 24774 14758 24791
rect 14786 24791 14791 24838
rect 14791 24791 14847 24838
rect 14847 24791 14850 24838
rect 14786 24774 14850 24791
rect 14878 24791 14885 24838
rect 14885 24791 14941 24838
rect 14941 24791 14942 24838
rect 14878 24774 14942 24791
rect 14970 24791 14979 24838
rect 14979 24791 15034 24838
rect 14970 24774 15034 24791
rect 14510 24709 14565 24757
rect 14565 24709 14574 24757
rect 14510 24693 14574 24709
rect 14602 24709 14603 24757
rect 14603 24709 14659 24757
rect 14659 24709 14666 24757
rect 14602 24693 14666 24709
rect 14694 24709 14697 24757
rect 14697 24709 14753 24757
rect 14753 24709 14758 24757
rect 14694 24693 14758 24709
rect 14786 24709 14791 24757
rect 14791 24709 14847 24757
rect 14847 24709 14850 24757
rect 14786 24693 14850 24709
rect 14878 24709 14885 24757
rect 14885 24709 14941 24757
rect 14941 24709 14942 24757
rect 14878 24693 14942 24709
rect 14970 24709 14979 24757
rect 14979 24709 15034 24757
rect 14970 24693 15034 24709
rect 14510 24627 14565 24676
rect 14565 24627 14574 24676
rect 14510 24612 14574 24627
rect 14602 24627 14603 24676
rect 14603 24627 14659 24676
rect 14659 24627 14666 24676
rect 14602 24612 14666 24627
rect 14694 24627 14697 24676
rect 14697 24627 14753 24676
rect 14753 24627 14758 24676
rect 14694 24612 14758 24627
rect 14786 24627 14791 24676
rect 14791 24627 14847 24676
rect 14847 24627 14850 24676
rect 14786 24612 14850 24627
rect 14878 24627 14885 24676
rect 14885 24627 14941 24676
rect 14941 24627 14942 24676
rect 14878 24612 14942 24627
rect 14970 24627 14979 24676
rect 14979 24627 15034 24676
rect 14970 24612 15034 24627
rect 14510 24545 14565 24595
rect 14565 24545 14574 24595
rect 14510 24531 14574 24545
rect 14602 24545 14603 24595
rect 14603 24545 14659 24595
rect 14659 24545 14666 24595
rect 14602 24531 14666 24545
rect 14694 24545 14697 24595
rect 14697 24545 14753 24595
rect 14753 24545 14758 24595
rect 14694 24531 14758 24545
rect 14786 24545 14791 24595
rect 14791 24545 14847 24595
rect 14847 24545 14850 24595
rect 14786 24531 14850 24545
rect 14878 24545 14885 24595
rect 14885 24545 14941 24595
rect 14941 24545 14942 24595
rect 14878 24531 14942 24545
rect 14970 24545 14979 24595
rect 14979 24545 15034 24595
rect 14970 24531 15034 24545
rect 14510 24463 14565 24514
rect 14565 24463 14574 24514
rect 14510 24450 14574 24463
rect 14602 24463 14603 24514
rect 14603 24463 14659 24514
rect 14659 24463 14666 24514
rect 14602 24450 14666 24463
rect 14694 24463 14697 24514
rect 14697 24463 14753 24514
rect 14753 24463 14758 24514
rect 14694 24450 14758 24463
rect 14786 24463 14791 24514
rect 14791 24463 14847 24514
rect 14847 24463 14850 24514
rect 14786 24450 14850 24463
rect 14878 24463 14885 24514
rect 14885 24463 14941 24514
rect 14941 24463 14942 24514
rect 14878 24450 14942 24463
rect 14970 24463 14979 24514
rect 14979 24463 15034 24514
rect 14970 24450 15034 24463
rect 14510 24381 14565 24433
rect 14565 24381 14574 24433
rect 14510 24369 14574 24381
rect 14602 24381 14603 24433
rect 14603 24381 14659 24433
rect 14659 24381 14666 24433
rect 14602 24369 14666 24381
rect 14694 24381 14697 24433
rect 14697 24381 14753 24433
rect 14753 24381 14758 24433
rect 14694 24369 14758 24381
rect 14786 24381 14791 24433
rect 14791 24381 14847 24433
rect 14847 24381 14850 24433
rect 14786 24369 14850 24381
rect 14878 24381 14885 24433
rect 14885 24381 14941 24433
rect 14941 24381 14942 24433
rect 14878 24369 14942 24381
rect 14970 24381 14979 24433
rect 14979 24381 15034 24433
rect 14970 24369 15034 24381
rect 14510 24299 14565 24352
rect 14565 24299 14574 24352
rect 14510 24288 14574 24299
rect 14602 24299 14603 24352
rect 14603 24299 14659 24352
rect 14659 24299 14666 24352
rect 14602 24288 14666 24299
rect 14694 24299 14697 24352
rect 14697 24299 14753 24352
rect 14753 24299 14758 24352
rect 14694 24288 14758 24299
rect 14786 24299 14791 24352
rect 14791 24299 14847 24352
rect 14847 24299 14850 24352
rect 14786 24288 14850 24299
rect 14878 24299 14885 24352
rect 14885 24299 14941 24352
rect 14941 24299 14942 24352
rect 14878 24288 14942 24299
rect 14970 24299 14979 24352
rect 14979 24299 15034 24352
rect 14970 24288 15034 24299
rect 14510 24217 14565 24271
rect 14565 24217 14574 24271
rect 14510 24207 14574 24217
rect 14602 24217 14603 24271
rect 14603 24217 14659 24271
rect 14659 24217 14666 24271
rect 14602 24207 14666 24217
rect 14694 24217 14697 24271
rect 14697 24217 14753 24271
rect 14753 24217 14758 24271
rect 14694 24207 14758 24217
rect 14786 24217 14791 24271
rect 14791 24217 14847 24271
rect 14847 24217 14850 24271
rect 14786 24207 14850 24217
rect 14878 24217 14885 24271
rect 14885 24217 14941 24271
rect 14941 24217 14942 24271
rect 14878 24207 14942 24217
rect 14970 24217 14979 24271
rect 14979 24217 15034 24271
rect 14970 24207 15034 24217
rect 14510 24135 14565 24190
rect 14565 24135 14574 24190
rect 14510 24126 14574 24135
rect 14602 24135 14603 24190
rect 14603 24135 14659 24190
rect 14659 24135 14666 24190
rect 14602 24126 14666 24135
rect 14694 24135 14697 24190
rect 14697 24135 14753 24190
rect 14753 24135 14758 24190
rect 14694 24126 14758 24135
rect 14786 24135 14791 24190
rect 14791 24135 14847 24190
rect 14847 24135 14850 24190
rect 14786 24126 14850 24135
rect 14878 24135 14885 24190
rect 14885 24135 14941 24190
rect 14941 24135 14942 24190
rect 14878 24126 14942 24135
rect 14970 24135 14979 24190
rect 14979 24135 15034 24190
rect 14970 24126 15034 24135
rect 14510 24053 14565 24109
rect 14565 24053 14574 24109
rect 14510 24045 14574 24053
rect 14602 24053 14603 24109
rect 14603 24053 14659 24109
rect 14659 24053 14666 24109
rect 14602 24045 14666 24053
rect 14694 24053 14697 24109
rect 14697 24053 14753 24109
rect 14753 24053 14758 24109
rect 14694 24045 14758 24053
rect 14786 24053 14791 24109
rect 14791 24053 14847 24109
rect 14847 24053 14850 24109
rect 14786 24045 14850 24053
rect 14878 24053 14885 24109
rect 14885 24053 14941 24109
rect 14941 24053 14942 24109
rect 14878 24045 14942 24053
rect 14970 24053 14979 24109
rect 14979 24053 15034 24109
rect 14970 24045 15034 24053
rect 14510 24027 14574 24028
rect 14510 23971 14565 24027
rect 14565 23971 14574 24027
rect 14510 23964 14574 23971
rect 14602 24027 14666 24028
rect 14602 23971 14603 24027
rect 14603 23971 14659 24027
rect 14659 23971 14666 24027
rect 14602 23964 14666 23971
rect 14694 24027 14758 24028
rect 14694 23971 14697 24027
rect 14697 23971 14753 24027
rect 14753 23971 14758 24027
rect 14694 23964 14758 23971
rect 14786 24027 14850 24028
rect 14786 23971 14791 24027
rect 14791 23971 14847 24027
rect 14847 23971 14850 24027
rect 14786 23964 14850 23971
rect 14878 24027 14942 24028
rect 14878 23971 14885 24027
rect 14885 23971 14941 24027
rect 14941 23971 14942 24027
rect 14878 23964 14942 23971
rect 14970 24027 15034 24028
rect 14970 23971 14979 24027
rect 14979 23971 15034 24027
rect 14970 23964 15034 23971
rect 14510 23945 14574 23947
rect 14510 23889 14565 23945
rect 14565 23889 14574 23945
rect 14510 23883 14574 23889
rect 14602 23945 14666 23947
rect 14602 23889 14603 23945
rect 14603 23889 14659 23945
rect 14659 23889 14666 23945
rect 14602 23883 14666 23889
rect 14694 23945 14758 23947
rect 14694 23889 14697 23945
rect 14697 23889 14753 23945
rect 14753 23889 14758 23945
rect 14694 23883 14758 23889
rect 14786 23945 14850 23947
rect 14786 23889 14791 23945
rect 14791 23889 14847 23945
rect 14847 23889 14850 23945
rect 14786 23883 14850 23889
rect 14878 23945 14942 23947
rect 14878 23889 14885 23945
rect 14885 23889 14941 23945
rect 14941 23889 14942 23945
rect 14878 23883 14942 23889
rect 14970 23945 15034 23947
rect 14970 23889 14979 23945
rect 14979 23889 15034 23945
rect 14970 23883 15034 23889
rect 14510 23863 14574 23866
rect 14510 23807 14565 23863
rect 14565 23807 14574 23863
rect 14510 23802 14574 23807
rect 14602 23863 14666 23866
rect 14602 23807 14603 23863
rect 14603 23807 14659 23863
rect 14659 23807 14666 23863
rect 14602 23802 14666 23807
rect 14694 23863 14758 23866
rect 14694 23807 14697 23863
rect 14697 23807 14753 23863
rect 14753 23807 14758 23863
rect 14694 23802 14758 23807
rect 14786 23863 14850 23866
rect 14786 23807 14791 23863
rect 14791 23807 14847 23863
rect 14847 23807 14850 23863
rect 14786 23802 14850 23807
rect 14878 23863 14942 23866
rect 14878 23807 14885 23863
rect 14885 23807 14941 23863
rect 14941 23807 14942 23863
rect 14878 23802 14942 23807
rect 14970 23863 15034 23866
rect 14970 23807 14979 23863
rect 14979 23807 15034 23863
rect 14970 23802 15034 23807
rect 14510 23781 14574 23785
rect 14510 23725 14565 23781
rect 14565 23725 14574 23781
rect 14510 23721 14574 23725
rect 14602 23781 14666 23785
rect 14602 23725 14603 23781
rect 14603 23725 14659 23781
rect 14659 23725 14666 23781
rect 14602 23721 14666 23725
rect 14694 23781 14758 23785
rect 14694 23725 14697 23781
rect 14697 23725 14753 23781
rect 14753 23725 14758 23781
rect 14694 23721 14758 23725
rect 14786 23781 14850 23785
rect 14786 23725 14791 23781
rect 14791 23725 14847 23781
rect 14847 23725 14850 23781
rect 14786 23721 14850 23725
rect 14878 23781 14942 23785
rect 14878 23725 14885 23781
rect 14885 23725 14941 23781
rect 14941 23725 14942 23781
rect 14878 23721 14942 23725
rect 14970 23781 15034 23785
rect 14970 23725 14979 23781
rect 14979 23725 15034 23781
rect 14970 23721 15034 23725
rect 14510 23699 14574 23704
rect 14510 23643 14565 23699
rect 14565 23643 14574 23699
rect 14510 23640 14574 23643
rect 14602 23699 14666 23704
rect 14602 23643 14603 23699
rect 14603 23643 14659 23699
rect 14659 23643 14666 23699
rect 14602 23640 14666 23643
rect 14694 23699 14758 23704
rect 14694 23643 14697 23699
rect 14697 23643 14753 23699
rect 14753 23643 14758 23699
rect 14694 23640 14758 23643
rect 14786 23699 14850 23704
rect 14786 23643 14791 23699
rect 14791 23643 14847 23699
rect 14847 23643 14850 23699
rect 14786 23640 14850 23643
rect 14878 23699 14942 23704
rect 14878 23643 14885 23699
rect 14885 23643 14941 23699
rect 14941 23643 14942 23699
rect 14878 23640 14942 23643
rect 14970 23699 15034 23704
rect 14970 23643 14979 23699
rect 14979 23643 15034 23699
rect 14970 23640 15034 23643
rect 14510 23617 14574 23623
rect 14510 23561 14565 23617
rect 14565 23561 14574 23617
rect 14510 23559 14574 23561
rect 14602 23617 14666 23623
rect 14602 23561 14603 23617
rect 14603 23561 14659 23617
rect 14659 23561 14666 23617
rect 14602 23559 14666 23561
rect 14694 23617 14758 23623
rect 14694 23561 14697 23617
rect 14697 23561 14753 23617
rect 14753 23561 14758 23617
rect 14694 23559 14758 23561
rect 14786 23617 14850 23623
rect 14786 23561 14791 23617
rect 14791 23561 14847 23617
rect 14847 23561 14850 23617
rect 14786 23559 14850 23561
rect 14878 23617 14942 23623
rect 14878 23561 14885 23617
rect 14885 23561 14941 23617
rect 14941 23561 14942 23617
rect 14878 23559 14942 23561
rect 14970 23617 15034 23623
rect 14970 23561 14979 23617
rect 14979 23561 15034 23617
rect 14970 23559 15034 23561
rect 14510 23535 14574 23542
rect 14510 23479 14565 23535
rect 14565 23479 14574 23535
rect 14510 23478 14574 23479
rect 14602 23535 14666 23542
rect 14602 23479 14603 23535
rect 14603 23479 14659 23535
rect 14659 23479 14666 23535
rect 14602 23478 14666 23479
rect 14694 23535 14758 23542
rect 14694 23479 14697 23535
rect 14697 23479 14753 23535
rect 14753 23479 14758 23535
rect 14694 23478 14758 23479
rect 14786 23535 14850 23542
rect 14786 23479 14791 23535
rect 14791 23479 14847 23535
rect 14847 23479 14850 23535
rect 14786 23478 14850 23479
rect 14878 23535 14942 23542
rect 14878 23479 14885 23535
rect 14885 23479 14941 23535
rect 14941 23479 14942 23535
rect 14878 23478 14942 23479
rect 14970 23535 15034 23542
rect 14970 23479 14979 23535
rect 14979 23479 15034 23535
rect 14970 23478 15034 23479
rect 14510 23453 14574 23461
rect 14510 23397 14565 23453
rect 14565 23397 14574 23453
rect 14602 23453 14666 23461
rect 14602 23397 14603 23453
rect 14603 23397 14659 23453
rect 14659 23397 14666 23453
rect 14694 23453 14758 23461
rect 14694 23397 14697 23453
rect 14697 23397 14753 23453
rect 14753 23397 14758 23453
rect 14786 23453 14850 23461
rect 14786 23397 14791 23453
rect 14791 23397 14847 23453
rect 14847 23397 14850 23453
rect 14878 23453 14942 23461
rect 14878 23397 14885 23453
rect 14885 23397 14941 23453
rect 14941 23397 14942 23453
rect 14970 23453 15034 23461
rect 14970 23397 14979 23453
rect 14979 23397 15034 23453
rect 14510 23371 14574 23380
rect 14510 23316 14565 23371
rect 14565 23316 14574 23371
rect 14602 23371 14666 23380
rect 14602 23316 14603 23371
rect 14603 23316 14659 23371
rect 14659 23316 14666 23371
rect 14694 23371 14758 23380
rect 14694 23316 14697 23371
rect 14697 23316 14753 23371
rect 14753 23316 14758 23371
rect 14786 23371 14850 23380
rect 14786 23316 14791 23371
rect 14791 23316 14847 23371
rect 14847 23316 14850 23371
rect 14878 23371 14942 23380
rect 14878 23316 14885 23371
rect 14885 23316 14941 23371
rect 14941 23316 14942 23371
rect 14970 23371 15034 23380
rect 14970 23316 14979 23371
rect 14979 23316 15034 23371
rect 14510 23289 14574 23299
rect 14510 23235 14565 23289
rect 14565 23235 14574 23289
rect 14602 23289 14666 23299
rect 14602 23235 14603 23289
rect 14603 23235 14659 23289
rect 14659 23235 14666 23289
rect 14694 23289 14758 23299
rect 14694 23235 14697 23289
rect 14697 23235 14753 23289
rect 14753 23235 14758 23289
rect 14786 23289 14850 23299
rect 14786 23235 14791 23289
rect 14791 23235 14847 23289
rect 14847 23235 14850 23289
rect 14878 23289 14942 23299
rect 14878 23235 14885 23289
rect 14885 23235 14941 23289
rect 14941 23235 14942 23289
rect 14970 23289 15034 23299
rect 14970 23235 14979 23289
rect 14979 23235 15034 23289
rect 14510 23207 14574 23218
rect 14510 23154 14565 23207
rect 14565 23154 14574 23207
rect 14602 23207 14666 23218
rect 14602 23154 14603 23207
rect 14603 23154 14659 23207
rect 14659 23154 14666 23207
rect 14694 23207 14758 23218
rect 14694 23154 14697 23207
rect 14697 23154 14753 23207
rect 14753 23154 14758 23207
rect 14786 23207 14850 23218
rect 14786 23154 14791 23207
rect 14791 23154 14847 23207
rect 14847 23154 14850 23207
rect 14878 23207 14942 23218
rect 14878 23154 14885 23207
rect 14885 23154 14941 23207
rect 14941 23154 14942 23207
rect 14970 23207 15034 23218
rect 14970 23154 14979 23207
rect 14979 23154 15034 23207
rect 292 18912 356 18976
rect 392 18912 456 18976
rect 492 18912 556 18976
rect 592 18912 656 18976
rect 292 18832 356 18896
rect 392 18832 456 18896
rect 492 18832 556 18896
rect 592 18832 656 18896
rect 292 18752 356 18816
rect 392 18752 456 18816
rect 492 18752 556 18816
rect 592 18752 656 18816
rect 292 18672 356 18736
rect 392 18672 456 18736
rect 492 18672 556 18736
rect 592 18672 656 18736
rect 292 18592 356 18656
rect 392 18592 456 18656
rect 492 18592 556 18656
rect 592 18592 656 18656
rect 292 18512 356 18576
rect 392 18512 456 18576
rect 492 18512 556 18576
rect 592 18512 656 18576
rect 292 18432 356 18496
rect 392 18432 456 18496
rect 492 18432 556 18496
rect 592 18432 656 18496
rect 292 18352 356 18416
rect 392 18352 456 18416
rect 492 18352 556 18416
rect 592 18352 656 18416
rect 292 18272 356 18336
rect 392 18272 456 18336
rect 492 18272 556 18336
rect 592 18272 656 18336
rect 292 18192 356 18256
rect 392 18192 456 18256
rect 492 18192 556 18256
rect 592 18192 656 18256
rect 292 18112 356 18176
rect 392 18112 456 18176
rect 492 18112 556 18176
rect 592 18112 656 18176
rect 292 18032 356 18096
rect 392 18032 456 18096
rect 492 18032 556 18096
rect 592 18032 656 18096
rect 292 17951 356 18015
rect 392 17951 456 18015
rect 492 17951 556 18015
rect 592 17951 656 18015
rect 292 17870 356 17934
rect 392 17870 456 17934
rect 492 17870 556 17934
rect 592 17870 656 17934
rect 292 17789 356 17853
rect 392 17789 456 17853
rect 492 17789 556 17853
rect 592 17789 656 17853
rect 292 17708 356 17772
rect 392 17708 456 17772
rect 492 17708 556 17772
rect 592 17708 656 17772
rect 292 17627 356 17691
rect 392 17627 456 17691
rect 492 17627 556 17691
rect 592 17627 656 17691
rect 292 17546 356 17610
rect 392 17546 456 17610
rect 492 17546 556 17610
rect 592 17546 656 17610
rect 292 17465 356 17529
rect 392 17465 456 17529
rect 492 17465 556 17529
rect 592 17465 656 17529
rect 292 17384 356 17448
rect 392 17384 456 17448
rect 492 17384 556 17448
rect 592 17384 656 17448
rect 292 17303 356 17367
rect 392 17303 456 17367
rect 492 17303 556 17367
rect 592 17303 656 17367
rect 292 17222 356 17286
rect 392 17222 456 17286
rect 492 17222 556 17286
rect 592 17222 656 17286
rect 292 17141 356 17205
rect 392 17141 456 17205
rect 492 17141 556 17205
rect 592 17141 656 17205
rect 292 17060 356 17124
rect 392 17060 456 17124
rect 492 17060 556 17124
rect 592 17060 656 17124
rect 292 16979 356 17043
rect 392 16979 456 17043
rect 492 16979 556 17043
rect 592 16979 656 17043
rect 292 16898 356 16962
rect 392 16898 456 16962
rect 492 16898 556 16962
rect 592 16898 656 16962
rect 292 16817 356 16881
rect 392 16817 456 16881
rect 492 16817 556 16881
rect 592 16817 656 16881
rect 292 16736 356 16800
rect 392 16736 456 16800
rect 492 16736 556 16800
rect 592 16736 656 16800
rect 292 16655 356 16719
rect 392 16655 456 16719
rect 492 16655 556 16719
rect 592 16655 656 16719
rect 292 16574 356 16638
rect 392 16574 456 16638
rect 492 16574 556 16638
rect 592 16574 656 16638
rect 292 16493 356 16557
rect 392 16493 456 16557
rect 492 16493 556 16557
rect 592 16493 656 16557
rect 292 16412 356 16476
rect 392 16412 456 16476
rect 492 16412 556 16476
rect 592 16412 656 16476
rect 292 16331 356 16395
rect 392 16331 456 16395
rect 492 16331 556 16395
rect 592 16331 656 16395
rect 292 16250 356 16314
rect 392 16250 456 16314
rect 492 16250 556 16314
rect 592 16250 656 16314
rect 292 16169 356 16233
rect 392 16169 456 16233
rect 492 16169 556 16233
rect 592 16169 656 16233
rect 292 16088 356 16152
rect 392 16088 456 16152
rect 492 16088 556 16152
rect 592 16088 656 16152
rect 292 16007 356 16071
rect 392 16007 456 16071
rect 492 16007 556 16071
rect 592 16007 656 16071
rect 292 15926 356 15990
rect 392 15926 456 15990
rect 492 15926 556 15990
rect 592 15926 656 15990
rect 292 15845 356 15909
rect 392 15845 456 15909
rect 492 15845 556 15909
rect 592 15845 656 15909
rect 292 15764 356 15828
rect 392 15764 456 15828
rect 492 15764 556 15828
rect 592 15764 656 15828
rect 292 15683 356 15747
rect 392 15683 456 15747
rect 492 15683 556 15747
rect 592 15683 656 15747
rect 292 15602 356 15666
rect 392 15602 456 15666
rect 492 15602 556 15666
rect 592 15602 656 15666
rect 292 15521 356 15585
rect 392 15521 456 15585
rect 492 15521 556 15585
rect 592 15521 656 15585
rect 292 15440 356 15504
rect 392 15440 456 15504
rect 492 15440 556 15504
rect 592 15440 656 15504
rect 292 15359 356 15423
rect 392 15359 456 15423
rect 492 15359 556 15423
rect 592 15359 656 15423
rect 292 15278 356 15342
rect 392 15278 456 15342
rect 492 15278 556 15342
rect 592 15278 656 15342
rect 292 15197 356 15261
rect 392 15197 456 15261
rect 492 15197 556 15261
rect 592 15197 656 15261
rect 292 15116 356 15180
rect 392 15116 456 15180
rect 492 15116 556 15180
rect 592 15116 656 15180
rect 292 15035 356 15099
rect 392 15035 456 15099
rect 492 15035 556 15099
rect 592 15035 656 15099
rect 292 14954 356 15018
rect 392 14954 456 15018
rect 492 14954 556 15018
rect 592 14954 656 15018
rect 292 14873 356 14937
rect 392 14873 456 14937
rect 492 14873 556 14937
rect 592 14873 656 14937
rect 292 14792 356 14856
rect 392 14792 456 14856
rect 492 14792 556 14856
rect 592 14792 656 14856
rect 292 14711 356 14775
rect 392 14711 456 14775
rect 492 14711 556 14775
rect 592 14711 656 14775
rect 292 14630 356 14694
rect 392 14630 456 14694
rect 492 14630 556 14694
rect 592 14630 656 14694
rect 292 14549 356 14613
rect 392 14549 456 14613
rect 492 14549 556 14613
rect 592 14549 656 14613
rect 292 14468 356 14532
rect 392 14468 456 14532
rect 492 14468 556 14532
rect 592 14468 656 14532
rect 292 14387 356 14451
rect 392 14387 456 14451
rect 492 14387 556 14451
rect 592 14387 656 14451
rect 292 14306 356 14370
rect 392 14306 456 14370
rect 492 14306 556 14370
rect 592 14306 656 14370
rect 292 14225 356 14289
rect 392 14225 456 14289
rect 492 14225 556 14289
rect 592 14225 656 14289
rect 292 14144 356 14208
rect 392 14144 456 14208
rect 492 14144 556 14208
rect 592 14144 656 14208
rect 292 14063 356 14127
rect 392 14063 456 14127
rect 492 14063 556 14127
rect 592 14063 656 14127
rect 522 11282 586 11346
rect 606 11282 670 11346
rect 690 11282 754 11346
rect 522 10499 586 10563
rect 606 10499 670 10563
rect 690 10499 754 10563
rect 522 10415 586 10479
rect 606 10415 670 10479
rect 690 10415 754 10479
rect 522 10331 586 10395
rect 606 10331 670 10395
rect 690 10331 754 10395
rect 522 9548 586 9612
rect 606 9548 670 9612
rect 690 9548 754 9612
rect 1372 13532 1436 13596
rect 1502 13532 1566 13596
rect 1372 13445 1436 13509
rect 1502 13445 1566 13509
rect 1372 13358 1436 13422
rect 1502 13358 1566 13422
rect 1372 13271 1436 13335
rect 1502 13271 1566 13335
rect 1372 13184 1436 13248
rect 1502 13184 1566 13248
rect 1372 13097 1436 13161
rect 1502 13097 1566 13161
rect 1372 13010 1436 13074
rect 1502 13010 1566 13074
rect 1372 12922 1436 12986
rect 1502 12922 1566 12986
rect 1372 12834 1436 12898
rect 1502 12834 1566 12898
rect 13738 20312 13802 20376
rect 13888 20312 13952 20376
rect 13738 20218 13802 20282
rect 13888 20218 13952 20282
rect 13738 20124 13802 20188
rect 13888 20124 13952 20188
rect 13738 20030 13802 20094
rect 13888 20030 13952 20094
rect 13738 19935 13802 19999
rect 13888 19935 13952 19999
rect 13738 19840 13802 19904
rect 13888 19840 13952 19904
rect 1138 9408 1202 9472
rect 1218 9408 1282 9472
rect 911 7174 975 7238
rect 991 7174 1055 7238
rect 1486 4822 1550 4886
rect 1570 4822 1634 4886
rect 1654 4852 1709 4886
rect 1709 4852 1718 4886
rect 1738 4852 1765 4886
rect 1765 4852 1797 4886
rect 1797 4852 1802 4886
rect 1822 4852 1853 4886
rect 1853 4852 1885 4886
rect 1885 4852 1886 4886
rect 1906 4852 1941 4886
rect 1941 4852 1970 4886
rect 1990 4852 2029 4886
rect 2029 4852 2054 4886
rect 2074 4852 2117 4886
rect 2117 4852 2138 4886
rect 1654 4828 1718 4852
rect 1738 4828 1802 4852
rect 1822 4828 1886 4852
rect 1906 4828 1970 4852
rect 1990 4828 2054 4852
rect 2074 4828 2138 4852
rect 1654 4822 1709 4828
rect 1709 4822 1718 4828
rect 1738 4822 1765 4828
rect 1765 4822 1797 4828
rect 1797 4822 1802 4828
rect 1822 4822 1853 4828
rect 1853 4822 1885 4828
rect 1885 4822 1886 4828
rect 1906 4822 1941 4828
rect 1941 4822 1970 4828
rect 1990 4822 2029 4828
rect 2029 4822 2054 4828
rect 2074 4822 2117 4828
rect 2117 4822 2138 4828
rect 1486 4736 1550 4800
rect 1570 4736 1634 4800
rect 1654 4772 1709 4800
rect 1709 4772 1718 4800
rect 1738 4772 1765 4800
rect 1765 4772 1797 4800
rect 1797 4772 1802 4800
rect 1822 4772 1853 4800
rect 1853 4772 1885 4800
rect 1885 4772 1886 4800
rect 1906 4772 1941 4800
rect 1941 4772 1970 4800
rect 1990 4772 2029 4800
rect 2029 4772 2054 4800
rect 2074 4772 2117 4800
rect 2117 4772 2138 4800
rect 1654 4747 1718 4772
rect 1738 4747 1802 4772
rect 1822 4747 1886 4772
rect 1906 4747 1970 4772
rect 1990 4747 2054 4772
rect 2074 4747 2138 4772
rect 1654 4736 1709 4747
rect 1709 4736 1718 4747
rect 1738 4736 1765 4747
rect 1765 4736 1797 4747
rect 1797 4736 1802 4747
rect 1822 4736 1853 4747
rect 1853 4736 1885 4747
rect 1885 4736 1886 4747
rect 1906 4736 1941 4747
rect 1941 4736 1970 4747
rect 1990 4736 2029 4747
rect 2029 4736 2054 4747
rect 2074 4736 2117 4747
rect 2117 4736 2138 4747
rect 1486 4650 1550 4714
rect 1570 4650 1634 4714
rect 1654 4691 1709 4714
rect 1709 4691 1718 4714
rect 1738 4691 1765 4714
rect 1765 4691 1797 4714
rect 1797 4691 1802 4714
rect 1822 4691 1853 4714
rect 1853 4691 1885 4714
rect 1885 4691 1886 4714
rect 1906 4691 1941 4714
rect 1941 4691 1970 4714
rect 1990 4691 2029 4714
rect 2029 4691 2054 4714
rect 2074 4691 2117 4714
rect 2117 4691 2138 4714
rect 1654 4666 1718 4691
rect 1738 4666 1802 4691
rect 1822 4666 1886 4691
rect 1906 4666 1970 4691
rect 1990 4666 2054 4691
rect 2074 4666 2138 4691
rect 1654 4650 1709 4666
rect 1709 4650 1718 4666
rect 1738 4650 1765 4666
rect 1765 4650 1797 4666
rect 1797 4650 1802 4666
rect 1822 4650 1853 4666
rect 1853 4650 1885 4666
rect 1885 4650 1886 4666
rect 1906 4650 1941 4666
rect 1941 4650 1970 4666
rect 1990 4650 2029 4666
rect 2029 4650 2054 4666
rect 2074 4650 2117 4666
rect 2117 4650 2138 4666
rect 1486 4564 1550 4628
rect 1570 4564 1634 4628
rect 1654 4610 1709 4628
rect 1709 4610 1718 4628
rect 1738 4610 1765 4628
rect 1765 4610 1797 4628
rect 1797 4610 1802 4628
rect 1822 4610 1853 4628
rect 1853 4610 1885 4628
rect 1885 4610 1886 4628
rect 1906 4610 1941 4628
rect 1941 4610 1970 4628
rect 1990 4610 2029 4628
rect 2029 4610 2054 4628
rect 2074 4610 2117 4628
rect 2117 4610 2138 4628
rect 1654 4585 1718 4610
rect 1738 4585 1802 4610
rect 1822 4585 1886 4610
rect 1906 4585 1970 4610
rect 1990 4585 2054 4610
rect 2074 4585 2138 4610
rect 1654 4564 1709 4585
rect 1709 4564 1718 4585
rect 1738 4564 1765 4585
rect 1765 4564 1797 4585
rect 1797 4564 1802 4585
rect 1822 4564 1853 4585
rect 1853 4564 1885 4585
rect 1885 4564 1886 4585
rect 1906 4564 1941 4585
rect 1941 4564 1970 4585
rect 1990 4564 2029 4585
rect 2029 4564 2054 4585
rect 2074 4564 2117 4585
rect 2117 4564 2138 4585
rect 1486 4478 1550 4542
rect 1570 4478 1634 4542
rect 1654 4529 1709 4542
rect 1709 4529 1718 4542
rect 1738 4529 1765 4542
rect 1765 4529 1797 4542
rect 1797 4529 1802 4542
rect 1822 4529 1853 4542
rect 1853 4529 1885 4542
rect 1885 4529 1886 4542
rect 1906 4529 1941 4542
rect 1941 4529 1970 4542
rect 1990 4529 2029 4542
rect 2029 4529 2054 4542
rect 2074 4529 2117 4542
rect 2117 4529 2138 4542
rect 1654 4504 1718 4529
rect 1738 4504 1802 4529
rect 1822 4504 1886 4529
rect 1906 4504 1970 4529
rect 1990 4504 2054 4529
rect 2074 4504 2138 4529
rect 1654 4478 1709 4504
rect 1709 4478 1718 4504
rect 1738 4478 1765 4504
rect 1765 4478 1797 4504
rect 1797 4478 1802 4504
rect 1822 4478 1853 4504
rect 1853 4478 1885 4504
rect 1885 4478 1886 4504
rect 1906 4478 1941 4504
rect 1941 4478 1970 4504
rect 1990 4478 2029 4504
rect 2029 4478 2054 4504
rect 2074 4478 2117 4504
rect 2117 4478 2138 4504
rect 1486 4392 1550 4456
rect 1570 4392 1634 4456
rect 1654 4448 1709 4456
rect 1709 4448 1718 4456
rect 1738 4448 1765 4456
rect 1765 4448 1797 4456
rect 1797 4448 1802 4456
rect 1822 4448 1853 4456
rect 1853 4448 1885 4456
rect 1885 4448 1886 4456
rect 1906 4448 1941 4456
rect 1941 4448 1970 4456
rect 1990 4448 2029 4456
rect 2029 4448 2054 4456
rect 2074 4448 2117 4456
rect 2117 4448 2138 4456
rect 1654 4423 1718 4448
rect 1738 4423 1802 4448
rect 1822 4423 1886 4448
rect 1906 4423 1970 4448
rect 1990 4423 2054 4448
rect 2074 4423 2138 4448
rect 1654 4392 1709 4423
rect 1709 4392 1718 4423
rect 1738 4392 1765 4423
rect 1765 4392 1797 4423
rect 1797 4392 1802 4423
rect 1822 4392 1853 4423
rect 1853 4392 1885 4423
rect 1885 4392 1886 4423
rect 1906 4392 1941 4423
rect 1941 4392 1970 4423
rect 1990 4392 2029 4423
rect 2029 4392 2054 4423
rect 2074 4392 2117 4423
rect 2117 4392 2138 4423
rect 1486 4306 1550 4370
rect 1570 4306 1634 4370
rect 1654 4367 1709 4370
rect 1709 4367 1718 4370
rect 1738 4367 1765 4370
rect 1765 4367 1797 4370
rect 1797 4367 1802 4370
rect 1822 4367 1853 4370
rect 1853 4367 1885 4370
rect 1885 4367 1886 4370
rect 1906 4367 1941 4370
rect 1941 4367 1970 4370
rect 1990 4367 2029 4370
rect 2029 4367 2054 4370
rect 2074 4367 2117 4370
rect 2117 4367 2138 4370
rect 1654 4342 1718 4367
rect 1738 4342 1802 4367
rect 1822 4342 1886 4367
rect 1906 4342 1970 4367
rect 1990 4342 2054 4367
rect 2074 4342 2138 4367
rect 1654 4306 1709 4342
rect 1709 4306 1718 4342
rect 1738 4306 1765 4342
rect 1765 4306 1797 4342
rect 1797 4306 1802 4342
rect 1822 4306 1853 4342
rect 1853 4306 1885 4342
rect 1885 4306 1886 4342
rect 1906 4306 1941 4342
rect 1941 4306 1970 4342
rect 1990 4306 2029 4342
rect 2029 4306 2054 4342
rect 2074 4306 2117 4342
rect 2117 4306 2138 4342
rect 1486 4219 1550 4283
rect 1570 4219 1634 4283
rect 1654 4261 1718 4283
rect 1738 4261 1802 4283
rect 1822 4261 1886 4283
rect 1906 4261 1970 4283
rect 1990 4261 2054 4283
rect 2074 4261 2138 4283
rect 1654 4219 1709 4261
rect 1709 4219 1718 4261
rect 1738 4219 1765 4261
rect 1765 4219 1797 4261
rect 1797 4219 1802 4261
rect 1822 4219 1853 4261
rect 1853 4219 1885 4261
rect 1885 4219 1886 4261
rect 1906 4219 1941 4261
rect 1941 4219 1970 4261
rect 1990 4219 2029 4261
rect 2029 4219 2054 4261
rect 2074 4219 2117 4261
rect 2117 4219 2138 4261
rect 1486 4132 1550 4196
rect 1570 4132 1634 4196
rect 1654 4180 1718 4196
rect 1738 4180 1802 4196
rect 1822 4180 1886 4196
rect 1906 4180 1970 4196
rect 1990 4180 2054 4196
rect 2074 4180 2138 4196
rect 1654 4132 1709 4180
rect 1709 4132 1718 4180
rect 1738 4132 1765 4180
rect 1765 4132 1797 4180
rect 1797 4132 1802 4180
rect 1822 4132 1853 4180
rect 1853 4132 1885 4180
rect 1885 4132 1886 4180
rect 1906 4132 1941 4180
rect 1941 4132 1970 4180
rect 1990 4132 2029 4180
rect 2029 4132 2054 4180
rect 2074 4132 2117 4180
rect 2117 4132 2138 4180
rect 1486 4045 1550 4109
rect 1570 4045 1634 4109
rect 1654 4099 1718 4109
rect 1738 4099 1802 4109
rect 1822 4099 1886 4109
rect 1906 4099 1970 4109
rect 1990 4099 2054 4109
rect 2074 4099 2138 4109
rect 1654 4045 1709 4099
rect 1709 4045 1718 4099
rect 1738 4045 1765 4099
rect 1765 4045 1797 4099
rect 1797 4045 1802 4099
rect 1822 4045 1853 4099
rect 1853 4045 1885 4099
rect 1885 4045 1886 4099
rect 1906 4045 1941 4099
rect 1941 4045 1970 4099
rect 1990 4045 2029 4099
rect 2029 4045 2054 4099
rect 2074 4045 2117 4099
rect 2117 4045 2138 4099
rect 1486 3958 1550 4022
rect 1570 3958 1634 4022
rect 1654 4018 1718 4022
rect 1738 4018 1802 4022
rect 1822 4018 1886 4022
rect 1906 4018 1970 4022
rect 1990 4018 2054 4022
rect 2074 4018 2138 4022
rect 1654 3962 1709 4018
rect 1709 3962 1718 4018
rect 1738 3962 1765 4018
rect 1765 3962 1797 4018
rect 1797 3962 1802 4018
rect 1822 3962 1853 4018
rect 1853 3962 1885 4018
rect 1885 3962 1886 4018
rect 1906 3962 1941 4018
rect 1941 3962 1970 4018
rect 1990 3962 2029 4018
rect 2029 3962 2054 4018
rect 2074 3962 2117 4018
rect 2117 3962 2138 4018
rect 1654 3958 1718 3962
rect 1738 3958 1802 3962
rect 1822 3958 1886 3962
rect 1906 3958 1970 3962
rect 1990 3958 2054 3962
rect 2074 3958 2138 3962
rect 291 274 344 298
rect 344 274 355 298
rect 291 250 355 274
rect 291 234 344 250
rect 344 234 355 250
rect 371 234 435 298
rect 2230 1432 2294 1496
rect 2310 1432 2374 1496
rect 2390 1432 2454 1496
rect 2470 1432 2534 1496
rect 2550 1432 2614 1496
rect 2630 1432 2694 1496
rect 2230 1348 2294 1412
rect 2310 1348 2374 1412
rect 2390 1348 2454 1412
rect 2470 1348 2534 1412
rect 2550 1348 2614 1412
rect 2630 1348 2694 1412
rect 2230 1264 2294 1328
rect 2310 1264 2374 1328
rect 2390 1264 2454 1328
rect 2470 1264 2534 1328
rect 2550 1264 2614 1328
rect 2630 1264 2694 1328
rect 2230 1180 2294 1244
rect 2310 1180 2374 1244
rect 2390 1180 2454 1244
rect 2470 1180 2534 1244
rect 2550 1180 2614 1244
rect 2630 1180 2694 1244
rect 2230 1096 2294 1160
rect 2310 1096 2374 1160
rect 2390 1096 2454 1160
rect 2470 1096 2534 1160
rect 2550 1096 2614 1160
rect 2630 1096 2694 1160
rect 2230 1012 2294 1076
rect 2310 1012 2374 1076
rect 2390 1012 2454 1076
rect 2470 1012 2534 1076
rect 2550 1012 2614 1076
rect 2630 1012 2694 1076
rect 2230 928 2294 992
rect 2310 928 2374 992
rect 2390 928 2454 992
rect 2470 928 2534 992
rect 2550 928 2614 992
rect 2630 928 2694 992
rect 2230 844 2294 908
rect 2310 844 2374 908
rect 2390 844 2454 908
rect 2470 844 2534 908
rect 2550 844 2614 908
rect 2630 844 2694 908
rect 2230 759 2294 823
rect 2310 759 2374 823
rect 2390 759 2454 823
rect 2470 759 2534 823
rect 2550 759 2614 823
rect 2630 759 2694 823
rect 2230 674 2294 738
rect 2310 674 2374 738
rect 2390 674 2454 738
rect 2470 674 2534 738
rect 2550 674 2614 738
rect 2630 674 2694 738
rect 2230 589 2294 653
rect 2310 589 2374 653
rect 2390 589 2454 653
rect 2470 589 2534 653
rect 2550 589 2614 653
rect 2630 589 2694 653
rect 2782 9204 2789 9246
rect 2789 9204 2845 9246
rect 2845 9204 2846 9246
rect 2782 9182 2846 9204
rect 2866 9204 2921 9246
rect 2921 9204 2930 9246
rect 2950 9204 2977 9246
rect 2977 9204 3014 9246
rect 2866 9182 2930 9204
rect 2950 9182 3014 9204
rect 3034 9204 3053 9246
rect 3053 9204 3098 9246
rect 3034 9182 3098 9204
rect 3118 9182 3182 9246
rect 3202 9204 3241 9246
rect 3241 9204 3266 9246
rect 3202 9182 3266 9204
rect 3286 9204 3317 9246
rect 3317 9204 3350 9246
rect 3370 9204 3373 9246
rect 3373 9204 3434 9246
rect 3454 9204 3505 9246
rect 3505 9204 3518 9246
rect 3286 9182 3350 9204
rect 3370 9182 3434 9204
rect 3454 9182 3518 9204
rect 3538 9204 3581 9246
rect 3581 9204 3602 9246
rect 3622 9204 3637 9246
rect 3637 9204 3686 9246
rect 3538 9182 3602 9204
rect 3622 9182 3686 9204
rect 3706 9204 3713 9246
rect 3713 9204 3769 9246
rect 3769 9204 3770 9246
rect 3706 9182 3770 9204
rect 2782 9120 2846 9160
rect 2782 9096 2789 9120
rect 2789 9096 2845 9120
rect 2845 9096 2846 9120
rect 2866 9120 2930 9160
rect 2950 9120 3014 9160
rect 2866 9096 2921 9120
rect 2921 9096 2930 9120
rect 2950 9096 2977 9120
rect 2977 9096 3014 9120
rect 3034 9120 3098 9160
rect 3034 9096 3053 9120
rect 3053 9096 3098 9120
rect 3118 9096 3182 9160
rect 3202 9120 3266 9160
rect 3202 9096 3241 9120
rect 3241 9096 3266 9120
rect 3286 9120 3350 9160
rect 3370 9120 3434 9160
rect 3454 9120 3518 9160
rect 3286 9096 3317 9120
rect 3317 9096 3350 9120
rect 3370 9096 3373 9120
rect 3373 9096 3434 9120
rect 3454 9096 3505 9120
rect 3505 9096 3518 9120
rect 3538 9120 3602 9160
rect 3622 9120 3686 9160
rect 3538 9096 3581 9120
rect 3581 9096 3602 9120
rect 3622 9096 3637 9120
rect 3637 9096 3686 9120
rect 3706 9120 3770 9160
rect 3706 9096 3713 9120
rect 3713 9096 3769 9120
rect 3769 9096 3770 9120
rect 2782 9064 2789 9074
rect 2789 9064 2845 9074
rect 2845 9064 2846 9074
rect 2782 9010 2846 9064
rect 2866 9064 2921 9074
rect 2921 9064 2930 9074
rect 2950 9064 2977 9074
rect 2977 9064 3014 9074
rect 2866 9010 2930 9064
rect 2950 9010 3014 9064
rect 3034 9064 3053 9074
rect 3053 9064 3098 9074
rect 3034 9010 3098 9064
rect 3118 9010 3182 9074
rect 3202 9064 3241 9074
rect 3241 9064 3266 9074
rect 3202 9010 3266 9064
rect 3286 9064 3317 9074
rect 3317 9064 3350 9074
rect 3370 9064 3373 9074
rect 3373 9064 3434 9074
rect 3454 9064 3505 9074
rect 3505 9064 3518 9074
rect 3286 9010 3350 9064
rect 3370 9010 3434 9064
rect 3454 9010 3518 9064
rect 3538 9064 3581 9074
rect 3581 9064 3602 9074
rect 3622 9064 3637 9074
rect 3637 9064 3686 9074
rect 3538 9010 3602 9064
rect 3622 9010 3686 9064
rect 3706 9064 3713 9074
rect 3713 9064 3769 9074
rect 3769 9064 3770 9074
rect 3706 9010 3770 9064
rect 2782 8924 2846 8988
rect 2866 8924 2930 8988
rect 2950 8924 3014 8988
rect 3034 8924 3098 8988
rect 3118 8924 3182 8988
rect 3202 8924 3266 8988
rect 3286 8924 3350 8988
rect 3370 8924 3434 8988
rect 3454 8924 3518 8988
rect 3538 8924 3602 8988
rect 3622 8924 3686 8988
rect 3706 8924 3770 8988
rect 2782 8838 2846 8902
rect 2866 8838 2930 8902
rect 2950 8838 3014 8902
rect 3034 8838 3098 8902
rect 3118 8838 3182 8902
rect 3202 8838 3266 8902
rect 3286 8838 3350 8902
rect 3370 8838 3434 8902
rect 3454 8838 3518 8902
rect 3538 8838 3602 8902
rect 3622 8838 3686 8902
rect 3706 8838 3770 8902
rect 2782 8752 2846 8816
rect 2866 8752 2930 8816
rect 2950 8752 3014 8816
rect 3034 8752 3098 8816
rect 3118 8752 3182 8816
rect 3202 8752 3266 8816
rect 3286 8752 3350 8816
rect 3370 8752 3434 8816
rect 3454 8752 3518 8816
rect 3538 8752 3602 8816
rect 3622 8752 3686 8816
rect 3706 8752 3770 8816
rect 2782 8666 2846 8730
rect 2866 8666 2930 8730
rect 2950 8666 3014 8730
rect 3034 8666 3098 8730
rect 3118 8666 3182 8730
rect 3202 8666 3266 8730
rect 3286 8666 3350 8730
rect 3370 8666 3434 8730
rect 3454 8666 3518 8730
rect 3538 8666 3602 8730
rect 3622 8666 3686 8730
rect 3706 8666 3770 8730
rect 2782 8579 2846 8643
rect 2866 8579 2930 8643
rect 2950 8579 3014 8643
rect 3034 8579 3098 8643
rect 3118 8579 3182 8643
rect 3202 8579 3266 8643
rect 3286 8579 3350 8643
rect 3370 8579 3434 8643
rect 3454 8579 3518 8643
rect 3538 8579 3602 8643
rect 3622 8579 3686 8643
rect 3706 8579 3770 8643
rect 2782 8492 2846 8556
rect 2866 8492 2930 8556
rect 2950 8492 3014 8556
rect 3034 8492 3098 8556
rect 3118 8492 3182 8556
rect 3202 8492 3266 8556
rect 3286 8492 3350 8556
rect 3370 8492 3434 8556
rect 3454 8492 3518 8556
rect 3538 8492 3602 8556
rect 3622 8492 3686 8556
rect 3706 8492 3770 8556
rect 2782 8405 2846 8469
rect 2866 8405 2930 8469
rect 2950 8405 3014 8469
rect 3034 8405 3098 8469
rect 3118 8405 3182 8469
rect 3202 8405 3266 8469
rect 3286 8405 3350 8469
rect 3370 8405 3434 8469
rect 3454 8405 3518 8469
rect 3538 8405 3602 8469
rect 3622 8405 3686 8469
rect 3706 8405 3770 8469
rect 2782 8318 2846 8382
rect 2866 8318 2930 8382
rect 2950 8318 3014 8382
rect 3034 8318 3098 8382
rect 3118 8318 3182 8382
rect 3202 8318 3266 8382
rect 3286 8318 3350 8382
rect 3370 8318 3434 8382
rect 3454 8318 3518 8382
rect 3538 8318 3602 8382
rect 3622 8318 3686 8382
rect 3706 8318 3770 8382
rect 4626 11528 4690 11533
rect 4626 11472 4681 11528
rect 4681 11472 4690 11528
rect 4626 11469 4690 11472
rect 4706 11528 4770 11533
rect 4706 11472 4715 11528
rect 4715 11472 4770 11528
rect 4706 11469 4770 11472
rect 4550 11282 4614 11346
rect 4634 11282 4698 11346
rect 4718 11282 4782 11346
rect 4550 10499 4614 10563
rect 4634 10499 4698 10563
rect 4718 10499 4782 10563
rect 4550 10415 4614 10479
rect 4634 10415 4698 10479
rect 4718 10415 4782 10479
rect 4550 10331 4614 10395
rect 4634 10331 4698 10395
rect 4718 10331 4782 10395
rect 4550 9548 4614 9612
rect 4634 9548 4698 9612
rect 4718 9548 4782 9612
rect 4332 7925 4396 7989
rect 4416 7925 4480 7989
rect 4499 7925 4563 7989
rect 4582 7925 4646 7989
rect 4665 7925 4729 7989
rect 4415 7840 4479 7904
rect 4499 7840 4563 7904
rect 4582 7840 4646 7904
rect 4665 7840 4729 7904
rect 4496 7754 4560 7818
rect 4581 7754 4645 7818
rect 4665 7754 4729 7818
rect 4578 7634 4642 7698
rect 4665 7634 4729 7698
rect 4454 7002 4518 7066
rect 4538 7002 4602 7066
rect 4622 7002 4686 7066
rect 4706 7002 4770 7066
rect 4454 6916 4518 6980
rect 4538 6916 4602 6980
rect 4622 6916 4686 6980
rect 4706 6916 4770 6980
rect 4454 6830 4518 6894
rect 4538 6830 4602 6894
rect 4622 6830 4686 6894
rect 4706 6830 4770 6894
rect 4454 6743 4518 6807
rect 4538 6743 4602 6807
rect 4622 6743 4686 6807
rect 4706 6743 4770 6807
rect 4454 6656 4518 6720
rect 4538 6656 4602 6720
rect 4622 6656 4686 6720
rect 4706 6656 4770 6720
rect 4454 6569 4518 6633
rect 4538 6569 4602 6633
rect 4622 6569 4686 6633
rect 4706 6569 4770 6633
rect 4454 6482 4518 6546
rect 4538 6482 4602 6546
rect 4622 6482 4686 6546
rect 4706 6482 4770 6546
rect 4454 6395 4518 6459
rect 4538 6395 4602 6459
rect 4622 6395 4686 6459
rect 4706 6395 4770 6459
rect 4918 3612 4982 3676
rect 5008 3612 5072 3676
rect 5098 3612 5162 3676
rect 5188 3612 5252 3676
rect 5278 3612 5342 3676
rect 5368 3612 5432 3676
rect 5458 3612 5522 3676
rect 4918 3526 4982 3590
rect 5008 3526 5072 3590
rect 5098 3526 5162 3590
rect 5188 3526 5252 3590
rect 5278 3526 5342 3590
rect 5368 3526 5432 3590
rect 5458 3526 5522 3590
rect 4918 3439 4982 3503
rect 5008 3439 5072 3503
rect 5098 3439 5162 3503
rect 5188 3439 5252 3503
rect 5278 3439 5342 3503
rect 5368 3439 5432 3503
rect 5458 3439 5522 3503
rect 4918 3352 4982 3416
rect 5008 3352 5072 3416
rect 5098 3352 5162 3416
rect 5188 3352 5252 3416
rect 5278 3352 5342 3416
rect 5368 3352 5432 3416
rect 5458 3352 5522 3416
rect 4918 3265 4982 3329
rect 5008 3265 5072 3329
rect 5098 3265 5162 3329
rect 5188 3265 5252 3329
rect 5278 3265 5342 3329
rect 5368 3265 5432 3329
rect 5458 3265 5522 3329
rect 4918 3178 4982 3242
rect 5008 3178 5072 3242
rect 5098 3178 5162 3242
rect 5188 3178 5252 3242
rect 5278 3178 5342 3242
rect 5368 3178 5432 3242
rect 5458 3178 5522 3242
rect 4918 3091 4982 3155
rect 5008 3091 5072 3155
rect 5098 3091 5162 3155
rect 5188 3091 5252 3155
rect 5278 3091 5342 3155
rect 5368 3091 5432 3155
rect 5458 3091 5522 3155
rect 4918 3004 4982 3068
rect 5008 3004 5072 3068
rect 5098 3004 5162 3068
rect 5188 3004 5252 3068
rect 5278 3004 5342 3068
rect 5368 3004 5432 3068
rect 5458 3004 5522 3068
rect 5648 13634 5712 13698
rect 5731 13634 5795 13698
rect 5814 13634 5878 13698
rect 5897 13634 5961 13698
rect 5980 13634 6044 13698
rect 6063 13634 6127 13698
rect 6146 13634 6210 13698
rect 6229 13634 6293 13698
rect 6312 13634 6376 13698
rect 6395 13634 6459 13698
rect 6478 13634 6542 13698
rect 6561 13634 6625 13698
rect 5648 13554 5712 13618
rect 5731 13554 5795 13618
rect 5814 13554 5878 13618
rect 5897 13554 5961 13618
rect 5980 13554 6044 13618
rect 6063 13554 6127 13618
rect 6146 13554 6210 13618
rect 6229 13554 6293 13618
rect 6312 13554 6376 13618
rect 6395 13554 6459 13618
rect 6478 13554 6542 13618
rect 6561 13554 6625 13618
rect 5648 13474 5712 13538
rect 5731 13474 5795 13538
rect 5814 13474 5878 13538
rect 5897 13474 5961 13538
rect 5980 13474 6044 13538
rect 6063 13474 6127 13538
rect 6146 13474 6210 13538
rect 6229 13474 6293 13538
rect 6312 13474 6376 13538
rect 6395 13474 6459 13538
rect 6478 13474 6542 13538
rect 6561 13474 6625 13538
rect 5648 13394 5712 13458
rect 5731 13394 5795 13458
rect 5814 13394 5878 13458
rect 5897 13394 5961 13458
rect 5980 13394 6044 13458
rect 6063 13394 6127 13458
rect 6146 13394 6210 13458
rect 6229 13394 6293 13458
rect 6312 13394 6376 13458
rect 6395 13394 6459 13458
rect 6478 13394 6542 13458
rect 6561 13394 6625 13458
rect 5648 13314 5712 13378
rect 5731 13314 5795 13378
rect 5814 13314 5878 13378
rect 5897 13314 5961 13378
rect 5980 13314 6044 13378
rect 6063 13314 6127 13378
rect 6146 13314 6210 13378
rect 6229 13314 6293 13378
rect 6312 13314 6376 13378
rect 6395 13314 6459 13378
rect 6478 13314 6542 13378
rect 6561 13314 6625 13378
rect 5648 13234 5712 13298
rect 5731 13234 5795 13298
rect 5814 13234 5878 13298
rect 5897 13234 5961 13298
rect 5980 13234 6044 13298
rect 6063 13234 6127 13298
rect 6146 13234 6210 13298
rect 6229 13234 6293 13298
rect 6312 13234 6376 13298
rect 6395 13234 6459 13298
rect 6478 13234 6542 13298
rect 6561 13234 6625 13298
rect 5648 13154 5712 13218
rect 5731 13154 5795 13218
rect 5814 13154 5878 13218
rect 5897 13154 5961 13218
rect 5980 13154 6044 13218
rect 6063 13154 6127 13218
rect 6146 13154 6210 13218
rect 6229 13154 6293 13218
rect 6312 13154 6376 13218
rect 6395 13154 6459 13218
rect 6478 13154 6542 13218
rect 6561 13154 6625 13218
rect 5648 13074 5712 13138
rect 5731 13074 5795 13138
rect 5814 13074 5878 13138
rect 5897 13074 5961 13138
rect 5980 13074 6044 13138
rect 6063 13074 6127 13138
rect 6146 13074 6210 13138
rect 6229 13074 6293 13138
rect 6312 13074 6376 13138
rect 6395 13074 6459 13138
rect 6478 13074 6542 13138
rect 6561 13074 6625 13138
rect 5648 12994 5712 13058
rect 5731 12994 5795 13058
rect 5814 12994 5878 13058
rect 5897 12994 5961 13058
rect 5980 12994 6044 13058
rect 6063 12994 6127 13058
rect 6146 12994 6210 13058
rect 6229 12994 6293 13058
rect 6312 12994 6376 13058
rect 6395 12994 6459 13058
rect 6478 12994 6542 13058
rect 6561 12994 6625 13058
rect 5648 12914 5712 12978
rect 5731 12914 5795 12978
rect 5814 12914 5878 12978
rect 5897 12914 5961 12978
rect 5980 12914 6044 12978
rect 6063 12914 6127 12978
rect 6146 12914 6210 12978
rect 6229 12914 6293 12978
rect 6312 12914 6376 12978
rect 6395 12914 6459 12978
rect 6478 12914 6542 12978
rect 6561 12914 6625 12978
rect 5648 12834 5712 12898
rect 5731 12834 5795 12898
rect 5814 12834 5878 12898
rect 5897 12834 5961 12898
rect 5980 12834 6044 12898
rect 6063 12834 6127 12898
rect 6146 12834 6210 12898
rect 6229 12834 6293 12898
rect 6312 12834 6376 12898
rect 6395 12834 6459 12898
rect 6478 12834 6542 12898
rect 6561 12834 6625 12898
rect 6705 11530 6760 11533
rect 6760 11530 6769 11533
rect 6705 11506 6769 11530
rect 6705 11469 6760 11506
rect 6760 11469 6769 11506
rect 6785 11469 6849 11533
rect 8171 11282 8235 11346
rect 8255 11282 8319 11346
rect 8339 11282 8403 11346
rect 9186 11282 9250 11346
rect 9270 11282 9334 11346
rect 9354 11282 9418 11346
rect 8171 10499 8235 10563
rect 8255 10499 8319 10563
rect 8339 10499 8403 10563
rect 8171 10415 8235 10479
rect 8255 10415 8319 10479
rect 8339 10415 8403 10479
rect 8171 10331 8235 10395
rect 8255 10331 8319 10395
rect 8339 10331 8403 10395
rect 8171 9548 8235 9612
rect 8255 9548 8319 9612
rect 8339 9548 8403 9612
rect 6916 9174 6980 9238
rect 7014 9174 7078 9238
rect 7112 9174 7176 9238
rect 6916 9089 6980 9153
rect 7014 9089 7078 9153
rect 7112 9089 7176 9153
rect 6916 9004 6980 9068
rect 7014 9004 7078 9068
rect 7112 9004 7176 9068
rect 6916 8919 6980 8983
rect 7014 8919 7078 8983
rect 7112 8919 7176 8983
rect 6916 8834 6980 8898
rect 7014 8834 7078 8898
rect 7112 8834 7176 8898
rect 6916 8749 6980 8813
rect 7014 8749 7078 8813
rect 7112 8749 7176 8813
rect 6916 8664 6980 8728
rect 7014 8664 7078 8728
rect 7112 8664 7176 8728
rect 6916 8579 6980 8643
rect 7014 8579 7078 8643
rect 7112 8579 7176 8643
rect 6916 8494 6980 8558
rect 7014 8494 7078 8558
rect 7112 8494 7176 8558
rect 6916 8408 6980 8472
rect 7014 8408 7078 8472
rect 7112 8408 7176 8472
rect 6916 8322 6980 8386
rect 7014 8322 7078 8386
rect 7112 8322 7176 8386
rect 9186 10499 9250 10563
rect 9270 10499 9334 10563
rect 9354 10499 9418 10563
rect 9186 10415 9250 10479
rect 9270 10415 9334 10479
rect 9354 10415 9418 10479
rect 9186 10331 9250 10395
rect 9270 10331 9334 10395
rect 9354 10331 9418 10395
rect 9186 9548 9250 9612
rect 9270 9548 9334 9612
rect 9354 9548 9418 9612
rect 8601 9177 8665 9241
rect 8699 9177 8763 9241
rect 8797 9177 8861 9241
rect 8601 9092 8665 9156
rect 8699 9092 8763 9156
rect 8797 9092 8861 9156
rect 8601 9006 8665 9070
rect 8699 9006 8763 9070
rect 8797 9006 8861 9070
rect 8601 8920 8665 8984
rect 8699 8920 8763 8984
rect 8797 8920 8861 8984
rect 8601 8834 8665 8898
rect 8699 8834 8763 8898
rect 8797 8834 8861 8898
rect 8601 8748 8665 8812
rect 8699 8748 8763 8812
rect 8797 8748 8861 8812
rect 8601 8662 8665 8726
rect 8699 8662 8763 8726
rect 8797 8662 8861 8726
rect 8601 8576 8665 8640
rect 8699 8576 8763 8640
rect 8797 8576 8861 8640
rect 8601 8490 8665 8554
rect 8699 8490 8763 8554
rect 8797 8490 8861 8554
rect 8601 8404 8665 8468
rect 8699 8404 8763 8468
rect 8797 8404 8861 8468
rect 8601 8318 8665 8382
rect 8699 8318 8763 8382
rect 8797 8318 8861 8382
rect 9114 9209 9121 9241
rect 9121 9209 9177 9241
rect 9177 9209 9178 9241
rect 9114 9178 9178 9209
rect 9114 9177 9121 9178
rect 9121 9177 9177 9178
rect 9177 9177 9178 9178
rect 9198 9209 9217 9241
rect 9217 9209 9262 9241
rect 9282 9209 9313 9241
rect 9313 9209 9346 9241
rect 9366 9209 9369 9241
rect 9369 9209 9409 9241
rect 9409 9209 9430 9241
rect 9450 9209 9465 9241
rect 9465 9209 9505 9241
rect 9505 9209 9514 9241
rect 9534 9209 9561 9241
rect 9561 9209 9598 9241
rect 9198 9178 9262 9209
rect 9282 9178 9346 9209
rect 9366 9178 9430 9209
rect 9450 9178 9514 9209
rect 9534 9178 9598 9209
rect 9198 9177 9217 9178
rect 9217 9177 9262 9178
rect 9282 9177 9313 9178
rect 9313 9177 9346 9178
rect 9366 9177 9369 9178
rect 9369 9177 9409 9178
rect 9409 9177 9430 9178
rect 9450 9177 9465 9178
rect 9465 9177 9505 9178
rect 9505 9177 9514 9178
rect 9534 9177 9561 9178
rect 9561 9177 9598 9178
rect 9618 9177 9682 9241
rect 9114 9122 9121 9156
rect 9121 9122 9177 9156
rect 9177 9122 9178 9156
rect 9114 9092 9178 9122
rect 9198 9122 9217 9156
rect 9217 9122 9262 9156
rect 9282 9122 9313 9156
rect 9313 9122 9346 9156
rect 9366 9122 9369 9156
rect 9369 9122 9409 9156
rect 9409 9122 9430 9156
rect 9450 9122 9465 9156
rect 9465 9122 9505 9156
rect 9505 9122 9514 9156
rect 9534 9122 9561 9156
rect 9561 9122 9598 9156
rect 9198 9092 9262 9122
rect 9282 9092 9346 9122
rect 9366 9092 9430 9122
rect 9450 9092 9514 9122
rect 9534 9092 9598 9122
rect 9618 9092 9682 9156
rect 9114 9035 9121 9071
rect 9121 9035 9177 9071
rect 9177 9035 9178 9071
rect 9114 9007 9178 9035
rect 9198 9035 9217 9071
rect 9217 9035 9262 9071
rect 9282 9035 9313 9071
rect 9313 9035 9346 9071
rect 9366 9035 9369 9071
rect 9369 9035 9409 9071
rect 9409 9035 9430 9071
rect 9450 9035 9465 9071
rect 9465 9035 9505 9071
rect 9505 9035 9514 9071
rect 9534 9035 9561 9071
rect 9561 9035 9598 9071
rect 9198 9007 9262 9035
rect 9282 9007 9346 9035
rect 9366 9007 9430 9035
rect 9450 9007 9514 9035
rect 9534 9007 9598 9035
rect 9618 9007 9682 9071
rect 9114 8948 9121 8986
rect 9121 8948 9177 8986
rect 9177 8948 9178 8986
rect 9114 8922 9178 8948
rect 9198 8948 9217 8986
rect 9217 8948 9262 8986
rect 9282 8948 9313 8986
rect 9313 8948 9346 8986
rect 9366 8948 9369 8986
rect 9369 8948 9409 8986
rect 9409 8948 9430 8986
rect 9450 8948 9465 8986
rect 9465 8948 9505 8986
rect 9505 8948 9514 8986
rect 9534 8948 9561 8986
rect 9561 8948 9598 8986
rect 9198 8922 9262 8948
rect 9282 8922 9346 8948
rect 9366 8922 9430 8948
rect 9450 8922 9514 8948
rect 9534 8922 9598 8948
rect 9618 8922 9682 8986
rect 9114 8861 9121 8901
rect 9121 8861 9177 8901
rect 9177 8861 9178 8901
rect 9114 8837 9178 8861
rect 9198 8861 9217 8901
rect 9217 8861 9262 8901
rect 9282 8861 9313 8901
rect 9313 8861 9346 8901
rect 9366 8861 9369 8901
rect 9369 8861 9409 8901
rect 9409 8861 9430 8901
rect 9450 8861 9465 8901
rect 9465 8861 9505 8901
rect 9505 8861 9514 8901
rect 9534 8861 9561 8901
rect 9561 8861 9598 8901
rect 9198 8837 9262 8861
rect 9282 8837 9346 8861
rect 9366 8837 9430 8861
rect 9450 8837 9514 8861
rect 9534 8837 9598 8861
rect 9618 8837 9682 8901
rect 9114 8774 9121 8816
rect 9121 8774 9177 8816
rect 9177 8774 9178 8816
rect 9114 8752 9178 8774
rect 9198 8774 9217 8816
rect 9217 8774 9262 8816
rect 9282 8774 9313 8816
rect 9313 8774 9346 8816
rect 9366 8774 9369 8816
rect 9369 8774 9409 8816
rect 9409 8774 9430 8816
rect 9450 8774 9465 8816
rect 9465 8774 9505 8816
rect 9505 8774 9514 8816
rect 9534 8774 9561 8816
rect 9561 8774 9598 8816
rect 9198 8752 9262 8774
rect 9282 8752 9346 8774
rect 9366 8752 9430 8774
rect 9450 8752 9514 8774
rect 9534 8752 9598 8774
rect 9618 8752 9682 8816
rect 9114 8686 9121 8731
rect 9121 8686 9177 8731
rect 9177 8686 9178 8731
rect 9114 8667 9178 8686
rect 9198 8686 9217 8731
rect 9217 8686 9262 8731
rect 9282 8686 9313 8731
rect 9313 8686 9346 8731
rect 9366 8686 9369 8731
rect 9369 8686 9409 8731
rect 9409 8686 9430 8731
rect 9450 8686 9465 8731
rect 9465 8686 9505 8731
rect 9505 8686 9514 8731
rect 9534 8686 9561 8731
rect 9561 8686 9598 8731
rect 9198 8667 9262 8686
rect 9282 8667 9346 8686
rect 9366 8667 9430 8686
rect 9450 8667 9514 8686
rect 9534 8667 9598 8686
rect 9618 8667 9682 8731
rect 9114 8598 9121 8645
rect 9121 8598 9177 8645
rect 9177 8598 9178 8645
rect 9114 8581 9178 8598
rect 9198 8598 9217 8645
rect 9217 8598 9262 8645
rect 9282 8598 9313 8645
rect 9313 8598 9346 8645
rect 9366 8598 9369 8645
rect 9369 8598 9409 8645
rect 9409 8598 9430 8645
rect 9450 8598 9465 8645
rect 9465 8598 9505 8645
rect 9505 8598 9514 8645
rect 9534 8598 9561 8645
rect 9561 8598 9598 8645
rect 9198 8581 9262 8598
rect 9282 8581 9346 8598
rect 9366 8581 9430 8598
rect 9450 8581 9514 8598
rect 9534 8581 9598 8598
rect 9618 8581 9682 8645
rect 9114 8510 9121 8559
rect 9121 8510 9177 8559
rect 9177 8510 9178 8559
rect 9114 8495 9178 8510
rect 9198 8510 9217 8559
rect 9217 8510 9262 8559
rect 9282 8510 9313 8559
rect 9313 8510 9346 8559
rect 9366 8510 9369 8559
rect 9369 8510 9409 8559
rect 9409 8510 9430 8559
rect 9450 8510 9465 8559
rect 9465 8510 9505 8559
rect 9505 8510 9514 8559
rect 9534 8510 9561 8559
rect 9561 8510 9598 8559
rect 9198 8495 9262 8510
rect 9282 8495 9346 8510
rect 9366 8495 9430 8510
rect 9450 8495 9514 8510
rect 9534 8495 9598 8510
rect 9618 8495 9682 8559
rect 9114 8422 9121 8473
rect 9121 8422 9177 8473
rect 9177 8422 9178 8473
rect 9114 8409 9178 8422
rect 9198 8422 9217 8473
rect 9217 8422 9262 8473
rect 9282 8422 9313 8473
rect 9313 8422 9346 8473
rect 9366 8422 9369 8473
rect 9369 8422 9409 8473
rect 9409 8422 9430 8473
rect 9450 8422 9465 8473
rect 9465 8422 9505 8473
rect 9505 8422 9514 8473
rect 9534 8422 9561 8473
rect 9561 8422 9598 8473
rect 9198 8409 9262 8422
rect 9282 8409 9346 8422
rect 9366 8409 9430 8422
rect 9450 8409 9514 8422
rect 9534 8409 9598 8422
rect 9618 8409 9682 8473
rect 9114 8334 9121 8387
rect 9121 8334 9177 8387
rect 9177 8334 9178 8387
rect 9114 8323 9178 8334
rect 9198 8334 9217 8387
rect 9217 8334 9262 8387
rect 9282 8334 9313 8387
rect 9313 8334 9346 8387
rect 9366 8334 9369 8387
rect 9369 8334 9409 8387
rect 9409 8334 9430 8387
rect 9450 8334 9465 8387
rect 9465 8334 9505 8387
rect 9505 8334 9514 8387
rect 9534 8334 9561 8387
rect 9561 8334 9598 8387
rect 9198 8323 9262 8334
rect 9282 8323 9346 8334
rect 9366 8323 9430 8334
rect 9450 8323 9514 8334
rect 9534 8323 9598 8334
rect 9618 8323 9682 8387
rect 6847 2653 6911 2706
rect 6847 2642 6903 2653
rect 6903 2642 6911 2653
rect 6927 2653 6991 2706
rect 6927 2642 6931 2653
rect 6931 2642 6987 2653
rect 6987 2642 6991 2653
rect 7007 2653 7071 2706
rect 7007 2642 7015 2653
rect 7015 2642 7071 2653
rect 6847 2597 6903 2620
rect 6903 2597 6911 2620
rect 6847 2556 6911 2597
rect 6927 2597 6931 2620
rect 6931 2597 6987 2620
rect 6987 2597 6991 2620
rect 6927 2556 6991 2597
rect 7007 2597 7015 2620
rect 7015 2597 7071 2620
rect 7007 2556 7071 2597
rect 6847 2530 6911 2534
rect 6847 2474 6903 2530
rect 6903 2474 6911 2530
rect 6847 2470 6911 2474
rect 6927 2530 6991 2534
rect 6927 2474 6931 2530
rect 6931 2474 6987 2530
rect 6987 2474 6991 2530
rect 6927 2470 6991 2474
rect 7007 2530 7071 2534
rect 7007 2474 7015 2530
rect 7015 2474 7071 2530
rect 7007 2470 7071 2474
rect 6847 2407 6911 2448
rect 6847 2384 6903 2407
rect 6903 2384 6911 2407
rect 6927 2407 6991 2448
rect 6927 2384 6931 2407
rect 6931 2384 6987 2407
rect 6987 2384 6991 2407
rect 7007 2407 7071 2448
rect 7007 2384 7015 2407
rect 7015 2384 7071 2407
rect 6847 2351 6903 2362
rect 6903 2351 6911 2362
rect 6847 2298 6911 2351
rect 6927 2351 6931 2362
rect 6931 2351 6987 2362
rect 6987 2351 6991 2362
rect 6927 2298 6991 2351
rect 7007 2351 7015 2362
rect 7015 2351 7071 2362
rect 7007 2298 7071 2351
rect 6847 2228 6903 2276
rect 6903 2228 6911 2276
rect 6847 2212 6911 2228
rect 6927 2228 6931 2276
rect 6931 2228 6987 2276
rect 6987 2228 6991 2276
rect 6927 2212 6991 2228
rect 7007 2228 7015 2276
rect 7015 2228 7071 2276
rect 7007 2212 7071 2228
rect 6847 2161 6911 2190
rect 6847 2126 6903 2161
rect 6903 2126 6911 2161
rect 6927 2161 6991 2190
rect 6927 2126 6931 2161
rect 6931 2126 6987 2161
rect 6987 2126 6991 2161
rect 7007 2161 7071 2190
rect 7007 2126 7015 2161
rect 7015 2126 7071 2161
rect 6847 2039 6911 2103
rect 6927 2039 6991 2103
rect 7007 2039 7071 2103
rect 6847 1982 6903 2016
rect 6903 1982 6911 2016
rect 6847 1952 6911 1982
rect 6927 1982 6931 2016
rect 6931 1982 6987 2016
rect 6987 1982 6991 2016
rect 6927 1952 6991 1982
rect 7007 1982 7015 2016
rect 7015 1982 7071 2016
rect 7007 1952 7071 1982
rect 6847 1915 6911 1929
rect 6847 1865 6903 1915
rect 6903 1865 6911 1915
rect 6927 1915 6991 1929
rect 6927 1865 6931 1915
rect 6931 1865 6987 1915
rect 6987 1865 6991 1915
rect 7007 1915 7071 1929
rect 7007 1865 7015 1915
rect 7015 1865 7071 1915
rect 6847 1778 6911 1842
rect 6927 1778 6991 1842
rect 7007 1778 7071 1842
rect 8610 2657 8674 2706
rect 8610 2642 8615 2657
rect 8615 2642 8671 2657
rect 8671 2642 8674 2657
rect 8716 2657 8780 2706
rect 8716 2642 8719 2657
rect 8719 2642 8775 2657
rect 8775 2642 8780 2657
rect 8610 2601 8615 2621
rect 8615 2601 8671 2621
rect 8671 2601 8674 2621
rect 8610 2557 8674 2601
rect 8716 2601 8719 2621
rect 8719 2601 8775 2621
rect 8775 2601 8780 2621
rect 8716 2557 8780 2601
rect 8610 2535 8674 2536
rect 8610 2479 8615 2535
rect 8615 2479 8671 2535
rect 8671 2479 8674 2535
rect 8610 2472 8674 2479
rect 8716 2535 8780 2536
rect 8716 2479 8719 2535
rect 8719 2479 8775 2535
rect 8775 2479 8780 2535
rect 8716 2472 8780 2479
rect 8610 2412 8674 2450
rect 8610 2386 8615 2412
rect 8615 2386 8671 2412
rect 8671 2386 8674 2412
rect 8716 2412 8780 2450
rect 8716 2386 8719 2412
rect 8719 2386 8775 2412
rect 8775 2386 8780 2412
rect 8610 2356 8615 2364
rect 8615 2356 8671 2364
rect 8671 2356 8674 2364
rect 8610 2300 8674 2356
rect 8716 2356 8719 2364
rect 8719 2356 8775 2364
rect 8775 2356 8780 2364
rect 8716 2300 8780 2356
rect 8610 2233 8615 2278
rect 8615 2233 8671 2278
rect 8671 2233 8674 2278
rect 8610 2214 8674 2233
rect 8716 2233 8719 2278
rect 8719 2233 8775 2278
rect 8775 2233 8780 2278
rect 8716 2214 8780 2233
rect 8610 2166 8674 2192
rect 8610 2128 8615 2166
rect 8615 2128 8671 2166
rect 8671 2128 8674 2166
rect 8716 2166 8780 2192
rect 8716 2128 8719 2166
rect 8719 2128 8775 2166
rect 8775 2128 8780 2166
rect 8610 2043 8674 2106
rect 8610 2042 8615 2043
rect 8615 2042 8671 2043
rect 8671 2042 8674 2043
rect 8716 2043 8780 2106
rect 8716 2042 8719 2043
rect 8719 2042 8775 2043
rect 8775 2042 8780 2043
rect 8610 1987 8615 2020
rect 8615 1987 8671 2020
rect 8671 1987 8674 2020
rect 8610 1956 8674 1987
rect 8716 1987 8719 2020
rect 8719 1987 8775 2020
rect 8775 1987 8780 2020
rect 8716 1956 8780 1987
rect 8610 1870 8674 1934
rect 8716 1870 8780 1934
rect 8610 1784 8674 1848
rect 8716 1784 8780 1848
rect 2230 504 2294 568
rect 2310 504 2374 568
rect 2390 504 2454 568
rect 2470 504 2534 568
rect 2550 504 2614 568
rect 2630 504 2694 568
rect 2230 419 2294 483
rect 2310 419 2374 483
rect 2390 419 2454 483
rect 2470 419 2534 483
rect 2550 419 2614 483
rect 2630 419 2694 483
rect 9382 7174 9446 7238
rect 9462 7174 9526 7238
rect 9598 7174 9662 7238
rect 9678 7174 9742 7238
rect 9815 7174 9879 7238
rect 9895 7174 9959 7238
rect 12128 9408 12192 9472
rect 12209 9408 12273 9472
rect 10026 3612 10090 3676
rect 10138 3612 10202 3676
rect 10250 3612 10314 3676
rect 10026 3526 10090 3590
rect 10138 3526 10202 3590
rect 10250 3526 10314 3590
rect 10026 3439 10090 3503
rect 10138 3439 10202 3503
rect 10250 3439 10314 3503
rect 10026 3352 10090 3416
rect 10138 3352 10202 3416
rect 10250 3352 10314 3416
rect 10026 3265 10090 3329
rect 10138 3265 10202 3329
rect 10250 3265 10314 3329
rect 10026 3178 10090 3242
rect 10138 3178 10202 3242
rect 10250 3178 10314 3242
rect 10026 3091 10090 3155
rect 10138 3091 10202 3155
rect 10250 3091 10314 3155
rect 10026 3004 10090 3068
rect 10138 3004 10202 3068
rect 10250 3004 10314 3068
rect 10503 9174 10567 9238
rect 10585 9174 10649 9238
rect 10667 9174 10731 9238
rect 10749 9174 10813 9238
rect 10831 9174 10895 9238
rect 10913 9174 10977 9238
rect 10995 9174 11059 9238
rect 11077 9174 11141 9238
rect 10503 9090 10567 9154
rect 10585 9090 10649 9154
rect 10667 9090 10731 9154
rect 10749 9090 10813 9154
rect 10831 9090 10895 9154
rect 10913 9090 10977 9154
rect 10995 9090 11059 9154
rect 11077 9090 11141 9154
rect 10503 9006 10567 9070
rect 10585 9006 10649 9070
rect 10667 9006 10731 9070
rect 10749 9006 10813 9070
rect 10831 9006 10895 9070
rect 10913 9006 10977 9070
rect 10995 9006 11059 9070
rect 11077 9006 11141 9070
rect 10503 8922 10567 8986
rect 10585 8922 10649 8986
rect 10667 8922 10731 8986
rect 10749 8922 10813 8986
rect 10831 8922 10895 8986
rect 10913 8922 10977 8986
rect 10995 8922 11059 8986
rect 11077 8922 11141 8986
rect 10503 8838 10567 8902
rect 10585 8838 10649 8902
rect 10667 8838 10731 8902
rect 10749 8838 10813 8902
rect 10831 8838 10895 8902
rect 10913 8838 10977 8902
rect 10995 8838 11059 8902
rect 11077 8838 11141 8902
rect 10503 8754 10567 8818
rect 10585 8754 10649 8818
rect 10667 8754 10731 8818
rect 10749 8754 10813 8818
rect 10831 8754 10895 8818
rect 10913 8754 10977 8818
rect 10995 8754 11059 8818
rect 11077 8754 11141 8818
rect 10503 8670 10567 8734
rect 10585 8670 10649 8734
rect 10667 8670 10731 8734
rect 10749 8670 10813 8734
rect 10831 8670 10895 8734
rect 10913 8670 10977 8734
rect 10995 8670 11059 8734
rect 11077 8670 11141 8734
rect 10503 8586 10567 8650
rect 10585 8586 10649 8650
rect 10667 8586 10731 8650
rect 10749 8586 10813 8650
rect 10831 8586 10895 8650
rect 10913 8586 10977 8650
rect 10995 8586 11059 8650
rect 11077 8586 11141 8650
rect 10503 8502 10567 8566
rect 10585 8502 10649 8566
rect 10667 8502 10731 8566
rect 10749 8502 10813 8566
rect 10831 8502 10895 8566
rect 10913 8502 10977 8566
rect 10995 8502 11059 8566
rect 11077 8502 11141 8566
rect 10503 8418 10567 8482
rect 10585 8418 10649 8482
rect 10667 8418 10731 8482
rect 10749 8418 10813 8482
rect 10831 8418 10895 8482
rect 10913 8418 10977 8482
rect 10995 8418 11059 8482
rect 11077 8418 11141 8482
rect 10503 8333 10567 8397
rect 10585 8333 10649 8397
rect 10667 8333 10731 8397
rect 10749 8333 10813 8397
rect 10831 8333 10895 8397
rect 10913 8333 10977 8397
rect 10995 8333 11059 8397
rect 11077 8333 11141 8397
rect 12674 7966 12738 8030
rect 12755 7966 12819 8030
rect 12836 7966 12900 8030
rect 12917 7966 12981 8030
rect 12998 7966 13062 8030
rect 13078 7966 13142 8030
rect 13158 7966 13222 8030
rect 13238 7966 13302 8030
rect 13318 7966 13382 8030
rect 13398 7966 13462 8030
rect 12674 7880 12738 7944
rect 12755 7880 12819 7944
rect 12836 7880 12900 7944
rect 12917 7880 12981 7944
rect 12998 7880 13062 7944
rect 13078 7880 13142 7944
rect 13158 7880 13222 7944
rect 13238 7880 13302 7944
rect 13318 7880 13382 7944
rect 13398 7880 13462 7944
rect 12674 7794 12738 7858
rect 12755 7794 12819 7858
rect 12836 7794 12900 7858
rect 12917 7794 12981 7858
rect 12998 7794 13062 7858
rect 13078 7794 13142 7858
rect 13158 7794 13222 7858
rect 13238 7794 13302 7858
rect 13318 7794 13382 7858
rect 13398 7794 13462 7858
rect 12674 7708 12738 7772
rect 12755 7708 12819 7772
rect 12836 7708 12900 7772
rect 12917 7708 12981 7772
rect 12998 7708 13062 7772
rect 13078 7708 13142 7772
rect 13158 7708 13222 7772
rect 13238 7708 13302 7772
rect 13318 7708 13382 7772
rect 13398 7708 13462 7772
rect 12674 7622 12738 7686
rect 12755 7622 12819 7686
rect 12836 7622 12900 7686
rect 12917 7622 12981 7686
rect 12998 7622 13062 7686
rect 13078 7622 13142 7686
rect 13158 7622 13222 7686
rect 13238 7622 13302 7686
rect 13318 7622 13382 7686
rect 13398 7622 13462 7686
rect 12674 7536 12738 7600
rect 12755 7536 12819 7600
rect 12836 7536 12900 7600
rect 12917 7536 12981 7600
rect 12998 7536 13062 7600
rect 13078 7536 13142 7600
rect 13158 7536 13222 7600
rect 13238 7536 13302 7600
rect 13318 7536 13382 7600
rect 13398 7536 13462 7600
rect 12674 7450 12738 7514
rect 12755 7450 12819 7514
rect 12836 7450 12900 7514
rect 12917 7450 12981 7514
rect 12998 7450 13062 7514
rect 13078 7450 13142 7514
rect 13158 7450 13222 7514
rect 13238 7450 13302 7514
rect 13318 7450 13382 7514
rect 13398 7450 13462 7514
rect 12674 7364 12738 7428
rect 12755 7364 12819 7428
rect 12836 7364 12900 7428
rect 12917 7364 12981 7428
rect 12998 7364 13062 7428
rect 13078 7364 13142 7428
rect 13158 7364 13222 7428
rect 13238 7364 13302 7428
rect 13318 7364 13382 7428
rect 13398 7364 13462 7428
rect 11342 2642 11406 2706
rect 11442 2642 11506 2706
rect 11542 2642 11606 2706
rect 11642 2642 11706 2706
rect 11342 2557 11406 2621
rect 11442 2557 11506 2621
rect 11542 2557 11606 2621
rect 11642 2557 11706 2621
rect 11342 2472 11406 2536
rect 11442 2472 11506 2536
rect 11542 2472 11606 2536
rect 11642 2472 11706 2536
rect 11342 2387 11406 2451
rect 11442 2387 11506 2451
rect 11542 2387 11606 2451
rect 11642 2387 11706 2451
rect 11342 2302 11406 2366
rect 11442 2302 11506 2366
rect 11542 2302 11606 2366
rect 11642 2302 11706 2366
rect 11342 2216 11406 2280
rect 11442 2216 11506 2280
rect 11542 2216 11606 2280
rect 11642 2216 11706 2280
rect 11342 2130 11406 2194
rect 11442 2130 11506 2194
rect 11542 2130 11606 2194
rect 11642 2130 11706 2194
rect 11342 2044 11406 2108
rect 11442 2044 11506 2108
rect 11542 2044 11606 2108
rect 11642 2044 11706 2108
rect 11342 1958 11406 2022
rect 11442 1958 11506 2022
rect 11542 1958 11606 2022
rect 11642 1958 11706 2022
rect 11342 1872 11406 1936
rect 11442 1872 11506 1936
rect 11542 1872 11606 1936
rect 11642 1872 11706 1936
rect 11342 1786 11406 1850
rect 11442 1786 11506 1850
rect 11542 1786 11606 1850
rect 11642 1786 11706 1850
rect 14139 4817 14203 4881
rect 14283 4817 14347 4881
rect 14139 4732 14203 4796
rect 14283 4732 14347 4796
rect 14139 4647 14203 4711
rect 14283 4647 14347 4711
rect 14139 4562 14203 4626
rect 14283 4562 14347 4626
rect 14139 4477 14203 4541
rect 14283 4477 14347 4541
rect 14139 4392 14203 4456
rect 14283 4392 14347 4456
rect 14139 4307 14203 4371
rect 14283 4307 14347 4371
rect 14139 4222 14203 4286
rect 14283 4222 14347 4286
rect 14139 4137 14203 4201
rect 14283 4137 14347 4201
rect 14139 4051 14203 4115
rect 14283 4051 14347 4115
rect 14139 3965 14203 4029
rect 14283 3965 14347 4029
rect 13569 2642 13633 2706
rect 13653 2642 13717 2706
rect 13737 2642 13801 2706
rect 13821 2642 13885 2706
rect 13905 2642 13969 2706
rect 13989 2642 14053 2706
rect 13569 2557 13633 2621
rect 13653 2557 13717 2621
rect 13737 2557 13801 2621
rect 13821 2557 13885 2621
rect 13905 2557 13969 2621
rect 13989 2557 14053 2621
rect 13569 2471 13633 2535
rect 13653 2471 13717 2535
rect 13737 2471 13801 2535
rect 13821 2471 13885 2535
rect 13905 2471 13969 2535
rect 13989 2471 14053 2535
rect 13569 2385 13633 2449
rect 13653 2385 13717 2449
rect 13737 2385 13801 2449
rect 13821 2385 13885 2449
rect 13905 2385 13969 2449
rect 13989 2385 14053 2449
rect 13569 2299 13633 2363
rect 13653 2299 13717 2363
rect 13737 2299 13801 2363
rect 13821 2299 13885 2363
rect 13905 2299 13969 2363
rect 13989 2299 14053 2363
rect 13569 2213 13633 2277
rect 13653 2213 13717 2277
rect 13737 2213 13801 2277
rect 13821 2213 13885 2277
rect 13905 2213 13969 2277
rect 13989 2213 14053 2277
rect 13569 2127 13633 2191
rect 13653 2127 13717 2191
rect 13737 2127 13801 2191
rect 13821 2127 13885 2191
rect 13905 2127 13969 2191
rect 13989 2127 14053 2191
rect 13569 2041 13633 2105
rect 13653 2041 13717 2105
rect 13737 2041 13801 2105
rect 13821 2041 13885 2105
rect 13905 2041 13969 2105
rect 13989 2041 14053 2105
rect 13569 1955 13633 2019
rect 13653 1955 13717 2019
rect 13737 1955 13801 2019
rect 13821 1955 13885 2019
rect 13905 1955 13969 2019
rect 13989 1955 14053 2019
rect 13569 1869 13633 1933
rect 13653 1869 13717 1933
rect 13737 1869 13801 1933
rect 13821 1869 13885 1933
rect 13905 1869 13969 1933
rect 13989 1869 14053 1933
rect 13569 1783 13633 1847
rect 13653 1783 13717 1847
rect 13737 1783 13801 1847
rect 13821 1783 13885 1847
rect 13905 1783 13969 1847
rect 13989 1783 14053 1847
rect 10343 293 10407 298
rect 10343 237 10347 293
rect 10347 237 10403 293
rect 10403 237 10407 293
rect 10343 234 10407 237
rect 10423 293 10487 298
rect 10423 237 10427 293
rect 10427 237 10483 293
rect 10483 237 10487 293
rect 10423 234 10487 237
rect 10714 234 10778 298
rect 10794 234 10858 298
rect 11207 234 11271 298
rect 11287 234 11351 298
rect 14438 1422 14502 1486
rect 14524 1422 14588 1486
rect 14610 1422 14674 1486
rect 14696 1422 14760 1486
rect 14782 1422 14846 1486
rect 14868 1422 14932 1486
rect 14954 1422 15018 1486
rect 15040 1422 15104 1486
rect 15126 1422 15190 1486
rect 15212 1422 15276 1486
rect 15298 1422 15362 1486
rect 14438 1337 14502 1401
rect 14524 1337 14588 1401
rect 14610 1337 14674 1401
rect 14696 1337 14760 1401
rect 14782 1337 14846 1401
rect 14868 1337 14932 1401
rect 14954 1337 15018 1401
rect 15040 1337 15104 1401
rect 15126 1337 15190 1401
rect 15212 1337 15276 1401
rect 15298 1337 15362 1401
rect 14438 1252 14502 1316
rect 14524 1252 14588 1316
rect 14610 1252 14674 1316
rect 14696 1252 14760 1316
rect 14782 1252 14846 1316
rect 14868 1252 14932 1316
rect 14954 1252 15018 1316
rect 15040 1252 15104 1316
rect 15126 1252 15190 1316
rect 15212 1252 15276 1316
rect 15298 1252 15362 1316
rect 14438 1166 14502 1230
rect 14524 1166 14588 1230
rect 14610 1166 14674 1230
rect 14696 1166 14760 1230
rect 14782 1166 14846 1230
rect 14868 1166 14932 1230
rect 14954 1166 15018 1230
rect 15040 1166 15104 1230
rect 15126 1166 15190 1230
rect 15212 1166 15276 1230
rect 15298 1166 15362 1230
rect 14438 1080 14502 1144
rect 14524 1080 14588 1144
rect 14610 1080 14674 1144
rect 14696 1080 14760 1144
rect 14782 1080 14846 1144
rect 14868 1080 14932 1144
rect 14954 1080 15018 1144
rect 15040 1080 15104 1144
rect 15126 1080 15190 1144
rect 15212 1080 15276 1144
rect 15298 1080 15362 1144
rect 14438 994 14502 1058
rect 14524 994 14588 1058
rect 14610 994 14674 1058
rect 14696 994 14760 1058
rect 14782 994 14846 1058
rect 14868 994 14932 1058
rect 14954 994 15018 1058
rect 15040 994 15104 1058
rect 15126 994 15190 1058
rect 15212 994 15276 1058
rect 15298 994 15362 1058
rect 14438 908 14502 972
rect 14524 908 14588 972
rect 14610 908 14674 972
rect 14696 908 14760 972
rect 14782 908 14846 972
rect 14868 908 14932 972
rect 14954 908 15018 972
rect 15040 908 15104 972
rect 15126 908 15190 972
rect 15212 908 15276 972
rect 15298 908 15362 972
rect 14438 822 14502 886
rect 14524 822 14588 886
rect 14610 822 14674 886
rect 14696 822 14760 886
rect 14782 822 14846 886
rect 14868 822 14932 886
rect 14954 822 15018 886
rect 15040 822 15104 886
rect 15126 822 15190 886
rect 15212 822 15276 886
rect 15298 822 15362 886
rect 14438 736 14502 800
rect 14524 736 14588 800
rect 14610 736 14674 800
rect 14696 736 14760 800
rect 14782 736 14846 800
rect 14868 736 14932 800
rect 14954 736 15018 800
rect 15040 736 15104 800
rect 15126 736 15190 800
rect 15212 736 15276 800
rect 15298 736 15362 800
rect 14438 650 14502 714
rect 14524 650 14588 714
rect 14610 650 14674 714
rect 14696 650 14760 714
rect 14782 650 14846 714
rect 14868 650 14932 714
rect 14954 650 15018 714
rect 15040 650 15104 714
rect 15126 650 15190 714
rect 15212 650 15276 714
rect 15298 650 15362 714
rect 14438 564 14502 628
rect 14524 564 14588 628
rect 14610 564 14674 628
rect 14696 564 14760 628
rect 14782 564 14846 628
rect 14868 564 14932 628
rect 14954 564 15018 628
rect 15040 564 15104 628
rect 15126 564 15190 628
rect 15212 564 15276 628
rect 15298 564 15362 628
rect 13013 234 13077 298
rect 13093 234 13157 298
rect 13318 295 13382 298
rect 13318 239 13373 295
rect 13373 239 13382 295
rect 13318 234 13382 239
rect 13398 295 13462 298
rect 13398 239 13407 295
rect 13407 239 13462 295
rect 13398 234 13462 239
rect 15030 234 15094 298
rect 15110 234 15174 298
rect 15488 293 15552 298
rect 15488 237 15543 293
rect 15543 237 15552 293
rect 15488 234 15552 237
rect 15568 293 15632 298
rect 15568 237 15577 293
rect 15577 237 15632 293
rect 15568 234 15632 237
<< metal4 >>
rect 0 35157 254 40000
rect 12586 39372 13006 39373
rect 5105 39365 6299 39366
rect 5105 39301 5110 39365
rect 5174 39301 5190 39365
rect 5254 39301 5270 39365
rect 5334 39301 5350 39365
rect 5414 39301 5430 39365
rect 5494 39301 5510 39365
rect 5574 39301 5590 39365
rect 5654 39301 5670 39365
rect 5734 39301 5750 39365
rect 5814 39301 5830 39365
rect 5894 39301 5910 39365
rect 5974 39301 5990 39365
rect 6054 39301 6070 39365
rect 6134 39301 6150 39365
rect 6214 39301 6230 39365
rect 6294 39301 6299 39365
rect 5105 39284 6299 39301
rect 5105 39220 5110 39284
rect 5174 39220 5190 39284
rect 5254 39220 5270 39284
rect 5334 39220 5350 39284
rect 5414 39220 5430 39284
rect 5494 39220 5510 39284
rect 5574 39220 5590 39284
rect 5654 39220 5670 39284
rect 5734 39220 5750 39284
rect 5814 39220 5830 39284
rect 5894 39220 5910 39284
rect 5974 39220 5990 39284
rect 6054 39220 6070 39284
rect 6134 39220 6150 39284
rect 6214 39220 6230 39284
rect 6294 39220 6299 39284
rect 5105 39203 6299 39220
rect 5105 39139 5110 39203
rect 5174 39139 5190 39203
rect 5254 39139 5270 39203
rect 5334 39139 5350 39203
rect 5414 39139 5430 39203
rect 5494 39139 5510 39203
rect 5574 39139 5590 39203
rect 5654 39139 5670 39203
rect 5734 39139 5750 39203
rect 5814 39139 5830 39203
rect 5894 39139 5910 39203
rect 5974 39139 5990 39203
rect 6054 39139 6070 39203
rect 6134 39139 6150 39203
rect 6214 39139 6230 39203
rect 6294 39139 6299 39203
rect 5105 39122 6299 39139
rect 5105 39058 5110 39122
rect 5174 39058 5190 39122
rect 5254 39058 5270 39122
rect 5334 39058 5350 39122
rect 5414 39058 5430 39122
rect 5494 39058 5510 39122
rect 5574 39058 5590 39122
rect 5654 39058 5670 39122
rect 5734 39058 5750 39122
rect 5814 39058 5830 39122
rect 5894 39058 5910 39122
rect 5974 39058 5990 39122
rect 6054 39058 6070 39122
rect 6134 39058 6150 39122
rect 6214 39058 6230 39122
rect 6294 39058 6299 39122
rect 5105 39041 6299 39058
rect 5105 38977 5110 39041
rect 5174 38977 5190 39041
rect 5254 38977 5270 39041
rect 5334 38977 5350 39041
rect 5414 38977 5430 39041
rect 5494 38977 5510 39041
rect 5574 38977 5590 39041
rect 5654 38977 5670 39041
rect 5734 38977 5750 39041
rect 5814 38977 5830 39041
rect 5894 38977 5910 39041
rect 5974 38977 5990 39041
rect 6054 38977 6070 39041
rect 6134 38977 6150 39041
rect 6214 38977 6230 39041
rect 6294 38977 6299 39041
rect 5105 38960 6299 38977
rect 5105 38896 5110 38960
rect 5174 38896 5190 38960
rect 5254 38896 5270 38960
rect 5334 38896 5350 38960
rect 5414 38896 5430 38960
rect 5494 38896 5510 38960
rect 5574 38896 5590 38960
rect 5654 38896 5670 38960
rect 5734 38896 5750 38960
rect 5814 38896 5830 38960
rect 5894 38896 5910 38960
rect 5974 38896 5990 38960
rect 6054 38896 6070 38960
rect 6134 38896 6150 38960
rect 6214 38896 6230 38960
rect 6294 38896 6299 38960
rect 5105 38879 6299 38896
rect 5105 38815 5110 38879
rect 5174 38815 5190 38879
rect 5254 38815 5270 38879
rect 5334 38815 5350 38879
rect 5414 38815 5430 38879
rect 5494 38815 5510 38879
rect 5574 38815 5590 38879
rect 5654 38815 5670 38879
rect 5734 38815 5750 38879
rect 5814 38815 5830 38879
rect 5894 38815 5910 38879
rect 5974 38815 5990 38879
rect 6054 38815 6070 38879
rect 6134 38815 6150 38879
rect 6214 38815 6230 38879
rect 6294 38815 6299 38879
rect 5105 38798 6299 38815
rect 5105 38734 5110 38798
rect 5174 38734 5190 38798
rect 5254 38734 5270 38798
rect 5334 38734 5350 38798
rect 5414 38734 5430 38798
rect 5494 38734 5510 38798
rect 5574 38734 5590 38798
rect 5654 38734 5670 38798
rect 5734 38734 5750 38798
rect 5814 38734 5830 38798
rect 5894 38734 5910 38798
rect 5974 38734 5990 38798
rect 6054 38734 6070 38798
rect 6134 38734 6150 38798
rect 6214 38734 6230 38798
rect 6294 38734 6299 38798
rect 5105 38717 6299 38734
rect 5105 38653 5110 38717
rect 5174 38653 5190 38717
rect 5254 38653 5270 38717
rect 5334 38653 5350 38717
rect 5414 38653 5430 38717
rect 5494 38653 5510 38717
rect 5574 38653 5590 38717
rect 5654 38653 5670 38717
rect 5734 38653 5750 38717
rect 5814 38653 5830 38717
rect 5894 38653 5910 38717
rect 5974 38653 5990 38717
rect 6054 38653 6070 38717
rect 6134 38653 6150 38717
rect 6214 38653 6230 38717
rect 6294 38653 6299 38717
rect 5105 38636 6299 38653
rect 5105 38572 5110 38636
rect 5174 38572 5190 38636
rect 5254 38572 5270 38636
rect 5334 38572 5350 38636
rect 5414 38572 5430 38636
rect 5494 38572 5510 38636
rect 5574 38572 5590 38636
rect 5654 38572 5670 38636
rect 5734 38572 5750 38636
rect 5814 38572 5830 38636
rect 5894 38572 5910 38636
rect 5974 38572 5990 38636
rect 6054 38572 6070 38636
rect 6134 38572 6150 38636
rect 6214 38572 6230 38636
rect 6294 38572 6299 38636
rect 5105 38555 6299 38572
rect 5105 38491 5110 38555
rect 5174 38491 5190 38555
rect 5254 38491 5270 38555
rect 5334 38491 5350 38555
rect 5414 38491 5430 38555
rect 5494 38491 5510 38555
rect 5574 38491 5590 38555
rect 5654 38491 5670 38555
rect 5734 38491 5750 38555
rect 5814 38491 5830 38555
rect 5894 38491 5910 38555
rect 5974 38491 5990 38555
rect 6054 38491 6070 38555
rect 6134 38491 6150 38555
rect 6214 38491 6230 38555
rect 6294 38491 6299 38555
rect 5105 38474 6299 38491
rect 5105 38410 5110 38474
rect 5174 38410 5190 38474
rect 5254 38410 5270 38474
rect 5334 38410 5350 38474
rect 5414 38410 5430 38474
rect 5494 38410 5510 38474
rect 5574 38410 5590 38474
rect 5654 38410 5670 38474
rect 5734 38410 5750 38474
rect 5814 38410 5830 38474
rect 5894 38410 5910 38474
rect 5974 38410 5990 38474
rect 6054 38410 6070 38474
rect 6134 38410 6150 38474
rect 6214 38410 6230 38474
rect 6294 38410 6299 38474
rect 5105 38393 6299 38410
rect 5105 38329 5110 38393
rect 5174 38329 5190 38393
rect 5254 38329 5270 38393
rect 5334 38329 5350 38393
rect 5414 38329 5430 38393
rect 5494 38329 5510 38393
rect 5574 38329 5590 38393
rect 5654 38329 5670 38393
rect 5734 38329 5750 38393
rect 5814 38329 5830 38393
rect 5894 38329 5910 38393
rect 5974 38329 5990 38393
rect 6054 38329 6070 38393
rect 6134 38329 6150 38393
rect 6214 38329 6230 38393
rect 6294 38329 6299 38393
rect 5105 38312 6299 38329
rect 5105 38248 5110 38312
rect 5174 38248 5190 38312
rect 5254 38248 5270 38312
rect 5334 38248 5350 38312
rect 5414 38248 5430 38312
rect 5494 38248 5510 38312
rect 5574 38248 5590 38312
rect 5654 38248 5670 38312
rect 5734 38248 5750 38312
rect 5814 38248 5830 38312
rect 5894 38248 5910 38312
rect 5974 38248 5990 38312
rect 6054 38248 6070 38312
rect 6134 38248 6150 38312
rect 6214 38248 6230 38312
rect 6294 38248 6299 38312
rect 5105 38231 6299 38248
rect 5105 38167 5110 38231
rect 5174 38167 5190 38231
rect 5254 38167 5270 38231
rect 5334 38167 5350 38231
rect 5414 38167 5430 38231
rect 5494 38167 5510 38231
rect 5574 38167 5590 38231
rect 5654 38167 5670 38231
rect 5734 38167 5750 38231
rect 5814 38167 5830 38231
rect 5894 38167 5910 38231
rect 5974 38167 5990 38231
rect 6054 38167 6070 38231
rect 6134 38167 6150 38231
rect 6214 38167 6230 38231
rect 6294 38167 6299 38231
rect 5105 38150 6299 38167
rect 5105 38086 5110 38150
rect 5174 38086 5190 38150
rect 5254 38086 5270 38150
rect 5334 38086 5350 38150
rect 5414 38086 5430 38150
rect 5494 38086 5510 38150
rect 5574 38086 5590 38150
rect 5654 38086 5670 38150
rect 5734 38086 5750 38150
rect 5814 38086 5830 38150
rect 5894 38086 5910 38150
rect 5974 38086 5990 38150
rect 6054 38086 6070 38150
rect 6134 38086 6150 38150
rect 6214 38086 6230 38150
rect 6294 38086 6299 38150
rect 5105 38069 6299 38086
rect 5105 38005 5110 38069
rect 5174 38005 5190 38069
rect 5254 38005 5270 38069
rect 5334 38005 5350 38069
rect 5414 38005 5430 38069
rect 5494 38005 5510 38069
rect 5574 38005 5590 38069
rect 5654 38005 5670 38069
rect 5734 38005 5750 38069
rect 5814 38005 5830 38069
rect 5894 38005 5910 38069
rect 5974 38005 5990 38069
rect 6054 38005 6070 38069
rect 6134 38005 6150 38069
rect 6214 38005 6230 38069
rect 6294 38005 6299 38069
rect 5105 37988 6299 38005
rect 5105 37924 5110 37988
rect 5174 37924 5190 37988
rect 5254 37924 5270 37988
rect 5334 37924 5350 37988
rect 5414 37924 5430 37988
rect 5494 37924 5510 37988
rect 5574 37924 5590 37988
rect 5654 37924 5670 37988
rect 5734 37924 5750 37988
rect 5814 37924 5830 37988
rect 5894 37924 5910 37988
rect 5974 37924 5990 37988
rect 6054 37924 6070 37988
rect 6134 37924 6150 37988
rect 6214 37924 6230 37988
rect 6294 37924 6299 37988
rect 5105 37907 6299 37924
rect 5105 37843 5110 37907
rect 5174 37843 5190 37907
rect 5254 37843 5270 37907
rect 5334 37843 5350 37907
rect 5414 37843 5430 37907
rect 5494 37843 5510 37907
rect 5574 37843 5590 37907
rect 5654 37843 5670 37907
rect 5734 37843 5750 37907
rect 5814 37843 5830 37907
rect 5894 37843 5910 37907
rect 5974 37843 5990 37907
rect 6054 37843 6070 37907
rect 6134 37843 6150 37907
rect 6214 37843 6230 37907
rect 6294 37843 6299 37907
rect 5105 37826 6299 37843
rect 5105 37762 5110 37826
rect 5174 37762 5190 37826
rect 5254 37762 5270 37826
rect 5334 37762 5350 37826
rect 5414 37762 5430 37826
rect 5494 37762 5510 37826
rect 5574 37762 5590 37826
rect 5654 37762 5670 37826
rect 5734 37762 5750 37826
rect 5814 37762 5830 37826
rect 5894 37762 5910 37826
rect 5974 37762 5990 37826
rect 6054 37762 6070 37826
rect 6134 37762 6150 37826
rect 6214 37762 6230 37826
rect 6294 37762 6299 37826
rect 5105 37745 6299 37762
rect 5105 37681 5110 37745
rect 5174 37681 5190 37745
rect 5254 37681 5270 37745
rect 5334 37681 5350 37745
rect 5414 37681 5430 37745
rect 5494 37681 5510 37745
rect 5574 37681 5590 37745
rect 5654 37681 5670 37745
rect 5734 37681 5750 37745
rect 5814 37681 5830 37745
rect 5894 37681 5910 37745
rect 5974 37681 5990 37745
rect 6054 37681 6070 37745
rect 6134 37681 6150 37745
rect 6214 37681 6230 37745
rect 6294 37681 6299 37745
rect 5105 37664 6299 37681
rect 5105 37600 5110 37664
rect 5174 37600 5190 37664
rect 5254 37600 5270 37664
rect 5334 37600 5350 37664
rect 5414 37600 5430 37664
rect 5494 37600 5510 37664
rect 5574 37600 5590 37664
rect 5654 37600 5670 37664
rect 5734 37600 5750 37664
rect 5814 37600 5830 37664
rect 5894 37600 5910 37664
rect 5974 37600 5990 37664
rect 6054 37600 6070 37664
rect 6134 37600 6150 37664
rect 6214 37600 6230 37664
rect 6294 37600 6299 37664
rect 5105 37583 6299 37600
rect 5105 37519 5110 37583
rect 5174 37519 5190 37583
rect 5254 37519 5270 37583
rect 5334 37519 5350 37583
rect 5414 37519 5430 37583
rect 5494 37519 5510 37583
rect 5574 37519 5590 37583
rect 5654 37519 5670 37583
rect 5734 37519 5750 37583
rect 5814 37519 5830 37583
rect 5894 37519 5910 37583
rect 5974 37519 5990 37583
rect 6054 37519 6070 37583
rect 6134 37519 6150 37583
rect 6214 37519 6230 37583
rect 6294 37519 6299 37583
rect 5105 37502 6299 37519
rect 5105 37438 5110 37502
rect 5174 37438 5190 37502
rect 5254 37438 5270 37502
rect 5334 37438 5350 37502
rect 5414 37438 5430 37502
rect 5494 37438 5510 37502
rect 5574 37438 5590 37502
rect 5654 37438 5670 37502
rect 5734 37438 5750 37502
rect 5814 37438 5830 37502
rect 5894 37438 5910 37502
rect 5974 37438 5990 37502
rect 6054 37438 6070 37502
rect 6134 37438 6150 37502
rect 6214 37438 6230 37502
rect 6294 37438 6299 37502
rect 5105 37421 6299 37438
rect 5105 37357 5110 37421
rect 5174 37357 5190 37421
rect 5254 37357 5270 37421
rect 5334 37357 5350 37421
rect 5414 37357 5430 37421
rect 5494 37357 5510 37421
rect 5574 37357 5590 37421
rect 5654 37357 5670 37421
rect 5734 37357 5750 37421
rect 5814 37357 5830 37421
rect 5894 37357 5910 37421
rect 5974 37357 5990 37421
rect 6054 37357 6070 37421
rect 6134 37357 6150 37421
rect 6214 37357 6230 37421
rect 6294 37357 6299 37421
rect 5105 37340 6299 37357
rect 5105 37276 5110 37340
rect 5174 37276 5190 37340
rect 5254 37276 5270 37340
rect 5334 37276 5350 37340
rect 5414 37276 5430 37340
rect 5494 37276 5510 37340
rect 5574 37276 5590 37340
rect 5654 37276 5670 37340
rect 5734 37276 5750 37340
rect 5814 37276 5830 37340
rect 5894 37276 5910 37340
rect 5974 37276 5990 37340
rect 6054 37276 6070 37340
rect 6134 37276 6150 37340
rect 6214 37276 6230 37340
rect 6294 37276 6299 37340
rect 5105 37259 6299 37276
rect 5105 37195 5110 37259
rect 5174 37195 5190 37259
rect 5254 37195 5270 37259
rect 5334 37195 5350 37259
rect 5414 37195 5430 37259
rect 5494 37195 5510 37259
rect 5574 37195 5590 37259
rect 5654 37195 5670 37259
rect 5734 37195 5750 37259
rect 5814 37195 5830 37259
rect 5894 37195 5910 37259
rect 5974 37195 5990 37259
rect 6054 37195 6070 37259
rect 6134 37195 6150 37259
rect 6214 37195 6230 37259
rect 6294 37195 6299 37259
rect 5105 37178 6299 37195
rect 5105 37114 5110 37178
rect 5174 37114 5190 37178
rect 5254 37114 5270 37178
rect 5334 37114 5350 37178
rect 5414 37114 5430 37178
rect 5494 37114 5510 37178
rect 5574 37114 5590 37178
rect 5654 37114 5670 37178
rect 5734 37114 5750 37178
rect 5814 37114 5830 37178
rect 5894 37114 5910 37178
rect 5974 37114 5990 37178
rect 6054 37114 6070 37178
rect 6134 37114 6150 37178
rect 6214 37114 6230 37178
rect 6294 37114 6299 37178
rect 5105 37097 6299 37114
rect 5105 37033 5110 37097
rect 5174 37033 5190 37097
rect 5254 37033 5270 37097
rect 5334 37033 5350 37097
rect 5414 37033 5430 37097
rect 5494 37033 5510 37097
rect 5574 37033 5590 37097
rect 5654 37033 5670 37097
rect 5734 37033 5750 37097
rect 5814 37033 5830 37097
rect 5894 37033 5910 37097
rect 5974 37033 5990 37097
rect 6054 37033 6070 37097
rect 6134 37033 6150 37097
rect 6214 37033 6230 37097
rect 6294 37033 6299 37097
rect 5105 37016 6299 37033
rect 5105 36952 5110 37016
rect 5174 36952 5190 37016
rect 5254 36952 5270 37016
rect 5334 36952 5350 37016
rect 5414 36952 5430 37016
rect 5494 36952 5510 37016
rect 5574 36952 5590 37016
rect 5654 36952 5670 37016
rect 5734 36952 5750 37016
rect 5814 36952 5830 37016
rect 5894 36952 5910 37016
rect 5974 36952 5990 37016
rect 6054 36952 6070 37016
rect 6134 36952 6150 37016
rect 6214 36952 6230 37016
rect 6294 36952 6299 37016
rect 5105 36935 6299 36952
rect 5105 36871 5110 36935
rect 5174 36871 5190 36935
rect 5254 36871 5270 36935
rect 5334 36871 5350 36935
rect 5414 36871 5430 36935
rect 5494 36871 5510 36935
rect 5574 36871 5590 36935
rect 5654 36871 5670 36935
rect 5734 36871 5750 36935
rect 5814 36871 5830 36935
rect 5894 36871 5910 36935
rect 5974 36871 5990 36935
rect 6054 36871 6070 36935
rect 6134 36871 6150 36935
rect 6214 36871 6230 36935
rect 6294 36871 6299 36935
rect 5105 36854 6299 36871
rect 5105 36790 5110 36854
rect 5174 36790 5190 36854
rect 5254 36790 5270 36854
rect 5334 36790 5350 36854
rect 5414 36790 5430 36854
rect 5494 36790 5510 36854
rect 5574 36790 5590 36854
rect 5654 36790 5670 36854
rect 5734 36790 5750 36854
rect 5814 36790 5830 36854
rect 5894 36790 5910 36854
rect 5974 36790 5990 36854
rect 6054 36790 6070 36854
rect 6134 36790 6150 36854
rect 6214 36790 6230 36854
rect 6294 36790 6299 36854
rect 5105 36773 6299 36790
rect 5105 36709 5110 36773
rect 5174 36709 5190 36773
rect 5254 36709 5270 36773
rect 5334 36709 5350 36773
rect 5414 36709 5430 36773
rect 5494 36709 5510 36773
rect 5574 36709 5590 36773
rect 5654 36709 5670 36773
rect 5734 36709 5750 36773
rect 5814 36709 5830 36773
rect 5894 36709 5910 36773
rect 5974 36709 5990 36773
rect 6054 36709 6070 36773
rect 6134 36709 6150 36773
rect 6214 36709 6230 36773
rect 6294 36709 6299 36773
rect 5105 36692 6299 36709
rect 5105 36628 5110 36692
rect 5174 36628 5190 36692
rect 5254 36628 5270 36692
rect 5334 36628 5350 36692
rect 5414 36628 5430 36692
rect 5494 36628 5510 36692
rect 5574 36628 5590 36692
rect 5654 36628 5670 36692
rect 5734 36628 5750 36692
rect 5814 36628 5830 36692
rect 5894 36628 5910 36692
rect 5974 36628 5990 36692
rect 6054 36628 6070 36692
rect 6134 36628 6150 36692
rect 6214 36628 6230 36692
rect 6294 36628 6299 36692
rect 5105 36611 6299 36628
rect 5105 36547 5110 36611
rect 5174 36547 5190 36611
rect 5254 36547 5270 36611
rect 5334 36547 5350 36611
rect 5414 36547 5430 36611
rect 5494 36547 5510 36611
rect 5574 36547 5590 36611
rect 5654 36547 5670 36611
rect 5734 36547 5750 36611
rect 5814 36547 5830 36611
rect 5894 36547 5910 36611
rect 5974 36547 5990 36611
rect 6054 36547 6070 36611
rect 6134 36547 6150 36611
rect 6214 36547 6230 36611
rect 6294 36547 6299 36611
rect 5105 36530 6299 36547
rect 5105 36466 5110 36530
rect 5174 36466 5190 36530
rect 5254 36466 5270 36530
rect 5334 36466 5350 36530
rect 5414 36466 5430 36530
rect 5494 36466 5510 36530
rect 5574 36466 5590 36530
rect 5654 36466 5670 36530
rect 5734 36466 5750 36530
rect 5814 36466 5830 36530
rect 5894 36466 5910 36530
rect 5974 36466 5990 36530
rect 6054 36466 6070 36530
rect 6134 36466 6150 36530
rect 6214 36466 6230 36530
rect 6294 36466 6299 36530
rect 5105 36449 6299 36466
rect 5105 36385 5110 36449
rect 5174 36385 5190 36449
rect 5254 36385 5270 36449
rect 5334 36385 5350 36449
rect 5414 36385 5430 36449
rect 5494 36385 5510 36449
rect 5574 36385 5590 36449
rect 5654 36385 5670 36449
rect 5734 36385 5750 36449
rect 5814 36385 5830 36449
rect 5894 36385 5910 36449
rect 5974 36385 5990 36449
rect 6054 36385 6070 36449
rect 6134 36385 6150 36449
rect 6214 36385 6230 36449
rect 6294 36385 6299 36449
rect 5105 36368 6299 36385
rect 5105 36304 5110 36368
rect 5174 36304 5190 36368
rect 5254 36304 5270 36368
rect 5334 36304 5350 36368
rect 5414 36304 5430 36368
rect 5494 36304 5510 36368
rect 5574 36304 5590 36368
rect 5654 36304 5670 36368
rect 5734 36304 5750 36368
rect 5814 36304 5830 36368
rect 5894 36304 5910 36368
rect 5974 36304 5990 36368
rect 6054 36304 6070 36368
rect 6134 36304 6150 36368
rect 6214 36304 6230 36368
rect 6294 36304 6299 36368
rect 5105 36287 6299 36304
rect 5105 36223 5110 36287
rect 5174 36223 5190 36287
rect 5254 36223 5270 36287
rect 5334 36223 5350 36287
rect 5414 36223 5430 36287
rect 5494 36223 5510 36287
rect 5574 36223 5590 36287
rect 5654 36223 5670 36287
rect 5734 36223 5750 36287
rect 5814 36223 5830 36287
rect 5894 36223 5910 36287
rect 5974 36223 5990 36287
rect 6054 36223 6070 36287
rect 6134 36223 6150 36287
rect 6214 36223 6230 36287
rect 6294 36223 6299 36287
rect 5105 36206 6299 36223
rect 5105 36142 5110 36206
rect 5174 36142 5190 36206
rect 5254 36142 5270 36206
rect 5334 36142 5350 36206
rect 5414 36142 5430 36206
rect 5494 36142 5510 36206
rect 5574 36142 5590 36206
rect 5654 36142 5670 36206
rect 5734 36142 5750 36206
rect 5814 36142 5830 36206
rect 5894 36142 5910 36206
rect 5974 36142 5990 36206
rect 6054 36142 6070 36206
rect 6134 36142 6150 36206
rect 6214 36142 6230 36206
rect 6294 36142 6299 36206
rect 5105 36124 6299 36142
rect 5105 36060 5110 36124
rect 5174 36060 5190 36124
rect 5254 36060 5270 36124
rect 5334 36060 5350 36124
rect 5414 36060 5430 36124
rect 5494 36060 5510 36124
rect 5574 36060 5590 36124
rect 5654 36060 5670 36124
rect 5734 36060 5750 36124
rect 5814 36060 5830 36124
rect 5894 36060 5910 36124
rect 5974 36060 5990 36124
rect 6054 36060 6070 36124
rect 6134 36060 6150 36124
rect 6214 36060 6230 36124
rect 6294 36060 6299 36124
rect 5105 36042 6299 36060
rect 5105 35978 5110 36042
rect 5174 35978 5190 36042
rect 5254 35978 5270 36042
rect 5334 35978 5350 36042
rect 5414 35978 5430 36042
rect 5494 35978 5510 36042
rect 5574 35978 5590 36042
rect 5654 35978 5670 36042
rect 5734 35978 5750 36042
rect 5814 35978 5830 36042
rect 5894 35978 5910 36042
rect 5974 35978 5990 36042
rect 6054 35978 6070 36042
rect 6134 35978 6150 36042
rect 6214 35978 6230 36042
rect 6294 35978 6299 36042
rect 5105 35960 6299 35978
rect 5105 35896 5110 35960
rect 5174 35896 5190 35960
rect 5254 35896 5270 35960
rect 5334 35896 5350 35960
rect 5414 35896 5430 35960
rect 5494 35896 5510 35960
rect 5574 35896 5590 35960
rect 5654 35896 5670 35960
rect 5734 35896 5750 35960
rect 5814 35896 5830 35960
rect 5894 35896 5910 35960
rect 5974 35896 5990 35960
rect 6054 35896 6070 35960
rect 6134 35896 6150 35960
rect 6214 35896 6230 35960
rect 6294 35896 6299 35960
rect 5105 35878 6299 35896
rect 5105 35814 5110 35878
rect 5174 35814 5190 35878
rect 5254 35814 5270 35878
rect 5334 35814 5350 35878
rect 5414 35814 5430 35878
rect 5494 35814 5510 35878
rect 5574 35814 5590 35878
rect 5654 35814 5670 35878
rect 5734 35814 5750 35878
rect 5814 35814 5830 35878
rect 5894 35814 5910 35878
rect 5974 35814 5990 35878
rect 6054 35814 6070 35878
rect 6134 35814 6150 35878
rect 6214 35814 6230 35878
rect 6294 35814 6299 35878
rect 5105 35796 6299 35814
rect 5105 35732 5110 35796
rect 5174 35732 5190 35796
rect 5254 35732 5270 35796
rect 5334 35732 5350 35796
rect 5414 35732 5430 35796
rect 5494 35732 5510 35796
rect 5574 35732 5590 35796
rect 5654 35732 5670 35796
rect 5734 35732 5750 35796
rect 5814 35732 5830 35796
rect 5894 35732 5910 35796
rect 5974 35732 5990 35796
rect 6054 35732 6070 35796
rect 6134 35732 6150 35796
rect 6214 35732 6230 35796
rect 6294 35732 6299 35796
rect 5105 35714 6299 35732
rect 5105 35650 5110 35714
rect 5174 35650 5190 35714
rect 5254 35650 5270 35714
rect 5334 35650 5350 35714
rect 5414 35650 5430 35714
rect 5494 35650 5510 35714
rect 5574 35650 5590 35714
rect 5654 35650 5670 35714
rect 5734 35650 5750 35714
rect 5814 35650 5830 35714
rect 5894 35650 5910 35714
rect 5974 35650 5990 35714
rect 6054 35650 6070 35714
rect 6134 35650 6150 35714
rect 6214 35650 6230 35714
rect 6294 35650 6299 35714
rect 5105 35632 6299 35650
rect 5105 35568 5110 35632
rect 5174 35568 5190 35632
rect 5254 35568 5270 35632
rect 5334 35568 5350 35632
rect 5414 35568 5430 35632
rect 5494 35568 5510 35632
rect 5574 35568 5590 35632
rect 5654 35568 5670 35632
rect 5734 35568 5750 35632
rect 5814 35568 5830 35632
rect 5894 35568 5910 35632
rect 5974 35568 5990 35632
rect 6054 35568 6070 35632
rect 6134 35568 6150 35632
rect 6214 35568 6230 35632
rect 6294 35568 6299 35632
rect 5105 35550 6299 35568
rect 5105 35486 5110 35550
rect 5174 35486 5190 35550
rect 5254 35486 5270 35550
rect 5334 35486 5350 35550
rect 5414 35486 5430 35550
rect 5494 35486 5510 35550
rect 5574 35486 5590 35550
rect 5654 35486 5670 35550
rect 5734 35486 5750 35550
rect 5814 35486 5830 35550
rect 5894 35486 5910 35550
rect 5974 35486 5990 35550
rect 6054 35486 6070 35550
rect 6134 35486 6150 35550
rect 6214 35486 6230 35550
rect 6294 35486 6299 35550
rect 5105 35468 6299 35486
rect 5105 35404 5110 35468
rect 5174 35404 5190 35468
rect 5254 35404 5270 35468
rect 5334 35404 5350 35468
rect 5414 35404 5430 35468
rect 5494 35404 5510 35468
rect 5574 35404 5590 35468
rect 5654 35404 5670 35468
rect 5734 35404 5750 35468
rect 5814 35404 5830 35468
rect 5894 35404 5910 35468
rect 5974 35404 5990 35468
rect 6054 35404 6070 35468
rect 6134 35404 6150 35468
rect 6214 35404 6230 35468
rect 6294 35404 6299 35468
rect 5105 35386 6299 35404
rect 5105 35322 5110 35386
rect 5174 35322 5190 35386
rect 5254 35322 5270 35386
rect 5334 35322 5350 35386
rect 5414 35322 5430 35386
rect 5494 35322 5510 35386
rect 5574 35322 5590 35386
rect 5654 35322 5670 35386
rect 5734 35322 5750 35386
rect 5814 35322 5830 35386
rect 5894 35322 5910 35386
rect 5974 35322 5990 35386
rect 6054 35322 6070 35386
rect 6134 35322 6150 35386
rect 6214 35322 6230 35386
rect 6294 35322 6299 35386
rect 5105 35304 6299 35322
rect 5105 35240 5110 35304
rect 5174 35240 5190 35304
rect 5254 35240 5270 35304
rect 5334 35240 5350 35304
rect 5414 35240 5430 35304
rect 5494 35240 5510 35304
rect 5574 35240 5590 35304
rect 5654 35240 5670 35304
rect 5734 35240 5750 35304
rect 5814 35240 5830 35304
rect 5894 35240 5910 35304
rect 5974 35240 5990 35304
rect 6054 35240 6070 35304
rect 6134 35240 6150 35304
rect 6214 35240 6230 35304
rect 6294 35240 6299 35304
rect 5105 35222 6299 35240
rect 5105 35158 5110 35222
rect 5174 35158 5190 35222
rect 5254 35158 5270 35222
rect 5334 35158 5350 35222
rect 5414 35158 5430 35222
rect 5494 35158 5510 35222
rect 5574 35158 5590 35222
rect 5654 35158 5670 35222
rect 5734 35158 5750 35222
rect 5814 35158 5830 35222
rect 5894 35158 5910 35222
rect 5974 35158 5990 35222
rect 6054 35158 6070 35222
rect 6134 35158 6150 35222
rect 6214 35158 6230 35222
rect 6294 35158 6299 35222
rect 5105 35157 6299 35158
rect 6602 39365 7796 39366
rect 6602 39301 6607 39365
rect 6671 39301 6687 39365
rect 6751 39301 6767 39365
rect 6831 39301 6847 39365
rect 6911 39301 6927 39365
rect 6991 39301 7007 39365
rect 7071 39301 7087 39365
rect 7151 39301 7167 39365
rect 7231 39301 7247 39365
rect 7311 39301 7327 39365
rect 7391 39301 7407 39365
rect 7471 39301 7487 39365
rect 7551 39301 7567 39365
rect 7631 39301 7647 39365
rect 7711 39301 7727 39365
rect 7791 39301 7796 39365
rect 6602 39284 7796 39301
rect 6602 39220 6607 39284
rect 6671 39220 6687 39284
rect 6751 39220 6767 39284
rect 6831 39220 6847 39284
rect 6911 39220 6927 39284
rect 6991 39220 7007 39284
rect 7071 39220 7087 39284
rect 7151 39220 7167 39284
rect 7231 39220 7247 39284
rect 7311 39220 7327 39284
rect 7391 39220 7407 39284
rect 7471 39220 7487 39284
rect 7551 39220 7567 39284
rect 7631 39220 7647 39284
rect 7711 39220 7727 39284
rect 7791 39220 7796 39284
rect 6602 39203 7796 39220
rect 6602 39139 6607 39203
rect 6671 39139 6687 39203
rect 6751 39139 6767 39203
rect 6831 39139 6847 39203
rect 6911 39139 6927 39203
rect 6991 39139 7007 39203
rect 7071 39139 7087 39203
rect 7151 39139 7167 39203
rect 7231 39139 7247 39203
rect 7311 39139 7327 39203
rect 7391 39139 7407 39203
rect 7471 39139 7487 39203
rect 7551 39139 7567 39203
rect 7631 39139 7647 39203
rect 7711 39139 7727 39203
rect 7791 39139 7796 39203
rect 6602 39122 7796 39139
rect 6602 39058 6607 39122
rect 6671 39058 6687 39122
rect 6751 39058 6767 39122
rect 6831 39058 6847 39122
rect 6911 39058 6927 39122
rect 6991 39058 7007 39122
rect 7071 39058 7087 39122
rect 7151 39058 7167 39122
rect 7231 39058 7247 39122
rect 7311 39058 7327 39122
rect 7391 39058 7407 39122
rect 7471 39058 7487 39122
rect 7551 39058 7567 39122
rect 7631 39058 7647 39122
rect 7711 39058 7727 39122
rect 7791 39058 7796 39122
rect 6602 39041 7796 39058
rect 6602 38977 6607 39041
rect 6671 38977 6687 39041
rect 6751 38977 6767 39041
rect 6831 38977 6847 39041
rect 6911 38977 6927 39041
rect 6991 38977 7007 39041
rect 7071 38977 7087 39041
rect 7151 38977 7167 39041
rect 7231 38977 7247 39041
rect 7311 38977 7327 39041
rect 7391 38977 7407 39041
rect 7471 38977 7487 39041
rect 7551 38977 7567 39041
rect 7631 38977 7647 39041
rect 7711 38977 7727 39041
rect 7791 38977 7796 39041
rect 6602 38960 7796 38977
rect 6602 38896 6607 38960
rect 6671 38896 6687 38960
rect 6751 38896 6767 38960
rect 6831 38896 6847 38960
rect 6911 38896 6927 38960
rect 6991 38896 7007 38960
rect 7071 38896 7087 38960
rect 7151 38896 7167 38960
rect 7231 38896 7247 38960
rect 7311 38896 7327 38960
rect 7391 38896 7407 38960
rect 7471 38896 7487 38960
rect 7551 38896 7567 38960
rect 7631 38896 7647 38960
rect 7711 38896 7727 38960
rect 7791 38896 7796 38960
rect 6602 38879 7796 38896
rect 6602 38815 6607 38879
rect 6671 38815 6687 38879
rect 6751 38815 6767 38879
rect 6831 38815 6847 38879
rect 6911 38815 6927 38879
rect 6991 38815 7007 38879
rect 7071 38815 7087 38879
rect 7151 38815 7167 38879
rect 7231 38815 7247 38879
rect 7311 38815 7327 38879
rect 7391 38815 7407 38879
rect 7471 38815 7487 38879
rect 7551 38815 7567 38879
rect 7631 38815 7647 38879
rect 7711 38815 7727 38879
rect 7791 38815 7796 38879
rect 6602 38798 7796 38815
rect 6602 38734 6607 38798
rect 6671 38734 6687 38798
rect 6751 38734 6767 38798
rect 6831 38734 6847 38798
rect 6911 38734 6927 38798
rect 6991 38734 7007 38798
rect 7071 38734 7087 38798
rect 7151 38734 7167 38798
rect 7231 38734 7247 38798
rect 7311 38734 7327 38798
rect 7391 38734 7407 38798
rect 7471 38734 7487 38798
rect 7551 38734 7567 38798
rect 7631 38734 7647 38798
rect 7711 38734 7727 38798
rect 7791 38734 7796 38798
rect 6602 38717 7796 38734
rect 6602 38653 6607 38717
rect 6671 38653 6687 38717
rect 6751 38653 6767 38717
rect 6831 38653 6847 38717
rect 6911 38653 6927 38717
rect 6991 38653 7007 38717
rect 7071 38653 7087 38717
rect 7151 38653 7167 38717
rect 7231 38653 7247 38717
rect 7311 38653 7327 38717
rect 7391 38653 7407 38717
rect 7471 38653 7487 38717
rect 7551 38653 7567 38717
rect 7631 38653 7647 38717
rect 7711 38653 7727 38717
rect 7791 38653 7796 38717
rect 6602 38636 7796 38653
rect 6602 38572 6607 38636
rect 6671 38572 6687 38636
rect 6751 38572 6767 38636
rect 6831 38572 6847 38636
rect 6911 38572 6927 38636
rect 6991 38572 7007 38636
rect 7071 38572 7087 38636
rect 7151 38572 7167 38636
rect 7231 38572 7247 38636
rect 7311 38572 7327 38636
rect 7391 38572 7407 38636
rect 7471 38572 7487 38636
rect 7551 38572 7567 38636
rect 7631 38572 7647 38636
rect 7711 38572 7727 38636
rect 7791 38572 7796 38636
rect 6602 38555 7796 38572
rect 6602 38491 6607 38555
rect 6671 38491 6687 38555
rect 6751 38491 6767 38555
rect 6831 38491 6847 38555
rect 6911 38491 6927 38555
rect 6991 38491 7007 38555
rect 7071 38491 7087 38555
rect 7151 38491 7167 38555
rect 7231 38491 7247 38555
rect 7311 38491 7327 38555
rect 7391 38491 7407 38555
rect 7471 38491 7487 38555
rect 7551 38491 7567 38555
rect 7631 38491 7647 38555
rect 7711 38491 7727 38555
rect 7791 38491 7796 38555
rect 6602 38474 7796 38491
rect 6602 38410 6607 38474
rect 6671 38410 6687 38474
rect 6751 38410 6767 38474
rect 6831 38410 6847 38474
rect 6911 38410 6927 38474
rect 6991 38410 7007 38474
rect 7071 38410 7087 38474
rect 7151 38410 7167 38474
rect 7231 38410 7247 38474
rect 7311 38410 7327 38474
rect 7391 38410 7407 38474
rect 7471 38410 7487 38474
rect 7551 38410 7567 38474
rect 7631 38410 7647 38474
rect 7711 38410 7727 38474
rect 7791 38410 7796 38474
rect 6602 38393 7796 38410
rect 6602 38329 6607 38393
rect 6671 38329 6687 38393
rect 6751 38329 6767 38393
rect 6831 38329 6847 38393
rect 6911 38329 6927 38393
rect 6991 38329 7007 38393
rect 7071 38329 7087 38393
rect 7151 38329 7167 38393
rect 7231 38329 7247 38393
rect 7311 38329 7327 38393
rect 7391 38329 7407 38393
rect 7471 38329 7487 38393
rect 7551 38329 7567 38393
rect 7631 38329 7647 38393
rect 7711 38329 7727 38393
rect 7791 38329 7796 38393
rect 6602 38312 7796 38329
rect 6602 38248 6607 38312
rect 6671 38248 6687 38312
rect 6751 38248 6767 38312
rect 6831 38248 6847 38312
rect 6911 38248 6927 38312
rect 6991 38248 7007 38312
rect 7071 38248 7087 38312
rect 7151 38248 7167 38312
rect 7231 38248 7247 38312
rect 7311 38248 7327 38312
rect 7391 38248 7407 38312
rect 7471 38248 7487 38312
rect 7551 38248 7567 38312
rect 7631 38248 7647 38312
rect 7711 38248 7727 38312
rect 7791 38248 7796 38312
rect 6602 38231 7796 38248
rect 6602 38167 6607 38231
rect 6671 38167 6687 38231
rect 6751 38167 6767 38231
rect 6831 38167 6847 38231
rect 6911 38167 6927 38231
rect 6991 38167 7007 38231
rect 7071 38167 7087 38231
rect 7151 38167 7167 38231
rect 7231 38167 7247 38231
rect 7311 38167 7327 38231
rect 7391 38167 7407 38231
rect 7471 38167 7487 38231
rect 7551 38167 7567 38231
rect 7631 38167 7647 38231
rect 7711 38167 7727 38231
rect 7791 38167 7796 38231
rect 6602 38150 7796 38167
rect 6602 38086 6607 38150
rect 6671 38086 6687 38150
rect 6751 38086 6767 38150
rect 6831 38086 6847 38150
rect 6911 38086 6927 38150
rect 6991 38086 7007 38150
rect 7071 38086 7087 38150
rect 7151 38086 7167 38150
rect 7231 38086 7247 38150
rect 7311 38086 7327 38150
rect 7391 38086 7407 38150
rect 7471 38086 7487 38150
rect 7551 38086 7567 38150
rect 7631 38086 7647 38150
rect 7711 38086 7727 38150
rect 7791 38086 7796 38150
rect 6602 38069 7796 38086
rect 6602 38005 6607 38069
rect 6671 38005 6687 38069
rect 6751 38005 6767 38069
rect 6831 38005 6847 38069
rect 6911 38005 6927 38069
rect 6991 38005 7007 38069
rect 7071 38005 7087 38069
rect 7151 38005 7167 38069
rect 7231 38005 7247 38069
rect 7311 38005 7327 38069
rect 7391 38005 7407 38069
rect 7471 38005 7487 38069
rect 7551 38005 7567 38069
rect 7631 38005 7647 38069
rect 7711 38005 7727 38069
rect 7791 38005 7796 38069
rect 6602 37988 7796 38005
rect 6602 37924 6607 37988
rect 6671 37924 6687 37988
rect 6751 37924 6767 37988
rect 6831 37924 6847 37988
rect 6911 37924 6927 37988
rect 6991 37924 7007 37988
rect 7071 37924 7087 37988
rect 7151 37924 7167 37988
rect 7231 37924 7247 37988
rect 7311 37924 7327 37988
rect 7391 37924 7407 37988
rect 7471 37924 7487 37988
rect 7551 37924 7567 37988
rect 7631 37924 7647 37988
rect 7711 37924 7727 37988
rect 7791 37924 7796 37988
rect 6602 37907 7796 37924
rect 6602 37843 6607 37907
rect 6671 37843 6687 37907
rect 6751 37843 6767 37907
rect 6831 37843 6847 37907
rect 6911 37843 6927 37907
rect 6991 37843 7007 37907
rect 7071 37843 7087 37907
rect 7151 37843 7167 37907
rect 7231 37843 7247 37907
rect 7311 37843 7327 37907
rect 7391 37843 7407 37907
rect 7471 37843 7487 37907
rect 7551 37843 7567 37907
rect 7631 37843 7647 37907
rect 7711 37843 7727 37907
rect 7791 37843 7796 37907
rect 6602 37826 7796 37843
rect 6602 37762 6607 37826
rect 6671 37762 6687 37826
rect 6751 37762 6767 37826
rect 6831 37762 6847 37826
rect 6911 37762 6927 37826
rect 6991 37762 7007 37826
rect 7071 37762 7087 37826
rect 7151 37762 7167 37826
rect 7231 37762 7247 37826
rect 7311 37762 7327 37826
rect 7391 37762 7407 37826
rect 7471 37762 7487 37826
rect 7551 37762 7567 37826
rect 7631 37762 7647 37826
rect 7711 37762 7727 37826
rect 7791 37762 7796 37826
rect 6602 37745 7796 37762
rect 6602 37681 6607 37745
rect 6671 37681 6687 37745
rect 6751 37681 6767 37745
rect 6831 37681 6847 37745
rect 6911 37681 6927 37745
rect 6991 37681 7007 37745
rect 7071 37681 7087 37745
rect 7151 37681 7167 37745
rect 7231 37681 7247 37745
rect 7311 37681 7327 37745
rect 7391 37681 7407 37745
rect 7471 37681 7487 37745
rect 7551 37681 7567 37745
rect 7631 37681 7647 37745
rect 7711 37681 7727 37745
rect 7791 37681 7796 37745
rect 6602 37664 7796 37681
rect 6602 37600 6607 37664
rect 6671 37600 6687 37664
rect 6751 37600 6767 37664
rect 6831 37600 6847 37664
rect 6911 37600 6927 37664
rect 6991 37600 7007 37664
rect 7071 37600 7087 37664
rect 7151 37600 7167 37664
rect 7231 37600 7247 37664
rect 7311 37600 7327 37664
rect 7391 37600 7407 37664
rect 7471 37600 7487 37664
rect 7551 37600 7567 37664
rect 7631 37600 7647 37664
rect 7711 37600 7727 37664
rect 7791 37600 7796 37664
rect 6602 37583 7796 37600
rect 6602 37519 6607 37583
rect 6671 37519 6687 37583
rect 6751 37519 6767 37583
rect 6831 37519 6847 37583
rect 6911 37519 6927 37583
rect 6991 37519 7007 37583
rect 7071 37519 7087 37583
rect 7151 37519 7167 37583
rect 7231 37519 7247 37583
rect 7311 37519 7327 37583
rect 7391 37519 7407 37583
rect 7471 37519 7487 37583
rect 7551 37519 7567 37583
rect 7631 37519 7647 37583
rect 7711 37519 7727 37583
rect 7791 37519 7796 37583
rect 6602 37502 7796 37519
rect 6602 37438 6607 37502
rect 6671 37438 6687 37502
rect 6751 37438 6767 37502
rect 6831 37438 6847 37502
rect 6911 37438 6927 37502
rect 6991 37438 7007 37502
rect 7071 37438 7087 37502
rect 7151 37438 7167 37502
rect 7231 37438 7247 37502
rect 7311 37438 7327 37502
rect 7391 37438 7407 37502
rect 7471 37438 7487 37502
rect 7551 37438 7567 37502
rect 7631 37438 7647 37502
rect 7711 37438 7727 37502
rect 7791 37438 7796 37502
rect 6602 37421 7796 37438
rect 6602 37357 6607 37421
rect 6671 37357 6687 37421
rect 6751 37357 6767 37421
rect 6831 37357 6847 37421
rect 6911 37357 6927 37421
rect 6991 37357 7007 37421
rect 7071 37357 7087 37421
rect 7151 37357 7167 37421
rect 7231 37357 7247 37421
rect 7311 37357 7327 37421
rect 7391 37357 7407 37421
rect 7471 37357 7487 37421
rect 7551 37357 7567 37421
rect 7631 37357 7647 37421
rect 7711 37357 7727 37421
rect 7791 37357 7796 37421
rect 6602 37340 7796 37357
rect 6602 37276 6607 37340
rect 6671 37276 6687 37340
rect 6751 37276 6767 37340
rect 6831 37276 6847 37340
rect 6911 37276 6927 37340
rect 6991 37276 7007 37340
rect 7071 37276 7087 37340
rect 7151 37276 7167 37340
rect 7231 37276 7247 37340
rect 7311 37276 7327 37340
rect 7391 37276 7407 37340
rect 7471 37276 7487 37340
rect 7551 37276 7567 37340
rect 7631 37276 7647 37340
rect 7711 37276 7727 37340
rect 7791 37276 7796 37340
rect 6602 37259 7796 37276
rect 6602 37195 6607 37259
rect 6671 37195 6687 37259
rect 6751 37195 6767 37259
rect 6831 37195 6847 37259
rect 6911 37195 6927 37259
rect 6991 37195 7007 37259
rect 7071 37195 7087 37259
rect 7151 37195 7167 37259
rect 7231 37195 7247 37259
rect 7311 37195 7327 37259
rect 7391 37195 7407 37259
rect 7471 37195 7487 37259
rect 7551 37195 7567 37259
rect 7631 37195 7647 37259
rect 7711 37195 7727 37259
rect 7791 37195 7796 37259
rect 6602 37178 7796 37195
rect 6602 37114 6607 37178
rect 6671 37114 6687 37178
rect 6751 37114 6767 37178
rect 6831 37114 6847 37178
rect 6911 37114 6927 37178
rect 6991 37114 7007 37178
rect 7071 37114 7087 37178
rect 7151 37114 7167 37178
rect 7231 37114 7247 37178
rect 7311 37114 7327 37178
rect 7391 37114 7407 37178
rect 7471 37114 7487 37178
rect 7551 37114 7567 37178
rect 7631 37114 7647 37178
rect 7711 37114 7727 37178
rect 7791 37114 7796 37178
rect 6602 37097 7796 37114
rect 6602 37033 6607 37097
rect 6671 37033 6687 37097
rect 6751 37033 6767 37097
rect 6831 37033 6847 37097
rect 6911 37033 6927 37097
rect 6991 37033 7007 37097
rect 7071 37033 7087 37097
rect 7151 37033 7167 37097
rect 7231 37033 7247 37097
rect 7311 37033 7327 37097
rect 7391 37033 7407 37097
rect 7471 37033 7487 37097
rect 7551 37033 7567 37097
rect 7631 37033 7647 37097
rect 7711 37033 7727 37097
rect 7791 37033 7796 37097
rect 6602 37016 7796 37033
rect 6602 36952 6607 37016
rect 6671 36952 6687 37016
rect 6751 36952 6767 37016
rect 6831 36952 6847 37016
rect 6911 36952 6927 37016
rect 6991 36952 7007 37016
rect 7071 36952 7087 37016
rect 7151 36952 7167 37016
rect 7231 36952 7247 37016
rect 7311 36952 7327 37016
rect 7391 36952 7407 37016
rect 7471 36952 7487 37016
rect 7551 36952 7567 37016
rect 7631 36952 7647 37016
rect 7711 36952 7727 37016
rect 7791 36952 7796 37016
rect 6602 36935 7796 36952
rect 6602 36871 6607 36935
rect 6671 36871 6687 36935
rect 6751 36871 6767 36935
rect 6831 36871 6847 36935
rect 6911 36871 6927 36935
rect 6991 36871 7007 36935
rect 7071 36871 7087 36935
rect 7151 36871 7167 36935
rect 7231 36871 7247 36935
rect 7311 36871 7327 36935
rect 7391 36871 7407 36935
rect 7471 36871 7487 36935
rect 7551 36871 7567 36935
rect 7631 36871 7647 36935
rect 7711 36871 7727 36935
rect 7791 36871 7796 36935
rect 6602 36854 7796 36871
rect 6602 36790 6607 36854
rect 6671 36790 6687 36854
rect 6751 36790 6767 36854
rect 6831 36790 6847 36854
rect 6911 36790 6927 36854
rect 6991 36790 7007 36854
rect 7071 36790 7087 36854
rect 7151 36790 7167 36854
rect 7231 36790 7247 36854
rect 7311 36790 7327 36854
rect 7391 36790 7407 36854
rect 7471 36790 7487 36854
rect 7551 36790 7567 36854
rect 7631 36790 7647 36854
rect 7711 36790 7727 36854
rect 7791 36790 7796 36854
rect 6602 36773 7796 36790
rect 6602 36709 6607 36773
rect 6671 36709 6687 36773
rect 6751 36709 6767 36773
rect 6831 36709 6847 36773
rect 6911 36709 6927 36773
rect 6991 36709 7007 36773
rect 7071 36709 7087 36773
rect 7151 36709 7167 36773
rect 7231 36709 7247 36773
rect 7311 36709 7327 36773
rect 7391 36709 7407 36773
rect 7471 36709 7487 36773
rect 7551 36709 7567 36773
rect 7631 36709 7647 36773
rect 7711 36709 7727 36773
rect 7791 36709 7796 36773
rect 6602 36692 7796 36709
rect 6602 36628 6607 36692
rect 6671 36628 6687 36692
rect 6751 36628 6767 36692
rect 6831 36628 6847 36692
rect 6911 36628 6927 36692
rect 6991 36628 7007 36692
rect 7071 36628 7087 36692
rect 7151 36628 7167 36692
rect 7231 36628 7247 36692
rect 7311 36628 7327 36692
rect 7391 36628 7407 36692
rect 7471 36628 7487 36692
rect 7551 36628 7567 36692
rect 7631 36628 7647 36692
rect 7711 36628 7727 36692
rect 7791 36628 7796 36692
rect 6602 36611 7796 36628
rect 6602 36547 6607 36611
rect 6671 36547 6687 36611
rect 6751 36547 6767 36611
rect 6831 36547 6847 36611
rect 6911 36547 6927 36611
rect 6991 36547 7007 36611
rect 7071 36547 7087 36611
rect 7151 36547 7167 36611
rect 7231 36547 7247 36611
rect 7311 36547 7327 36611
rect 7391 36547 7407 36611
rect 7471 36547 7487 36611
rect 7551 36547 7567 36611
rect 7631 36547 7647 36611
rect 7711 36547 7727 36611
rect 7791 36547 7796 36611
rect 6602 36530 7796 36547
rect 6602 36466 6607 36530
rect 6671 36466 6687 36530
rect 6751 36466 6767 36530
rect 6831 36466 6847 36530
rect 6911 36466 6927 36530
rect 6991 36466 7007 36530
rect 7071 36466 7087 36530
rect 7151 36466 7167 36530
rect 7231 36466 7247 36530
rect 7311 36466 7327 36530
rect 7391 36466 7407 36530
rect 7471 36466 7487 36530
rect 7551 36466 7567 36530
rect 7631 36466 7647 36530
rect 7711 36466 7727 36530
rect 7791 36466 7796 36530
rect 6602 36449 7796 36466
rect 6602 36385 6607 36449
rect 6671 36385 6687 36449
rect 6751 36385 6767 36449
rect 6831 36385 6847 36449
rect 6911 36385 6927 36449
rect 6991 36385 7007 36449
rect 7071 36385 7087 36449
rect 7151 36385 7167 36449
rect 7231 36385 7247 36449
rect 7311 36385 7327 36449
rect 7391 36385 7407 36449
rect 7471 36385 7487 36449
rect 7551 36385 7567 36449
rect 7631 36385 7647 36449
rect 7711 36385 7727 36449
rect 7791 36385 7796 36449
rect 6602 36368 7796 36385
rect 6602 36304 6607 36368
rect 6671 36304 6687 36368
rect 6751 36304 6767 36368
rect 6831 36304 6847 36368
rect 6911 36304 6927 36368
rect 6991 36304 7007 36368
rect 7071 36304 7087 36368
rect 7151 36304 7167 36368
rect 7231 36304 7247 36368
rect 7311 36304 7327 36368
rect 7391 36304 7407 36368
rect 7471 36304 7487 36368
rect 7551 36304 7567 36368
rect 7631 36304 7647 36368
rect 7711 36304 7727 36368
rect 7791 36304 7796 36368
rect 6602 36287 7796 36304
rect 6602 36223 6607 36287
rect 6671 36223 6687 36287
rect 6751 36223 6767 36287
rect 6831 36223 6847 36287
rect 6911 36223 6927 36287
rect 6991 36223 7007 36287
rect 7071 36223 7087 36287
rect 7151 36223 7167 36287
rect 7231 36223 7247 36287
rect 7311 36223 7327 36287
rect 7391 36223 7407 36287
rect 7471 36223 7487 36287
rect 7551 36223 7567 36287
rect 7631 36223 7647 36287
rect 7711 36223 7727 36287
rect 7791 36223 7796 36287
rect 6602 36206 7796 36223
rect 6602 36142 6607 36206
rect 6671 36142 6687 36206
rect 6751 36142 6767 36206
rect 6831 36142 6847 36206
rect 6911 36142 6927 36206
rect 6991 36142 7007 36206
rect 7071 36142 7087 36206
rect 7151 36142 7167 36206
rect 7231 36142 7247 36206
rect 7311 36142 7327 36206
rect 7391 36142 7407 36206
rect 7471 36142 7487 36206
rect 7551 36142 7567 36206
rect 7631 36142 7647 36206
rect 7711 36142 7727 36206
rect 7791 36142 7796 36206
rect 6602 36124 7796 36142
rect 6602 36060 6607 36124
rect 6671 36060 6687 36124
rect 6751 36060 6767 36124
rect 6831 36060 6847 36124
rect 6911 36060 6927 36124
rect 6991 36060 7007 36124
rect 7071 36060 7087 36124
rect 7151 36060 7167 36124
rect 7231 36060 7247 36124
rect 7311 36060 7327 36124
rect 7391 36060 7407 36124
rect 7471 36060 7487 36124
rect 7551 36060 7567 36124
rect 7631 36060 7647 36124
rect 7711 36060 7727 36124
rect 7791 36060 7796 36124
rect 6602 36042 7796 36060
rect 6602 35978 6607 36042
rect 6671 35978 6687 36042
rect 6751 35978 6767 36042
rect 6831 35978 6847 36042
rect 6911 35978 6927 36042
rect 6991 35978 7007 36042
rect 7071 35978 7087 36042
rect 7151 35978 7167 36042
rect 7231 35978 7247 36042
rect 7311 35978 7327 36042
rect 7391 35978 7407 36042
rect 7471 35978 7487 36042
rect 7551 35978 7567 36042
rect 7631 35978 7647 36042
rect 7711 35978 7727 36042
rect 7791 35978 7796 36042
rect 6602 35960 7796 35978
rect 6602 35896 6607 35960
rect 6671 35896 6687 35960
rect 6751 35896 6767 35960
rect 6831 35896 6847 35960
rect 6911 35896 6927 35960
rect 6991 35896 7007 35960
rect 7071 35896 7087 35960
rect 7151 35896 7167 35960
rect 7231 35896 7247 35960
rect 7311 35896 7327 35960
rect 7391 35896 7407 35960
rect 7471 35896 7487 35960
rect 7551 35896 7567 35960
rect 7631 35896 7647 35960
rect 7711 35896 7727 35960
rect 7791 35896 7796 35960
rect 6602 35878 7796 35896
rect 6602 35814 6607 35878
rect 6671 35814 6687 35878
rect 6751 35814 6767 35878
rect 6831 35814 6847 35878
rect 6911 35814 6927 35878
rect 6991 35814 7007 35878
rect 7071 35814 7087 35878
rect 7151 35814 7167 35878
rect 7231 35814 7247 35878
rect 7311 35814 7327 35878
rect 7391 35814 7407 35878
rect 7471 35814 7487 35878
rect 7551 35814 7567 35878
rect 7631 35814 7647 35878
rect 7711 35814 7727 35878
rect 7791 35814 7796 35878
rect 6602 35796 7796 35814
rect 6602 35732 6607 35796
rect 6671 35732 6687 35796
rect 6751 35732 6767 35796
rect 6831 35732 6847 35796
rect 6911 35732 6927 35796
rect 6991 35732 7007 35796
rect 7071 35732 7087 35796
rect 7151 35732 7167 35796
rect 7231 35732 7247 35796
rect 7311 35732 7327 35796
rect 7391 35732 7407 35796
rect 7471 35732 7487 35796
rect 7551 35732 7567 35796
rect 7631 35732 7647 35796
rect 7711 35732 7727 35796
rect 7791 35732 7796 35796
rect 6602 35714 7796 35732
rect 6602 35650 6607 35714
rect 6671 35650 6687 35714
rect 6751 35650 6767 35714
rect 6831 35650 6847 35714
rect 6911 35650 6927 35714
rect 6991 35650 7007 35714
rect 7071 35650 7087 35714
rect 7151 35650 7167 35714
rect 7231 35650 7247 35714
rect 7311 35650 7327 35714
rect 7391 35650 7407 35714
rect 7471 35650 7487 35714
rect 7551 35650 7567 35714
rect 7631 35650 7647 35714
rect 7711 35650 7727 35714
rect 7791 35650 7796 35714
rect 6602 35632 7796 35650
rect 6602 35568 6607 35632
rect 6671 35568 6687 35632
rect 6751 35568 6767 35632
rect 6831 35568 6847 35632
rect 6911 35568 6927 35632
rect 6991 35568 7007 35632
rect 7071 35568 7087 35632
rect 7151 35568 7167 35632
rect 7231 35568 7247 35632
rect 7311 35568 7327 35632
rect 7391 35568 7407 35632
rect 7471 35568 7487 35632
rect 7551 35568 7567 35632
rect 7631 35568 7647 35632
rect 7711 35568 7727 35632
rect 7791 35568 7796 35632
rect 6602 35550 7796 35568
rect 6602 35486 6607 35550
rect 6671 35486 6687 35550
rect 6751 35486 6767 35550
rect 6831 35486 6847 35550
rect 6911 35486 6927 35550
rect 6991 35486 7007 35550
rect 7071 35486 7087 35550
rect 7151 35486 7167 35550
rect 7231 35486 7247 35550
rect 7311 35486 7327 35550
rect 7391 35486 7407 35550
rect 7471 35486 7487 35550
rect 7551 35486 7567 35550
rect 7631 35486 7647 35550
rect 7711 35486 7727 35550
rect 7791 35486 7796 35550
rect 6602 35468 7796 35486
rect 6602 35404 6607 35468
rect 6671 35404 6687 35468
rect 6751 35404 6767 35468
rect 6831 35404 6847 35468
rect 6911 35404 6927 35468
rect 6991 35404 7007 35468
rect 7071 35404 7087 35468
rect 7151 35404 7167 35468
rect 7231 35404 7247 35468
rect 7311 35404 7327 35468
rect 7391 35404 7407 35468
rect 7471 35404 7487 35468
rect 7551 35404 7567 35468
rect 7631 35404 7647 35468
rect 7711 35404 7727 35468
rect 7791 35404 7796 35468
rect 6602 35386 7796 35404
rect 6602 35322 6607 35386
rect 6671 35322 6687 35386
rect 6751 35322 6767 35386
rect 6831 35322 6847 35386
rect 6911 35322 6927 35386
rect 6991 35322 7007 35386
rect 7071 35322 7087 35386
rect 7151 35322 7167 35386
rect 7231 35322 7247 35386
rect 7311 35322 7327 35386
rect 7391 35322 7407 35386
rect 7471 35322 7487 35386
rect 7551 35322 7567 35386
rect 7631 35322 7647 35386
rect 7711 35322 7727 35386
rect 7791 35322 7796 35386
rect 6602 35304 7796 35322
rect 6602 35240 6607 35304
rect 6671 35240 6687 35304
rect 6751 35240 6767 35304
rect 6831 35240 6847 35304
rect 6911 35240 6927 35304
rect 6991 35240 7007 35304
rect 7071 35240 7087 35304
rect 7151 35240 7167 35304
rect 7231 35240 7247 35304
rect 7311 35240 7327 35304
rect 7391 35240 7407 35304
rect 7471 35240 7487 35304
rect 7551 35240 7567 35304
rect 7631 35240 7647 35304
rect 7711 35240 7727 35304
rect 7791 35240 7796 35304
rect 6602 35222 7796 35240
rect 6602 35158 6607 35222
rect 6671 35158 6687 35222
rect 6751 35158 6767 35222
rect 6831 35158 6847 35222
rect 6911 35158 6927 35222
rect 6991 35158 7007 35222
rect 7071 35158 7087 35222
rect 7151 35158 7167 35222
rect 7231 35158 7247 35222
rect 7311 35158 7327 35222
rect 7391 35158 7407 35222
rect 7471 35158 7487 35222
rect 7551 35158 7567 35222
rect 7631 35158 7647 35222
rect 7711 35158 7727 35222
rect 7791 35158 7796 35222
rect 6602 35157 7796 35158
rect 8095 39365 9289 39366
rect 8095 39301 8100 39365
rect 8164 39301 8180 39365
rect 8244 39301 8260 39365
rect 8324 39301 8340 39365
rect 8404 39301 8420 39365
rect 8484 39301 8500 39365
rect 8564 39301 8580 39365
rect 8644 39301 8660 39365
rect 8724 39301 8740 39365
rect 8804 39301 8820 39365
rect 8884 39301 8900 39365
rect 8964 39301 8980 39365
rect 9044 39301 9060 39365
rect 9124 39301 9140 39365
rect 9204 39301 9220 39365
rect 9284 39301 9289 39365
rect 8095 39284 9289 39301
rect 8095 39220 8100 39284
rect 8164 39220 8180 39284
rect 8244 39220 8260 39284
rect 8324 39220 8340 39284
rect 8404 39220 8420 39284
rect 8484 39220 8500 39284
rect 8564 39220 8580 39284
rect 8644 39220 8660 39284
rect 8724 39220 8740 39284
rect 8804 39220 8820 39284
rect 8884 39220 8900 39284
rect 8964 39220 8980 39284
rect 9044 39220 9060 39284
rect 9124 39220 9140 39284
rect 9204 39220 9220 39284
rect 9284 39220 9289 39284
rect 8095 39203 9289 39220
rect 8095 39139 8100 39203
rect 8164 39139 8180 39203
rect 8244 39139 8260 39203
rect 8324 39139 8340 39203
rect 8404 39139 8420 39203
rect 8484 39139 8500 39203
rect 8564 39139 8580 39203
rect 8644 39139 8660 39203
rect 8724 39139 8740 39203
rect 8804 39139 8820 39203
rect 8884 39139 8900 39203
rect 8964 39139 8980 39203
rect 9044 39139 9060 39203
rect 9124 39139 9140 39203
rect 9204 39139 9220 39203
rect 9284 39139 9289 39203
rect 8095 39122 9289 39139
rect 8095 39058 8100 39122
rect 8164 39058 8180 39122
rect 8244 39058 8260 39122
rect 8324 39058 8340 39122
rect 8404 39058 8420 39122
rect 8484 39058 8500 39122
rect 8564 39058 8580 39122
rect 8644 39058 8660 39122
rect 8724 39058 8740 39122
rect 8804 39058 8820 39122
rect 8884 39058 8900 39122
rect 8964 39058 8980 39122
rect 9044 39058 9060 39122
rect 9124 39058 9140 39122
rect 9204 39058 9220 39122
rect 9284 39058 9289 39122
rect 8095 39041 9289 39058
rect 8095 38977 8100 39041
rect 8164 38977 8180 39041
rect 8244 38977 8260 39041
rect 8324 38977 8340 39041
rect 8404 38977 8420 39041
rect 8484 38977 8500 39041
rect 8564 38977 8580 39041
rect 8644 38977 8660 39041
rect 8724 38977 8740 39041
rect 8804 38977 8820 39041
rect 8884 38977 8900 39041
rect 8964 38977 8980 39041
rect 9044 38977 9060 39041
rect 9124 38977 9140 39041
rect 9204 38977 9220 39041
rect 9284 38977 9289 39041
rect 8095 38960 9289 38977
rect 8095 38896 8100 38960
rect 8164 38896 8180 38960
rect 8244 38896 8260 38960
rect 8324 38896 8340 38960
rect 8404 38896 8420 38960
rect 8484 38896 8500 38960
rect 8564 38896 8580 38960
rect 8644 38896 8660 38960
rect 8724 38896 8740 38960
rect 8804 38896 8820 38960
rect 8884 38896 8900 38960
rect 8964 38896 8980 38960
rect 9044 38896 9060 38960
rect 9124 38896 9140 38960
rect 9204 38896 9220 38960
rect 9284 38896 9289 38960
rect 8095 38879 9289 38896
rect 8095 38815 8100 38879
rect 8164 38815 8180 38879
rect 8244 38815 8260 38879
rect 8324 38815 8340 38879
rect 8404 38815 8420 38879
rect 8484 38815 8500 38879
rect 8564 38815 8580 38879
rect 8644 38815 8660 38879
rect 8724 38815 8740 38879
rect 8804 38815 8820 38879
rect 8884 38815 8900 38879
rect 8964 38815 8980 38879
rect 9044 38815 9060 38879
rect 9124 38815 9140 38879
rect 9204 38815 9220 38879
rect 9284 38815 9289 38879
rect 8095 38798 9289 38815
rect 8095 38734 8100 38798
rect 8164 38734 8180 38798
rect 8244 38734 8260 38798
rect 8324 38734 8340 38798
rect 8404 38734 8420 38798
rect 8484 38734 8500 38798
rect 8564 38734 8580 38798
rect 8644 38734 8660 38798
rect 8724 38734 8740 38798
rect 8804 38734 8820 38798
rect 8884 38734 8900 38798
rect 8964 38734 8980 38798
rect 9044 38734 9060 38798
rect 9124 38734 9140 38798
rect 9204 38734 9220 38798
rect 9284 38734 9289 38798
rect 8095 38717 9289 38734
rect 8095 38653 8100 38717
rect 8164 38653 8180 38717
rect 8244 38653 8260 38717
rect 8324 38653 8340 38717
rect 8404 38653 8420 38717
rect 8484 38653 8500 38717
rect 8564 38653 8580 38717
rect 8644 38653 8660 38717
rect 8724 38653 8740 38717
rect 8804 38653 8820 38717
rect 8884 38653 8900 38717
rect 8964 38653 8980 38717
rect 9044 38653 9060 38717
rect 9124 38653 9140 38717
rect 9204 38653 9220 38717
rect 9284 38653 9289 38717
rect 8095 38636 9289 38653
rect 8095 38572 8100 38636
rect 8164 38572 8180 38636
rect 8244 38572 8260 38636
rect 8324 38572 8340 38636
rect 8404 38572 8420 38636
rect 8484 38572 8500 38636
rect 8564 38572 8580 38636
rect 8644 38572 8660 38636
rect 8724 38572 8740 38636
rect 8804 38572 8820 38636
rect 8884 38572 8900 38636
rect 8964 38572 8980 38636
rect 9044 38572 9060 38636
rect 9124 38572 9140 38636
rect 9204 38572 9220 38636
rect 9284 38572 9289 38636
rect 8095 38555 9289 38572
rect 8095 38491 8100 38555
rect 8164 38491 8180 38555
rect 8244 38491 8260 38555
rect 8324 38491 8340 38555
rect 8404 38491 8420 38555
rect 8484 38491 8500 38555
rect 8564 38491 8580 38555
rect 8644 38491 8660 38555
rect 8724 38491 8740 38555
rect 8804 38491 8820 38555
rect 8884 38491 8900 38555
rect 8964 38491 8980 38555
rect 9044 38491 9060 38555
rect 9124 38491 9140 38555
rect 9204 38491 9220 38555
rect 9284 38491 9289 38555
rect 8095 38474 9289 38491
rect 8095 38410 8100 38474
rect 8164 38410 8180 38474
rect 8244 38410 8260 38474
rect 8324 38410 8340 38474
rect 8404 38410 8420 38474
rect 8484 38410 8500 38474
rect 8564 38410 8580 38474
rect 8644 38410 8660 38474
rect 8724 38410 8740 38474
rect 8804 38410 8820 38474
rect 8884 38410 8900 38474
rect 8964 38410 8980 38474
rect 9044 38410 9060 38474
rect 9124 38410 9140 38474
rect 9204 38410 9220 38474
rect 9284 38410 9289 38474
rect 8095 38393 9289 38410
rect 8095 38329 8100 38393
rect 8164 38329 8180 38393
rect 8244 38329 8260 38393
rect 8324 38329 8340 38393
rect 8404 38329 8420 38393
rect 8484 38329 8500 38393
rect 8564 38329 8580 38393
rect 8644 38329 8660 38393
rect 8724 38329 8740 38393
rect 8804 38329 8820 38393
rect 8884 38329 8900 38393
rect 8964 38329 8980 38393
rect 9044 38329 9060 38393
rect 9124 38329 9140 38393
rect 9204 38329 9220 38393
rect 9284 38329 9289 38393
rect 8095 38312 9289 38329
rect 8095 38248 8100 38312
rect 8164 38248 8180 38312
rect 8244 38248 8260 38312
rect 8324 38248 8340 38312
rect 8404 38248 8420 38312
rect 8484 38248 8500 38312
rect 8564 38248 8580 38312
rect 8644 38248 8660 38312
rect 8724 38248 8740 38312
rect 8804 38248 8820 38312
rect 8884 38248 8900 38312
rect 8964 38248 8980 38312
rect 9044 38248 9060 38312
rect 9124 38248 9140 38312
rect 9204 38248 9220 38312
rect 9284 38248 9289 38312
rect 8095 38231 9289 38248
rect 8095 38167 8100 38231
rect 8164 38167 8180 38231
rect 8244 38167 8260 38231
rect 8324 38167 8340 38231
rect 8404 38167 8420 38231
rect 8484 38167 8500 38231
rect 8564 38167 8580 38231
rect 8644 38167 8660 38231
rect 8724 38167 8740 38231
rect 8804 38167 8820 38231
rect 8884 38167 8900 38231
rect 8964 38167 8980 38231
rect 9044 38167 9060 38231
rect 9124 38167 9140 38231
rect 9204 38167 9220 38231
rect 9284 38167 9289 38231
rect 8095 38150 9289 38167
rect 8095 38086 8100 38150
rect 8164 38086 8180 38150
rect 8244 38086 8260 38150
rect 8324 38086 8340 38150
rect 8404 38086 8420 38150
rect 8484 38086 8500 38150
rect 8564 38086 8580 38150
rect 8644 38086 8660 38150
rect 8724 38086 8740 38150
rect 8804 38086 8820 38150
rect 8884 38086 8900 38150
rect 8964 38086 8980 38150
rect 9044 38086 9060 38150
rect 9124 38086 9140 38150
rect 9204 38086 9220 38150
rect 9284 38086 9289 38150
rect 8095 38069 9289 38086
rect 8095 38005 8100 38069
rect 8164 38005 8180 38069
rect 8244 38005 8260 38069
rect 8324 38005 8340 38069
rect 8404 38005 8420 38069
rect 8484 38005 8500 38069
rect 8564 38005 8580 38069
rect 8644 38005 8660 38069
rect 8724 38005 8740 38069
rect 8804 38005 8820 38069
rect 8884 38005 8900 38069
rect 8964 38005 8980 38069
rect 9044 38005 9060 38069
rect 9124 38005 9140 38069
rect 9204 38005 9220 38069
rect 9284 38005 9289 38069
rect 8095 37988 9289 38005
rect 8095 37924 8100 37988
rect 8164 37924 8180 37988
rect 8244 37924 8260 37988
rect 8324 37924 8340 37988
rect 8404 37924 8420 37988
rect 8484 37924 8500 37988
rect 8564 37924 8580 37988
rect 8644 37924 8660 37988
rect 8724 37924 8740 37988
rect 8804 37924 8820 37988
rect 8884 37924 8900 37988
rect 8964 37924 8980 37988
rect 9044 37924 9060 37988
rect 9124 37924 9140 37988
rect 9204 37924 9220 37988
rect 9284 37924 9289 37988
rect 8095 37907 9289 37924
rect 8095 37843 8100 37907
rect 8164 37843 8180 37907
rect 8244 37843 8260 37907
rect 8324 37843 8340 37907
rect 8404 37843 8420 37907
rect 8484 37843 8500 37907
rect 8564 37843 8580 37907
rect 8644 37843 8660 37907
rect 8724 37843 8740 37907
rect 8804 37843 8820 37907
rect 8884 37843 8900 37907
rect 8964 37843 8980 37907
rect 9044 37843 9060 37907
rect 9124 37843 9140 37907
rect 9204 37843 9220 37907
rect 9284 37843 9289 37907
rect 8095 37826 9289 37843
rect 8095 37762 8100 37826
rect 8164 37762 8180 37826
rect 8244 37762 8260 37826
rect 8324 37762 8340 37826
rect 8404 37762 8420 37826
rect 8484 37762 8500 37826
rect 8564 37762 8580 37826
rect 8644 37762 8660 37826
rect 8724 37762 8740 37826
rect 8804 37762 8820 37826
rect 8884 37762 8900 37826
rect 8964 37762 8980 37826
rect 9044 37762 9060 37826
rect 9124 37762 9140 37826
rect 9204 37762 9220 37826
rect 9284 37762 9289 37826
rect 8095 37745 9289 37762
rect 8095 37681 8100 37745
rect 8164 37681 8180 37745
rect 8244 37681 8260 37745
rect 8324 37681 8340 37745
rect 8404 37681 8420 37745
rect 8484 37681 8500 37745
rect 8564 37681 8580 37745
rect 8644 37681 8660 37745
rect 8724 37681 8740 37745
rect 8804 37681 8820 37745
rect 8884 37681 8900 37745
rect 8964 37681 8980 37745
rect 9044 37681 9060 37745
rect 9124 37681 9140 37745
rect 9204 37681 9220 37745
rect 9284 37681 9289 37745
rect 8095 37664 9289 37681
rect 8095 37600 8100 37664
rect 8164 37600 8180 37664
rect 8244 37600 8260 37664
rect 8324 37600 8340 37664
rect 8404 37600 8420 37664
rect 8484 37600 8500 37664
rect 8564 37600 8580 37664
rect 8644 37600 8660 37664
rect 8724 37600 8740 37664
rect 8804 37600 8820 37664
rect 8884 37600 8900 37664
rect 8964 37600 8980 37664
rect 9044 37600 9060 37664
rect 9124 37600 9140 37664
rect 9204 37600 9220 37664
rect 9284 37600 9289 37664
rect 8095 37583 9289 37600
rect 8095 37519 8100 37583
rect 8164 37519 8180 37583
rect 8244 37519 8260 37583
rect 8324 37519 8340 37583
rect 8404 37519 8420 37583
rect 8484 37519 8500 37583
rect 8564 37519 8580 37583
rect 8644 37519 8660 37583
rect 8724 37519 8740 37583
rect 8804 37519 8820 37583
rect 8884 37519 8900 37583
rect 8964 37519 8980 37583
rect 9044 37519 9060 37583
rect 9124 37519 9140 37583
rect 9204 37519 9220 37583
rect 9284 37519 9289 37583
rect 8095 37502 9289 37519
rect 8095 37438 8100 37502
rect 8164 37438 8180 37502
rect 8244 37438 8260 37502
rect 8324 37438 8340 37502
rect 8404 37438 8420 37502
rect 8484 37438 8500 37502
rect 8564 37438 8580 37502
rect 8644 37438 8660 37502
rect 8724 37438 8740 37502
rect 8804 37438 8820 37502
rect 8884 37438 8900 37502
rect 8964 37438 8980 37502
rect 9044 37438 9060 37502
rect 9124 37438 9140 37502
rect 9204 37438 9220 37502
rect 9284 37438 9289 37502
rect 8095 37421 9289 37438
rect 8095 37357 8100 37421
rect 8164 37357 8180 37421
rect 8244 37357 8260 37421
rect 8324 37357 8340 37421
rect 8404 37357 8420 37421
rect 8484 37357 8500 37421
rect 8564 37357 8580 37421
rect 8644 37357 8660 37421
rect 8724 37357 8740 37421
rect 8804 37357 8820 37421
rect 8884 37357 8900 37421
rect 8964 37357 8980 37421
rect 9044 37357 9060 37421
rect 9124 37357 9140 37421
rect 9204 37357 9220 37421
rect 9284 37357 9289 37421
rect 8095 37340 9289 37357
rect 8095 37276 8100 37340
rect 8164 37276 8180 37340
rect 8244 37276 8260 37340
rect 8324 37276 8340 37340
rect 8404 37276 8420 37340
rect 8484 37276 8500 37340
rect 8564 37276 8580 37340
rect 8644 37276 8660 37340
rect 8724 37276 8740 37340
rect 8804 37276 8820 37340
rect 8884 37276 8900 37340
rect 8964 37276 8980 37340
rect 9044 37276 9060 37340
rect 9124 37276 9140 37340
rect 9204 37276 9220 37340
rect 9284 37276 9289 37340
rect 8095 37259 9289 37276
rect 8095 37195 8100 37259
rect 8164 37195 8180 37259
rect 8244 37195 8260 37259
rect 8324 37195 8340 37259
rect 8404 37195 8420 37259
rect 8484 37195 8500 37259
rect 8564 37195 8580 37259
rect 8644 37195 8660 37259
rect 8724 37195 8740 37259
rect 8804 37195 8820 37259
rect 8884 37195 8900 37259
rect 8964 37195 8980 37259
rect 9044 37195 9060 37259
rect 9124 37195 9140 37259
rect 9204 37195 9220 37259
rect 9284 37195 9289 37259
rect 8095 37178 9289 37195
rect 8095 37114 8100 37178
rect 8164 37114 8180 37178
rect 8244 37114 8260 37178
rect 8324 37114 8340 37178
rect 8404 37114 8420 37178
rect 8484 37114 8500 37178
rect 8564 37114 8580 37178
rect 8644 37114 8660 37178
rect 8724 37114 8740 37178
rect 8804 37114 8820 37178
rect 8884 37114 8900 37178
rect 8964 37114 8980 37178
rect 9044 37114 9060 37178
rect 9124 37114 9140 37178
rect 9204 37114 9220 37178
rect 9284 37114 9289 37178
rect 8095 37097 9289 37114
rect 8095 37033 8100 37097
rect 8164 37033 8180 37097
rect 8244 37033 8260 37097
rect 8324 37033 8340 37097
rect 8404 37033 8420 37097
rect 8484 37033 8500 37097
rect 8564 37033 8580 37097
rect 8644 37033 8660 37097
rect 8724 37033 8740 37097
rect 8804 37033 8820 37097
rect 8884 37033 8900 37097
rect 8964 37033 8980 37097
rect 9044 37033 9060 37097
rect 9124 37033 9140 37097
rect 9204 37033 9220 37097
rect 9284 37033 9289 37097
rect 8095 37016 9289 37033
rect 8095 36952 8100 37016
rect 8164 36952 8180 37016
rect 8244 36952 8260 37016
rect 8324 36952 8340 37016
rect 8404 36952 8420 37016
rect 8484 36952 8500 37016
rect 8564 36952 8580 37016
rect 8644 36952 8660 37016
rect 8724 36952 8740 37016
rect 8804 36952 8820 37016
rect 8884 36952 8900 37016
rect 8964 36952 8980 37016
rect 9044 36952 9060 37016
rect 9124 36952 9140 37016
rect 9204 36952 9220 37016
rect 9284 36952 9289 37016
rect 8095 36935 9289 36952
rect 8095 36871 8100 36935
rect 8164 36871 8180 36935
rect 8244 36871 8260 36935
rect 8324 36871 8340 36935
rect 8404 36871 8420 36935
rect 8484 36871 8500 36935
rect 8564 36871 8580 36935
rect 8644 36871 8660 36935
rect 8724 36871 8740 36935
rect 8804 36871 8820 36935
rect 8884 36871 8900 36935
rect 8964 36871 8980 36935
rect 9044 36871 9060 36935
rect 9124 36871 9140 36935
rect 9204 36871 9220 36935
rect 9284 36871 9289 36935
rect 8095 36854 9289 36871
rect 8095 36790 8100 36854
rect 8164 36790 8180 36854
rect 8244 36790 8260 36854
rect 8324 36790 8340 36854
rect 8404 36790 8420 36854
rect 8484 36790 8500 36854
rect 8564 36790 8580 36854
rect 8644 36790 8660 36854
rect 8724 36790 8740 36854
rect 8804 36790 8820 36854
rect 8884 36790 8900 36854
rect 8964 36790 8980 36854
rect 9044 36790 9060 36854
rect 9124 36790 9140 36854
rect 9204 36790 9220 36854
rect 9284 36790 9289 36854
rect 8095 36773 9289 36790
rect 8095 36709 8100 36773
rect 8164 36709 8180 36773
rect 8244 36709 8260 36773
rect 8324 36709 8340 36773
rect 8404 36709 8420 36773
rect 8484 36709 8500 36773
rect 8564 36709 8580 36773
rect 8644 36709 8660 36773
rect 8724 36709 8740 36773
rect 8804 36709 8820 36773
rect 8884 36709 8900 36773
rect 8964 36709 8980 36773
rect 9044 36709 9060 36773
rect 9124 36709 9140 36773
rect 9204 36709 9220 36773
rect 9284 36709 9289 36773
rect 8095 36692 9289 36709
rect 8095 36628 8100 36692
rect 8164 36628 8180 36692
rect 8244 36628 8260 36692
rect 8324 36628 8340 36692
rect 8404 36628 8420 36692
rect 8484 36628 8500 36692
rect 8564 36628 8580 36692
rect 8644 36628 8660 36692
rect 8724 36628 8740 36692
rect 8804 36628 8820 36692
rect 8884 36628 8900 36692
rect 8964 36628 8980 36692
rect 9044 36628 9060 36692
rect 9124 36628 9140 36692
rect 9204 36628 9220 36692
rect 9284 36628 9289 36692
rect 8095 36611 9289 36628
rect 8095 36547 8100 36611
rect 8164 36547 8180 36611
rect 8244 36547 8260 36611
rect 8324 36547 8340 36611
rect 8404 36547 8420 36611
rect 8484 36547 8500 36611
rect 8564 36547 8580 36611
rect 8644 36547 8660 36611
rect 8724 36547 8740 36611
rect 8804 36547 8820 36611
rect 8884 36547 8900 36611
rect 8964 36547 8980 36611
rect 9044 36547 9060 36611
rect 9124 36547 9140 36611
rect 9204 36547 9220 36611
rect 9284 36547 9289 36611
rect 8095 36530 9289 36547
rect 8095 36466 8100 36530
rect 8164 36466 8180 36530
rect 8244 36466 8260 36530
rect 8324 36466 8340 36530
rect 8404 36466 8420 36530
rect 8484 36466 8500 36530
rect 8564 36466 8580 36530
rect 8644 36466 8660 36530
rect 8724 36466 8740 36530
rect 8804 36466 8820 36530
rect 8884 36466 8900 36530
rect 8964 36466 8980 36530
rect 9044 36466 9060 36530
rect 9124 36466 9140 36530
rect 9204 36466 9220 36530
rect 9284 36466 9289 36530
rect 8095 36449 9289 36466
rect 8095 36385 8100 36449
rect 8164 36385 8180 36449
rect 8244 36385 8260 36449
rect 8324 36385 8340 36449
rect 8404 36385 8420 36449
rect 8484 36385 8500 36449
rect 8564 36385 8580 36449
rect 8644 36385 8660 36449
rect 8724 36385 8740 36449
rect 8804 36385 8820 36449
rect 8884 36385 8900 36449
rect 8964 36385 8980 36449
rect 9044 36385 9060 36449
rect 9124 36385 9140 36449
rect 9204 36385 9220 36449
rect 9284 36385 9289 36449
rect 8095 36368 9289 36385
rect 8095 36304 8100 36368
rect 8164 36304 8180 36368
rect 8244 36304 8260 36368
rect 8324 36304 8340 36368
rect 8404 36304 8420 36368
rect 8484 36304 8500 36368
rect 8564 36304 8580 36368
rect 8644 36304 8660 36368
rect 8724 36304 8740 36368
rect 8804 36304 8820 36368
rect 8884 36304 8900 36368
rect 8964 36304 8980 36368
rect 9044 36304 9060 36368
rect 9124 36304 9140 36368
rect 9204 36304 9220 36368
rect 9284 36304 9289 36368
rect 8095 36287 9289 36304
rect 8095 36223 8100 36287
rect 8164 36223 8180 36287
rect 8244 36223 8260 36287
rect 8324 36223 8340 36287
rect 8404 36223 8420 36287
rect 8484 36223 8500 36287
rect 8564 36223 8580 36287
rect 8644 36223 8660 36287
rect 8724 36223 8740 36287
rect 8804 36223 8820 36287
rect 8884 36223 8900 36287
rect 8964 36223 8980 36287
rect 9044 36223 9060 36287
rect 9124 36223 9140 36287
rect 9204 36223 9220 36287
rect 9284 36223 9289 36287
rect 8095 36206 9289 36223
rect 8095 36142 8100 36206
rect 8164 36142 8180 36206
rect 8244 36142 8260 36206
rect 8324 36142 8340 36206
rect 8404 36142 8420 36206
rect 8484 36142 8500 36206
rect 8564 36142 8580 36206
rect 8644 36142 8660 36206
rect 8724 36142 8740 36206
rect 8804 36142 8820 36206
rect 8884 36142 8900 36206
rect 8964 36142 8980 36206
rect 9044 36142 9060 36206
rect 9124 36142 9140 36206
rect 9204 36142 9220 36206
rect 9284 36142 9289 36206
rect 8095 36124 9289 36142
rect 8095 36060 8100 36124
rect 8164 36060 8180 36124
rect 8244 36060 8260 36124
rect 8324 36060 8340 36124
rect 8404 36060 8420 36124
rect 8484 36060 8500 36124
rect 8564 36060 8580 36124
rect 8644 36060 8660 36124
rect 8724 36060 8740 36124
rect 8804 36060 8820 36124
rect 8884 36060 8900 36124
rect 8964 36060 8980 36124
rect 9044 36060 9060 36124
rect 9124 36060 9140 36124
rect 9204 36060 9220 36124
rect 9284 36060 9289 36124
rect 8095 36042 9289 36060
rect 8095 35978 8100 36042
rect 8164 35978 8180 36042
rect 8244 35978 8260 36042
rect 8324 35978 8340 36042
rect 8404 35978 8420 36042
rect 8484 35978 8500 36042
rect 8564 35978 8580 36042
rect 8644 35978 8660 36042
rect 8724 35978 8740 36042
rect 8804 35978 8820 36042
rect 8884 35978 8900 36042
rect 8964 35978 8980 36042
rect 9044 35978 9060 36042
rect 9124 35978 9140 36042
rect 9204 35978 9220 36042
rect 9284 35978 9289 36042
rect 8095 35960 9289 35978
rect 8095 35896 8100 35960
rect 8164 35896 8180 35960
rect 8244 35896 8260 35960
rect 8324 35896 8340 35960
rect 8404 35896 8420 35960
rect 8484 35896 8500 35960
rect 8564 35896 8580 35960
rect 8644 35896 8660 35960
rect 8724 35896 8740 35960
rect 8804 35896 8820 35960
rect 8884 35896 8900 35960
rect 8964 35896 8980 35960
rect 9044 35896 9060 35960
rect 9124 35896 9140 35960
rect 9204 35896 9220 35960
rect 9284 35896 9289 35960
rect 8095 35878 9289 35896
rect 8095 35814 8100 35878
rect 8164 35814 8180 35878
rect 8244 35814 8260 35878
rect 8324 35814 8340 35878
rect 8404 35814 8420 35878
rect 8484 35814 8500 35878
rect 8564 35814 8580 35878
rect 8644 35814 8660 35878
rect 8724 35814 8740 35878
rect 8804 35814 8820 35878
rect 8884 35814 8900 35878
rect 8964 35814 8980 35878
rect 9044 35814 9060 35878
rect 9124 35814 9140 35878
rect 9204 35814 9220 35878
rect 9284 35814 9289 35878
rect 8095 35796 9289 35814
rect 8095 35732 8100 35796
rect 8164 35732 8180 35796
rect 8244 35732 8260 35796
rect 8324 35732 8340 35796
rect 8404 35732 8420 35796
rect 8484 35732 8500 35796
rect 8564 35732 8580 35796
rect 8644 35732 8660 35796
rect 8724 35732 8740 35796
rect 8804 35732 8820 35796
rect 8884 35732 8900 35796
rect 8964 35732 8980 35796
rect 9044 35732 9060 35796
rect 9124 35732 9140 35796
rect 9204 35732 9220 35796
rect 9284 35732 9289 35796
rect 8095 35714 9289 35732
rect 8095 35650 8100 35714
rect 8164 35650 8180 35714
rect 8244 35650 8260 35714
rect 8324 35650 8340 35714
rect 8404 35650 8420 35714
rect 8484 35650 8500 35714
rect 8564 35650 8580 35714
rect 8644 35650 8660 35714
rect 8724 35650 8740 35714
rect 8804 35650 8820 35714
rect 8884 35650 8900 35714
rect 8964 35650 8980 35714
rect 9044 35650 9060 35714
rect 9124 35650 9140 35714
rect 9204 35650 9220 35714
rect 9284 35650 9289 35714
rect 8095 35632 9289 35650
rect 8095 35568 8100 35632
rect 8164 35568 8180 35632
rect 8244 35568 8260 35632
rect 8324 35568 8340 35632
rect 8404 35568 8420 35632
rect 8484 35568 8500 35632
rect 8564 35568 8580 35632
rect 8644 35568 8660 35632
rect 8724 35568 8740 35632
rect 8804 35568 8820 35632
rect 8884 35568 8900 35632
rect 8964 35568 8980 35632
rect 9044 35568 9060 35632
rect 9124 35568 9140 35632
rect 9204 35568 9220 35632
rect 9284 35568 9289 35632
rect 8095 35550 9289 35568
rect 8095 35486 8100 35550
rect 8164 35486 8180 35550
rect 8244 35486 8260 35550
rect 8324 35486 8340 35550
rect 8404 35486 8420 35550
rect 8484 35486 8500 35550
rect 8564 35486 8580 35550
rect 8644 35486 8660 35550
rect 8724 35486 8740 35550
rect 8804 35486 8820 35550
rect 8884 35486 8900 35550
rect 8964 35486 8980 35550
rect 9044 35486 9060 35550
rect 9124 35486 9140 35550
rect 9204 35486 9220 35550
rect 9284 35486 9289 35550
rect 8095 35468 9289 35486
rect 8095 35404 8100 35468
rect 8164 35404 8180 35468
rect 8244 35404 8260 35468
rect 8324 35404 8340 35468
rect 8404 35404 8420 35468
rect 8484 35404 8500 35468
rect 8564 35404 8580 35468
rect 8644 35404 8660 35468
rect 8724 35404 8740 35468
rect 8804 35404 8820 35468
rect 8884 35404 8900 35468
rect 8964 35404 8980 35468
rect 9044 35404 9060 35468
rect 9124 35404 9140 35468
rect 9204 35404 9220 35468
rect 9284 35404 9289 35468
rect 8095 35386 9289 35404
rect 8095 35322 8100 35386
rect 8164 35322 8180 35386
rect 8244 35322 8260 35386
rect 8324 35322 8340 35386
rect 8404 35322 8420 35386
rect 8484 35322 8500 35386
rect 8564 35322 8580 35386
rect 8644 35322 8660 35386
rect 8724 35322 8740 35386
rect 8804 35322 8820 35386
rect 8884 35322 8900 35386
rect 8964 35322 8980 35386
rect 9044 35322 9060 35386
rect 9124 35322 9140 35386
rect 9204 35322 9220 35386
rect 9284 35322 9289 35386
rect 8095 35304 9289 35322
rect 8095 35240 8100 35304
rect 8164 35240 8180 35304
rect 8244 35240 8260 35304
rect 8324 35240 8340 35304
rect 8404 35240 8420 35304
rect 8484 35240 8500 35304
rect 8564 35240 8580 35304
rect 8644 35240 8660 35304
rect 8724 35240 8740 35304
rect 8804 35240 8820 35304
rect 8884 35240 8900 35304
rect 8964 35240 8980 35304
rect 9044 35240 9060 35304
rect 9124 35240 9140 35304
rect 9204 35240 9220 35304
rect 9284 35240 9289 35304
rect 8095 35222 9289 35240
rect 8095 35158 8100 35222
rect 8164 35158 8180 35222
rect 8244 35158 8260 35222
rect 8324 35158 8340 35222
rect 8404 35158 8420 35222
rect 8484 35158 8500 35222
rect 8564 35158 8580 35222
rect 8644 35158 8660 35222
rect 8724 35158 8740 35222
rect 8804 35158 8820 35222
rect 8884 35158 8900 35222
rect 8964 35158 8980 35222
rect 9044 35158 9060 35222
rect 9124 35158 9140 35222
rect 9204 35158 9220 35222
rect 9284 35158 9289 35222
rect 8095 35157 9289 35158
rect 9592 39365 10786 39366
rect 9592 39301 9597 39365
rect 9661 39301 9677 39365
rect 9741 39301 9757 39365
rect 9821 39301 9837 39365
rect 9901 39301 9917 39365
rect 9981 39301 9997 39365
rect 10061 39301 10077 39365
rect 10141 39301 10157 39365
rect 10221 39301 10237 39365
rect 10301 39301 10317 39365
rect 10381 39301 10397 39365
rect 10461 39301 10477 39365
rect 10541 39301 10557 39365
rect 10621 39301 10637 39365
rect 10701 39301 10717 39365
rect 10781 39301 10786 39365
rect 9592 39284 10786 39301
rect 9592 39220 9597 39284
rect 9661 39220 9677 39284
rect 9741 39220 9757 39284
rect 9821 39220 9837 39284
rect 9901 39220 9917 39284
rect 9981 39220 9997 39284
rect 10061 39220 10077 39284
rect 10141 39220 10157 39284
rect 10221 39220 10237 39284
rect 10301 39220 10317 39284
rect 10381 39220 10397 39284
rect 10461 39220 10477 39284
rect 10541 39220 10557 39284
rect 10621 39220 10637 39284
rect 10701 39220 10717 39284
rect 10781 39220 10786 39284
rect 9592 39203 10786 39220
rect 9592 39139 9597 39203
rect 9661 39139 9677 39203
rect 9741 39139 9757 39203
rect 9821 39139 9837 39203
rect 9901 39139 9917 39203
rect 9981 39139 9997 39203
rect 10061 39139 10077 39203
rect 10141 39139 10157 39203
rect 10221 39139 10237 39203
rect 10301 39139 10317 39203
rect 10381 39139 10397 39203
rect 10461 39139 10477 39203
rect 10541 39139 10557 39203
rect 10621 39139 10637 39203
rect 10701 39139 10717 39203
rect 10781 39139 10786 39203
rect 9592 39122 10786 39139
rect 9592 39058 9597 39122
rect 9661 39058 9677 39122
rect 9741 39058 9757 39122
rect 9821 39058 9837 39122
rect 9901 39058 9917 39122
rect 9981 39058 9997 39122
rect 10061 39058 10077 39122
rect 10141 39058 10157 39122
rect 10221 39058 10237 39122
rect 10301 39058 10317 39122
rect 10381 39058 10397 39122
rect 10461 39058 10477 39122
rect 10541 39058 10557 39122
rect 10621 39058 10637 39122
rect 10701 39058 10717 39122
rect 10781 39058 10786 39122
rect 9592 39041 10786 39058
rect 9592 38977 9597 39041
rect 9661 38977 9677 39041
rect 9741 38977 9757 39041
rect 9821 38977 9837 39041
rect 9901 38977 9917 39041
rect 9981 38977 9997 39041
rect 10061 38977 10077 39041
rect 10141 38977 10157 39041
rect 10221 38977 10237 39041
rect 10301 38977 10317 39041
rect 10381 38977 10397 39041
rect 10461 38977 10477 39041
rect 10541 38977 10557 39041
rect 10621 38977 10637 39041
rect 10701 38977 10717 39041
rect 10781 38977 10786 39041
rect 9592 38960 10786 38977
rect 9592 38896 9597 38960
rect 9661 38896 9677 38960
rect 9741 38896 9757 38960
rect 9821 38896 9837 38960
rect 9901 38896 9917 38960
rect 9981 38896 9997 38960
rect 10061 38896 10077 38960
rect 10141 38896 10157 38960
rect 10221 38896 10237 38960
rect 10301 38896 10317 38960
rect 10381 38896 10397 38960
rect 10461 38896 10477 38960
rect 10541 38896 10557 38960
rect 10621 38896 10637 38960
rect 10701 38896 10717 38960
rect 10781 38896 10786 38960
rect 9592 38879 10786 38896
rect 9592 38815 9597 38879
rect 9661 38815 9677 38879
rect 9741 38815 9757 38879
rect 9821 38815 9837 38879
rect 9901 38815 9917 38879
rect 9981 38815 9997 38879
rect 10061 38815 10077 38879
rect 10141 38815 10157 38879
rect 10221 38815 10237 38879
rect 10301 38815 10317 38879
rect 10381 38815 10397 38879
rect 10461 38815 10477 38879
rect 10541 38815 10557 38879
rect 10621 38815 10637 38879
rect 10701 38815 10717 38879
rect 10781 38815 10786 38879
rect 9592 38798 10786 38815
rect 9592 38734 9597 38798
rect 9661 38734 9677 38798
rect 9741 38734 9757 38798
rect 9821 38734 9837 38798
rect 9901 38734 9917 38798
rect 9981 38734 9997 38798
rect 10061 38734 10077 38798
rect 10141 38734 10157 38798
rect 10221 38734 10237 38798
rect 10301 38734 10317 38798
rect 10381 38734 10397 38798
rect 10461 38734 10477 38798
rect 10541 38734 10557 38798
rect 10621 38734 10637 38798
rect 10701 38734 10717 38798
rect 10781 38734 10786 38798
rect 9592 38717 10786 38734
rect 9592 38653 9597 38717
rect 9661 38653 9677 38717
rect 9741 38653 9757 38717
rect 9821 38653 9837 38717
rect 9901 38653 9917 38717
rect 9981 38653 9997 38717
rect 10061 38653 10077 38717
rect 10141 38653 10157 38717
rect 10221 38653 10237 38717
rect 10301 38653 10317 38717
rect 10381 38653 10397 38717
rect 10461 38653 10477 38717
rect 10541 38653 10557 38717
rect 10621 38653 10637 38717
rect 10701 38653 10717 38717
rect 10781 38653 10786 38717
rect 9592 38636 10786 38653
rect 9592 38572 9597 38636
rect 9661 38572 9677 38636
rect 9741 38572 9757 38636
rect 9821 38572 9837 38636
rect 9901 38572 9917 38636
rect 9981 38572 9997 38636
rect 10061 38572 10077 38636
rect 10141 38572 10157 38636
rect 10221 38572 10237 38636
rect 10301 38572 10317 38636
rect 10381 38572 10397 38636
rect 10461 38572 10477 38636
rect 10541 38572 10557 38636
rect 10621 38572 10637 38636
rect 10701 38572 10717 38636
rect 10781 38572 10786 38636
rect 9592 38555 10786 38572
rect 9592 38491 9597 38555
rect 9661 38491 9677 38555
rect 9741 38491 9757 38555
rect 9821 38491 9837 38555
rect 9901 38491 9917 38555
rect 9981 38491 9997 38555
rect 10061 38491 10077 38555
rect 10141 38491 10157 38555
rect 10221 38491 10237 38555
rect 10301 38491 10317 38555
rect 10381 38491 10397 38555
rect 10461 38491 10477 38555
rect 10541 38491 10557 38555
rect 10621 38491 10637 38555
rect 10701 38491 10717 38555
rect 10781 38491 10786 38555
rect 9592 38474 10786 38491
rect 9592 38410 9597 38474
rect 9661 38410 9677 38474
rect 9741 38410 9757 38474
rect 9821 38410 9837 38474
rect 9901 38410 9917 38474
rect 9981 38410 9997 38474
rect 10061 38410 10077 38474
rect 10141 38410 10157 38474
rect 10221 38410 10237 38474
rect 10301 38410 10317 38474
rect 10381 38410 10397 38474
rect 10461 38410 10477 38474
rect 10541 38410 10557 38474
rect 10621 38410 10637 38474
rect 10701 38410 10717 38474
rect 10781 38410 10786 38474
rect 9592 38393 10786 38410
rect 9592 38329 9597 38393
rect 9661 38329 9677 38393
rect 9741 38329 9757 38393
rect 9821 38329 9837 38393
rect 9901 38329 9917 38393
rect 9981 38329 9997 38393
rect 10061 38329 10077 38393
rect 10141 38329 10157 38393
rect 10221 38329 10237 38393
rect 10301 38329 10317 38393
rect 10381 38329 10397 38393
rect 10461 38329 10477 38393
rect 10541 38329 10557 38393
rect 10621 38329 10637 38393
rect 10701 38329 10717 38393
rect 10781 38329 10786 38393
rect 9592 38312 10786 38329
rect 9592 38248 9597 38312
rect 9661 38248 9677 38312
rect 9741 38248 9757 38312
rect 9821 38248 9837 38312
rect 9901 38248 9917 38312
rect 9981 38248 9997 38312
rect 10061 38248 10077 38312
rect 10141 38248 10157 38312
rect 10221 38248 10237 38312
rect 10301 38248 10317 38312
rect 10381 38248 10397 38312
rect 10461 38248 10477 38312
rect 10541 38248 10557 38312
rect 10621 38248 10637 38312
rect 10701 38248 10717 38312
rect 10781 38248 10786 38312
rect 9592 38231 10786 38248
rect 9592 38167 9597 38231
rect 9661 38167 9677 38231
rect 9741 38167 9757 38231
rect 9821 38167 9837 38231
rect 9901 38167 9917 38231
rect 9981 38167 9997 38231
rect 10061 38167 10077 38231
rect 10141 38167 10157 38231
rect 10221 38167 10237 38231
rect 10301 38167 10317 38231
rect 10381 38167 10397 38231
rect 10461 38167 10477 38231
rect 10541 38167 10557 38231
rect 10621 38167 10637 38231
rect 10701 38167 10717 38231
rect 10781 38167 10786 38231
rect 9592 38150 10786 38167
rect 9592 38086 9597 38150
rect 9661 38086 9677 38150
rect 9741 38086 9757 38150
rect 9821 38086 9837 38150
rect 9901 38086 9917 38150
rect 9981 38086 9997 38150
rect 10061 38086 10077 38150
rect 10141 38086 10157 38150
rect 10221 38086 10237 38150
rect 10301 38086 10317 38150
rect 10381 38086 10397 38150
rect 10461 38086 10477 38150
rect 10541 38086 10557 38150
rect 10621 38086 10637 38150
rect 10701 38086 10717 38150
rect 10781 38086 10786 38150
rect 9592 38069 10786 38086
rect 9592 38005 9597 38069
rect 9661 38005 9677 38069
rect 9741 38005 9757 38069
rect 9821 38005 9837 38069
rect 9901 38005 9917 38069
rect 9981 38005 9997 38069
rect 10061 38005 10077 38069
rect 10141 38005 10157 38069
rect 10221 38005 10237 38069
rect 10301 38005 10317 38069
rect 10381 38005 10397 38069
rect 10461 38005 10477 38069
rect 10541 38005 10557 38069
rect 10621 38005 10637 38069
rect 10701 38005 10717 38069
rect 10781 38005 10786 38069
rect 9592 37988 10786 38005
rect 9592 37924 9597 37988
rect 9661 37924 9677 37988
rect 9741 37924 9757 37988
rect 9821 37924 9837 37988
rect 9901 37924 9917 37988
rect 9981 37924 9997 37988
rect 10061 37924 10077 37988
rect 10141 37924 10157 37988
rect 10221 37924 10237 37988
rect 10301 37924 10317 37988
rect 10381 37924 10397 37988
rect 10461 37924 10477 37988
rect 10541 37924 10557 37988
rect 10621 37924 10637 37988
rect 10701 37924 10717 37988
rect 10781 37924 10786 37988
rect 9592 37907 10786 37924
rect 9592 37843 9597 37907
rect 9661 37843 9677 37907
rect 9741 37843 9757 37907
rect 9821 37843 9837 37907
rect 9901 37843 9917 37907
rect 9981 37843 9997 37907
rect 10061 37843 10077 37907
rect 10141 37843 10157 37907
rect 10221 37843 10237 37907
rect 10301 37843 10317 37907
rect 10381 37843 10397 37907
rect 10461 37843 10477 37907
rect 10541 37843 10557 37907
rect 10621 37843 10637 37907
rect 10701 37843 10717 37907
rect 10781 37843 10786 37907
rect 9592 37826 10786 37843
rect 9592 37762 9597 37826
rect 9661 37762 9677 37826
rect 9741 37762 9757 37826
rect 9821 37762 9837 37826
rect 9901 37762 9917 37826
rect 9981 37762 9997 37826
rect 10061 37762 10077 37826
rect 10141 37762 10157 37826
rect 10221 37762 10237 37826
rect 10301 37762 10317 37826
rect 10381 37762 10397 37826
rect 10461 37762 10477 37826
rect 10541 37762 10557 37826
rect 10621 37762 10637 37826
rect 10701 37762 10717 37826
rect 10781 37762 10786 37826
rect 9592 37745 10786 37762
rect 9592 37681 9597 37745
rect 9661 37681 9677 37745
rect 9741 37681 9757 37745
rect 9821 37681 9837 37745
rect 9901 37681 9917 37745
rect 9981 37681 9997 37745
rect 10061 37681 10077 37745
rect 10141 37681 10157 37745
rect 10221 37681 10237 37745
rect 10301 37681 10317 37745
rect 10381 37681 10397 37745
rect 10461 37681 10477 37745
rect 10541 37681 10557 37745
rect 10621 37681 10637 37745
rect 10701 37681 10717 37745
rect 10781 37681 10786 37745
rect 9592 37664 10786 37681
rect 9592 37600 9597 37664
rect 9661 37600 9677 37664
rect 9741 37600 9757 37664
rect 9821 37600 9837 37664
rect 9901 37600 9917 37664
rect 9981 37600 9997 37664
rect 10061 37600 10077 37664
rect 10141 37600 10157 37664
rect 10221 37600 10237 37664
rect 10301 37600 10317 37664
rect 10381 37600 10397 37664
rect 10461 37600 10477 37664
rect 10541 37600 10557 37664
rect 10621 37600 10637 37664
rect 10701 37600 10717 37664
rect 10781 37600 10786 37664
rect 9592 37583 10786 37600
rect 9592 37519 9597 37583
rect 9661 37519 9677 37583
rect 9741 37519 9757 37583
rect 9821 37519 9837 37583
rect 9901 37519 9917 37583
rect 9981 37519 9997 37583
rect 10061 37519 10077 37583
rect 10141 37519 10157 37583
rect 10221 37519 10237 37583
rect 10301 37519 10317 37583
rect 10381 37519 10397 37583
rect 10461 37519 10477 37583
rect 10541 37519 10557 37583
rect 10621 37519 10637 37583
rect 10701 37519 10717 37583
rect 10781 37519 10786 37583
rect 9592 37502 10786 37519
rect 9592 37438 9597 37502
rect 9661 37438 9677 37502
rect 9741 37438 9757 37502
rect 9821 37438 9837 37502
rect 9901 37438 9917 37502
rect 9981 37438 9997 37502
rect 10061 37438 10077 37502
rect 10141 37438 10157 37502
rect 10221 37438 10237 37502
rect 10301 37438 10317 37502
rect 10381 37438 10397 37502
rect 10461 37438 10477 37502
rect 10541 37438 10557 37502
rect 10621 37438 10637 37502
rect 10701 37438 10717 37502
rect 10781 37438 10786 37502
rect 9592 37421 10786 37438
rect 9592 37357 9597 37421
rect 9661 37357 9677 37421
rect 9741 37357 9757 37421
rect 9821 37357 9837 37421
rect 9901 37357 9917 37421
rect 9981 37357 9997 37421
rect 10061 37357 10077 37421
rect 10141 37357 10157 37421
rect 10221 37357 10237 37421
rect 10301 37357 10317 37421
rect 10381 37357 10397 37421
rect 10461 37357 10477 37421
rect 10541 37357 10557 37421
rect 10621 37357 10637 37421
rect 10701 37357 10717 37421
rect 10781 37357 10786 37421
rect 9592 37340 10786 37357
rect 9592 37276 9597 37340
rect 9661 37276 9677 37340
rect 9741 37276 9757 37340
rect 9821 37276 9837 37340
rect 9901 37276 9917 37340
rect 9981 37276 9997 37340
rect 10061 37276 10077 37340
rect 10141 37276 10157 37340
rect 10221 37276 10237 37340
rect 10301 37276 10317 37340
rect 10381 37276 10397 37340
rect 10461 37276 10477 37340
rect 10541 37276 10557 37340
rect 10621 37276 10637 37340
rect 10701 37276 10717 37340
rect 10781 37276 10786 37340
rect 9592 37259 10786 37276
rect 9592 37195 9597 37259
rect 9661 37195 9677 37259
rect 9741 37195 9757 37259
rect 9821 37195 9837 37259
rect 9901 37195 9917 37259
rect 9981 37195 9997 37259
rect 10061 37195 10077 37259
rect 10141 37195 10157 37259
rect 10221 37195 10237 37259
rect 10301 37195 10317 37259
rect 10381 37195 10397 37259
rect 10461 37195 10477 37259
rect 10541 37195 10557 37259
rect 10621 37195 10637 37259
rect 10701 37195 10717 37259
rect 10781 37195 10786 37259
rect 9592 37178 10786 37195
rect 9592 37114 9597 37178
rect 9661 37114 9677 37178
rect 9741 37114 9757 37178
rect 9821 37114 9837 37178
rect 9901 37114 9917 37178
rect 9981 37114 9997 37178
rect 10061 37114 10077 37178
rect 10141 37114 10157 37178
rect 10221 37114 10237 37178
rect 10301 37114 10317 37178
rect 10381 37114 10397 37178
rect 10461 37114 10477 37178
rect 10541 37114 10557 37178
rect 10621 37114 10637 37178
rect 10701 37114 10717 37178
rect 10781 37114 10786 37178
rect 9592 37097 10786 37114
rect 9592 37033 9597 37097
rect 9661 37033 9677 37097
rect 9741 37033 9757 37097
rect 9821 37033 9837 37097
rect 9901 37033 9917 37097
rect 9981 37033 9997 37097
rect 10061 37033 10077 37097
rect 10141 37033 10157 37097
rect 10221 37033 10237 37097
rect 10301 37033 10317 37097
rect 10381 37033 10397 37097
rect 10461 37033 10477 37097
rect 10541 37033 10557 37097
rect 10621 37033 10637 37097
rect 10701 37033 10717 37097
rect 10781 37033 10786 37097
rect 9592 37016 10786 37033
rect 9592 36952 9597 37016
rect 9661 36952 9677 37016
rect 9741 36952 9757 37016
rect 9821 36952 9837 37016
rect 9901 36952 9917 37016
rect 9981 36952 9997 37016
rect 10061 36952 10077 37016
rect 10141 36952 10157 37016
rect 10221 36952 10237 37016
rect 10301 36952 10317 37016
rect 10381 36952 10397 37016
rect 10461 36952 10477 37016
rect 10541 36952 10557 37016
rect 10621 36952 10637 37016
rect 10701 36952 10717 37016
rect 10781 36952 10786 37016
rect 9592 36935 10786 36952
rect 9592 36871 9597 36935
rect 9661 36871 9677 36935
rect 9741 36871 9757 36935
rect 9821 36871 9837 36935
rect 9901 36871 9917 36935
rect 9981 36871 9997 36935
rect 10061 36871 10077 36935
rect 10141 36871 10157 36935
rect 10221 36871 10237 36935
rect 10301 36871 10317 36935
rect 10381 36871 10397 36935
rect 10461 36871 10477 36935
rect 10541 36871 10557 36935
rect 10621 36871 10637 36935
rect 10701 36871 10717 36935
rect 10781 36871 10786 36935
rect 9592 36854 10786 36871
rect 9592 36790 9597 36854
rect 9661 36790 9677 36854
rect 9741 36790 9757 36854
rect 9821 36790 9837 36854
rect 9901 36790 9917 36854
rect 9981 36790 9997 36854
rect 10061 36790 10077 36854
rect 10141 36790 10157 36854
rect 10221 36790 10237 36854
rect 10301 36790 10317 36854
rect 10381 36790 10397 36854
rect 10461 36790 10477 36854
rect 10541 36790 10557 36854
rect 10621 36790 10637 36854
rect 10701 36790 10717 36854
rect 10781 36790 10786 36854
rect 9592 36773 10786 36790
rect 9592 36709 9597 36773
rect 9661 36709 9677 36773
rect 9741 36709 9757 36773
rect 9821 36709 9837 36773
rect 9901 36709 9917 36773
rect 9981 36709 9997 36773
rect 10061 36709 10077 36773
rect 10141 36709 10157 36773
rect 10221 36709 10237 36773
rect 10301 36709 10317 36773
rect 10381 36709 10397 36773
rect 10461 36709 10477 36773
rect 10541 36709 10557 36773
rect 10621 36709 10637 36773
rect 10701 36709 10717 36773
rect 10781 36709 10786 36773
rect 9592 36692 10786 36709
rect 9592 36628 9597 36692
rect 9661 36628 9677 36692
rect 9741 36628 9757 36692
rect 9821 36628 9837 36692
rect 9901 36628 9917 36692
rect 9981 36628 9997 36692
rect 10061 36628 10077 36692
rect 10141 36628 10157 36692
rect 10221 36628 10237 36692
rect 10301 36628 10317 36692
rect 10381 36628 10397 36692
rect 10461 36628 10477 36692
rect 10541 36628 10557 36692
rect 10621 36628 10637 36692
rect 10701 36628 10717 36692
rect 10781 36628 10786 36692
rect 9592 36611 10786 36628
rect 9592 36547 9597 36611
rect 9661 36547 9677 36611
rect 9741 36547 9757 36611
rect 9821 36547 9837 36611
rect 9901 36547 9917 36611
rect 9981 36547 9997 36611
rect 10061 36547 10077 36611
rect 10141 36547 10157 36611
rect 10221 36547 10237 36611
rect 10301 36547 10317 36611
rect 10381 36547 10397 36611
rect 10461 36547 10477 36611
rect 10541 36547 10557 36611
rect 10621 36547 10637 36611
rect 10701 36547 10717 36611
rect 10781 36547 10786 36611
rect 9592 36530 10786 36547
rect 9592 36466 9597 36530
rect 9661 36466 9677 36530
rect 9741 36466 9757 36530
rect 9821 36466 9837 36530
rect 9901 36466 9917 36530
rect 9981 36466 9997 36530
rect 10061 36466 10077 36530
rect 10141 36466 10157 36530
rect 10221 36466 10237 36530
rect 10301 36466 10317 36530
rect 10381 36466 10397 36530
rect 10461 36466 10477 36530
rect 10541 36466 10557 36530
rect 10621 36466 10637 36530
rect 10701 36466 10717 36530
rect 10781 36466 10786 36530
rect 9592 36449 10786 36466
rect 9592 36385 9597 36449
rect 9661 36385 9677 36449
rect 9741 36385 9757 36449
rect 9821 36385 9837 36449
rect 9901 36385 9917 36449
rect 9981 36385 9997 36449
rect 10061 36385 10077 36449
rect 10141 36385 10157 36449
rect 10221 36385 10237 36449
rect 10301 36385 10317 36449
rect 10381 36385 10397 36449
rect 10461 36385 10477 36449
rect 10541 36385 10557 36449
rect 10621 36385 10637 36449
rect 10701 36385 10717 36449
rect 10781 36385 10786 36449
rect 9592 36368 10786 36385
rect 9592 36304 9597 36368
rect 9661 36304 9677 36368
rect 9741 36304 9757 36368
rect 9821 36304 9837 36368
rect 9901 36304 9917 36368
rect 9981 36304 9997 36368
rect 10061 36304 10077 36368
rect 10141 36304 10157 36368
rect 10221 36304 10237 36368
rect 10301 36304 10317 36368
rect 10381 36304 10397 36368
rect 10461 36304 10477 36368
rect 10541 36304 10557 36368
rect 10621 36304 10637 36368
rect 10701 36304 10717 36368
rect 10781 36304 10786 36368
rect 9592 36287 10786 36304
rect 9592 36223 9597 36287
rect 9661 36223 9677 36287
rect 9741 36223 9757 36287
rect 9821 36223 9837 36287
rect 9901 36223 9917 36287
rect 9981 36223 9997 36287
rect 10061 36223 10077 36287
rect 10141 36223 10157 36287
rect 10221 36223 10237 36287
rect 10301 36223 10317 36287
rect 10381 36223 10397 36287
rect 10461 36223 10477 36287
rect 10541 36223 10557 36287
rect 10621 36223 10637 36287
rect 10701 36223 10717 36287
rect 10781 36223 10786 36287
rect 9592 36206 10786 36223
rect 9592 36142 9597 36206
rect 9661 36142 9677 36206
rect 9741 36142 9757 36206
rect 9821 36142 9837 36206
rect 9901 36142 9917 36206
rect 9981 36142 9997 36206
rect 10061 36142 10077 36206
rect 10141 36142 10157 36206
rect 10221 36142 10237 36206
rect 10301 36142 10317 36206
rect 10381 36142 10397 36206
rect 10461 36142 10477 36206
rect 10541 36142 10557 36206
rect 10621 36142 10637 36206
rect 10701 36142 10717 36206
rect 10781 36142 10786 36206
rect 9592 36124 10786 36142
rect 9592 36060 9597 36124
rect 9661 36060 9677 36124
rect 9741 36060 9757 36124
rect 9821 36060 9837 36124
rect 9901 36060 9917 36124
rect 9981 36060 9997 36124
rect 10061 36060 10077 36124
rect 10141 36060 10157 36124
rect 10221 36060 10237 36124
rect 10301 36060 10317 36124
rect 10381 36060 10397 36124
rect 10461 36060 10477 36124
rect 10541 36060 10557 36124
rect 10621 36060 10637 36124
rect 10701 36060 10717 36124
rect 10781 36060 10786 36124
rect 9592 36042 10786 36060
rect 9592 35978 9597 36042
rect 9661 35978 9677 36042
rect 9741 35978 9757 36042
rect 9821 35978 9837 36042
rect 9901 35978 9917 36042
rect 9981 35978 9997 36042
rect 10061 35978 10077 36042
rect 10141 35978 10157 36042
rect 10221 35978 10237 36042
rect 10301 35978 10317 36042
rect 10381 35978 10397 36042
rect 10461 35978 10477 36042
rect 10541 35978 10557 36042
rect 10621 35978 10637 36042
rect 10701 35978 10717 36042
rect 10781 35978 10786 36042
rect 9592 35960 10786 35978
rect 9592 35896 9597 35960
rect 9661 35896 9677 35960
rect 9741 35896 9757 35960
rect 9821 35896 9837 35960
rect 9901 35896 9917 35960
rect 9981 35896 9997 35960
rect 10061 35896 10077 35960
rect 10141 35896 10157 35960
rect 10221 35896 10237 35960
rect 10301 35896 10317 35960
rect 10381 35896 10397 35960
rect 10461 35896 10477 35960
rect 10541 35896 10557 35960
rect 10621 35896 10637 35960
rect 10701 35896 10717 35960
rect 10781 35896 10786 35960
rect 9592 35878 10786 35896
rect 9592 35814 9597 35878
rect 9661 35814 9677 35878
rect 9741 35814 9757 35878
rect 9821 35814 9837 35878
rect 9901 35814 9917 35878
rect 9981 35814 9997 35878
rect 10061 35814 10077 35878
rect 10141 35814 10157 35878
rect 10221 35814 10237 35878
rect 10301 35814 10317 35878
rect 10381 35814 10397 35878
rect 10461 35814 10477 35878
rect 10541 35814 10557 35878
rect 10621 35814 10637 35878
rect 10701 35814 10717 35878
rect 10781 35814 10786 35878
rect 9592 35796 10786 35814
rect 9592 35732 9597 35796
rect 9661 35732 9677 35796
rect 9741 35732 9757 35796
rect 9821 35732 9837 35796
rect 9901 35732 9917 35796
rect 9981 35732 9997 35796
rect 10061 35732 10077 35796
rect 10141 35732 10157 35796
rect 10221 35732 10237 35796
rect 10301 35732 10317 35796
rect 10381 35732 10397 35796
rect 10461 35732 10477 35796
rect 10541 35732 10557 35796
rect 10621 35732 10637 35796
rect 10701 35732 10717 35796
rect 10781 35732 10786 35796
rect 9592 35714 10786 35732
rect 9592 35650 9597 35714
rect 9661 35650 9677 35714
rect 9741 35650 9757 35714
rect 9821 35650 9837 35714
rect 9901 35650 9917 35714
rect 9981 35650 9997 35714
rect 10061 35650 10077 35714
rect 10141 35650 10157 35714
rect 10221 35650 10237 35714
rect 10301 35650 10317 35714
rect 10381 35650 10397 35714
rect 10461 35650 10477 35714
rect 10541 35650 10557 35714
rect 10621 35650 10637 35714
rect 10701 35650 10717 35714
rect 10781 35650 10786 35714
rect 9592 35632 10786 35650
rect 9592 35568 9597 35632
rect 9661 35568 9677 35632
rect 9741 35568 9757 35632
rect 9821 35568 9837 35632
rect 9901 35568 9917 35632
rect 9981 35568 9997 35632
rect 10061 35568 10077 35632
rect 10141 35568 10157 35632
rect 10221 35568 10237 35632
rect 10301 35568 10317 35632
rect 10381 35568 10397 35632
rect 10461 35568 10477 35632
rect 10541 35568 10557 35632
rect 10621 35568 10637 35632
rect 10701 35568 10717 35632
rect 10781 35568 10786 35632
rect 9592 35550 10786 35568
rect 9592 35486 9597 35550
rect 9661 35486 9677 35550
rect 9741 35486 9757 35550
rect 9821 35486 9837 35550
rect 9901 35486 9917 35550
rect 9981 35486 9997 35550
rect 10061 35486 10077 35550
rect 10141 35486 10157 35550
rect 10221 35486 10237 35550
rect 10301 35486 10317 35550
rect 10381 35486 10397 35550
rect 10461 35486 10477 35550
rect 10541 35486 10557 35550
rect 10621 35486 10637 35550
rect 10701 35486 10717 35550
rect 10781 35486 10786 35550
rect 9592 35468 10786 35486
rect 9592 35404 9597 35468
rect 9661 35404 9677 35468
rect 9741 35404 9757 35468
rect 9821 35404 9837 35468
rect 9901 35404 9917 35468
rect 9981 35404 9997 35468
rect 10061 35404 10077 35468
rect 10141 35404 10157 35468
rect 10221 35404 10237 35468
rect 10301 35404 10317 35468
rect 10381 35404 10397 35468
rect 10461 35404 10477 35468
rect 10541 35404 10557 35468
rect 10621 35404 10637 35468
rect 10701 35404 10717 35468
rect 10781 35404 10786 35468
rect 9592 35386 10786 35404
rect 9592 35322 9597 35386
rect 9661 35322 9677 35386
rect 9741 35322 9757 35386
rect 9821 35322 9837 35386
rect 9901 35322 9917 35386
rect 9981 35322 9997 35386
rect 10061 35322 10077 35386
rect 10141 35322 10157 35386
rect 10221 35322 10237 35386
rect 10301 35322 10317 35386
rect 10381 35322 10397 35386
rect 10461 35322 10477 35386
rect 10541 35322 10557 35386
rect 10621 35322 10637 35386
rect 10701 35322 10717 35386
rect 10781 35322 10786 35386
rect 9592 35304 10786 35322
rect 9592 35240 9597 35304
rect 9661 35240 9677 35304
rect 9741 35240 9757 35304
rect 9821 35240 9837 35304
rect 9901 35240 9917 35304
rect 9981 35240 9997 35304
rect 10061 35240 10077 35304
rect 10141 35240 10157 35304
rect 10221 35240 10237 35304
rect 10301 35240 10317 35304
rect 10381 35240 10397 35304
rect 10461 35240 10477 35304
rect 10541 35240 10557 35304
rect 10621 35240 10637 35304
rect 10701 35240 10717 35304
rect 10781 35240 10786 35304
rect 9592 35222 10786 35240
rect 9592 35158 9597 35222
rect 9661 35158 9677 35222
rect 9741 35158 9757 35222
rect 9821 35158 9837 35222
rect 9901 35158 9917 35222
rect 9981 35158 9997 35222
rect 10061 35158 10077 35222
rect 10141 35158 10157 35222
rect 10221 35158 10237 35222
rect 10301 35158 10317 35222
rect 10381 35158 10397 35222
rect 10461 35158 10477 35222
rect 10541 35158 10557 35222
rect 10621 35158 10637 35222
rect 10701 35158 10717 35222
rect 10781 35158 10786 35222
rect 9592 35157 10786 35158
rect 11093 39365 12287 39366
rect 11093 39301 11098 39365
rect 11162 39301 11178 39365
rect 11242 39301 11258 39365
rect 11322 39301 11338 39365
rect 11402 39301 11418 39365
rect 11482 39301 11498 39365
rect 11562 39301 11578 39365
rect 11642 39301 11658 39365
rect 11722 39301 11738 39365
rect 11802 39301 11818 39365
rect 11882 39301 11898 39365
rect 11962 39301 11978 39365
rect 12042 39301 12058 39365
rect 12122 39301 12138 39365
rect 12202 39301 12218 39365
rect 12282 39301 12287 39365
rect 11093 39284 12287 39301
rect 11093 39220 11098 39284
rect 11162 39220 11178 39284
rect 11242 39220 11258 39284
rect 11322 39220 11338 39284
rect 11402 39220 11418 39284
rect 11482 39220 11498 39284
rect 11562 39220 11578 39284
rect 11642 39220 11658 39284
rect 11722 39220 11738 39284
rect 11802 39220 11818 39284
rect 11882 39220 11898 39284
rect 11962 39220 11978 39284
rect 12042 39220 12058 39284
rect 12122 39220 12138 39284
rect 12202 39220 12218 39284
rect 12282 39220 12287 39284
rect 11093 39203 12287 39220
rect 11093 39139 11098 39203
rect 11162 39139 11178 39203
rect 11242 39139 11258 39203
rect 11322 39139 11338 39203
rect 11402 39139 11418 39203
rect 11482 39139 11498 39203
rect 11562 39139 11578 39203
rect 11642 39139 11658 39203
rect 11722 39139 11738 39203
rect 11802 39139 11818 39203
rect 11882 39139 11898 39203
rect 11962 39139 11978 39203
rect 12042 39139 12058 39203
rect 12122 39139 12138 39203
rect 12202 39139 12218 39203
rect 12282 39139 12287 39203
rect 11093 39122 12287 39139
rect 11093 39058 11098 39122
rect 11162 39058 11178 39122
rect 11242 39058 11258 39122
rect 11322 39058 11338 39122
rect 11402 39058 11418 39122
rect 11482 39058 11498 39122
rect 11562 39058 11578 39122
rect 11642 39058 11658 39122
rect 11722 39058 11738 39122
rect 11802 39058 11818 39122
rect 11882 39058 11898 39122
rect 11962 39058 11978 39122
rect 12042 39058 12058 39122
rect 12122 39058 12138 39122
rect 12202 39058 12218 39122
rect 12282 39058 12287 39122
rect 11093 39041 12287 39058
rect 11093 38977 11098 39041
rect 11162 38977 11178 39041
rect 11242 38977 11258 39041
rect 11322 38977 11338 39041
rect 11402 38977 11418 39041
rect 11482 38977 11498 39041
rect 11562 38977 11578 39041
rect 11642 38977 11658 39041
rect 11722 38977 11738 39041
rect 11802 38977 11818 39041
rect 11882 38977 11898 39041
rect 11962 38977 11978 39041
rect 12042 38977 12058 39041
rect 12122 38977 12138 39041
rect 12202 38977 12218 39041
rect 12282 38977 12287 39041
rect 11093 38960 12287 38977
rect 11093 38896 11098 38960
rect 11162 38896 11178 38960
rect 11242 38896 11258 38960
rect 11322 38896 11338 38960
rect 11402 38896 11418 38960
rect 11482 38896 11498 38960
rect 11562 38896 11578 38960
rect 11642 38896 11658 38960
rect 11722 38896 11738 38960
rect 11802 38896 11818 38960
rect 11882 38896 11898 38960
rect 11962 38896 11978 38960
rect 12042 38896 12058 38960
rect 12122 38896 12138 38960
rect 12202 38896 12218 38960
rect 12282 38896 12287 38960
rect 11093 38879 12287 38896
rect 11093 38815 11098 38879
rect 11162 38815 11178 38879
rect 11242 38815 11258 38879
rect 11322 38815 11338 38879
rect 11402 38815 11418 38879
rect 11482 38815 11498 38879
rect 11562 38815 11578 38879
rect 11642 38815 11658 38879
rect 11722 38815 11738 38879
rect 11802 38815 11818 38879
rect 11882 38815 11898 38879
rect 11962 38815 11978 38879
rect 12042 38815 12058 38879
rect 12122 38815 12138 38879
rect 12202 38815 12218 38879
rect 12282 38815 12287 38879
rect 11093 38798 12287 38815
rect 11093 38734 11098 38798
rect 11162 38734 11178 38798
rect 11242 38734 11258 38798
rect 11322 38734 11338 38798
rect 11402 38734 11418 38798
rect 11482 38734 11498 38798
rect 11562 38734 11578 38798
rect 11642 38734 11658 38798
rect 11722 38734 11738 38798
rect 11802 38734 11818 38798
rect 11882 38734 11898 38798
rect 11962 38734 11978 38798
rect 12042 38734 12058 38798
rect 12122 38734 12138 38798
rect 12202 38734 12218 38798
rect 12282 38734 12287 38798
rect 11093 38717 12287 38734
rect 11093 38653 11098 38717
rect 11162 38653 11178 38717
rect 11242 38653 11258 38717
rect 11322 38653 11338 38717
rect 11402 38653 11418 38717
rect 11482 38653 11498 38717
rect 11562 38653 11578 38717
rect 11642 38653 11658 38717
rect 11722 38653 11738 38717
rect 11802 38653 11818 38717
rect 11882 38653 11898 38717
rect 11962 38653 11978 38717
rect 12042 38653 12058 38717
rect 12122 38653 12138 38717
rect 12202 38653 12218 38717
rect 12282 38653 12287 38717
rect 11093 38636 12287 38653
rect 11093 38572 11098 38636
rect 11162 38572 11178 38636
rect 11242 38572 11258 38636
rect 11322 38572 11338 38636
rect 11402 38572 11418 38636
rect 11482 38572 11498 38636
rect 11562 38572 11578 38636
rect 11642 38572 11658 38636
rect 11722 38572 11738 38636
rect 11802 38572 11818 38636
rect 11882 38572 11898 38636
rect 11962 38572 11978 38636
rect 12042 38572 12058 38636
rect 12122 38572 12138 38636
rect 12202 38572 12218 38636
rect 12282 38572 12287 38636
rect 11093 38555 12287 38572
rect 11093 38491 11098 38555
rect 11162 38491 11178 38555
rect 11242 38491 11258 38555
rect 11322 38491 11338 38555
rect 11402 38491 11418 38555
rect 11482 38491 11498 38555
rect 11562 38491 11578 38555
rect 11642 38491 11658 38555
rect 11722 38491 11738 38555
rect 11802 38491 11818 38555
rect 11882 38491 11898 38555
rect 11962 38491 11978 38555
rect 12042 38491 12058 38555
rect 12122 38491 12138 38555
rect 12202 38491 12218 38555
rect 12282 38491 12287 38555
rect 11093 38474 12287 38491
rect 11093 38410 11098 38474
rect 11162 38410 11178 38474
rect 11242 38410 11258 38474
rect 11322 38410 11338 38474
rect 11402 38410 11418 38474
rect 11482 38410 11498 38474
rect 11562 38410 11578 38474
rect 11642 38410 11658 38474
rect 11722 38410 11738 38474
rect 11802 38410 11818 38474
rect 11882 38410 11898 38474
rect 11962 38410 11978 38474
rect 12042 38410 12058 38474
rect 12122 38410 12138 38474
rect 12202 38410 12218 38474
rect 12282 38410 12287 38474
rect 11093 38393 12287 38410
rect 11093 38329 11098 38393
rect 11162 38329 11178 38393
rect 11242 38329 11258 38393
rect 11322 38329 11338 38393
rect 11402 38329 11418 38393
rect 11482 38329 11498 38393
rect 11562 38329 11578 38393
rect 11642 38329 11658 38393
rect 11722 38329 11738 38393
rect 11802 38329 11818 38393
rect 11882 38329 11898 38393
rect 11962 38329 11978 38393
rect 12042 38329 12058 38393
rect 12122 38329 12138 38393
rect 12202 38329 12218 38393
rect 12282 38329 12287 38393
rect 11093 38312 12287 38329
rect 11093 38248 11098 38312
rect 11162 38248 11178 38312
rect 11242 38248 11258 38312
rect 11322 38248 11338 38312
rect 11402 38248 11418 38312
rect 11482 38248 11498 38312
rect 11562 38248 11578 38312
rect 11642 38248 11658 38312
rect 11722 38248 11738 38312
rect 11802 38248 11818 38312
rect 11882 38248 11898 38312
rect 11962 38248 11978 38312
rect 12042 38248 12058 38312
rect 12122 38248 12138 38312
rect 12202 38248 12218 38312
rect 12282 38248 12287 38312
rect 11093 38231 12287 38248
rect 11093 38167 11098 38231
rect 11162 38167 11178 38231
rect 11242 38167 11258 38231
rect 11322 38167 11338 38231
rect 11402 38167 11418 38231
rect 11482 38167 11498 38231
rect 11562 38167 11578 38231
rect 11642 38167 11658 38231
rect 11722 38167 11738 38231
rect 11802 38167 11818 38231
rect 11882 38167 11898 38231
rect 11962 38167 11978 38231
rect 12042 38167 12058 38231
rect 12122 38167 12138 38231
rect 12202 38167 12218 38231
rect 12282 38167 12287 38231
rect 11093 38150 12287 38167
rect 11093 38086 11098 38150
rect 11162 38086 11178 38150
rect 11242 38086 11258 38150
rect 11322 38086 11338 38150
rect 11402 38086 11418 38150
rect 11482 38086 11498 38150
rect 11562 38086 11578 38150
rect 11642 38086 11658 38150
rect 11722 38086 11738 38150
rect 11802 38086 11818 38150
rect 11882 38086 11898 38150
rect 11962 38086 11978 38150
rect 12042 38086 12058 38150
rect 12122 38086 12138 38150
rect 12202 38086 12218 38150
rect 12282 38086 12287 38150
rect 11093 38069 12287 38086
rect 11093 38005 11098 38069
rect 11162 38005 11178 38069
rect 11242 38005 11258 38069
rect 11322 38005 11338 38069
rect 11402 38005 11418 38069
rect 11482 38005 11498 38069
rect 11562 38005 11578 38069
rect 11642 38005 11658 38069
rect 11722 38005 11738 38069
rect 11802 38005 11818 38069
rect 11882 38005 11898 38069
rect 11962 38005 11978 38069
rect 12042 38005 12058 38069
rect 12122 38005 12138 38069
rect 12202 38005 12218 38069
rect 12282 38005 12287 38069
rect 11093 37988 12287 38005
rect 11093 37924 11098 37988
rect 11162 37924 11178 37988
rect 11242 37924 11258 37988
rect 11322 37924 11338 37988
rect 11402 37924 11418 37988
rect 11482 37924 11498 37988
rect 11562 37924 11578 37988
rect 11642 37924 11658 37988
rect 11722 37924 11738 37988
rect 11802 37924 11818 37988
rect 11882 37924 11898 37988
rect 11962 37924 11978 37988
rect 12042 37924 12058 37988
rect 12122 37924 12138 37988
rect 12202 37924 12218 37988
rect 12282 37924 12287 37988
rect 11093 37907 12287 37924
rect 11093 37843 11098 37907
rect 11162 37843 11178 37907
rect 11242 37843 11258 37907
rect 11322 37843 11338 37907
rect 11402 37843 11418 37907
rect 11482 37843 11498 37907
rect 11562 37843 11578 37907
rect 11642 37843 11658 37907
rect 11722 37843 11738 37907
rect 11802 37843 11818 37907
rect 11882 37843 11898 37907
rect 11962 37843 11978 37907
rect 12042 37843 12058 37907
rect 12122 37843 12138 37907
rect 12202 37843 12218 37907
rect 12282 37843 12287 37907
rect 11093 37826 12287 37843
rect 11093 37762 11098 37826
rect 11162 37762 11178 37826
rect 11242 37762 11258 37826
rect 11322 37762 11338 37826
rect 11402 37762 11418 37826
rect 11482 37762 11498 37826
rect 11562 37762 11578 37826
rect 11642 37762 11658 37826
rect 11722 37762 11738 37826
rect 11802 37762 11818 37826
rect 11882 37762 11898 37826
rect 11962 37762 11978 37826
rect 12042 37762 12058 37826
rect 12122 37762 12138 37826
rect 12202 37762 12218 37826
rect 12282 37762 12287 37826
rect 11093 37745 12287 37762
rect 11093 37681 11098 37745
rect 11162 37681 11178 37745
rect 11242 37681 11258 37745
rect 11322 37681 11338 37745
rect 11402 37681 11418 37745
rect 11482 37681 11498 37745
rect 11562 37681 11578 37745
rect 11642 37681 11658 37745
rect 11722 37681 11738 37745
rect 11802 37681 11818 37745
rect 11882 37681 11898 37745
rect 11962 37681 11978 37745
rect 12042 37681 12058 37745
rect 12122 37681 12138 37745
rect 12202 37681 12218 37745
rect 12282 37681 12287 37745
rect 11093 37664 12287 37681
rect 11093 37600 11098 37664
rect 11162 37600 11178 37664
rect 11242 37600 11258 37664
rect 11322 37600 11338 37664
rect 11402 37600 11418 37664
rect 11482 37600 11498 37664
rect 11562 37600 11578 37664
rect 11642 37600 11658 37664
rect 11722 37600 11738 37664
rect 11802 37600 11818 37664
rect 11882 37600 11898 37664
rect 11962 37600 11978 37664
rect 12042 37600 12058 37664
rect 12122 37600 12138 37664
rect 12202 37600 12218 37664
rect 12282 37600 12287 37664
rect 11093 37583 12287 37600
rect 11093 37519 11098 37583
rect 11162 37519 11178 37583
rect 11242 37519 11258 37583
rect 11322 37519 11338 37583
rect 11402 37519 11418 37583
rect 11482 37519 11498 37583
rect 11562 37519 11578 37583
rect 11642 37519 11658 37583
rect 11722 37519 11738 37583
rect 11802 37519 11818 37583
rect 11882 37519 11898 37583
rect 11962 37519 11978 37583
rect 12042 37519 12058 37583
rect 12122 37519 12138 37583
rect 12202 37519 12218 37583
rect 12282 37519 12287 37583
rect 11093 37502 12287 37519
rect 11093 37438 11098 37502
rect 11162 37438 11178 37502
rect 11242 37438 11258 37502
rect 11322 37438 11338 37502
rect 11402 37438 11418 37502
rect 11482 37438 11498 37502
rect 11562 37438 11578 37502
rect 11642 37438 11658 37502
rect 11722 37438 11738 37502
rect 11802 37438 11818 37502
rect 11882 37438 11898 37502
rect 11962 37438 11978 37502
rect 12042 37438 12058 37502
rect 12122 37438 12138 37502
rect 12202 37438 12218 37502
rect 12282 37438 12287 37502
rect 11093 37421 12287 37438
rect 11093 37357 11098 37421
rect 11162 37357 11178 37421
rect 11242 37357 11258 37421
rect 11322 37357 11338 37421
rect 11402 37357 11418 37421
rect 11482 37357 11498 37421
rect 11562 37357 11578 37421
rect 11642 37357 11658 37421
rect 11722 37357 11738 37421
rect 11802 37357 11818 37421
rect 11882 37357 11898 37421
rect 11962 37357 11978 37421
rect 12042 37357 12058 37421
rect 12122 37357 12138 37421
rect 12202 37357 12218 37421
rect 12282 37357 12287 37421
rect 11093 37340 12287 37357
rect 11093 37276 11098 37340
rect 11162 37276 11178 37340
rect 11242 37276 11258 37340
rect 11322 37276 11338 37340
rect 11402 37276 11418 37340
rect 11482 37276 11498 37340
rect 11562 37276 11578 37340
rect 11642 37276 11658 37340
rect 11722 37276 11738 37340
rect 11802 37276 11818 37340
rect 11882 37276 11898 37340
rect 11962 37276 11978 37340
rect 12042 37276 12058 37340
rect 12122 37276 12138 37340
rect 12202 37276 12218 37340
rect 12282 37276 12287 37340
rect 11093 37259 12287 37276
rect 11093 37195 11098 37259
rect 11162 37195 11178 37259
rect 11242 37195 11258 37259
rect 11322 37195 11338 37259
rect 11402 37195 11418 37259
rect 11482 37195 11498 37259
rect 11562 37195 11578 37259
rect 11642 37195 11658 37259
rect 11722 37195 11738 37259
rect 11802 37195 11818 37259
rect 11882 37195 11898 37259
rect 11962 37195 11978 37259
rect 12042 37195 12058 37259
rect 12122 37195 12138 37259
rect 12202 37195 12218 37259
rect 12282 37195 12287 37259
rect 11093 37178 12287 37195
rect 11093 37114 11098 37178
rect 11162 37114 11178 37178
rect 11242 37114 11258 37178
rect 11322 37114 11338 37178
rect 11402 37114 11418 37178
rect 11482 37114 11498 37178
rect 11562 37114 11578 37178
rect 11642 37114 11658 37178
rect 11722 37114 11738 37178
rect 11802 37114 11818 37178
rect 11882 37114 11898 37178
rect 11962 37114 11978 37178
rect 12042 37114 12058 37178
rect 12122 37114 12138 37178
rect 12202 37114 12218 37178
rect 12282 37114 12287 37178
rect 11093 37097 12287 37114
rect 11093 37033 11098 37097
rect 11162 37033 11178 37097
rect 11242 37033 11258 37097
rect 11322 37033 11338 37097
rect 11402 37033 11418 37097
rect 11482 37033 11498 37097
rect 11562 37033 11578 37097
rect 11642 37033 11658 37097
rect 11722 37033 11738 37097
rect 11802 37033 11818 37097
rect 11882 37033 11898 37097
rect 11962 37033 11978 37097
rect 12042 37033 12058 37097
rect 12122 37033 12138 37097
rect 12202 37033 12218 37097
rect 12282 37033 12287 37097
rect 11093 37016 12287 37033
rect 11093 36952 11098 37016
rect 11162 36952 11178 37016
rect 11242 36952 11258 37016
rect 11322 36952 11338 37016
rect 11402 36952 11418 37016
rect 11482 36952 11498 37016
rect 11562 36952 11578 37016
rect 11642 36952 11658 37016
rect 11722 36952 11738 37016
rect 11802 36952 11818 37016
rect 11882 36952 11898 37016
rect 11962 36952 11978 37016
rect 12042 36952 12058 37016
rect 12122 36952 12138 37016
rect 12202 36952 12218 37016
rect 12282 36952 12287 37016
rect 11093 36935 12287 36952
rect 11093 36871 11098 36935
rect 11162 36871 11178 36935
rect 11242 36871 11258 36935
rect 11322 36871 11338 36935
rect 11402 36871 11418 36935
rect 11482 36871 11498 36935
rect 11562 36871 11578 36935
rect 11642 36871 11658 36935
rect 11722 36871 11738 36935
rect 11802 36871 11818 36935
rect 11882 36871 11898 36935
rect 11962 36871 11978 36935
rect 12042 36871 12058 36935
rect 12122 36871 12138 36935
rect 12202 36871 12218 36935
rect 12282 36871 12287 36935
rect 11093 36854 12287 36871
rect 11093 36790 11098 36854
rect 11162 36790 11178 36854
rect 11242 36790 11258 36854
rect 11322 36790 11338 36854
rect 11402 36790 11418 36854
rect 11482 36790 11498 36854
rect 11562 36790 11578 36854
rect 11642 36790 11658 36854
rect 11722 36790 11738 36854
rect 11802 36790 11818 36854
rect 11882 36790 11898 36854
rect 11962 36790 11978 36854
rect 12042 36790 12058 36854
rect 12122 36790 12138 36854
rect 12202 36790 12218 36854
rect 12282 36790 12287 36854
rect 11093 36773 12287 36790
rect 11093 36709 11098 36773
rect 11162 36709 11178 36773
rect 11242 36709 11258 36773
rect 11322 36709 11338 36773
rect 11402 36709 11418 36773
rect 11482 36709 11498 36773
rect 11562 36709 11578 36773
rect 11642 36709 11658 36773
rect 11722 36709 11738 36773
rect 11802 36709 11818 36773
rect 11882 36709 11898 36773
rect 11962 36709 11978 36773
rect 12042 36709 12058 36773
rect 12122 36709 12138 36773
rect 12202 36709 12218 36773
rect 12282 36709 12287 36773
rect 11093 36692 12287 36709
rect 11093 36628 11098 36692
rect 11162 36628 11178 36692
rect 11242 36628 11258 36692
rect 11322 36628 11338 36692
rect 11402 36628 11418 36692
rect 11482 36628 11498 36692
rect 11562 36628 11578 36692
rect 11642 36628 11658 36692
rect 11722 36628 11738 36692
rect 11802 36628 11818 36692
rect 11882 36628 11898 36692
rect 11962 36628 11978 36692
rect 12042 36628 12058 36692
rect 12122 36628 12138 36692
rect 12202 36628 12218 36692
rect 12282 36628 12287 36692
rect 11093 36611 12287 36628
rect 11093 36547 11098 36611
rect 11162 36547 11178 36611
rect 11242 36547 11258 36611
rect 11322 36547 11338 36611
rect 11402 36547 11418 36611
rect 11482 36547 11498 36611
rect 11562 36547 11578 36611
rect 11642 36547 11658 36611
rect 11722 36547 11738 36611
rect 11802 36547 11818 36611
rect 11882 36547 11898 36611
rect 11962 36547 11978 36611
rect 12042 36547 12058 36611
rect 12122 36547 12138 36611
rect 12202 36547 12218 36611
rect 12282 36547 12287 36611
rect 11093 36530 12287 36547
rect 11093 36466 11098 36530
rect 11162 36466 11178 36530
rect 11242 36466 11258 36530
rect 11322 36466 11338 36530
rect 11402 36466 11418 36530
rect 11482 36466 11498 36530
rect 11562 36466 11578 36530
rect 11642 36466 11658 36530
rect 11722 36466 11738 36530
rect 11802 36466 11818 36530
rect 11882 36466 11898 36530
rect 11962 36466 11978 36530
rect 12042 36466 12058 36530
rect 12122 36466 12138 36530
rect 12202 36466 12218 36530
rect 12282 36466 12287 36530
rect 11093 36449 12287 36466
rect 11093 36385 11098 36449
rect 11162 36385 11178 36449
rect 11242 36385 11258 36449
rect 11322 36385 11338 36449
rect 11402 36385 11418 36449
rect 11482 36385 11498 36449
rect 11562 36385 11578 36449
rect 11642 36385 11658 36449
rect 11722 36385 11738 36449
rect 11802 36385 11818 36449
rect 11882 36385 11898 36449
rect 11962 36385 11978 36449
rect 12042 36385 12058 36449
rect 12122 36385 12138 36449
rect 12202 36385 12218 36449
rect 12282 36385 12287 36449
rect 11093 36368 12287 36385
rect 11093 36304 11098 36368
rect 11162 36304 11178 36368
rect 11242 36304 11258 36368
rect 11322 36304 11338 36368
rect 11402 36304 11418 36368
rect 11482 36304 11498 36368
rect 11562 36304 11578 36368
rect 11642 36304 11658 36368
rect 11722 36304 11738 36368
rect 11802 36304 11818 36368
rect 11882 36304 11898 36368
rect 11962 36304 11978 36368
rect 12042 36304 12058 36368
rect 12122 36304 12138 36368
rect 12202 36304 12218 36368
rect 12282 36304 12287 36368
rect 11093 36287 12287 36304
rect 11093 36223 11098 36287
rect 11162 36223 11178 36287
rect 11242 36223 11258 36287
rect 11322 36223 11338 36287
rect 11402 36223 11418 36287
rect 11482 36223 11498 36287
rect 11562 36223 11578 36287
rect 11642 36223 11658 36287
rect 11722 36223 11738 36287
rect 11802 36223 11818 36287
rect 11882 36223 11898 36287
rect 11962 36223 11978 36287
rect 12042 36223 12058 36287
rect 12122 36223 12138 36287
rect 12202 36223 12218 36287
rect 12282 36223 12287 36287
rect 11093 36206 12287 36223
rect 11093 36142 11098 36206
rect 11162 36142 11178 36206
rect 11242 36142 11258 36206
rect 11322 36142 11338 36206
rect 11402 36142 11418 36206
rect 11482 36142 11498 36206
rect 11562 36142 11578 36206
rect 11642 36142 11658 36206
rect 11722 36142 11738 36206
rect 11802 36142 11818 36206
rect 11882 36142 11898 36206
rect 11962 36142 11978 36206
rect 12042 36142 12058 36206
rect 12122 36142 12138 36206
rect 12202 36142 12218 36206
rect 12282 36142 12287 36206
rect 11093 36124 12287 36142
rect 11093 36060 11098 36124
rect 11162 36060 11178 36124
rect 11242 36060 11258 36124
rect 11322 36060 11338 36124
rect 11402 36060 11418 36124
rect 11482 36060 11498 36124
rect 11562 36060 11578 36124
rect 11642 36060 11658 36124
rect 11722 36060 11738 36124
rect 11802 36060 11818 36124
rect 11882 36060 11898 36124
rect 11962 36060 11978 36124
rect 12042 36060 12058 36124
rect 12122 36060 12138 36124
rect 12202 36060 12218 36124
rect 12282 36060 12287 36124
rect 11093 36042 12287 36060
rect 11093 35978 11098 36042
rect 11162 35978 11178 36042
rect 11242 35978 11258 36042
rect 11322 35978 11338 36042
rect 11402 35978 11418 36042
rect 11482 35978 11498 36042
rect 11562 35978 11578 36042
rect 11642 35978 11658 36042
rect 11722 35978 11738 36042
rect 11802 35978 11818 36042
rect 11882 35978 11898 36042
rect 11962 35978 11978 36042
rect 12042 35978 12058 36042
rect 12122 35978 12138 36042
rect 12202 35978 12218 36042
rect 12282 35978 12287 36042
rect 11093 35960 12287 35978
rect 11093 35896 11098 35960
rect 11162 35896 11178 35960
rect 11242 35896 11258 35960
rect 11322 35896 11338 35960
rect 11402 35896 11418 35960
rect 11482 35896 11498 35960
rect 11562 35896 11578 35960
rect 11642 35896 11658 35960
rect 11722 35896 11738 35960
rect 11802 35896 11818 35960
rect 11882 35896 11898 35960
rect 11962 35896 11978 35960
rect 12042 35896 12058 35960
rect 12122 35896 12138 35960
rect 12202 35896 12218 35960
rect 12282 35896 12287 35960
rect 12586 39308 12588 39372
rect 12652 39308 12676 39372
rect 12740 39308 12764 39372
rect 12828 39308 12852 39372
rect 12916 39308 12940 39372
rect 13004 39308 13006 39372
rect 12586 39292 13006 39308
rect 12586 39228 12588 39292
rect 12652 39228 12676 39292
rect 12740 39228 12764 39292
rect 12828 39228 12852 39292
rect 12916 39228 12940 39292
rect 13004 39228 13006 39292
rect 12586 39212 13006 39228
rect 12586 39148 12588 39212
rect 12652 39148 12676 39212
rect 12740 39148 12764 39212
rect 12828 39148 12852 39212
rect 12916 39148 12940 39212
rect 13004 39148 13006 39212
rect 12586 39132 13006 39148
rect 12586 39068 12588 39132
rect 12652 39068 12676 39132
rect 12740 39068 12764 39132
rect 12828 39068 12852 39132
rect 12916 39068 12940 39132
rect 13004 39068 13006 39132
rect 12586 39052 13006 39068
rect 12586 38988 12588 39052
rect 12652 38988 12676 39052
rect 12740 38988 12764 39052
rect 12828 38988 12852 39052
rect 12916 38988 12940 39052
rect 13004 38988 13006 39052
rect 12586 38972 13006 38988
rect 12586 38908 12588 38972
rect 12652 38908 12676 38972
rect 12740 38908 12764 38972
rect 12828 38908 12852 38972
rect 12916 38908 12940 38972
rect 13004 38908 13006 38972
rect 12586 38892 13006 38908
rect 12586 38828 12588 38892
rect 12652 38828 12676 38892
rect 12740 38828 12764 38892
rect 12828 38828 12852 38892
rect 12916 38828 12940 38892
rect 13004 38828 13006 38892
rect 12586 38812 13006 38828
rect 12586 38748 12588 38812
rect 12652 38748 12676 38812
rect 12740 38748 12764 38812
rect 12828 38748 12852 38812
rect 12916 38748 12940 38812
rect 13004 38748 13006 38812
rect 12586 38731 13006 38748
rect 12586 38667 12588 38731
rect 12652 38667 12676 38731
rect 12740 38667 12764 38731
rect 12828 38667 12852 38731
rect 12916 38667 12940 38731
rect 13004 38667 13006 38731
rect 12586 38650 13006 38667
rect 12586 38586 12588 38650
rect 12652 38586 12676 38650
rect 12740 38586 12764 38650
rect 12828 38586 12852 38650
rect 12916 38586 12940 38650
rect 13004 38586 13006 38650
rect 12586 38569 13006 38586
rect 12586 38505 12588 38569
rect 12652 38505 12676 38569
rect 12740 38505 12764 38569
rect 12828 38505 12852 38569
rect 12916 38505 12940 38569
rect 13004 38505 13006 38569
rect 12586 38488 13006 38505
rect 12586 38424 12588 38488
rect 12652 38424 12676 38488
rect 12740 38424 12764 38488
rect 12828 38424 12852 38488
rect 12916 38424 12940 38488
rect 13004 38424 13006 38488
rect 12586 38407 13006 38424
rect 12586 38343 12588 38407
rect 12652 38343 12676 38407
rect 12740 38343 12764 38407
rect 12828 38343 12852 38407
rect 12916 38343 12940 38407
rect 13004 38343 13006 38407
rect 12586 38326 13006 38343
rect 12586 38262 12588 38326
rect 12652 38262 12676 38326
rect 12740 38262 12764 38326
rect 12828 38262 12852 38326
rect 12916 38262 12940 38326
rect 13004 38262 13006 38326
rect 12586 38245 13006 38262
rect 12586 38181 12588 38245
rect 12652 38181 12676 38245
rect 12740 38181 12764 38245
rect 12828 38181 12852 38245
rect 12916 38181 12940 38245
rect 13004 38181 13006 38245
rect 12586 38164 13006 38181
rect 12586 38100 12588 38164
rect 12652 38100 12676 38164
rect 12740 38100 12764 38164
rect 12828 38100 12852 38164
rect 12916 38100 12940 38164
rect 13004 38100 13006 38164
rect 12586 38083 13006 38100
rect 12586 38019 12588 38083
rect 12652 38019 12676 38083
rect 12740 38019 12764 38083
rect 12828 38019 12852 38083
rect 12916 38019 12940 38083
rect 13004 38019 13006 38083
rect 12586 38002 13006 38019
rect 12586 37938 12588 38002
rect 12652 37938 12676 38002
rect 12740 37938 12764 38002
rect 12828 37938 12852 38002
rect 12916 37938 12940 38002
rect 13004 37938 13006 38002
rect 12586 37921 13006 37938
rect 12586 37857 12588 37921
rect 12652 37857 12676 37921
rect 12740 37857 12764 37921
rect 12828 37857 12852 37921
rect 12916 37857 12940 37921
rect 13004 37857 13006 37921
rect 12586 37840 13006 37857
rect 12586 37776 12588 37840
rect 12652 37776 12676 37840
rect 12740 37776 12764 37840
rect 12828 37776 12852 37840
rect 12916 37776 12940 37840
rect 13004 37776 13006 37840
rect 12586 37759 13006 37776
rect 12586 37695 12588 37759
rect 12652 37695 12676 37759
rect 12740 37695 12764 37759
rect 12828 37695 12852 37759
rect 12916 37695 12940 37759
rect 13004 37695 13006 37759
rect 12586 37678 13006 37695
rect 12586 37614 12588 37678
rect 12652 37614 12676 37678
rect 12740 37614 12764 37678
rect 12828 37614 12852 37678
rect 12916 37614 12940 37678
rect 13004 37614 13006 37678
rect 12586 37597 13006 37614
rect 12586 37533 12588 37597
rect 12652 37533 12676 37597
rect 12740 37533 12764 37597
rect 12828 37533 12852 37597
rect 12916 37533 12940 37597
rect 13004 37533 13006 37597
rect 12586 37516 13006 37533
rect 12586 37452 12588 37516
rect 12652 37452 12676 37516
rect 12740 37452 12764 37516
rect 12828 37452 12852 37516
rect 12916 37452 12940 37516
rect 13004 37452 13006 37516
rect 12586 37435 13006 37452
rect 12586 37371 12588 37435
rect 12652 37371 12676 37435
rect 12740 37371 12764 37435
rect 12828 37371 12852 37435
rect 12916 37371 12940 37435
rect 13004 37371 13006 37435
rect 12586 37354 13006 37371
rect 12586 37290 12588 37354
rect 12652 37290 12676 37354
rect 12740 37290 12764 37354
rect 12828 37290 12852 37354
rect 12916 37290 12940 37354
rect 13004 37290 13006 37354
rect 12586 37273 13006 37290
rect 12586 37209 12588 37273
rect 12652 37209 12676 37273
rect 12740 37209 12764 37273
rect 12828 37209 12852 37273
rect 12916 37209 12940 37273
rect 13004 37209 13006 37273
rect 12586 37192 13006 37209
rect 12586 37128 12588 37192
rect 12652 37128 12676 37192
rect 12740 37128 12764 37192
rect 12828 37128 12852 37192
rect 12916 37128 12940 37192
rect 13004 37128 13006 37192
rect 12586 37111 13006 37128
rect 12586 37047 12588 37111
rect 12652 37047 12676 37111
rect 12740 37047 12764 37111
rect 12828 37047 12852 37111
rect 12916 37047 12940 37111
rect 13004 37047 13006 37111
rect 12586 37030 13006 37047
rect 12586 36966 12588 37030
rect 12652 36966 12676 37030
rect 12740 36966 12764 37030
rect 12828 36966 12852 37030
rect 12916 36966 12940 37030
rect 13004 36966 13006 37030
rect 12586 36949 13006 36966
rect 12586 36885 12588 36949
rect 12652 36885 12676 36949
rect 12740 36885 12764 36949
rect 12828 36885 12852 36949
rect 12916 36885 12940 36949
rect 13004 36885 13006 36949
rect 12586 36868 13006 36885
rect 12586 36804 12588 36868
rect 12652 36804 12676 36868
rect 12740 36804 12764 36868
rect 12828 36804 12852 36868
rect 12916 36804 12940 36868
rect 13004 36804 13006 36868
rect 12586 36787 13006 36804
rect 12586 36723 12588 36787
rect 12652 36723 12676 36787
rect 12740 36723 12764 36787
rect 12828 36723 12852 36787
rect 12916 36723 12940 36787
rect 13004 36723 13006 36787
rect 12586 36706 13006 36723
rect 12586 36642 12588 36706
rect 12652 36642 12676 36706
rect 12740 36642 12764 36706
rect 12828 36642 12852 36706
rect 12916 36642 12940 36706
rect 13004 36642 13006 36706
rect 12586 36625 13006 36642
rect 12586 36561 12588 36625
rect 12652 36561 12676 36625
rect 12740 36561 12764 36625
rect 12828 36561 12852 36625
rect 12916 36561 12940 36625
rect 13004 36561 13006 36625
rect 12586 36544 13006 36561
rect 12586 36480 12588 36544
rect 12652 36480 12676 36544
rect 12740 36480 12764 36544
rect 12828 36480 12852 36544
rect 12916 36480 12940 36544
rect 13004 36480 13006 36544
rect 12586 36463 13006 36480
rect 12586 36399 12588 36463
rect 12652 36399 12676 36463
rect 12740 36399 12764 36463
rect 12828 36399 12852 36463
rect 12916 36399 12940 36463
rect 13004 36399 13006 36463
rect 12586 36382 13006 36399
rect 12586 36318 12588 36382
rect 12652 36318 12676 36382
rect 12740 36318 12764 36382
rect 12828 36318 12852 36382
rect 12916 36318 12940 36382
rect 13004 36318 13006 36382
rect 12586 36301 13006 36318
rect 12586 36237 12588 36301
rect 12652 36237 12676 36301
rect 12740 36237 12764 36301
rect 12828 36237 12852 36301
rect 12916 36237 12940 36301
rect 13004 36237 13006 36301
rect 12586 36220 13006 36237
rect 12586 36156 12588 36220
rect 12652 36156 12676 36220
rect 12740 36156 12764 36220
rect 12828 36156 12852 36220
rect 12916 36156 12940 36220
rect 13004 36156 13006 36220
rect 12586 36139 13006 36156
rect 12586 36075 12588 36139
rect 12652 36075 12676 36139
rect 12740 36075 12764 36139
rect 12828 36075 12852 36139
rect 12916 36075 12940 36139
rect 13004 36075 13006 36139
rect 12586 36058 13006 36075
rect 12586 35994 12588 36058
rect 12652 35994 12676 36058
rect 12740 35994 12764 36058
rect 12828 35994 12852 36058
rect 12916 35994 12940 36058
rect 13004 35994 13006 36058
rect 12586 35977 13006 35994
rect 12586 35913 12588 35977
rect 12652 35913 12676 35977
rect 12740 35913 12764 35977
rect 12828 35913 12852 35977
rect 12916 35913 12940 35977
rect 13004 35913 13006 35977
rect 12586 35912 13006 35913
rect 11093 35878 12287 35896
rect 11093 35814 11098 35878
rect 11162 35814 11178 35878
rect 11242 35814 11258 35878
rect 11322 35814 11338 35878
rect 11402 35814 11418 35878
rect 11482 35814 11498 35878
rect 11562 35814 11578 35878
rect 11642 35814 11658 35878
rect 11722 35814 11738 35878
rect 11802 35814 11818 35878
rect 11882 35814 11898 35878
rect 11962 35814 11978 35878
rect 12042 35814 12058 35878
rect 12122 35814 12138 35878
rect 12202 35814 12218 35878
rect 12282 35814 12287 35878
rect 11093 35796 12287 35814
rect 11093 35732 11098 35796
rect 11162 35732 11178 35796
rect 11242 35732 11258 35796
rect 11322 35732 11338 35796
rect 11402 35732 11418 35796
rect 11482 35732 11498 35796
rect 11562 35732 11578 35796
rect 11642 35732 11658 35796
rect 11722 35732 11738 35796
rect 11802 35732 11818 35796
rect 11882 35732 11898 35796
rect 11962 35732 11978 35796
rect 12042 35732 12058 35796
rect 12122 35732 12138 35796
rect 12202 35732 12218 35796
rect 12282 35732 12287 35796
rect 11093 35714 12287 35732
rect 11093 35650 11098 35714
rect 11162 35650 11178 35714
rect 11242 35650 11258 35714
rect 11322 35650 11338 35714
rect 11402 35650 11418 35714
rect 11482 35650 11498 35714
rect 11562 35650 11578 35714
rect 11642 35650 11658 35714
rect 11722 35650 11738 35714
rect 11802 35650 11818 35714
rect 11882 35650 11898 35714
rect 11962 35650 11978 35714
rect 12042 35650 12058 35714
rect 12122 35650 12138 35714
rect 12202 35650 12218 35714
rect 12282 35650 12287 35714
rect 11093 35632 12287 35650
rect 11093 35568 11098 35632
rect 11162 35568 11178 35632
rect 11242 35568 11258 35632
rect 11322 35568 11338 35632
rect 11402 35568 11418 35632
rect 11482 35568 11498 35632
rect 11562 35568 11578 35632
rect 11642 35568 11658 35632
rect 11722 35568 11738 35632
rect 11802 35568 11818 35632
rect 11882 35568 11898 35632
rect 11962 35568 11978 35632
rect 12042 35568 12058 35632
rect 12122 35568 12138 35632
rect 12202 35568 12218 35632
rect 12282 35568 12287 35632
rect 11093 35550 12287 35568
rect 11093 35486 11098 35550
rect 11162 35486 11178 35550
rect 11242 35486 11258 35550
rect 11322 35486 11338 35550
rect 11402 35486 11418 35550
rect 11482 35486 11498 35550
rect 11562 35486 11578 35550
rect 11642 35486 11658 35550
rect 11722 35486 11738 35550
rect 11802 35486 11818 35550
rect 11882 35486 11898 35550
rect 11962 35486 11978 35550
rect 12042 35486 12058 35550
rect 12122 35486 12138 35550
rect 12202 35486 12218 35550
rect 12282 35486 12287 35550
rect 11093 35468 12287 35486
rect 11093 35404 11098 35468
rect 11162 35404 11178 35468
rect 11242 35404 11258 35468
rect 11322 35404 11338 35468
rect 11402 35404 11418 35468
rect 11482 35404 11498 35468
rect 11562 35404 11578 35468
rect 11642 35404 11658 35468
rect 11722 35404 11738 35468
rect 11802 35404 11818 35468
rect 11882 35404 11898 35468
rect 11962 35404 11978 35468
rect 12042 35404 12058 35468
rect 12122 35404 12138 35468
rect 12202 35404 12218 35468
rect 12282 35404 12287 35468
rect 11093 35386 12287 35404
rect 11093 35322 11098 35386
rect 11162 35322 11178 35386
rect 11242 35322 11258 35386
rect 11322 35322 11338 35386
rect 11402 35322 11418 35386
rect 11482 35322 11498 35386
rect 11562 35322 11578 35386
rect 11642 35322 11658 35386
rect 11722 35322 11738 35386
rect 11802 35322 11818 35386
rect 11882 35322 11898 35386
rect 11962 35322 11978 35386
rect 12042 35322 12058 35386
rect 12122 35322 12138 35386
rect 12202 35322 12218 35386
rect 12282 35322 12287 35386
rect 12597 35851 13247 35852
rect 12597 35787 12598 35851
rect 12662 35787 12682 35851
rect 12746 35787 12766 35851
rect 12830 35787 12850 35851
rect 12914 35787 12933 35851
rect 12997 35787 13016 35851
rect 13080 35787 13099 35851
rect 13163 35787 13182 35851
rect 13246 35787 13247 35851
rect 12597 35767 13247 35787
rect 12597 35703 12598 35767
rect 12662 35703 12682 35767
rect 12746 35703 12766 35767
rect 12830 35703 12850 35767
rect 12914 35703 12933 35767
rect 12997 35703 13016 35767
rect 13080 35703 13099 35767
rect 13163 35703 13182 35767
rect 13246 35703 13247 35767
rect 12597 35683 13247 35703
rect 12597 35619 12598 35683
rect 12662 35619 12682 35683
rect 12746 35619 12766 35683
rect 12830 35619 12850 35683
rect 12914 35619 12933 35683
rect 12997 35619 13016 35683
rect 13080 35619 13099 35683
rect 13163 35619 13182 35683
rect 13246 35619 13247 35683
rect 12597 35599 13247 35619
rect 12597 35535 12598 35599
rect 12662 35535 12682 35599
rect 12746 35535 12766 35599
rect 12830 35535 12850 35599
rect 12914 35535 12933 35599
rect 12997 35535 13016 35599
rect 13080 35535 13099 35599
rect 13163 35535 13182 35599
rect 13246 35535 13247 35599
rect 12597 35515 13247 35535
rect 12597 35451 12598 35515
rect 12662 35451 12682 35515
rect 12746 35451 12766 35515
rect 12830 35451 12850 35515
rect 12914 35451 12933 35515
rect 12997 35451 13016 35515
rect 13080 35451 13099 35515
rect 13163 35451 13182 35515
rect 13246 35451 13247 35515
rect 12597 35431 13247 35451
rect 12597 35367 12598 35431
rect 12662 35367 12682 35431
rect 12746 35367 12766 35431
rect 12830 35367 12850 35431
rect 12914 35367 12933 35431
rect 12997 35367 13016 35431
rect 13080 35367 13099 35431
rect 13163 35367 13182 35431
rect 13246 35367 13247 35431
rect 12597 35366 13247 35367
rect 11093 35304 12287 35322
rect 11093 35240 11098 35304
rect 11162 35240 11178 35304
rect 11242 35240 11258 35304
rect 11322 35240 11338 35304
rect 11402 35240 11418 35304
rect 11482 35240 11498 35304
rect 11562 35240 11578 35304
rect 11642 35240 11658 35304
rect 11722 35240 11738 35304
rect 11802 35240 11818 35304
rect 11882 35240 11898 35304
rect 11962 35240 11978 35304
rect 12042 35240 12058 35304
rect 12122 35240 12138 35304
rect 12202 35240 12218 35304
rect 12282 35240 12287 35304
rect 11093 35222 12287 35240
rect 11093 35158 11098 35222
rect 11162 35158 11178 35222
rect 11242 35158 11258 35222
rect 11322 35158 11338 35222
rect 11402 35158 11418 35222
rect 11482 35158 11498 35222
rect 11562 35158 11578 35222
rect 11642 35158 11658 35222
rect 11722 35158 11738 35222
rect 11802 35158 11818 35222
rect 11882 35158 11898 35222
rect 11962 35158 11978 35222
rect 12042 35158 12058 35222
rect 12122 35158 12138 35222
rect 12202 35158 12218 35222
rect 12282 35158 12287 35222
rect 11093 35157 12287 35158
rect 15746 35157 16000 40000
rect 4082 34681 4718 34684
rect 4082 34617 4083 34681
rect 4147 34617 4165 34681
rect 4229 34617 4247 34681
rect 4311 34617 4329 34681
rect 4393 34617 4410 34681
rect 4474 34617 4491 34681
rect 4555 34617 4572 34681
rect 4636 34617 4653 34681
rect 4717 34617 4718 34681
rect 4082 34593 4718 34617
rect 4082 34529 4083 34593
rect 4147 34529 4165 34593
rect 4229 34529 4247 34593
rect 4311 34529 4329 34593
rect 4393 34529 4410 34593
rect 4474 34529 4491 34593
rect 4555 34529 4572 34593
rect 4636 34529 4653 34593
rect 4717 34529 4718 34593
rect 4082 34505 4718 34529
rect 4082 34441 4083 34505
rect 4147 34441 4165 34505
rect 4229 34441 4247 34505
rect 4311 34441 4329 34505
rect 4393 34441 4410 34505
rect 4474 34441 4491 34505
rect 4555 34441 4572 34505
rect 4636 34441 4653 34505
rect 4717 34441 4718 34505
rect 4082 34417 4718 34441
rect 4082 34353 4083 34417
rect 4147 34353 4165 34417
rect 4229 34353 4247 34417
rect 4311 34353 4329 34417
rect 4393 34353 4410 34417
rect 4474 34353 4491 34417
rect 4555 34353 4572 34417
rect 4636 34353 4653 34417
rect 4717 34353 4718 34417
rect 4082 34329 4718 34353
rect 4082 34265 4083 34329
rect 4147 34265 4165 34329
rect 4229 34265 4247 34329
rect 4311 34265 4329 34329
rect 4393 34265 4410 34329
rect 4474 34265 4491 34329
rect 4555 34265 4572 34329
rect 4636 34265 4653 34329
rect 4717 34265 4718 34329
rect 4082 34241 4718 34265
rect 4082 34177 4083 34241
rect 4147 34177 4165 34241
rect 4229 34177 4247 34241
rect 4311 34177 4329 34241
rect 4393 34177 4410 34241
rect 4474 34177 4491 34241
rect 4555 34177 4572 34241
rect 4636 34177 4653 34241
rect 4717 34177 4718 34241
rect 4082 34174 4718 34177
tri 15029 31179 15299 31449 sw
rect 14501 31178 15299 31179
rect 2131 31167 2497 31168
rect 2131 31103 2132 31167
rect 2196 31103 2232 31167
rect 2296 31103 2332 31167
rect 2396 31103 2432 31167
rect 2496 31103 2497 31167
rect 2131 31085 2497 31103
rect 2131 31021 2132 31085
rect 2196 31021 2232 31085
rect 2296 31021 2332 31085
rect 2396 31021 2432 31085
rect 2496 31021 2497 31085
rect 2131 31003 2497 31021
rect 2131 30939 2132 31003
rect 2196 30939 2232 31003
rect 2296 30939 2332 31003
rect 2396 30939 2432 31003
rect 2496 30939 2497 31003
rect 2131 30921 2497 30939
rect 2131 30857 2132 30921
rect 2196 30857 2232 30921
rect 2296 30857 2332 30921
rect 2396 30857 2432 30921
rect 2496 30857 2497 30921
rect 2131 30839 2497 30857
rect 2131 30775 2132 30839
rect 2196 30775 2232 30839
rect 2296 30775 2332 30839
rect 2396 30775 2432 30839
rect 2496 30775 2497 30839
rect 2131 30757 2497 30775
rect 2131 30693 2132 30757
rect 2196 30693 2232 30757
rect 2296 30693 2332 30757
rect 2396 30693 2432 30757
rect 2496 30693 2497 30757
rect 2131 30675 2497 30693
rect 2131 30611 2132 30675
rect 2196 30611 2232 30675
rect 2296 30611 2332 30675
rect 2396 30611 2432 30675
rect 2496 30611 2497 30675
rect 2131 30593 2497 30611
rect 2131 30529 2132 30593
rect 2196 30529 2232 30593
rect 2296 30529 2332 30593
rect 2396 30529 2432 30593
rect 2496 30529 2497 30593
rect 2131 30511 2497 30529
rect 2131 30447 2132 30511
rect 2196 30447 2232 30511
rect 2296 30447 2332 30511
rect 2396 30447 2432 30511
rect 2496 30447 2497 30511
rect 2131 30429 2497 30447
rect 2131 30365 2132 30429
rect 2196 30365 2232 30429
rect 2296 30365 2332 30429
rect 2396 30365 2432 30429
rect 2496 30365 2497 30429
rect 2131 30347 2497 30365
rect 2131 30283 2132 30347
rect 2196 30283 2232 30347
rect 2296 30283 2332 30347
rect 2396 30283 2432 30347
rect 2496 30283 2497 30347
rect 2131 30264 2497 30283
rect 2131 30200 2132 30264
rect 2196 30200 2232 30264
rect 2296 30200 2332 30264
rect 2396 30200 2432 30264
rect 2496 30200 2497 30264
rect 2131 30181 2497 30200
rect 2131 30117 2132 30181
rect 2196 30117 2232 30181
rect 2296 30117 2332 30181
rect 2396 30117 2432 30181
rect 2496 30117 2497 30181
rect 2131 30098 2497 30117
rect 2131 30034 2132 30098
rect 2196 30034 2232 30098
rect 2296 30034 2332 30098
rect 2396 30034 2432 30098
rect 2496 30034 2497 30098
rect 2131 30015 2497 30034
rect 2131 29951 2132 30015
rect 2196 29951 2232 30015
rect 2296 29951 2332 30015
rect 2396 29951 2432 30015
rect 2496 29951 2497 30015
rect 2131 29932 2497 29951
rect 2131 29868 2132 29932
rect 2196 29868 2232 29932
rect 2296 29868 2332 29932
rect 2396 29868 2432 29932
rect 2496 29868 2497 29932
rect 2131 29849 2497 29868
rect 2131 29785 2132 29849
rect 2196 29785 2232 29849
rect 2296 29785 2332 29849
rect 2396 29785 2432 29849
rect 2496 29785 2497 29849
rect 2131 29766 2497 29785
rect 2131 29702 2132 29766
rect 2196 29702 2232 29766
rect 2296 29702 2332 29766
rect 2396 29702 2432 29766
rect 2496 29702 2497 29766
rect 2131 29683 2497 29702
rect 2131 29619 2132 29683
rect 2196 29619 2232 29683
rect 2296 29619 2332 29683
rect 2396 29619 2432 29683
rect 2496 29619 2497 29683
rect 2131 29600 2497 29619
rect 2131 29536 2132 29600
rect 2196 29536 2232 29600
rect 2296 29536 2332 29600
rect 2396 29536 2432 29600
rect 2496 29536 2497 29600
rect 2131 29517 2497 29536
rect 2131 29453 2132 29517
rect 2196 29453 2232 29517
rect 2296 29453 2332 29517
rect 2396 29453 2432 29517
rect 2496 29453 2497 29517
rect 2131 29434 2497 29453
rect 2131 29370 2132 29434
rect 2196 29370 2232 29434
rect 2296 29370 2332 29434
rect 2396 29370 2432 29434
rect 2496 29370 2497 29434
rect 2131 29351 2497 29370
rect 2131 29287 2132 29351
rect 2196 29287 2232 29351
rect 2296 29287 2332 29351
rect 2396 29287 2432 29351
rect 2496 29287 2497 29351
rect 2131 29268 2497 29287
rect 2131 29204 2132 29268
rect 2196 29204 2232 29268
rect 2296 29204 2332 29268
rect 2396 29204 2432 29268
rect 2496 29204 2497 29268
rect 2131 29185 2497 29204
rect 2131 29121 2132 29185
rect 2196 29121 2232 29185
rect 2296 29121 2332 29185
rect 2396 29121 2432 29185
rect 2496 29121 2497 29185
rect 2131 29102 2497 29121
rect 2131 29038 2132 29102
rect 2196 29038 2232 29102
rect 2296 29038 2332 29102
rect 2396 29038 2432 29102
rect 2496 29038 2497 29102
rect 2131 29019 2497 29038
rect 2131 28955 2132 29019
rect 2196 28955 2232 29019
rect 2296 28955 2332 29019
rect 2396 28955 2432 29019
rect 2496 28955 2497 29019
rect 2131 28936 2497 28955
rect 2131 28872 2132 28936
rect 2196 28872 2232 28936
rect 2296 28872 2332 28936
rect 2396 28872 2432 28936
rect 2496 28872 2497 28936
rect 2131 28871 2497 28872
rect 14501 29034 14508 31178
rect 15292 29034 15299 31178
rect 14501 29017 15299 29034
rect 14501 28953 14508 29017
rect 14572 28953 14588 29017
rect 14652 28953 14668 29017
rect 14732 28953 14748 29017
rect 14812 28953 14828 29017
rect 14892 28953 14908 29017
rect 14972 28953 14988 29017
rect 15052 28953 15068 29017
rect 15132 28953 15148 29017
rect 15212 28953 15228 29017
rect 15292 28953 15299 29017
rect 14501 28936 15299 28953
rect 14501 28872 14508 28936
rect 14572 28872 14588 28936
rect 14652 28872 14668 28936
rect 14732 28872 14748 28936
rect 14812 28872 14828 28936
rect 14892 28872 14908 28936
rect 14972 28872 14988 28936
rect 15052 28872 15068 28936
rect 15132 28872 15148 28936
rect 15212 28872 15228 28936
rect 15292 28872 15299 28936
rect 14501 28871 15299 28872
tri 15029 28601 15299 28871 nw
rect 14516 27593 15040 27594
rect 14516 27529 14521 27593
rect 14585 27529 14611 27593
rect 14675 27529 14701 27593
rect 14765 27529 14791 27593
rect 14855 27529 14881 27593
rect 14945 27529 14971 27593
rect 15035 27529 15040 27593
rect 14516 27512 15040 27529
rect 14516 27448 14521 27512
rect 14585 27448 14611 27512
rect 14675 27448 14701 27512
rect 14765 27448 14791 27512
rect 14855 27448 14881 27512
rect 14945 27448 14971 27512
rect 15035 27448 15040 27512
rect 14516 27431 15040 27448
rect 14516 27367 14521 27431
rect 14585 27367 14611 27431
rect 14675 27367 14701 27431
rect 14765 27367 14791 27431
rect 14855 27367 14881 27431
rect 14945 27367 14971 27431
rect 15035 27367 15040 27431
rect 14516 27350 15040 27367
rect 14516 27286 14521 27350
rect 14585 27286 14611 27350
rect 14675 27286 14701 27350
rect 14765 27286 14791 27350
rect 14855 27286 14881 27350
rect 14945 27286 14971 27350
rect 15035 27286 15040 27350
rect 14516 27268 15040 27286
rect 14516 27204 14521 27268
rect 14585 27204 14611 27268
rect 14675 27204 14701 27268
rect 14765 27204 14791 27268
rect 14855 27204 14881 27268
rect 14945 27204 14971 27268
rect 15035 27204 15040 27268
rect 14516 27186 15040 27204
rect 14516 27122 14521 27186
rect 14585 27122 14611 27186
rect 14675 27122 14701 27186
rect 14765 27122 14791 27186
rect 14855 27122 14881 27186
rect 14945 27122 14971 27186
rect 15035 27122 15040 27186
rect 14516 27104 15040 27122
rect 14516 27040 14521 27104
rect 14585 27040 14611 27104
rect 14675 27040 14701 27104
rect 14765 27040 14791 27104
rect 14855 27040 14881 27104
rect 14945 27040 14971 27104
rect 15035 27040 15040 27104
rect 14516 27039 15040 27040
rect 1976 25853 2492 25854
rect 1976 25789 1977 25853
rect 2041 25789 2067 25853
rect 2131 25789 2157 25853
rect 2221 25789 2247 25853
rect 2311 25789 2337 25853
rect 2401 25789 2427 25853
rect 2491 25789 2492 25853
rect 1976 25770 2492 25789
rect 1976 25706 1977 25770
rect 2041 25706 2067 25770
rect 2131 25706 2157 25770
rect 2221 25706 2247 25770
rect 2311 25706 2337 25770
rect 2401 25706 2427 25770
rect 2491 25706 2492 25770
rect 1976 25687 2492 25706
rect 1976 25623 1977 25687
rect 2041 25623 2067 25687
rect 2131 25623 2157 25687
rect 2221 25623 2247 25687
rect 2311 25623 2337 25687
rect 2401 25623 2427 25687
rect 2491 25623 2492 25687
rect 1976 25604 2492 25623
rect 1976 25540 1977 25604
rect 2041 25540 2067 25604
rect 2131 25540 2157 25604
rect 2221 25540 2247 25604
rect 2311 25540 2337 25604
rect 2401 25540 2427 25604
rect 2491 25540 2492 25604
rect 1976 25521 2492 25540
rect 1976 25457 1977 25521
rect 2041 25457 2067 25521
rect 2131 25457 2157 25521
rect 2221 25457 2247 25521
rect 2311 25457 2337 25521
rect 2401 25457 2427 25521
rect 2491 25457 2492 25521
rect 1976 25437 2492 25457
rect 1976 25373 1977 25437
rect 2041 25373 2067 25437
rect 2131 25373 2157 25437
rect 2221 25373 2247 25437
rect 2311 25373 2337 25437
rect 2401 25373 2427 25437
rect 2491 25373 2492 25437
rect 1976 25353 2492 25373
rect 1976 25289 1977 25353
rect 2041 25289 2067 25353
rect 2131 25289 2157 25353
rect 2221 25289 2247 25353
rect 2311 25289 2337 25353
rect 2401 25289 2427 25353
rect 2491 25289 2492 25353
rect 1976 25269 2492 25289
rect 1976 25205 1977 25269
rect 2041 25205 2067 25269
rect 2131 25205 2157 25269
rect 2221 25205 2247 25269
rect 2311 25205 2337 25269
rect 2401 25205 2427 25269
rect 2491 25205 2492 25269
rect 1976 25185 2492 25205
rect 1976 25121 1977 25185
rect 2041 25121 2067 25185
rect 2131 25121 2157 25185
rect 2221 25121 2247 25185
rect 2311 25121 2337 25185
rect 2401 25121 2427 25185
rect 2491 25121 2492 25185
rect 1976 25101 2492 25121
rect 1976 25037 1977 25101
rect 2041 25037 2067 25101
rect 2131 25037 2157 25101
rect 2221 25037 2247 25101
rect 2311 25037 2337 25101
rect 2401 25037 2427 25101
rect 2491 25037 2492 25101
rect 1976 25017 2492 25037
rect 1976 24953 1977 25017
rect 2041 24953 2067 25017
rect 2131 24953 2157 25017
rect 2221 24953 2247 25017
rect 2311 24953 2337 25017
rect 2401 24953 2427 25017
rect 2491 24953 2492 25017
rect 1976 24933 2492 24953
rect 1976 24869 1977 24933
rect 2041 24869 2067 24933
rect 2131 24869 2157 24933
rect 2221 24869 2247 24933
rect 2311 24869 2337 24933
rect 2401 24869 2427 24933
rect 2491 24869 2492 24933
rect 1976 24849 2492 24869
rect 1976 24785 1977 24849
rect 2041 24785 2067 24849
rect 2131 24785 2157 24849
rect 2221 24785 2247 24849
rect 2311 24785 2337 24849
rect 2401 24785 2427 24849
rect 2491 24785 2492 24849
rect 1976 24765 2492 24785
rect 1976 24701 1977 24765
rect 2041 24701 2067 24765
rect 2131 24701 2157 24765
rect 2221 24701 2247 24765
rect 2311 24701 2337 24765
rect 2401 24701 2427 24765
rect 2491 24701 2492 24765
rect 1976 24681 2492 24701
rect 1976 24617 1977 24681
rect 2041 24617 2067 24681
rect 2131 24617 2157 24681
rect 2221 24617 2247 24681
rect 2311 24617 2337 24681
rect 2401 24617 2427 24681
rect 2491 24617 2492 24681
rect 1976 24597 2492 24617
rect 1976 24533 1977 24597
rect 2041 24533 2067 24597
rect 2131 24533 2157 24597
rect 2221 24533 2247 24597
rect 2311 24533 2337 24597
rect 2401 24533 2427 24597
rect 2491 24533 2492 24597
rect 1976 24513 2492 24533
rect 1976 24449 1977 24513
rect 2041 24449 2067 24513
rect 2131 24449 2157 24513
rect 2221 24449 2247 24513
rect 2311 24449 2337 24513
rect 2401 24449 2427 24513
rect 2491 24449 2492 24513
rect 1976 24429 2492 24449
rect 1976 24365 1977 24429
rect 2041 24365 2067 24429
rect 2131 24365 2157 24429
rect 2221 24365 2247 24429
rect 2311 24365 2337 24429
rect 2401 24365 2427 24429
rect 2491 24365 2492 24429
rect 1976 24345 2492 24365
rect 1976 24281 1977 24345
rect 2041 24281 2067 24345
rect 2131 24281 2157 24345
rect 2221 24281 2247 24345
rect 2311 24281 2337 24345
rect 2401 24281 2427 24345
rect 2491 24281 2492 24345
rect 1976 24280 2492 24281
rect 14506 25809 15038 25810
rect 14506 25745 14510 25809
rect 14574 25745 14602 25809
rect 14666 25745 14694 25809
rect 14758 25745 14786 25809
rect 14850 25745 14878 25809
rect 14942 25745 14970 25809
rect 15034 25745 15038 25809
rect 14506 25729 15038 25745
rect 14506 25665 14510 25729
rect 14574 25665 14602 25729
rect 14666 25665 14694 25729
rect 14758 25665 14786 25729
rect 14850 25665 14878 25729
rect 14942 25665 14970 25729
rect 15034 25665 15038 25729
rect 14506 25648 15038 25665
rect 14506 25584 14510 25648
rect 14574 25584 14602 25648
rect 14666 25584 14694 25648
rect 14758 25584 14786 25648
rect 14850 25584 14878 25648
rect 14942 25584 14970 25648
rect 15034 25584 15038 25648
rect 14506 25567 15038 25584
rect 14506 25503 14510 25567
rect 14574 25503 14602 25567
rect 14666 25503 14694 25567
rect 14758 25503 14786 25567
rect 14850 25503 14878 25567
rect 14942 25503 14970 25567
rect 15034 25503 15038 25567
rect 14506 25486 15038 25503
rect 14506 25422 14510 25486
rect 14574 25422 14602 25486
rect 14666 25422 14694 25486
rect 14758 25422 14786 25486
rect 14850 25422 14878 25486
rect 14942 25422 14970 25486
rect 15034 25422 15038 25486
rect 14506 25405 15038 25422
rect 14506 25341 14510 25405
rect 14574 25341 14602 25405
rect 14666 25341 14694 25405
rect 14758 25341 14786 25405
rect 14850 25341 14878 25405
rect 14942 25341 14970 25405
rect 15034 25341 15038 25405
rect 14506 25324 15038 25341
rect 14506 25260 14510 25324
rect 14574 25260 14602 25324
rect 14666 25260 14694 25324
rect 14758 25260 14786 25324
rect 14850 25260 14878 25324
rect 14942 25260 14970 25324
rect 15034 25260 15038 25324
rect 14506 25243 15038 25260
rect 14506 25179 14510 25243
rect 14574 25179 14602 25243
rect 14666 25179 14694 25243
rect 14758 25179 14786 25243
rect 14850 25179 14878 25243
rect 14942 25179 14970 25243
rect 15034 25179 15038 25243
rect 14506 25162 15038 25179
rect 14506 25098 14510 25162
rect 14574 25098 14602 25162
rect 14666 25098 14694 25162
rect 14758 25098 14786 25162
rect 14850 25098 14878 25162
rect 14942 25098 14970 25162
rect 15034 25098 15038 25162
rect 14506 25081 15038 25098
rect 14506 25017 14510 25081
rect 14574 25017 14602 25081
rect 14666 25017 14694 25081
rect 14758 25017 14786 25081
rect 14850 25017 14878 25081
rect 14942 25017 14970 25081
rect 15034 25017 15038 25081
rect 14506 25000 15038 25017
rect 14506 24936 14510 25000
rect 14574 24936 14602 25000
rect 14666 24936 14694 25000
rect 14758 24936 14786 25000
rect 14850 24936 14878 25000
rect 14942 24936 14970 25000
rect 15034 24936 15038 25000
rect 14506 24919 15038 24936
rect 14506 24855 14510 24919
rect 14574 24855 14602 24919
rect 14666 24855 14694 24919
rect 14758 24855 14786 24919
rect 14850 24855 14878 24919
rect 14942 24855 14970 24919
rect 15034 24855 15038 24919
rect 14506 24838 15038 24855
rect 14506 24774 14510 24838
rect 14574 24774 14602 24838
rect 14666 24774 14694 24838
rect 14758 24774 14786 24838
rect 14850 24774 14878 24838
rect 14942 24774 14970 24838
rect 15034 24774 15038 24838
rect 14506 24757 15038 24774
rect 14506 24693 14510 24757
rect 14574 24693 14602 24757
rect 14666 24693 14694 24757
rect 14758 24693 14786 24757
rect 14850 24693 14878 24757
rect 14942 24693 14970 24757
rect 15034 24693 15038 24757
rect 14506 24676 15038 24693
rect 14506 24612 14510 24676
rect 14574 24612 14602 24676
rect 14666 24612 14694 24676
rect 14758 24612 14786 24676
rect 14850 24612 14878 24676
rect 14942 24612 14970 24676
rect 15034 24612 15038 24676
rect 14506 24595 15038 24612
rect 14506 24531 14510 24595
rect 14574 24531 14602 24595
rect 14666 24531 14694 24595
rect 14758 24531 14786 24595
rect 14850 24531 14878 24595
rect 14942 24531 14970 24595
rect 15034 24531 15038 24595
rect 14506 24514 15038 24531
rect 14506 24450 14510 24514
rect 14574 24450 14602 24514
rect 14666 24450 14694 24514
rect 14758 24450 14786 24514
rect 14850 24450 14878 24514
rect 14942 24450 14970 24514
rect 15034 24450 15038 24514
rect 14506 24433 15038 24450
rect 14506 24369 14510 24433
rect 14574 24369 14602 24433
rect 14666 24369 14694 24433
rect 14758 24369 14786 24433
rect 14850 24369 14878 24433
rect 14942 24369 14970 24433
rect 15034 24369 15038 24433
rect 14506 24352 15038 24369
rect 14506 24288 14510 24352
rect 14574 24288 14602 24352
rect 14666 24288 14694 24352
rect 14758 24288 14786 24352
rect 14850 24288 14878 24352
rect 14942 24288 14970 24352
rect 15034 24288 15038 24352
rect 14506 24271 15038 24288
tri 1960 24248 1962 24250 se
rect 1962 24248 2500 24250
rect 1714 24240 2500 24248
rect 1714 24176 1977 24240
rect 2041 24176 2065 24240
rect 2129 24176 2153 24240
rect 2217 24176 2241 24240
rect 2305 24176 2328 24240
rect 2392 24176 2415 24240
rect 2479 24176 2500 24240
rect 1714 24144 2500 24176
rect 1714 24080 1977 24144
rect 2041 24080 2065 24144
rect 2129 24080 2153 24144
rect 2217 24080 2241 24144
rect 2305 24080 2328 24144
rect 2392 24080 2415 24144
rect 2479 24080 2500 24144
rect 1714 24048 2500 24080
rect 1714 24002 1977 24048
rect 1503 24001 1977 24002
rect 1503 23937 1739 24001
rect 1803 23937 1875 24001
rect 1939 23984 1977 24001
rect 2041 23984 2065 24048
rect 2129 23984 2153 24048
rect 2217 23984 2241 24048
rect 2305 23984 2328 24048
rect 2392 23984 2415 24048
rect 2479 23984 2500 24048
rect 1939 23952 2500 23984
rect 1939 23937 1977 23952
rect 1503 23888 1977 23937
rect 2041 23888 2065 23952
rect 2129 23888 2153 23952
rect 2217 23888 2241 23952
rect 2305 23888 2328 23952
rect 2392 23888 2415 23952
rect 2479 23888 2500 23952
rect 1503 23865 2500 23888
rect 1503 23801 1739 23865
rect 1803 23801 1875 23865
rect 1939 23856 2500 23865
rect 1939 23801 1977 23856
rect 1503 23792 1977 23801
rect 2041 23792 2065 23856
rect 2129 23792 2153 23856
rect 2217 23792 2241 23856
rect 2305 23792 2328 23856
rect 2392 23792 2415 23856
rect 2479 23792 2500 23856
rect 1503 23791 2500 23792
rect 400 23785 1460 23791
rect 400 23721 1094 23785
rect 1158 23721 1188 23785
rect 1252 23721 1282 23785
rect 1346 23721 1376 23785
rect 1440 23721 1460 23785
rect 400 23703 1460 23721
rect 400 23639 1094 23703
rect 1158 23639 1188 23703
rect 1252 23639 1282 23703
rect 1346 23639 1376 23703
rect 1440 23639 1460 23703
rect 400 23621 1460 23639
rect 400 23557 1094 23621
rect 1158 23557 1188 23621
rect 1252 23557 1282 23621
rect 1346 23557 1376 23621
rect 1440 23557 1460 23621
rect 400 23539 1460 23557
rect 400 23475 1094 23539
rect 1158 23475 1188 23539
rect 1252 23475 1282 23539
rect 1346 23475 1376 23539
rect 1440 23475 1460 23539
rect 400 23457 1460 23475
rect 400 23393 1094 23457
rect 1158 23393 1188 23457
rect 1252 23393 1282 23457
rect 1346 23393 1376 23457
rect 1440 23393 1460 23457
rect 400 23375 1460 23393
rect 400 23311 1094 23375
rect 1158 23311 1188 23375
rect 1252 23311 1282 23375
rect 1346 23311 1376 23375
rect 1440 23311 1460 23375
rect 400 23293 1460 23311
rect 400 23229 1094 23293
rect 1158 23229 1188 23293
rect 1252 23229 1282 23293
rect 1346 23229 1376 23293
rect 1440 23229 1460 23293
rect 400 23211 1460 23229
rect 400 23147 1094 23211
rect 1158 23147 1188 23211
rect 1252 23147 1282 23211
rect 1346 23147 1376 23211
rect 1440 23147 1460 23211
rect 400 23129 1460 23147
rect 400 23065 1094 23129
rect 1158 23065 1188 23129
rect 1252 23065 1282 23129
rect 1346 23065 1376 23129
rect 1440 23065 1460 23129
rect 400 23047 1460 23065
rect 400 22983 1094 23047
rect 1158 22983 1188 23047
rect 1252 22983 1282 23047
rect 1346 22983 1376 23047
rect 1440 22983 1460 23047
rect 400 22964 1460 22983
rect 400 22900 1094 22964
rect 1158 22900 1188 22964
rect 1252 22900 1282 22964
rect 1346 22900 1376 22964
rect 1440 22900 1460 22964
rect 400 22881 1460 22900
rect 400 22817 1094 22881
rect 1158 22817 1188 22881
rect 1252 22817 1282 22881
rect 1346 22817 1376 22881
rect 1440 22817 1460 22881
rect 400 22798 1460 22817
rect 400 22734 1094 22798
rect 1158 22734 1188 22798
rect 1252 22734 1282 22798
rect 1346 22734 1376 22798
rect 1440 22734 1460 22798
rect 400 22715 1460 22734
rect 400 22651 1094 22715
rect 1158 22651 1188 22715
rect 1252 22651 1282 22715
rect 1346 22651 1376 22715
rect 1440 22651 1460 22715
rect 400 22632 1460 22651
rect 400 22568 1094 22632
rect 1158 22568 1188 22632
rect 1252 22568 1282 22632
rect 1346 22568 1376 22632
rect 1440 22568 1460 22632
rect 400 22549 1460 22568
rect 400 22485 1094 22549
rect 1158 22485 1188 22549
rect 1252 22485 1282 22549
rect 1346 22485 1376 22549
rect 1440 22485 1460 22549
rect 400 22466 1460 22485
rect 400 22402 1094 22466
rect 1158 22402 1188 22466
rect 1252 22402 1282 22466
rect 1346 22402 1376 22466
rect 1440 22402 1460 22466
rect 400 22383 1460 22402
rect 400 22319 1094 22383
rect 1158 22319 1188 22383
rect 1252 22319 1282 22383
rect 1346 22319 1376 22383
rect 1440 22319 1460 22383
rect 400 22300 1460 22319
rect 400 22236 1094 22300
rect 1158 22236 1188 22300
rect 1252 22236 1282 22300
rect 1346 22236 1376 22300
rect 1440 22236 1460 22300
rect 400 22217 1460 22236
rect 400 22153 1094 22217
rect 1158 22153 1188 22217
rect 1252 22153 1282 22217
rect 1346 22153 1376 22217
rect 1440 22153 1460 22217
rect 400 22134 1460 22153
rect 400 22070 1094 22134
rect 1158 22070 1188 22134
rect 1252 22070 1282 22134
rect 1346 22070 1376 22134
rect 1440 22070 1460 22134
rect 400 22051 1460 22070
rect 400 21987 1094 22051
rect 1158 21987 1188 22051
rect 1252 21987 1282 22051
rect 1346 21987 1376 22051
rect 1440 21987 1460 22051
rect 400 21968 1460 21987
rect 400 21904 1094 21968
rect 1158 21904 1188 21968
rect 1252 21904 1282 21968
rect 1346 21904 1376 21968
rect 1440 21904 1460 21968
rect 400 21885 1460 21904
rect 400 21821 1094 21885
rect 1158 21821 1188 21885
rect 1252 21821 1282 21885
rect 1346 21821 1376 21885
rect 1440 21821 1460 21885
rect 400 21802 1460 21821
rect 400 21738 1094 21802
rect 1158 21738 1188 21802
rect 1252 21738 1282 21802
rect 1346 21738 1376 21802
rect 1440 21738 1460 21802
rect 400 21719 1460 21738
rect 400 21655 1094 21719
rect 1158 21655 1188 21719
rect 1252 21655 1282 21719
rect 1346 21655 1376 21719
rect 1440 21655 1460 21719
rect 400 21636 1460 21655
rect 400 21572 1094 21636
rect 1158 21572 1188 21636
rect 1252 21572 1282 21636
rect 1346 21572 1376 21636
rect 1440 21572 1460 21636
rect 400 21553 1460 21572
rect 400 21489 1094 21553
rect 1158 21489 1188 21553
rect 1252 21489 1282 21553
rect 1346 21489 1376 21553
rect 1440 21489 1460 21553
rect 400 21470 1460 21489
rect 400 21406 1094 21470
rect 1158 21406 1188 21470
rect 1252 21406 1282 21470
rect 1346 21406 1376 21470
rect 1440 21406 1460 21470
rect 400 21387 1460 21406
rect 400 21323 1094 21387
rect 1158 21323 1188 21387
rect 1252 21323 1282 21387
rect 1346 21323 1376 21387
rect 1440 21323 1460 21387
rect 400 21317 1460 21323
rect 1467 23773 2500 23791
rect 1467 23709 1474 23773
rect 1538 23709 1554 23773
rect 1618 23709 1634 23773
rect 1698 23709 1714 23773
rect 1778 23709 1794 23773
rect 1858 23709 1874 23773
rect 1938 23709 1954 23773
rect 2018 23709 2034 23773
rect 2098 23709 2114 23773
rect 2178 23709 2194 23773
rect 2258 23709 2274 23773
rect 2338 23709 2354 23773
rect 2418 23709 2434 23773
rect 2498 23709 2500 23773
rect 1467 23691 2500 23709
rect 1467 23627 1474 23691
rect 1538 23627 1554 23691
rect 1618 23627 1634 23691
rect 1698 23627 1714 23691
rect 1778 23627 1794 23691
rect 1858 23627 1874 23691
rect 1938 23627 1954 23691
rect 2018 23627 2034 23691
rect 2098 23627 2114 23691
rect 2178 23627 2194 23691
rect 2258 23627 2274 23691
rect 2338 23627 2354 23691
rect 2418 23627 2434 23691
rect 2498 23627 2500 23691
rect 1467 23609 2500 23627
rect 1467 23545 1474 23609
rect 1538 23545 1554 23609
rect 1618 23545 1634 23609
rect 1698 23545 1714 23609
rect 1778 23545 1794 23609
rect 1858 23545 1874 23609
rect 1938 23545 1954 23609
rect 2018 23545 2034 23609
rect 2098 23545 2114 23609
rect 2178 23545 2194 23609
rect 2258 23545 2274 23609
rect 2338 23545 2354 23609
rect 2418 23545 2434 23609
rect 2498 23545 2500 23609
rect 1467 23527 2500 23545
rect 1467 23463 1474 23527
rect 1538 23463 1554 23527
rect 1618 23463 1634 23527
rect 1698 23463 1714 23527
rect 1778 23463 1794 23527
rect 1858 23463 1874 23527
rect 1938 23463 1954 23527
rect 2018 23463 2034 23527
rect 2098 23463 2114 23527
rect 2178 23463 2194 23527
rect 2258 23463 2274 23527
rect 2338 23463 2354 23527
rect 2418 23463 2434 23527
rect 2498 23463 2500 23527
rect 1467 23445 2500 23463
rect 1467 23381 1474 23445
rect 1538 23381 1554 23445
rect 1618 23381 1634 23445
rect 1698 23381 1714 23445
rect 1778 23381 1794 23445
rect 1858 23381 1874 23445
rect 1938 23381 1954 23445
rect 2018 23381 2034 23445
rect 2098 23381 2114 23445
rect 2178 23381 2194 23445
rect 2258 23381 2274 23445
rect 2338 23381 2354 23445
rect 2418 23381 2434 23445
rect 2498 23381 2500 23445
rect 1467 23363 2500 23381
rect 1467 23299 1474 23363
rect 1538 23299 1554 23363
rect 1618 23299 1634 23363
rect 1698 23299 1714 23363
rect 1778 23299 1794 23363
rect 1858 23299 1874 23363
rect 1938 23299 1954 23363
rect 2018 23299 2034 23363
rect 2098 23299 2114 23363
rect 2178 23299 2194 23363
rect 2258 23299 2274 23363
rect 2338 23299 2354 23363
rect 2418 23299 2434 23363
rect 2498 23299 2500 23363
rect 1467 23281 2500 23299
rect 1467 23217 1474 23281
rect 1538 23217 1554 23281
rect 1618 23217 1634 23281
rect 1698 23217 1714 23281
rect 1778 23217 1794 23281
rect 1858 23217 1874 23281
rect 1938 23217 1954 23281
rect 2018 23217 2034 23281
rect 2098 23217 2114 23281
rect 2178 23217 2194 23281
rect 2258 23217 2274 23281
rect 2338 23217 2354 23281
rect 2418 23217 2434 23281
rect 2498 23217 2500 23281
rect 1467 23199 2500 23217
rect 1467 23135 1474 23199
rect 1538 23135 1554 23199
rect 1618 23135 1634 23199
rect 1698 23135 1714 23199
rect 1778 23135 1794 23199
rect 1858 23135 1874 23199
rect 1938 23135 1954 23199
rect 2018 23135 2034 23199
rect 2098 23135 2114 23199
rect 2178 23135 2194 23199
rect 2258 23135 2274 23199
rect 2338 23135 2354 23199
rect 2418 23135 2434 23199
rect 2498 23135 2500 23199
rect 14506 24207 14510 24271
rect 14574 24207 14602 24271
rect 14666 24207 14694 24271
rect 14758 24207 14786 24271
rect 14850 24207 14878 24271
rect 14942 24207 14970 24271
rect 15034 24207 15038 24271
rect 14506 24190 15038 24207
rect 14506 24126 14510 24190
rect 14574 24126 14602 24190
rect 14666 24126 14694 24190
rect 14758 24126 14786 24190
rect 14850 24126 14878 24190
rect 14942 24126 14970 24190
rect 15034 24126 15038 24190
rect 14506 24109 15038 24126
rect 14506 24045 14510 24109
rect 14574 24045 14602 24109
rect 14666 24045 14694 24109
rect 14758 24045 14786 24109
rect 14850 24045 14878 24109
rect 14942 24045 14970 24109
rect 15034 24045 15038 24109
rect 14506 24028 15038 24045
rect 14506 23964 14510 24028
rect 14574 23964 14602 24028
rect 14666 23964 14694 24028
rect 14758 23964 14786 24028
rect 14850 23964 14878 24028
rect 14942 23964 14970 24028
rect 15034 23964 15038 24028
rect 14506 23947 15038 23964
rect 14506 23883 14510 23947
rect 14574 23883 14602 23947
rect 14666 23883 14694 23947
rect 14758 23883 14786 23947
rect 14850 23883 14878 23947
rect 14942 23883 14970 23947
rect 15034 23883 15038 23947
rect 14506 23866 15038 23883
rect 14506 23802 14510 23866
rect 14574 23802 14602 23866
rect 14666 23802 14694 23866
rect 14758 23802 14786 23866
rect 14850 23802 14878 23866
rect 14942 23802 14970 23866
rect 15034 23802 15038 23866
rect 14506 23785 15038 23802
rect 14506 23721 14510 23785
rect 14574 23721 14602 23785
rect 14666 23721 14694 23785
rect 14758 23721 14786 23785
rect 14850 23721 14878 23785
rect 14942 23721 14970 23785
rect 15034 23721 15038 23785
rect 14506 23704 15038 23721
rect 14506 23640 14510 23704
rect 14574 23640 14602 23704
rect 14666 23640 14694 23704
rect 14758 23640 14786 23704
rect 14850 23640 14878 23704
rect 14942 23640 14970 23704
rect 15034 23640 15038 23704
rect 14506 23623 15038 23640
rect 14506 23559 14510 23623
rect 14574 23559 14602 23623
rect 14666 23559 14694 23623
rect 14758 23559 14786 23623
rect 14850 23559 14878 23623
rect 14942 23559 14970 23623
rect 15034 23559 15038 23623
rect 14506 23542 15038 23559
rect 14506 23478 14510 23542
rect 14574 23478 14602 23542
rect 14666 23478 14694 23542
rect 14758 23478 14786 23542
rect 14850 23478 14878 23542
rect 14942 23478 14970 23542
rect 15034 23478 15038 23542
rect 14506 23461 15038 23478
rect 14506 23397 14510 23461
rect 14574 23397 14602 23461
rect 14666 23397 14694 23461
rect 14758 23397 14786 23461
rect 14850 23397 14878 23461
rect 14942 23397 14970 23461
rect 15034 23397 15038 23461
rect 14506 23380 15038 23397
rect 14506 23316 14510 23380
rect 14574 23316 14602 23380
rect 14666 23316 14694 23380
rect 14758 23316 14786 23380
rect 14850 23316 14878 23380
rect 14942 23316 14970 23380
rect 15034 23316 15038 23380
rect 14506 23299 15038 23316
rect 14506 23235 14510 23299
rect 14574 23235 14602 23299
rect 14666 23235 14694 23299
rect 14758 23235 14786 23299
rect 14850 23235 14878 23299
rect 14942 23235 14970 23299
rect 15034 23235 15038 23299
rect 14506 23218 15038 23235
rect 14506 23154 14510 23218
rect 14574 23154 14602 23218
rect 14666 23154 14694 23218
rect 14758 23154 14786 23218
rect 14850 23154 14878 23218
rect 14942 23154 14970 23218
rect 15034 23154 15038 23218
rect 14506 23153 15038 23154
rect 1467 23117 2500 23135
rect 1467 23053 1474 23117
rect 1538 23053 1554 23117
rect 1618 23053 1634 23117
rect 1698 23053 1714 23117
rect 1778 23053 1794 23117
rect 1858 23053 1874 23117
rect 1938 23053 1954 23117
rect 2018 23053 2034 23117
rect 2098 23053 2114 23117
rect 2178 23053 2194 23117
rect 2258 23053 2274 23117
rect 2338 23053 2354 23117
rect 2418 23053 2434 23117
rect 2498 23053 2500 23117
rect 1467 23035 2500 23053
rect 1467 22971 1474 23035
rect 1538 22971 1554 23035
rect 1618 22971 1634 23035
rect 1698 22971 1714 23035
rect 1778 22971 1794 23035
rect 1858 22971 1874 23035
rect 1938 22971 1954 23035
rect 2018 22971 2034 23035
rect 2098 22971 2114 23035
rect 2178 22971 2194 23035
rect 2258 22971 2274 23035
rect 2338 22971 2354 23035
rect 2418 22971 2434 23035
rect 2498 22971 2500 23035
rect 1467 22953 2500 22971
rect 1467 22889 1474 22953
rect 1538 22889 1554 22953
rect 1618 22889 1634 22953
rect 1698 22889 1714 22953
rect 1778 22889 1794 22953
rect 1858 22889 1874 22953
rect 1938 22889 1954 22953
rect 2018 22889 2034 22953
rect 2098 22889 2114 22953
rect 2178 22889 2194 22953
rect 2258 22889 2274 22953
rect 2338 22889 2354 22953
rect 2418 22889 2434 22953
rect 2498 22889 2500 22953
rect 1467 22871 2500 22889
rect 1467 22807 1474 22871
rect 1538 22807 1554 22871
rect 1618 22807 1634 22871
rect 1698 22807 1714 22871
rect 1778 22807 1794 22871
rect 1858 22807 1874 22871
rect 1938 22807 1954 22871
rect 2018 22807 2034 22871
rect 2098 22807 2114 22871
rect 2178 22807 2194 22871
rect 2258 22807 2274 22871
rect 2338 22807 2354 22871
rect 2418 22807 2434 22871
rect 2498 22807 2500 22871
rect 1467 22789 2500 22807
rect 1467 22725 1474 22789
rect 1538 22725 1554 22789
rect 1618 22725 1634 22789
rect 1698 22725 1714 22789
rect 1778 22725 1794 22789
rect 1858 22725 1874 22789
rect 1938 22725 1954 22789
rect 2018 22725 2034 22789
rect 2098 22725 2114 22789
rect 2178 22725 2194 22789
rect 2258 22725 2274 22789
rect 2338 22725 2354 22789
rect 2418 22725 2434 22789
rect 2498 22725 2500 22789
rect 1467 22707 2500 22725
rect 1467 22643 1474 22707
rect 1538 22643 1554 22707
rect 1618 22643 1634 22707
rect 1698 22643 1714 22707
rect 1778 22643 1794 22707
rect 1858 22643 1874 22707
rect 1938 22643 1954 22707
rect 2018 22643 2034 22707
rect 2098 22643 2114 22707
rect 2178 22643 2194 22707
rect 2258 22643 2274 22707
rect 2338 22643 2354 22707
rect 2418 22643 2434 22707
rect 2498 22643 2500 22707
rect 1467 22625 2500 22643
rect 1467 22561 1474 22625
rect 1538 22561 1554 22625
rect 1618 22561 1634 22625
rect 1698 22561 1714 22625
rect 1778 22561 1794 22625
rect 1858 22561 1874 22625
rect 1938 22561 1954 22625
rect 2018 22561 2034 22625
rect 2098 22561 2114 22625
rect 2178 22561 2194 22625
rect 2258 22561 2274 22625
rect 2338 22561 2354 22625
rect 2418 22561 2434 22625
rect 2498 22561 2500 22625
rect 1467 22543 2500 22561
rect 1467 22479 1474 22543
rect 1538 22479 1554 22543
rect 1618 22479 1634 22543
rect 1698 22479 1714 22543
rect 1778 22479 1794 22543
rect 1858 22479 1874 22543
rect 1938 22479 1954 22543
rect 2018 22479 2034 22543
rect 2098 22479 2114 22543
rect 2178 22479 2194 22543
rect 2258 22479 2274 22543
rect 2338 22479 2354 22543
rect 2418 22479 2434 22543
rect 2498 22479 2500 22543
rect 1467 22461 2500 22479
rect 1467 22397 1474 22461
rect 1538 22397 1554 22461
rect 1618 22397 1634 22461
rect 1698 22397 1714 22461
rect 1778 22397 1794 22461
rect 1858 22397 1874 22461
rect 1938 22397 1954 22461
rect 2018 22397 2034 22461
rect 2098 22397 2114 22461
rect 2178 22397 2194 22461
rect 2258 22397 2274 22461
rect 2338 22397 2354 22461
rect 2418 22397 2434 22461
rect 2498 22397 2500 22461
rect 1467 22379 2500 22397
rect 1467 22315 1474 22379
rect 1538 22315 1554 22379
rect 1618 22315 1634 22379
rect 1698 22315 1714 22379
rect 1778 22315 1794 22379
rect 1858 22315 1874 22379
rect 1938 22315 1954 22379
rect 2018 22315 2034 22379
rect 2098 22315 2114 22379
rect 2178 22315 2194 22379
rect 2258 22315 2274 22379
rect 2338 22315 2354 22379
rect 2418 22315 2434 22379
rect 2498 22315 2500 22379
rect 1467 22297 2500 22315
rect 1467 22233 1474 22297
rect 1538 22233 1554 22297
rect 1618 22233 1634 22297
rect 1698 22233 1714 22297
rect 1778 22233 1794 22297
rect 1858 22233 1874 22297
rect 1938 22233 1954 22297
rect 2018 22233 2034 22297
rect 2098 22233 2114 22297
rect 2178 22233 2194 22297
rect 2258 22233 2274 22297
rect 2338 22233 2354 22297
rect 2418 22233 2434 22297
rect 2498 22233 2500 22297
rect 1467 22215 2500 22233
rect 1467 22151 1474 22215
rect 1538 22151 1554 22215
rect 1618 22151 1634 22215
rect 1698 22151 1714 22215
rect 1778 22151 1794 22215
rect 1858 22151 1874 22215
rect 1938 22151 1954 22215
rect 2018 22151 2034 22215
rect 2098 22151 2114 22215
rect 2178 22151 2194 22215
rect 2258 22151 2274 22215
rect 2338 22151 2354 22215
rect 2418 22151 2434 22215
rect 2498 22151 2500 22215
rect 1467 22133 2500 22151
rect 1467 22069 1474 22133
rect 1538 22069 1554 22133
rect 1618 22069 1634 22133
rect 1698 22069 1714 22133
rect 1778 22069 1794 22133
rect 1858 22069 1874 22133
rect 1938 22069 1954 22133
rect 2018 22069 2034 22133
rect 2098 22069 2114 22133
rect 2178 22069 2194 22133
rect 2258 22069 2274 22133
rect 2338 22069 2354 22133
rect 2418 22069 2434 22133
rect 2498 22069 2500 22133
rect 1467 22051 2500 22069
rect 1467 21987 1474 22051
rect 1538 21987 1554 22051
rect 1618 21987 1634 22051
rect 1698 21987 1714 22051
rect 1778 21987 1794 22051
rect 1858 21987 1874 22051
rect 1938 21987 1954 22051
rect 2018 21987 2034 22051
rect 2098 21987 2114 22051
rect 2178 21987 2194 22051
rect 2258 21987 2274 22051
rect 2338 21987 2354 22051
rect 2418 21987 2434 22051
rect 2498 21987 2500 22051
rect 1467 21968 2500 21987
rect 1467 21904 1474 21968
rect 1538 21904 1554 21968
rect 1618 21904 1634 21968
rect 1698 21904 1714 21968
rect 1778 21904 1794 21968
rect 1858 21904 1874 21968
rect 1938 21904 1954 21968
rect 2018 21904 2034 21968
rect 2098 21904 2114 21968
rect 2178 21904 2194 21968
rect 2258 21904 2274 21968
rect 2338 21904 2354 21968
rect 2418 21904 2434 21968
rect 2498 21904 2500 21968
rect 1467 21885 2500 21904
rect 1467 21821 1474 21885
rect 1538 21821 1554 21885
rect 1618 21821 1634 21885
rect 1698 21821 1714 21885
rect 1778 21821 1794 21885
rect 1858 21821 1874 21885
rect 1938 21821 1954 21885
rect 2018 21821 2034 21885
rect 2098 21821 2114 21885
rect 2178 21821 2194 21885
rect 2258 21821 2274 21885
rect 2338 21821 2354 21885
rect 2418 21821 2434 21885
rect 2498 21821 2500 21885
rect 1467 21802 2500 21821
rect 1467 21738 1474 21802
rect 1538 21738 1554 21802
rect 1618 21738 1634 21802
rect 1698 21738 1714 21802
rect 1778 21738 1794 21802
rect 1858 21738 1874 21802
rect 1938 21738 1954 21802
rect 2018 21738 2034 21802
rect 2098 21738 2114 21802
rect 2178 21738 2194 21802
rect 2258 21738 2274 21802
rect 2338 21738 2354 21802
rect 2418 21738 2434 21802
rect 2498 21738 2500 21802
rect 1467 21719 2500 21738
rect 1467 21655 1474 21719
rect 1538 21655 1554 21719
rect 1618 21655 1634 21719
rect 1698 21655 1714 21719
rect 1778 21655 1794 21719
rect 1858 21655 1874 21719
rect 1938 21655 1954 21719
rect 2018 21655 2034 21719
rect 2098 21655 2114 21719
rect 2178 21655 2194 21719
rect 2258 21655 2274 21719
rect 2338 21655 2354 21719
rect 2418 21655 2434 21719
rect 2498 21655 2500 21719
rect 1467 21636 2500 21655
rect 1467 21572 1474 21636
rect 1538 21572 1554 21636
rect 1618 21572 1634 21636
rect 1698 21572 1714 21636
rect 1778 21572 1794 21636
rect 1858 21572 1874 21636
rect 1938 21572 1954 21636
rect 2018 21572 2034 21636
rect 2098 21572 2114 21636
rect 2178 21572 2194 21636
rect 2258 21572 2274 21636
rect 2338 21572 2354 21636
rect 2418 21572 2434 21636
rect 2498 21572 2500 21636
rect 1467 21553 2500 21572
rect 1467 21489 1474 21553
rect 1538 21489 1554 21553
rect 1618 21489 1634 21553
rect 1698 21489 1714 21553
rect 1778 21489 1794 21553
rect 1858 21489 1874 21553
rect 1938 21489 1954 21553
rect 2018 21489 2034 21553
rect 2098 21489 2114 21553
rect 2178 21489 2194 21553
rect 2258 21489 2274 21553
rect 2338 21489 2354 21553
rect 2418 21489 2434 21553
rect 2498 21489 2500 21553
rect 1467 21470 2500 21489
rect 1467 21406 1474 21470
rect 1538 21406 1554 21470
rect 1618 21406 1634 21470
rect 1698 21406 1714 21470
rect 1778 21406 1794 21470
rect 1858 21406 1874 21470
rect 1938 21406 1954 21470
rect 2018 21406 2034 21470
rect 2098 21406 2114 21470
rect 2178 21406 2194 21470
rect 2258 21406 2274 21470
rect 2338 21406 2354 21470
rect 2418 21406 2434 21470
rect 2498 21406 2500 21470
rect 1467 21387 2500 21406
rect 1467 21323 1474 21387
rect 1538 21323 1554 21387
rect 1618 21323 1634 21387
rect 1698 21323 1714 21387
rect 1778 21323 1794 21387
rect 1858 21323 1874 21387
rect 1938 21323 1954 21387
rect 2018 21323 2034 21387
rect 2098 21323 2114 21387
rect 2178 21323 2194 21387
rect 2258 21323 2274 21387
rect 2338 21323 2354 21387
rect 2418 21323 2434 21387
rect 2498 21323 2500 21387
rect 1467 21317 2500 21323
rect 1566 21242 2500 21317
rect 1641 21006 2500 21242
rect 1877 20923 2500 21006
rect 1877 20879 2004 20923
rect 13738 20376 13952 20382
rect 13802 20312 13888 20376
rect 13738 20282 13952 20312
rect 13802 20218 13888 20282
rect 13738 20188 13952 20218
rect 13802 20124 13888 20188
rect 13738 20094 13952 20124
rect 13802 20030 13888 20094
rect 13738 19999 13952 20030
rect 13802 19935 13888 19999
rect 13738 19904 13952 19935
rect 13802 19840 13888 19904
rect 13738 19834 13952 19840
rect 0 14007 254 19000
rect 291 18976 657 18977
rect 291 18912 292 18976
rect 356 18912 392 18976
rect 456 18912 492 18976
rect 556 18912 592 18976
rect 656 18912 657 18976
rect 291 18896 657 18912
rect 291 18832 292 18896
rect 356 18832 392 18896
rect 456 18832 492 18896
rect 556 18832 592 18896
rect 656 18832 657 18896
rect 291 18816 657 18832
rect 291 18752 292 18816
rect 356 18752 392 18816
rect 456 18752 492 18816
rect 556 18752 592 18816
rect 656 18752 657 18816
rect 291 18736 657 18752
rect 291 18672 292 18736
rect 356 18672 392 18736
rect 456 18672 492 18736
rect 556 18672 592 18736
rect 656 18672 657 18736
rect 291 18656 657 18672
rect 291 18592 292 18656
rect 356 18592 392 18656
rect 456 18592 492 18656
rect 556 18592 592 18656
rect 656 18592 657 18656
rect 291 18576 657 18592
rect 291 18512 292 18576
rect 356 18512 392 18576
rect 456 18512 492 18576
rect 556 18512 592 18576
rect 656 18512 657 18576
rect 291 18496 657 18512
rect 291 18432 292 18496
rect 356 18432 392 18496
rect 456 18432 492 18496
rect 556 18432 592 18496
rect 656 18432 657 18496
rect 291 18416 657 18432
rect 291 18352 292 18416
rect 356 18352 392 18416
rect 456 18352 492 18416
rect 556 18352 592 18416
rect 656 18352 657 18416
rect 291 18336 657 18352
rect 291 18272 292 18336
rect 356 18272 392 18336
rect 456 18272 492 18336
rect 556 18272 592 18336
rect 656 18272 657 18336
rect 291 18256 657 18272
rect 291 18192 292 18256
rect 356 18192 392 18256
rect 456 18192 492 18256
rect 556 18192 592 18256
rect 656 18192 657 18256
rect 291 18176 657 18192
rect 291 18112 292 18176
rect 356 18112 392 18176
rect 456 18112 492 18176
rect 556 18112 592 18176
rect 656 18112 657 18176
rect 291 18096 657 18112
rect 291 18032 292 18096
rect 356 18032 392 18096
rect 456 18032 492 18096
rect 556 18032 592 18096
rect 656 18032 657 18096
rect 291 18015 657 18032
rect 291 17951 292 18015
rect 356 17951 392 18015
rect 456 17951 492 18015
rect 556 17951 592 18015
rect 656 17951 657 18015
rect 291 17934 657 17951
rect 291 17870 292 17934
rect 356 17870 392 17934
rect 456 17870 492 17934
rect 556 17870 592 17934
rect 656 17870 657 17934
rect 291 17853 657 17870
rect 291 17789 292 17853
rect 356 17789 392 17853
rect 456 17789 492 17853
rect 556 17789 592 17853
rect 656 17789 657 17853
rect 291 17772 657 17789
rect 291 17708 292 17772
rect 356 17708 392 17772
rect 456 17708 492 17772
rect 556 17708 592 17772
rect 656 17708 657 17772
rect 291 17691 657 17708
rect 291 17627 292 17691
rect 356 17627 392 17691
rect 456 17627 492 17691
rect 556 17627 592 17691
rect 656 17627 657 17691
rect 291 17610 657 17627
rect 291 17546 292 17610
rect 356 17546 392 17610
rect 456 17546 492 17610
rect 556 17546 592 17610
rect 656 17546 657 17610
rect 291 17529 657 17546
rect 291 17465 292 17529
rect 356 17465 392 17529
rect 456 17465 492 17529
rect 556 17465 592 17529
rect 656 17465 657 17529
rect 291 17448 657 17465
rect 291 17384 292 17448
rect 356 17384 392 17448
rect 456 17384 492 17448
rect 556 17384 592 17448
rect 656 17384 657 17448
rect 291 17367 657 17384
rect 291 17303 292 17367
rect 356 17303 392 17367
rect 456 17303 492 17367
rect 556 17303 592 17367
rect 656 17303 657 17367
rect 291 17286 657 17303
rect 291 17222 292 17286
rect 356 17222 392 17286
rect 456 17222 492 17286
rect 556 17222 592 17286
rect 656 17222 657 17286
rect 291 17205 657 17222
rect 291 17141 292 17205
rect 356 17141 392 17205
rect 456 17141 492 17205
rect 556 17141 592 17205
rect 656 17141 657 17205
rect 291 17124 657 17141
rect 291 17060 292 17124
rect 356 17060 392 17124
rect 456 17060 492 17124
rect 556 17060 592 17124
rect 656 17060 657 17124
rect 291 17043 657 17060
rect 291 16979 292 17043
rect 356 16979 392 17043
rect 456 16979 492 17043
rect 556 16979 592 17043
rect 656 16979 657 17043
rect 291 16962 657 16979
rect 291 16898 292 16962
rect 356 16898 392 16962
rect 456 16898 492 16962
rect 556 16898 592 16962
rect 656 16898 657 16962
rect 291 16881 657 16898
rect 291 16817 292 16881
rect 356 16817 392 16881
rect 456 16817 492 16881
rect 556 16817 592 16881
rect 656 16817 657 16881
rect 291 16800 657 16817
rect 291 16736 292 16800
rect 356 16736 392 16800
rect 456 16736 492 16800
rect 556 16736 592 16800
rect 656 16736 657 16800
rect 291 16719 657 16736
rect 291 16655 292 16719
rect 356 16655 392 16719
rect 456 16655 492 16719
rect 556 16655 592 16719
rect 656 16655 657 16719
rect 291 16638 657 16655
rect 291 16574 292 16638
rect 356 16574 392 16638
rect 456 16574 492 16638
rect 556 16574 592 16638
rect 656 16574 657 16638
rect 291 16557 657 16574
rect 291 16493 292 16557
rect 356 16493 392 16557
rect 456 16493 492 16557
rect 556 16493 592 16557
rect 656 16493 657 16557
rect 291 16476 657 16493
rect 291 16412 292 16476
rect 356 16412 392 16476
rect 456 16412 492 16476
rect 556 16412 592 16476
rect 656 16412 657 16476
rect 291 16395 657 16412
rect 291 16331 292 16395
rect 356 16331 392 16395
rect 456 16331 492 16395
rect 556 16331 592 16395
rect 656 16331 657 16395
rect 291 16314 657 16331
rect 291 16250 292 16314
rect 356 16250 392 16314
rect 456 16250 492 16314
rect 556 16250 592 16314
rect 656 16250 657 16314
rect 291 16233 657 16250
rect 291 16169 292 16233
rect 356 16169 392 16233
rect 456 16169 492 16233
rect 556 16169 592 16233
rect 656 16169 657 16233
rect 291 16152 657 16169
rect 291 16088 292 16152
rect 356 16088 392 16152
rect 456 16088 492 16152
rect 556 16088 592 16152
rect 656 16088 657 16152
rect 291 16071 657 16088
rect 291 16007 292 16071
rect 356 16007 392 16071
rect 456 16007 492 16071
rect 556 16007 592 16071
rect 656 16007 657 16071
rect 291 15990 657 16007
rect 291 15926 292 15990
rect 356 15926 392 15990
rect 456 15926 492 15990
rect 556 15926 592 15990
rect 656 15926 657 15990
rect 291 15909 657 15926
rect 291 15845 292 15909
rect 356 15845 392 15909
rect 456 15845 492 15909
rect 556 15845 592 15909
rect 656 15845 657 15909
rect 291 15828 657 15845
rect 291 15764 292 15828
rect 356 15764 392 15828
rect 456 15764 492 15828
rect 556 15764 592 15828
rect 656 15764 657 15828
rect 291 15747 657 15764
rect 291 15683 292 15747
rect 356 15683 392 15747
rect 456 15683 492 15747
rect 556 15683 592 15747
rect 656 15683 657 15747
rect 291 15666 657 15683
rect 291 15602 292 15666
rect 356 15602 392 15666
rect 456 15602 492 15666
rect 556 15602 592 15666
rect 656 15602 657 15666
rect 291 15585 657 15602
rect 291 15521 292 15585
rect 356 15521 392 15585
rect 456 15521 492 15585
rect 556 15521 592 15585
rect 656 15521 657 15585
rect 291 15504 657 15521
rect 291 15440 292 15504
rect 356 15440 392 15504
rect 456 15440 492 15504
rect 556 15440 592 15504
rect 656 15440 657 15504
rect 291 15423 657 15440
rect 291 15359 292 15423
rect 356 15359 392 15423
rect 456 15359 492 15423
rect 556 15359 592 15423
rect 656 15359 657 15423
rect 291 15342 657 15359
rect 291 15278 292 15342
rect 356 15278 392 15342
rect 456 15278 492 15342
rect 556 15278 592 15342
rect 656 15278 657 15342
rect 291 15261 657 15278
rect 291 15197 292 15261
rect 356 15197 392 15261
rect 456 15197 492 15261
rect 556 15197 592 15261
rect 656 15197 657 15261
rect 291 15180 657 15197
rect 291 15116 292 15180
rect 356 15116 392 15180
rect 456 15116 492 15180
rect 556 15116 592 15180
rect 656 15116 657 15180
rect 291 15099 657 15116
rect 291 15035 292 15099
rect 356 15035 392 15099
rect 456 15035 492 15099
rect 556 15035 592 15099
rect 656 15035 657 15099
rect 291 15018 657 15035
rect 291 14954 292 15018
rect 356 14954 392 15018
rect 456 14954 492 15018
rect 556 14954 592 15018
rect 656 14954 657 15018
rect 291 14937 657 14954
rect 291 14873 292 14937
rect 356 14873 392 14937
rect 456 14873 492 14937
rect 556 14873 592 14937
rect 656 14873 657 14937
rect 291 14856 657 14873
rect 291 14792 292 14856
rect 356 14792 392 14856
rect 456 14792 492 14856
rect 556 14792 592 14856
rect 656 14792 657 14856
rect 291 14775 657 14792
rect 291 14711 292 14775
rect 356 14711 392 14775
rect 456 14711 492 14775
rect 556 14711 592 14775
rect 656 14711 657 14775
rect 291 14694 657 14711
rect 291 14630 292 14694
rect 356 14630 392 14694
rect 456 14630 492 14694
rect 556 14630 592 14694
rect 656 14630 657 14694
rect 291 14613 657 14630
rect 291 14549 292 14613
rect 356 14549 392 14613
rect 456 14549 492 14613
rect 556 14549 592 14613
rect 656 14549 657 14613
rect 291 14532 657 14549
rect 291 14468 292 14532
rect 356 14468 392 14532
rect 456 14468 492 14532
rect 556 14468 592 14532
rect 656 14468 657 14532
rect 291 14451 657 14468
rect 291 14387 292 14451
rect 356 14387 392 14451
rect 456 14387 492 14451
rect 556 14387 592 14451
rect 656 14387 657 14451
rect 291 14370 657 14387
rect 291 14306 292 14370
rect 356 14306 392 14370
rect 456 14306 492 14370
rect 556 14306 592 14370
rect 656 14306 657 14370
rect 291 14289 657 14306
rect 291 14225 292 14289
rect 356 14225 392 14289
rect 456 14225 492 14289
rect 556 14225 592 14289
rect 656 14225 657 14289
rect 291 14208 657 14225
rect 291 14144 292 14208
rect 356 14144 392 14208
rect 456 14144 492 14208
rect 556 14144 592 14208
rect 656 14144 657 14208
rect 291 14127 657 14144
rect 291 14063 292 14127
rect 356 14063 392 14127
rect 456 14063 492 14127
rect 556 14063 592 14127
rect 656 14063 657 14127
rect 291 14062 657 14063
rect 15746 14007 16000 19000
rect 0 12817 254 13707
rect 5647 13698 6626 13707
rect 5647 13634 5648 13698
rect 5712 13634 5731 13698
rect 5795 13634 5814 13698
rect 5878 13634 5897 13698
rect 5961 13634 5980 13698
rect 6044 13634 6063 13698
rect 6127 13634 6146 13698
rect 6210 13634 6229 13698
rect 6293 13634 6312 13698
rect 6376 13634 6395 13698
rect 6459 13634 6478 13698
rect 6542 13634 6561 13698
rect 6625 13634 6626 13698
rect 5647 13618 6626 13634
rect 1371 13596 1567 13597
rect 1371 13532 1372 13596
rect 1436 13532 1502 13596
rect 1566 13532 1567 13596
rect 1371 13509 1567 13532
rect 1371 13445 1372 13509
rect 1436 13445 1502 13509
rect 1566 13445 1567 13509
rect 1371 13422 1567 13445
rect 1371 13358 1372 13422
rect 1436 13358 1502 13422
rect 1566 13358 1567 13422
rect 1371 13335 1567 13358
rect 1371 13271 1372 13335
rect 1436 13271 1502 13335
rect 1566 13271 1567 13335
rect 1371 13248 1567 13271
rect 1371 13184 1372 13248
rect 1436 13184 1502 13248
rect 1566 13184 1567 13248
rect 1371 13161 1567 13184
rect 1371 13097 1372 13161
rect 1436 13097 1502 13161
rect 1566 13097 1567 13161
rect 1371 13074 1567 13097
rect 1371 13010 1372 13074
rect 1436 13010 1502 13074
rect 1566 13010 1567 13074
rect 1371 12986 1567 13010
rect 1371 12922 1372 12986
rect 1436 12922 1502 12986
rect 1566 12922 1567 12986
rect 1371 12898 1567 12922
rect 1371 12834 1372 12898
rect 1436 12834 1502 12898
rect 1566 12834 1567 12898
rect 1371 12833 1567 12834
rect 5647 13554 5648 13618
rect 5712 13554 5731 13618
rect 5795 13554 5814 13618
rect 5878 13554 5897 13618
rect 5961 13554 5980 13618
rect 6044 13554 6063 13618
rect 6127 13554 6146 13618
rect 6210 13554 6229 13618
rect 6293 13554 6312 13618
rect 6376 13554 6395 13618
rect 6459 13554 6478 13618
rect 6542 13554 6561 13618
rect 6625 13554 6626 13618
rect 5647 13538 6626 13554
rect 5647 13474 5648 13538
rect 5712 13474 5731 13538
rect 5795 13474 5814 13538
rect 5878 13474 5897 13538
rect 5961 13474 5980 13538
rect 6044 13474 6063 13538
rect 6127 13474 6146 13538
rect 6210 13474 6229 13538
rect 6293 13474 6312 13538
rect 6376 13474 6395 13538
rect 6459 13474 6478 13538
rect 6542 13474 6561 13538
rect 6625 13474 6626 13538
rect 5647 13458 6626 13474
rect 5647 13394 5648 13458
rect 5712 13394 5731 13458
rect 5795 13394 5814 13458
rect 5878 13394 5897 13458
rect 5961 13394 5980 13458
rect 6044 13394 6063 13458
rect 6127 13394 6146 13458
rect 6210 13394 6229 13458
rect 6293 13394 6312 13458
rect 6376 13394 6395 13458
rect 6459 13394 6478 13458
rect 6542 13394 6561 13458
rect 6625 13394 6626 13458
rect 5647 13378 6626 13394
rect 5647 13314 5648 13378
rect 5712 13314 5731 13378
rect 5795 13314 5814 13378
rect 5878 13314 5897 13378
rect 5961 13314 5980 13378
rect 6044 13314 6063 13378
rect 6127 13314 6146 13378
rect 6210 13314 6229 13378
rect 6293 13314 6312 13378
rect 6376 13314 6395 13378
rect 6459 13314 6478 13378
rect 6542 13314 6561 13378
rect 6625 13314 6626 13378
rect 5647 13298 6626 13314
rect 5647 13234 5648 13298
rect 5712 13234 5731 13298
rect 5795 13234 5814 13298
rect 5878 13234 5897 13298
rect 5961 13234 5980 13298
rect 6044 13234 6063 13298
rect 6127 13234 6146 13298
rect 6210 13234 6229 13298
rect 6293 13234 6312 13298
rect 6376 13234 6395 13298
rect 6459 13234 6478 13298
rect 6542 13234 6561 13298
rect 6625 13234 6626 13298
rect 5647 13218 6626 13234
rect 5647 13154 5648 13218
rect 5712 13154 5731 13218
rect 5795 13154 5814 13218
rect 5878 13154 5897 13218
rect 5961 13154 5980 13218
rect 6044 13154 6063 13218
rect 6127 13154 6146 13218
rect 6210 13154 6229 13218
rect 6293 13154 6312 13218
rect 6376 13154 6395 13218
rect 6459 13154 6478 13218
rect 6542 13154 6561 13218
rect 6625 13154 6626 13218
rect 5647 13138 6626 13154
rect 5647 13074 5648 13138
rect 5712 13074 5731 13138
rect 5795 13074 5814 13138
rect 5878 13074 5897 13138
rect 5961 13074 5980 13138
rect 6044 13074 6063 13138
rect 6127 13074 6146 13138
rect 6210 13074 6229 13138
rect 6293 13074 6312 13138
rect 6376 13074 6395 13138
rect 6459 13074 6478 13138
rect 6542 13074 6561 13138
rect 6625 13074 6626 13138
rect 5647 13058 6626 13074
rect 5647 12994 5648 13058
rect 5712 12994 5731 13058
rect 5795 12994 5814 13058
rect 5878 12994 5897 13058
rect 5961 12994 5980 13058
rect 6044 12994 6063 13058
rect 6127 12994 6146 13058
rect 6210 12994 6229 13058
rect 6293 12994 6312 13058
rect 6376 12994 6395 13058
rect 6459 12994 6478 13058
rect 6542 12994 6561 13058
rect 6625 12994 6626 13058
rect 5647 12978 6626 12994
rect 5647 12914 5648 12978
rect 5712 12914 5731 12978
rect 5795 12914 5814 12978
rect 5878 12914 5897 12978
rect 5961 12914 5980 12978
rect 6044 12914 6063 12978
rect 6127 12914 6146 12978
rect 6210 12914 6229 12978
rect 6293 12914 6312 12978
rect 6376 12914 6395 12978
rect 6459 12914 6478 12978
rect 6542 12914 6561 12978
rect 6625 12914 6626 12978
rect 5647 12898 6626 12914
rect 5647 12834 5648 12898
rect 5712 12834 5731 12898
rect 5795 12834 5814 12898
rect 5878 12834 5897 12898
rect 5961 12834 5980 12898
rect 6044 12834 6063 12898
rect 6127 12834 6146 12898
rect 6210 12834 6229 12898
rect 6293 12834 6312 12898
rect 6376 12834 6395 12898
rect 6459 12834 6478 12898
rect 6542 12834 6561 12898
rect 6625 12834 6626 12898
rect 5647 12825 6626 12834
rect 15746 12817 16000 13707
rect 0 11647 254 12537
rect 15746 11647 16000 12537
rect 4625 11533 6856 11534
rect 4625 11469 4626 11533
rect 4690 11469 4706 11533
rect 4770 11469 6705 11533
rect 6769 11469 6785 11533
rect 6849 11469 6856 11533
rect 4625 11468 6856 11469
rect 0 11281 254 11347
rect 521 11346 755 11347
rect 521 11282 522 11346
rect 586 11282 606 11346
rect 670 11282 690 11346
rect 754 11282 755 11346
rect 521 11281 755 11282
rect 4549 11346 4783 11347
rect 4549 11282 4550 11346
rect 4614 11282 4634 11346
rect 4698 11282 4718 11346
rect 4782 11282 4783 11346
rect 4549 11281 4783 11282
rect 8170 11346 8404 11347
rect 8170 11282 8171 11346
rect 8235 11282 8255 11346
rect 8319 11282 8339 11346
rect 8403 11282 8404 11346
rect 8170 11281 8404 11282
rect 9185 11346 9419 11347
rect 9185 11282 9186 11346
rect 9250 11282 9270 11346
rect 9334 11282 9354 11346
rect 9418 11282 9419 11346
rect 9185 11281 9419 11282
rect 15746 11281 16000 11347
rect 0 10625 254 11221
rect 15746 10625 16000 11221
rect 0 10329 254 10565
rect 521 10563 755 10565
rect 521 10499 522 10563
rect 586 10499 606 10563
rect 670 10499 690 10563
rect 754 10499 755 10563
rect 521 10479 755 10499
rect 521 10415 522 10479
rect 586 10415 606 10479
rect 670 10415 690 10479
rect 754 10415 755 10479
rect 521 10395 755 10415
rect 521 10331 522 10395
rect 586 10331 606 10395
rect 670 10331 690 10395
rect 754 10331 755 10395
rect 521 10329 755 10331
rect 4549 10563 4783 10565
rect 4549 10499 4550 10563
rect 4614 10499 4634 10563
rect 4698 10499 4718 10563
rect 4782 10499 4783 10563
rect 4549 10479 4783 10499
rect 4549 10415 4550 10479
rect 4614 10415 4634 10479
rect 4698 10415 4718 10479
rect 4782 10415 4783 10479
rect 4549 10395 4783 10415
rect 4549 10331 4550 10395
rect 4614 10331 4634 10395
rect 4698 10331 4718 10395
rect 4782 10331 4783 10395
rect 4549 10329 4783 10331
rect 8170 10563 8404 10565
rect 8170 10499 8171 10563
rect 8235 10499 8255 10563
rect 8319 10499 8339 10563
rect 8403 10499 8404 10563
rect 8170 10479 8404 10499
rect 8170 10415 8171 10479
rect 8235 10415 8255 10479
rect 8319 10415 8339 10479
rect 8403 10415 8404 10479
rect 8170 10395 8404 10415
rect 8170 10331 8171 10395
rect 8235 10331 8255 10395
rect 8319 10331 8339 10395
rect 8403 10331 8404 10395
rect 8170 10329 8404 10331
rect 9185 10563 9419 10565
rect 9185 10499 9186 10563
rect 9250 10499 9270 10563
rect 9334 10499 9354 10563
rect 9418 10499 9419 10563
rect 9185 10479 9419 10499
rect 9185 10415 9186 10479
rect 9250 10415 9270 10479
rect 9334 10415 9354 10479
rect 9418 10415 9419 10479
rect 9185 10395 9419 10415
rect 9185 10331 9186 10395
rect 9250 10331 9270 10395
rect 9334 10331 9354 10395
rect 9418 10331 9419 10395
rect 9185 10329 9419 10331
rect 15746 10329 16000 10565
rect 0 9673 254 10269
rect 15746 9673 16000 10269
rect 0 9547 254 9613
rect 521 9612 755 9613
rect 521 9548 522 9612
rect 586 9548 606 9612
rect 670 9548 690 9612
rect 754 9548 755 9612
rect 521 9547 755 9548
rect 4549 9612 4783 9613
rect 4549 9548 4550 9612
rect 4614 9548 4634 9612
rect 4698 9548 4718 9612
rect 4782 9548 4783 9612
rect 4549 9547 4783 9548
rect 8170 9612 8404 9613
rect 8170 9548 8171 9612
rect 8235 9548 8255 9612
rect 8319 9548 8339 9612
rect 8403 9548 8404 9612
rect 8170 9547 8404 9548
rect 9185 9612 9419 9613
rect 9185 9548 9186 9612
rect 9250 9548 9270 9612
rect 9334 9548 9354 9612
rect 9418 9548 9419 9612
rect 9185 9547 9419 9548
rect 15746 9547 16000 9613
rect 1137 9472 12274 9473
rect 1137 9408 1138 9472
rect 1202 9408 1218 9472
rect 1282 9408 12128 9472
rect 12192 9408 12209 9472
rect 12273 9408 12274 9472
rect 1137 9407 12274 9408
rect 0 8317 254 9247
rect 2780 9246 3772 9247
rect 2780 9182 2782 9246
rect 2846 9182 2866 9246
rect 2930 9182 2950 9246
rect 3014 9182 3034 9246
rect 3098 9182 3118 9246
rect 3182 9182 3202 9246
rect 3266 9182 3286 9246
rect 3350 9182 3370 9246
rect 3434 9182 3454 9246
rect 3518 9182 3538 9246
rect 3602 9182 3622 9246
rect 3686 9182 3706 9246
rect 3770 9182 3772 9246
rect 8600 9241 8862 9242
rect 2780 9160 3772 9182
rect 2780 9096 2782 9160
rect 2846 9096 2866 9160
rect 2930 9096 2950 9160
rect 3014 9096 3034 9160
rect 3098 9096 3118 9160
rect 3182 9096 3202 9160
rect 3266 9096 3286 9160
rect 3350 9096 3370 9160
rect 3434 9096 3454 9160
rect 3518 9096 3538 9160
rect 3602 9096 3622 9160
rect 3686 9096 3706 9160
rect 3770 9096 3772 9160
rect 2780 9074 3772 9096
rect 2780 9010 2782 9074
rect 2846 9010 2866 9074
rect 2930 9010 2950 9074
rect 3014 9010 3034 9074
rect 3098 9010 3118 9074
rect 3182 9010 3202 9074
rect 3266 9010 3286 9074
rect 3350 9010 3370 9074
rect 3434 9010 3454 9074
rect 3518 9010 3538 9074
rect 3602 9010 3622 9074
rect 3686 9010 3706 9074
rect 3770 9010 3772 9074
rect 2780 8988 3772 9010
rect 2780 8924 2782 8988
rect 2846 8924 2866 8988
rect 2930 8924 2950 8988
rect 3014 8924 3034 8988
rect 3098 8924 3118 8988
rect 3182 8924 3202 8988
rect 3266 8924 3286 8988
rect 3350 8924 3370 8988
rect 3434 8924 3454 8988
rect 3518 8924 3538 8988
rect 3602 8924 3622 8988
rect 3686 8924 3706 8988
rect 3770 8924 3772 8988
rect 2780 8902 3772 8924
rect 2780 8838 2782 8902
rect 2846 8838 2866 8902
rect 2930 8838 2950 8902
rect 3014 8838 3034 8902
rect 3098 8838 3118 8902
rect 3182 8838 3202 8902
rect 3266 8838 3286 8902
rect 3350 8838 3370 8902
rect 3434 8838 3454 8902
rect 3518 8838 3538 8902
rect 3602 8838 3622 8902
rect 3686 8838 3706 8902
rect 3770 8838 3772 8902
rect 2780 8816 3772 8838
rect 2780 8752 2782 8816
rect 2846 8752 2866 8816
rect 2930 8752 2950 8816
rect 3014 8752 3034 8816
rect 3098 8752 3118 8816
rect 3182 8752 3202 8816
rect 3266 8752 3286 8816
rect 3350 8752 3370 8816
rect 3434 8752 3454 8816
rect 3518 8752 3538 8816
rect 3602 8752 3622 8816
rect 3686 8752 3706 8816
rect 3770 8752 3772 8816
rect 2780 8730 3772 8752
rect 2780 8666 2782 8730
rect 2846 8666 2866 8730
rect 2930 8666 2950 8730
rect 3014 8666 3034 8730
rect 3098 8666 3118 8730
rect 3182 8666 3202 8730
rect 3266 8666 3286 8730
rect 3350 8666 3370 8730
rect 3434 8666 3454 8730
rect 3518 8666 3538 8730
rect 3602 8666 3622 8730
rect 3686 8666 3706 8730
rect 3770 8666 3772 8730
rect 2780 8643 3772 8666
rect 2780 8579 2782 8643
rect 2846 8579 2866 8643
rect 2930 8579 2950 8643
rect 3014 8579 3034 8643
rect 3098 8579 3118 8643
rect 3182 8579 3202 8643
rect 3266 8579 3286 8643
rect 3350 8579 3370 8643
rect 3434 8579 3454 8643
rect 3518 8579 3538 8643
rect 3602 8579 3622 8643
rect 3686 8579 3706 8643
rect 3770 8579 3772 8643
rect 2780 8556 3772 8579
rect 2780 8492 2782 8556
rect 2846 8492 2866 8556
rect 2930 8492 2950 8556
rect 3014 8492 3034 8556
rect 3098 8492 3118 8556
rect 3182 8492 3202 8556
rect 3266 8492 3286 8556
rect 3350 8492 3370 8556
rect 3434 8492 3454 8556
rect 3518 8492 3538 8556
rect 3602 8492 3622 8556
rect 3686 8492 3706 8556
rect 3770 8492 3772 8556
rect 2780 8469 3772 8492
rect 2780 8405 2782 8469
rect 2846 8405 2866 8469
rect 2930 8405 2950 8469
rect 3014 8405 3034 8469
rect 3098 8405 3118 8469
rect 3182 8405 3202 8469
rect 3266 8405 3286 8469
rect 3350 8405 3370 8469
rect 3434 8405 3454 8469
rect 3518 8405 3538 8469
rect 3602 8405 3622 8469
rect 3686 8405 3706 8469
rect 3770 8405 3772 8469
rect 2780 8382 3772 8405
rect 2780 8318 2782 8382
rect 2846 8318 2866 8382
rect 2930 8318 2950 8382
rect 3014 8318 3034 8382
rect 3098 8318 3118 8382
rect 3182 8318 3202 8382
rect 3266 8318 3286 8382
rect 3350 8318 3370 8382
rect 3434 8318 3454 8382
rect 3518 8318 3538 8382
rect 3602 8318 3622 8382
rect 3686 8318 3706 8382
rect 3770 8318 3772 8382
rect 6915 9238 7177 9239
rect 6915 9174 6916 9238
rect 6980 9174 7014 9238
rect 7078 9174 7112 9238
rect 7176 9174 7177 9238
rect 6915 9153 7177 9174
rect 6915 9089 6916 9153
rect 6980 9089 7014 9153
rect 7078 9089 7112 9153
rect 7176 9089 7177 9153
rect 6915 9068 7177 9089
rect 6915 9004 6916 9068
rect 6980 9004 7014 9068
rect 7078 9004 7112 9068
rect 7176 9004 7177 9068
rect 6915 8983 7177 9004
rect 6915 8919 6916 8983
rect 6980 8919 7014 8983
rect 7078 8919 7112 8983
rect 7176 8919 7177 8983
rect 6915 8898 7177 8919
rect 6915 8834 6916 8898
rect 6980 8834 7014 8898
rect 7078 8834 7112 8898
rect 7176 8834 7177 8898
rect 6915 8813 7177 8834
rect 6915 8749 6916 8813
rect 6980 8749 7014 8813
rect 7078 8749 7112 8813
rect 7176 8749 7177 8813
rect 6915 8728 7177 8749
rect 6915 8664 6916 8728
rect 6980 8664 7014 8728
rect 7078 8664 7112 8728
rect 7176 8664 7177 8728
rect 6915 8643 7177 8664
rect 6915 8579 6916 8643
rect 6980 8579 7014 8643
rect 7078 8579 7112 8643
rect 7176 8579 7177 8643
rect 6915 8558 7177 8579
rect 6915 8494 6916 8558
rect 6980 8494 7014 8558
rect 7078 8494 7112 8558
rect 7176 8494 7177 8558
rect 6915 8472 7177 8494
rect 6915 8408 6916 8472
rect 6980 8408 7014 8472
rect 7078 8408 7112 8472
rect 7176 8408 7177 8472
rect 6915 8386 7177 8408
rect 6915 8322 6916 8386
rect 6980 8322 7014 8386
rect 7078 8322 7112 8386
rect 7176 8322 7177 8386
rect 6915 8321 7177 8322
rect 8600 9177 8601 9241
rect 8665 9177 8699 9241
rect 8763 9177 8797 9241
rect 8861 9177 8862 9241
rect 8600 9156 8862 9177
rect 8600 9092 8601 9156
rect 8665 9092 8699 9156
rect 8763 9092 8797 9156
rect 8861 9092 8862 9156
rect 8600 9070 8862 9092
rect 8600 9006 8601 9070
rect 8665 9006 8699 9070
rect 8763 9006 8797 9070
rect 8861 9006 8862 9070
rect 8600 8984 8862 9006
rect 8600 8920 8601 8984
rect 8665 8920 8699 8984
rect 8763 8920 8797 8984
rect 8861 8920 8862 8984
rect 8600 8898 8862 8920
rect 8600 8834 8601 8898
rect 8665 8834 8699 8898
rect 8763 8834 8797 8898
rect 8861 8834 8862 8898
rect 8600 8812 8862 8834
rect 8600 8748 8601 8812
rect 8665 8748 8699 8812
rect 8763 8748 8797 8812
rect 8861 8748 8862 8812
rect 8600 8726 8862 8748
rect 8600 8662 8601 8726
rect 8665 8662 8699 8726
rect 8763 8662 8797 8726
rect 8861 8662 8862 8726
rect 8600 8640 8862 8662
rect 8600 8576 8601 8640
rect 8665 8576 8699 8640
rect 8763 8576 8797 8640
rect 8861 8576 8862 8640
rect 8600 8554 8862 8576
rect 8600 8490 8601 8554
rect 8665 8490 8699 8554
rect 8763 8490 8797 8554
rect 8861 8490 8862 8554
rect 8600 8468 8862 8490
rect 8600 8404 8601 8468
rect 8665 8404 8699 8468
rect 8763 8404 8797 8468
rect 8861 8404 8862 8468
rect 8600 8382 8862 8404
rect 2780 8317 3772 8318
rect 8600 8318 8601 8382
rect 8665 8318 8699 8382
rect 8763 8318 8797 8382
rect 8861 8318 8862 8382
rect 9108 9241 9688 9242
rect 9108 9177 9114 9241
rect 9178 9177 9198 9241
rect 9262 9177 9282 9241
rect 9346 9177 9366 9241
rect 9430 9177 9450 9241
rect 9514 9177 9534 9241
rect 9598 9177 9618 9241
rect 9682 9177 9688 9241
rect 9108 9156 9688 9177
rect 9108 9092 9114 9156
rect 9178 9092 9198 9156
rect 9262 9092 9282 9156
rect 9346 9092 9366 9156
rect 9430 9092 9450 9156
rect 9514 9092 9534 9156
rect 9598 9092 9618 9156
rect 9682 9092 9688 9156
rect 9108 9071 9688 9092
rect 9108 9007 9114 9071
rect 9178 9007 9198 9071
rect 9262 9007 9282 9071
rect 9346 9007 9366 9071
rect 9430 9007 9450 9071
rect 9514 9007 9534 9071
rect 9598 9007 9618 9071
rect 9682 9007 9688 9071
rect 9108 8986 9688 9007
rect 9108 8922 9114 8986
rect 9178 8922 9198 8986
rect 9262 8922 9282 8986
rect 9346 8922 9366 8986
rect 9430 8922 9450 8986
rect 9514 8922 9534 8986
rect 9598 8922 9618 8986
rect 9682 8922 9688 8986
rect 9108 8901 9688 8922
rect 9108 8837 9114 8901
rect 9178 8837 9198 8901
rect 9262 8837 9282 8901
rect 9346 8837 9366 8901
rect 9430 8837 9450 8901
rect 9514 8837 9534 8901
rect 9598 8837 9618 8901
rect 9682 8837 9688 8901
rect 9108 8816 9688 8837
rect 9108 8752 9114 8816
rect 9178 8752 9198 8816
rect 9262 8752 9282 8816
rect 9346 8752 9366 8816
rect 9430 8752 9450 8816
rect 9514 8752 9534 8816
rect 9598 8752 9618 8816
rect 9682 8752 9688 8816
rect 9108 8731 9688 8752
rect 9108 8667 9114 8731
rect 9178 8667 9198 8731
rect 9262 8667 9282 8731
rect 9346 8667 9366 8731
rect 9430 8667 9450 8731
rect 9514 8667 9534 8731
rect 9598 8667 9618 8731
rect 9682 8667 9688 8731
rect 9108 8645 9688 8667
rect 9108 8581 9114 8645
rect 9178 8581 9198 8645
rect 9262 8581 9282 8645
rect 9346 8581 9366 8645
rect 9430 8581 9450 8645
rect 9514 8581 9534 8645
rect 9598 8581 9618 8645
rect 9682 8581 9688 8645
rect 9108 8559 9688 8581
rect 9108 8495 9114 8559
rect 9178 8495 9198 8559
rect 9262 8495 9282 8559
rect 9346 8495 9366 8559
rect 9430 8495 9450 8559
rect 9514 8495 9534 8559
rect 9598 8495 9618 8559
rect 9682 8495 9688 8559
rect 9108 8473 9688 8495
rect 9108 8409 9114 8473
rect 9178 8409 9198 8473
rect 9262 8409 9282 8473
rect 9346 8409 9366 8473
rect 9430 8409 9450 8473
rect 9514 8409 9534 8473
rect 9598 8409 9618 8473
rect 9682 8409 9688 8473
rect 9108 8387 9688 8409
rect 9108 8323 9114 8387
rect 9178 8323 9198 8387
rect 9262 8323 9282 8387
rect 9346 8323 9366 8387
rect 9430 8323 9450 8387
rect 9514 8323 9534 8387
rect 9598 8323 9618 8387
rect 9682 8323 9688 8387
rect 10497 9238 11147 9239
rect 10497 9174 10503 9238
rect 10567 9174 10585 9238
rect 10649 9174 10667 9238
rect 10731 9174 10749 9238
rect 10813 9174 10831 9238
rect 10895 9174 10913 9238
rect 10977 9174 10995 9238
rect 11059 9174 11077 9238
rect 11141 9174 11147 9238
rect 10497 9154 11147 9174
rect 10497 9090 10503 9154
rect 10567 9090 10585 9154
rect 10649 9090 10667 9154
rect 10731 9090 10749 9154
rect 10813 9090 10831 9154
rect 10895 9090 10913 9154
rect 10977 9090 10995 9154
rect 11059 9090 11077 9154
rect 11141 9090 11147 9154
rect 10497 9070 11147 9090
rect 10497 9006 10503 9070
rect 10567 9006 10585 9070
rect 10649 9006 10667 9070
rect 10731 9006 10749 9070
rect 10813 9006 10831 9070
rect 10895 9006 10913 9070
rect 10977 9006 10995 9070
rect 11059 9006 11077 9070
rect 11141 9006 11147 9070
rect 10497 8986 11147 9006
rect 10497 8922 10503 8986
rect 10567 8922 10585 8986
rect 10649 8922 10667 8986
rect 10731 8922 10749 8986
rect 10813 8922 10831 8986
rect 10895 8922 10913 8986
rect 10977 8922 10995 8986
rect 11059 8922 11077 8986
rect 11141 8922 11147 8986
rect 10497 8902 11147 8922
rect 10497 8838 10503 8902
rect 10567 8838 10585 8902
rect 10649 8838 10667 8902
rect 10731 8838 10749 8902
rect 10813 8838 10831 8902
rect 10895 8838 10913 8902
rect 10977 8838 10995 8902
rect 11059 8838 11077 8902
rect 11141 8838 11147 8902
rect 10497 8818 11147 8838
rect 10497 8754 10503 8818
rect 10567 8754 10585 8818
rect 10649 8754 10667 8818
rect 10731 8754 10749 8818
rect 10813 8754 10831 8818
rect 10895 8754 10913 8818
rect 10977 8754 10995 8818
rect 11059 8754 11077 8818
rect 11141 8754 11147 8818
rect 10497 8734 11147 8754
rect 10497 8670 10503 8734
rect 10567 8670 10585 8734
rect 10649 8670 10667 8734
rect 10731 8670 10749 8734
rect 10813 8670 10831 8734
rect 10895 8670 10913 8734
rect 10977 8670 10995 8734
rect 11059 8670 11077 8734
rect 11141 8670 11147 8734
rect 10497 8650 11147 8670
rect 10497 8586 10503 8650
rect 10567 8586 10585 8650
rect 10649 8586 10667 8650
rect 10731 8586 10749 8650
rect 10813 8586 10831 8650
rect 10895 8586 10913 8650
rect 10977 8586 10995 8650
rect 11059 8586 11077 8650
rect 11141 8586 11147 8650
rect 10497 8566 11147 8586
rect 10497 8502 10503 8566
rect 10567 8502 10585 8566
rect 10649 8502 10667 8566
rect 10731 8502 10749 8566
rect 10813 8502 10831 8566
rect 10895 8502 10913 8566
rect 10977 8502 10995 8566
rect 11059 8502 11077 8566
rect 11141 8502 11147 8566
rect 10497 8482 11147 8502
rect 10497 8418 10503 8482
rect 10567 8418 10585 8482
rect 10649 8418 10667 8482
rect 10731 8418 10749 8482
rect 10813 8418 10831 8482
rect 10895 8418 10913 8482
rect 10977 8418 10995 8482
rect 11059 8418 11077 8482
rect 11141 8418 11147 8482
rect 10497 8397 11147 8418
rect 10497 8333 10503 8397
rect 10567 8333 10585 8397
rect 10649 8333 10667 8397
rect 10731 8333 10749 8397
rect 10813 8333 10831 8397
rect 10895 8333 10913 8397
rect 10977 8333 10995 8397
rect 11059 8333 11077 8397
rect 11141 8333 11147 8397
rect 10497 8332 11147 8333
rect 9108 8322 9688 8323
rect 8600 8317 8862 8318
rect 15746 8317 16000 9247
rect 0 7347 254 8037
rect 12673 8030 13463 8037
rect 4331 7989 4730 7992
rect 4331 7925 4332 7989
rect 4396 7925 4416 7989
rect 4480 7925 4499 7989
rect 4563 7925 4582 7989
rect 4646 7925 4665 7989
rect 4729 7925 4730 7989
rect 4331 7922 4730 7925
rect 12673 7966 12674 8030
rect 12738 7966 12755 8030
rect 12819 7966 12836 8030
rect 12900 7966 12917 8030
rect 12981 7966 12998 8030
rect 13062 7966 13078 8030
rect 13142 7966 13158 8030
rect 13222 7966 13238 8030
rect 13302 7966 13318 8030
rect 13382 7966 13398 8030
rect 13462 7966 13463 8030
rect 12673 7944 13463 7966
rect 4414 7904 4730 7907
rect 4414 7840 4415 7904
rect 4479 7840 4499 7904
rect 4563 7840 4582 7904
rect 4646 7840 4665 7904
rect 4729 7840 4730 7904
rect 4414 7837 4730 7840
rect 12673 7880 12674 7944
rect 12738 7880 12755 7944
rect 12819 7880 12836 7944
rect 12900 7880 12917 7944
rect 12981 7880 12998 7944
rect 13062 7880 13078 7944
rect 13142 7880 13158 7944
rect 13222 7880 13238 7944
rect 13302 7880 13318 7944
rect 13382 7880 13398 7944
rect 13462 7880 13463 7944
rect 12673 7858 13463 7880
rect 4495 7818 4730 7821
rect 4495 7754 4496 7818
rect 4560 7754 4581 7818
rect 4645 7754 4665 7818
rect 4729 7754 4730 7818
rect 4495 7751 4730 7754
rect 12673 7794 12674 7858
rect 12738 7794 12755 7858
rect 12819 7794 12836 7858
rect 12900 7794 12917 7858
rect 12981 7794 12998 7858
rect 13062 7794 13078 7858
rect 13142 7794 13158 7858
rect 13222 7794 13238 7858
rect 13302 7794 13318 7858
rect 13382 7794 13398 7858
rect 13462 7794 13463 7858
rect 12673 7772 13463 7794
rect 12673 7708 12674 7772
rect 12738 7708 12755 7772
rect 12819 7708 12836 7772
rect 12900 7708 12917 7772
rect 12981 7708 12998 7772
rect 13062 7708 13078 7772
rect 13142 7708 13158 7772
rect 13222 7708 13238 7772
rect 13302 7708 13318 7772
rect 13382 7708 13398 7772
rect 13462 7708 13463 7772
rect 4577 7698 4730 7701
rect 4577 7634 4578 7698
rect 4642 7634 4665 7698
rect 4729 7634 4730 7698
rect 4577 7631 4730 7634
rect 12673 7686 13463 7708
rect 12673 7622 12674 7686
rect 12738 7622 12755 7686
rect 12819 7622 12836 7686
rect 12900 7622 12917 7686
rect 12981 7622 12998 7686
rect 13062 7622 13078 7686
rect 13142 7622 13158 7686
rect 13222 7622 13238 7686
rect 13302 7622 13318 7686
rect 13382 7622 13398 7686
rect 13462 7622 13463 7686
rect 12673 7600 13463 7622
rect 12673 7536 12674 7600
rect 12738 7536 12755 7600
rect 12819 7536 12836 7600
rect 12900 7536 12917 7600
rect 12981 7536 12998 7600
rect 13062 7536 13078 7600
rect 13142 7536 13158 7600
rect 13222 7536 13238 7600
rect 13302 7536 13318 7600
rect 13382 7536 13398 7600
rect 13462 7536 13463 7600
rect 12673 7514 13463 7536
rect 12673 7450 12674 7514
rect 12738 7450 12755 7514
rect 12819 7450 12836 7514
rect 12900 7450 12917 7514
rect 12981 7450 12998 7514
rect 13062 7450 13078 7514
rect 13142 7450 13158 7514
rect 13222 7450 13238 7514
rect 13302 7450 13318 7514
rect 13382 7450 13398 7514
rect 13462 7450 13463 7514
rect 12673 7428 13463 7450
rect 12673 7364 12674 7428
rect 12738 7364 12755 7428
rect 12819 7364 12836 7428
rect 12900 7364 12917 7428
rect 12981 7364 12998 7428
rect 13062 7364 13078 7428
rect 13142 7364 13158 7428
rect 13222 7364 13238 7428
rect 13302 7364 13318 7428
rect 13382 7364 13398 7428
rect 13462 7364 13463 7428
rect 12673 7357 13463 7364
rect 15746 7347 16000 8037
rect 910 7238 9527 7239
rect 910 7174 911 7238
rect 975 7174 991 7238
rect 1055 7174 9382 7238
rect 9446 7174 9462 7238
rect 9526 7174 9527 7238
rect 910 7173 9527 7174
rect 9597 7238 9960 7239
rect 9597 7174 9598 7238
rect 9662 7174 9678 7238
rect 9742 7174 9815 7238
rect 9879 7174 9895 7238
rect 9959 7174 9960 7238
rect 9597 7173 9960 7174
rect 0 6377 254 7067
rect 4451 7066 4773 7067
rect 4451 7002 4454 7066
rect 4518 7002 4538 7066
rect 4602 7002 4622 7066
rect 4686 7002 4706 7066
rect 4770 7002 4773 7066
rect 4451 6980 4773 7002
rect 4451 6916 4454 6980
rect 4518 6916 4538 6980
rect 4602 6916 4622 6980
rect 4686 6916 4706 6980
rect 4770 6916 4773 6980
rect 4451 6894 4773 6916
rect 4451 6830 4454 6894
rect 4518 6830 4538 6894
rect 4602 6830 4622 6894
rect 4686 6830 4706 6894
rect 4770 6830 4773 6894
rect 4451 6807 4773 6830
rect 4451 6743 4454 6807
rect 4518 6743 4538 6807
rect 4602 6743 4622 6807
rect 4686 6743 4706 6807
rect 4770 6743 4773 6807
rect 4451 6720 4773 6743
rect 4451 6656 4454 6720
rect 4518 6656 4538 6720
rect 4602 6656 4622 6720
rect 4686 6656 4706 6720
rect 4770 6656 4773 6720
rect 4451 6633 4773 6656
rect 4451 6569 4454 6633
rect 4518 6569 4538 6633
rect 4602 6569 4622 6633
rect 4686 6569 4706 6633
rect 4770 6569 4773 6633
rect 4451 6546 4773 6569
rect 4451 6482 4454 6546
rect 4518 6482 4538 6546
rect 4602 6482 4622 6546
rect 4686 6482 4706 6546
rect 4770 6482 4773 6546
rect 4451 6459 4773 6482
rect 4451 6395 4454 6459
rect 4518 6395 4538 6459
rect 4602 6395 4622 6459
rect 4686 6395 4706 6459
rect 4770 6395 4773 6459
rect 4451 6394 4773 6395
rect 15746 6377 16000 7067
rect 0 5167 254 6097
rect 15746 5167 16000 6097
rect 0 3957 254 4887
rect 1484 4886 2140 4887
rect 1484 4822 1486 4886
rect 1550 4822 1570 4886
rect 1634 4822 1654 4886
rect 1718 4822 1738 4886
rect 1802 4822 1822 4886
rect 1886 4822 1906 4886
rect 1970 4822 1990 4886
rect 2054 4822 2074 4886
rect 2138 4822 2140 4886
rect 1484 4800 2140 4822
rect 1484 4736 1486 4800
rect 1550 4736 1570 4800
rect 1634 4736 1654 4800
rect 1718 4736 1738 4800
rect 1802 4736 1822 4800
rect 1886 4736 1906 4800
rect 1970 4736 1990 4800
rect 2054 4736 2074 4800
rect 2138 4736 2140 4800
rect 1484 4714 2140 4736
rect 1484 4650 1486 4714
rect 1550 4650 1570 4714
rect 1634 4650 1654 4714
rect 1718 4650 1738 4714
rect 1802 4650 1822 4714
rect 1886 4650 1906 4714
rect 1970 4650 1990 4714
rect 2054 4650 2074 4714
rect 2138 4650 2140 4714
rect 1484 4628 2140 4650
rect 1484 4564 1486 4628
rect 1550 4564 1570 4628
rect 1634 4564 1654 4628
rect 1718 4564 1738 4628
rect 1802 4564 1822 4628
rect 1886 4564 1906 4628
rect 1970 4564 1990 4628
rect 2054 4564 2074 4628
rect 2138 4564 2140 4628
rect 1484 4542 2140 4564
rect 1484 4478 1486 4542
rect 1550 4478 1570 4542
rect 1634 4478 1654 4542
rect 1718 4478 1738 4542
rect 1802 4478 1822 4542
rect 1886 4478 1906 4542
rect 1970 4478 1990 4542
rect 2054 4478 2074 4542
rect 2138 4478 2140 4542
rect 1484 4456 2140 4478
rect 1484 4392 1486 4456
rect 1550 4392 1570 4456
rect 1634 4392 1654 4456
rect 1718 4392 1738 4456
rect 1802 4392 1822 4456
rect 1886 4392 1906 4456
rect 1970 4392 1990 4456
rect 2054 4392 2074 4456
rect 2138 4392 2140 4456
rect 1484 4370 2140 4392
rect 1484 4306 1486 4370
rect 1550 4306 1570 4370
rect 1634 4306 1654 4370
rect 1718 4306 1738 4370
rect 1802 4306 1822 4370
rect 1886 4306 1906 4370
rect 1970 4306 1990 4370
rect 2054 4306 2074 4370
rect 2138 4306 2140 4370
rect 1484 4283 2140 4306
rect 1484 4219 1486 4283
rect 1550 4219 1570 4283
rect 1634 4219 1654 4283
rect 1718 4219 1738 4283
rect 1802 4219 1822 4283
rect 1886 4219 1906 4283
rect 1970 4219 1990 4283
rect 2054 4219 2074 4283
rect 2138 4219 2140 4283
rect 1484 4196 2140 4219
rect 1484 4132 1486 4196
rect 1550 4132 1570 4196
rect 1634 4132 1654 4196
rect 1718 4132 1738 4196
rect 1802 4132 1822 4196
rect 1886 4132 1906 4196
rect 1970 4132 1990 4196
rect 2054 4132 2074 4196
rect 2138 4132 2140 4196
rect 1484 4109 2140 4132
rect 1484 4045 1486 4109
rect 1550 4045 1570 4109
rect 1634 4045 1654 4109
rect 1718 4045 1738 4109
rect 1802 4045 1822 4109
rect 1886 4045 1906 4109
rect 1970 4045 1990 4109
rect 2054 4045 2074 4109
rect 2138 4045 2140 4109
rect 1484 4022 2140 4045
rect 1484 3958 1486 4022
rect 1550 3958 1570 4022
rect 1634 3958 1654 4022
rect 1718 3958 1738 4022
rect 1802 3958 1822 4022
rect 1886 3958 1906 4022
rect 1970 3958 1990 4022
rect 2054 3958 2074 4022
rect 2138 3958 2140 4022
rect 14138 4881 14348 4882
rect 14138 4817 14139 4881
rect 14203 4817 14283 4881
rect 14347 4817 14348 4881
rect 14138 4796 14348 4817
rect 14138 4732 14139 4796
rect 14203 4732 14283 4796
rect 14347 4732 14348 4796
rect 14138 4711 14348 4732
rect 14138 4647 14139 4711
rect 14203 4647 14283 4711
rect 14347 4647 14348 4711
rect 14138 4626 14348 4647
rect 14138 4562 14139 4626
rect 14203 4562 14283 4626
rect 14347 4562 14348 4626
rect 14138 4541 14348 4562
rect 14138 4477 14139 4541
rect 14203 4477 14283 4541
rect 14347 4477 14348 4541
rect 14138 4456 14348 4477
rect 14138 4392 14139 4456
rect 14203 4392 14283 4456
rect 14347 4392 14348 4456
rect 14138 4371 14348 4392
rect 14138 4307 14139 4371
rect 14203 4307 14283 4371
rect 14347 4307 14348 4371
rect 14138 4286 14348 4307
rect 14138 4222 14139 4286
rect 14203 4222 14283 4286
rect 14347 4222 14348 4286
rect 14138 4201 14348 4222
rect 14138 4137 14139 4201
rect 14203 4137 14283 4201
rect 14347 4137 14348 4201
rect 14138 4115 14348 4137
rect 14138 4051 14139 4115
rect 14203 4051 14283 4115
rect 14347 4051 14348 4115
rect 14138 4029 14348 4051
rect 14138 3965 14139 4029
rect 14203 3965 14283 4029
rect 14347 3965 14348 4029
rect 14138 3964 14348 3965
rect 1484 3957 2140 3958
rect 15746 3957 16000 4887
rect 0 2987 193 3677
rect 4912 3676 5528 3677
rect 4912 3612 4918 3676
rect 4982 3612 5008 3676
rect 5072 3612 5098 3676
rect 5162 3612 5188 3676
rect 5252 3612 5278 3676
rect 5342 3612 5368 3676
rect 5432 3612 5458 3676
rect 5522 3612 5528 3676
rect 4912 3590 5528 3612
rect 4912 3526 4918 3590
rect 4982 3526 5008 3590
rect 5072 3526 5098 3590
rect 5162 3526 5188 3590
rect 5252 3526 5278 3590
rect 5342 3526 5368 3590
rect 5432 3526 5458 3590
rect 5522 3526 5528 3590
rect 4912 3503 5528 3526
rect 4912 3439 4918 3503
rect 4982 3439 5008 3503
rect 5072 3439 5098 3503
rect 5162 3439 5188 3503
rect 5252 3439 5278 3503
rect 5342 3439 5368 3503
rect 5432 3439 5458 3503
rect 5522 3439 5528 3503
rect 4912 3416 5528 3439
rect 4912 3352 4918 3416
rect 4982 3352 5008 3416
rect 5072 3352 5098 3416
rect 5162 3352 5188 3416
rect 5252 3352 5278 3416
rect 5342 3352 5368 3416
rect 5432 3352 5458 3416
rect 5522 3352 5528 3416
rect 4912 3329 5528 3352
rect 4912 3265 4918 3329
rect 4982 3265 5008 3329
rect 5072 3265 5098 3329
rect 5162 3265 5188 3329
rect 5252 3265 5278 3329
rect 5342 3265 5368 3329
rect 5432 3265 5458 3329
rect 5522 3265 5528 3329
rect 4912 3242 5528 3265
rect 4912 3178 4918 3242
rect 4982 3178 5008 3242
rect 5072 3178 5098 3242
rect 5162 3178 5188 3242
rect 5252 3178 5278 3242
rect 5342 3178 5368 3242
rect 5432 3178 5458 3242
rect 5522 3178 5528 3242
rect 4912 3155 5528 3178
rect 4912 3091 4918 3155
rect 4982 3091 5008 3155
rect 5072 3091 5098 3155
rect 5162 3091 5188 3155
rect 5252 3091 5278 3155
rect 5342 3091 5368 3155
rect 5432 3091 5458 3155
rect 5522 3091 5528 3155
rect 4912 3068 5528 3091
rect 4912 3004 4918 3068
rect 4982 3004 5008 3068
rect 5072 3004 5098 3068
rect 5162 3004 5188 3068
rect 5252 3004 5278 3068
rect 5342 3004 5368 3068
rect 5432 3004 5458 3068
rect 5522 3004 5528 3068
rect 4912 3003 5528 3004
rect 10024 3676 10316 3677
rect 10024 3612 10026 3676
rect 10090 3612 10138 3676
rect 10202 3612 10250 3676
rect 10314 3612 10316 3676
rect 10024 3590 10316 3612
rect 10024 3526 10026 3590
rect 10090 3526 10138 3590
rect 10202 3526 10250 3590
rect 10314 3526 10316 3590
rect 10024 3503 10316 3526
rect 10024 3439 10026 3503
rect 10090 3439 10138 3503
rect 10202 3439 10250 3503
rect 10314 3439 10316 3503
rect 10024 3416 10316 3439
rect 10024 3352 10026 3416
rect 10090 3352 10138 3416
rect 10202 3352 10250 3416
rect 10314 3352 10316 3416
rect 10024 3329 10316 3352
rect 10024 3265 10026 3329
rect 10090 3265 10138 3329
rect 10202 3265 10250 3329
rect 10314 3265 10316 3329
rect 10024 3242 10316 3265
rect 10024 3178 10026 3242
rect 10090 3178 10138 3242
rect 10202 3178 10250 3242
rect 10314 3178 10316 3242
rect 10024 3155 10316 3178
rect 10024 3091 10026 3155
rect 10090 3091 10138 3155
rect 10202 3091 10250 3155
rect 10314 3091 10316 3155
rect 10024 3068 10316 3091
rect 10024 3004 10026 3068
rect 10090 3004 10138 3068
rect 10202 3004 10250 3068
rect 10314 3004 10316 3068
rect 10024 3003 10316 3004
rect 15807 2987 16000 3677
rect 0 1777 254 2707
rect 6846 2706 7072 2707
rect 6846 2642 6847 2706
rect 6911 2642 6927 2706
rect 6991 2642 7007 2706
rect 7071 2642 7072 2706
rect 6846 2620 7072 2642
rect 6846 2556 6847 2620
rect 6911 2556 6927 2620
rect 6991 2556 7007 2620
rect 7071 2556 7072 2620
rect 6846 2534 7072 2556
rect 6846 2470 6847 2534
rect 6911 2470 6927 2534
rect 6991 2470 7007 2534
rect 7071 2470 7072 2534
rect 6846 2448 7072 2470
rect 6846 2384 6847 2448
rect 6911 2384 6927 2448
rect 6991 2384 7007 2448
rect 7071 2384 7072 2448
rect 6846 2362 7072 2384
rect 6846 2298 6847 2362
rect 6911 2298 6927 2362
rect 6991 2298 7007 2362
rect 7071 2298 7072 2362
rect 6846 2276 7072 2298
rect 6846 2212 6847 2276
rect 6911 2212 6927 2276
rect 6991 2212 7007 2276
rect 7071 2212 7072 2276
rect 6846 2190 7072 2212
rect 6846 2126 6847 2190
rect 6911 2126 6927 2190
rect 6991 2126 7007 2190
rect 7071 2126 7072 2190
rect 6846 2103 7072 2126
rect 6846 2039 6847 2103
rect 6911 2039 6927 2103
rect 6991 2039 7007 2103
rect 7071 2039 7072 2103
rect 6846 2016 7072 2039
rect 6846 1952 6847 2016
rect 6911 1952 6927 2016
rect 6991 1952 7007 2016
rect 7071 1952 7072 2016
rect 6846 1929 7072 1952
rect 6846 1865 6847 1929
rect 6911 1865 6927 1929
rect 6991 1865 7007 1929
rect 7071 1865 7072 1929
rect 6846 1842 7072 1865
rect 6846 1778 6847 1842
rect 6911 1778 6927 1842
rect 6991 1778 7007 1842
rect 7071 1778 7072 1842
rect 8609 2706 8781 2707
rect 8609 2642 8610 2706
rect 8674 2642 8716 2706
rect 8780 2642 8781 2706
rect 8609 2621 8781 2642
rect 8609 2557 8610 2621
rect 8674 2557 8716 2621
rect 8780 2557 8781 2621
rect 8609 2536 8781 2557
rect 8609 2472 8610 2536
rect 8674 2472 8716 2536
rect 8780 2472 8781 2536
rect 8609 2450 8781 2472
rect 8609 2386 8610 2450
rect 8674 2386 8716 2450
rect 8780 2386 8781 2450
rect 8609 2364 8781 2386
rect 8609 2300 8610 2364
rect 8674 2300 8716 2364
rect 8780 2300 8781 2364
rect 8609 2278 8781 2300
rect 8609 2214 8610 2278
rect 8674 2214 8716 2278
rect 8780 2214 8781 2278
rect 8609 2192 8781 2214
rect 8609 2128 8610 2192
rect 8674 2128 8716 2192
rect 8780 2128 8781 2192
rect 8609 2106 8781 2128
rect 8609 2042 8610 2106
rect 8674 2042 8716 2106
rect 8780 2042 8781 2106
rect 8609 2020 8781 2042
rect 8609 1956 8610 2020
rect 8674 1956 8716 2020
rect 8780 1956 8781 2020
rect 8609 1934 8781 1956
rect 8609 1870 8610 1934
rect 8674 1870 8716 1934
rect 8780 1870 8781 1934
rect 8609 1848 8781 1870
rect 8609 1784 8610 1848
rect 8674 1784 8716 1848
rect 8780 1784 8781 1848
rect 11340 2706 11708 2707
rect 11340 2642 11342 2706
rect 11406 2642 11442 2706
rect 11506 2642 11542 2706
rect 11606 2642 11642 2706
rect 11706 2642 11708 2706
rect 11340 2621 11708 2642
rect 11340 2557 11342 2621
rect 11406 2557 11442 2621
rect 11506 2557 11542 2621
rect 11606 2557 11642 2621
rect 11706 2557 11708 2621
rect 11340 2536 11708 2557
rect 11340 2472 11342 2536
rect 11406 2472 11442 2536
rect 11506 2472 11542 2536
rect 11606 2472 11642 2536
rect 11706 2472 11708 2536
rect 11340 2451 11708 2472
rect 11340 2387 11342 2451
rect 11406 2387 11442 2451
rect 11506 2387 11542 2451
rect 11606 2387 11642 2451
rect 11706 2387 11708 2451
rect 11340 2366 11708 2387
rect 11340 2302 11342 2366
rect 11406 2302 11442 2366
rect 11506 2302 11542 2366
rect 11606 2302 11642 2366
rect 11706 2302 11708 2366
rect 11340 2280 11708 2302
rect 11340 2216 11342 2280
rect 11406 2216 11442 2280
rect 11506 2216 11542 2280
rect 11606 2216 11642 2280
rect 11706 2216 11708 2280
rect 11340 2194 11708 2216
rect 11340 2130 11342 2194
rect 11406 2130 11442 2194
rect 11506 2130 11542 2194
rect 11606 2130 11642 2194
rect 11706 2130 11708 2194
rect 11340 2108 11708 2130
rect 11340 2044 11342 2108
rect 11406 2044 11442 2108
rect 11506 2044 11542 2108
rect 11606 2044 11642 2108
rect 11706 2044 11708 2108
rect 11340 2022 11708 2044
rect 11340 1958 11342 2022
rect 11406 1958 11442 2022
rect 11506 1958 11542 2022
rect 11606 1958 11642 2022
rect 11706 1958 11708 2022
rect 11340 1936 11708 1958
rect 11340 1872 11342 1936
rect 11406 1872 11442 1936
rect 11506 1872 11542 1936
rect 11606 1872 11642 1936
rect 11706 1872 11708 1936
rect 11340 1850 11708 1872
rect 11340 1786 11342 1850
rect 11406 1786 11442 1850
rect 11506 1786 11542 1850
rect 11606 1786 11642 1850
rect 11706 1786 11708 1850
rect 11340 1785 11708 1786
rect 13565 2706 14057 2707
rect 13565 2642 13569 2706
rect 13633 2642 13653 2706
rect 13717 2642 13737 2706
rect 13801 2642 13821 2706
rect 13885 2642 13905 2706
rect 13969 2642 13989 2706
rect 14053 2642 14057 2706
rect 13565 2621 14057 2642
rect 13565 2557 13569 2621
rect 13633 2557 13653 2621
rect 13717 2557 13737 2621
rect 13801 2557 13821 2621
rect 13885 2557 13905 2621
rect 13969 2557 13989 2621
rect 14053 2557 14057 2621
rect 13565 2535 14057 2557
rect 13565 2471 13569 2535
rect 13633 2471 13653 2535
rect 13717 2471 13737 2535
rect 13801 2471 13821 2535
rect 13885 2471 13905 2535
rect 13969 2471 13989 2535
rect 14053 2471 14057 2535
rect 13565 2449 14057 2471
rect 13565 2385 13569 2449
rect 13633 2385 13653 2449
rect 13717 2385 13737 2449
rect 13801 2385 13821 2449
rect 13885 2385 13905 2449
rect 13969 2385 13989 2449
rect 14053 2385 14057 2449
rect 13565 2363 14057 2385
rect 13565 2299 13569 2363
rect 13633 2299 13653 2363
rect 13717 2299 13737 2363
rect 13801 2299 13821 2363
rect 13885 2299 13905 2363
rect 13969 2299 13989 2363
rect 14053 2299 14057 2363
rect 13565 2277 14057 2299
rect 13565 2213 13569 2277
rect 13633 2213 13653 2277
rect 13717 2213 13737 2277
rect 13801 2213 13821 2277
rect 13885 2213 13905 2277
rect 13969 2213 13989 2277
rect 14053 2213 14057 2277
rect 13565 2191 14057 2213
rect 13565 2127 13569 2191
rect 13633 2127 13653 2191
rect 13717 2127 13737 2191
rect 13801 2127 13821 2191
rect 13885 2127 13905 2191
rect 13969 2127 13989 2191
rect 14053 2127 14057 2191
rect 13565 2105 14057 2127
rect 13565 2041 13569 2105
rect 13633 2041 13653 2105
rect 13717 2041 13737 2105
rect 13801 2041 13821 2105
rect 13885 2041 13905 2105
rect 13969 2041 13989 2105
rect 14053 2041 14057 2105
rect 13565 2019 14057 2041
rect 13565 1955 13569 2019
rect 13633 1955 13653 2019
rect 13717 1955 13737 2019
rect 13801 1955 13821 2019
rect 13885 1955 13905 2019
rect 13969 1955 13989 2019
rect 14053 1955 14057 2019
rect 13565 1933 14057 1955
rect 13565 1869 13569 1933
rect 13633 1869 13653 1933
rect 13717 1869 13737 1933
rect 13801 1869 13821 1933
rect 13885 1869 13905 1933
rect 13969 1869 13989 1933
rect 14053 1869 14057 1933
rect 13565 1847 14057 1869
rect 8609 1783 8781 1784
rect 13565 1783 13569 1847
rect 13633 1783 13653 1847
rect 13717 1783 13737 1847
rect 13801 1783 13821 1847
rect 13885 1783 13905 1847
rect 13969 1783 13989 1847
rect 14053 1783 14057 1847
rect 13565 1782 14057 1783
rect 6846 1777 7072 1778
rect 15746 1777 16000 2707
rect 0 407 254 1497
rect 2225 1496 2699 1497
rect 2225 1432 2230 1496
rect 2294 1432 2310 1496
rect 2374 1432 2390 1496
rect 2454 1432 2470 1496
rect 2534 1432 2550 1496
rect 2614 1432 2630 1496
rect 2694 1432 2699 1496
rect 2225 1412 2699 1432
rect 2225 1348 2230 1412
rect 2294 1348 2310 1412
rect 2374 1348 2390 1412
rect 2454 1348 2470 1412
rect 2534 1348 2550 1412
rect 2614 1348 2630 1412
rect 2694 1348 2699 1412
rect 2225 1328 2699 1348
rect 2225 1264 2230 1328
rect 2294 1264 2310 1328
rect 2374 1264 2390 1328
rect 2454 1264 2470 1328
rect 2534 1264 2550 1328
rect 2614 1264 2630 1328
rect 2694 1264 2699 1328
rect 2225 1244 2699 1264
rect 2225 1180 2230 1244
rect 2294 1180 2310 1244
rect 2374 1180 2390 1244
rect 2454 1180 2470 1244
rect 2534 1180 2550 1244
rect 2614 1180 2630 1244
rect 2694 1180 2699 1244
rect 2225 1160 2699 1180
rect 2225 1096 2230 1160
rect 2294 1096 2310 1160
rect 2374 1096 2390 1160
rect 2454 1096 2470 1160
rect 2534 1096 2550 1160
rect 2614 1096 2630 1160
rect 2694 1096 2699 1160
rect 2225 1076 2699 1096
rect 2225 1012 2230 1076
rect 2294 1012 2310 1076
rect 2374 1012 2390 1076
rect 2454 1012 2470 1076
rect 2534 1012 2550 1076
rect 2614 1012 2630 1076
rect 2694 1012 2699 1076
rect 2225 992 2699 1012
rect 2225 928 2230 992
rect 2294 928 2310 992
rect 2374 928 2390 992
rect 2454 928 2470 992
rect 2534 928 2550 992
rect 2614 928 2630 992
rect 2694 928 2699 992
rect 2225 908 2699 928
rect 2225 844 2230 908
rect 2294 844 2310 908
rect 2374 844 2390 908
rect 2454 844 2470 908
rect 2534 844 2550 908
rect 2614 844 2630 908
rect 2694 844 2699 908
rect 2225 823 2699 844
rect 2225 759 2230 823
rect 2294 759 2310 823
rect 2374 759 2390 823
rect 2454 759 2470 823
rect 2534 759 2550 823
rect 2614 759 2630 823
rect 2694 759 2699 823
rect 2225 738 2699 759
rect 2225 674 2230 738
rect 2294 674 2310 738
rect 2374 674 2390 738
rect 2454 674 2470 738
rect 2534 674 2550 738
rect 2614 674 2630 738
rect 2694 674 2699 738
rect 2225 653 2699 674
rect 2225 589 2230 653
rect 2294 589 2310 653
rect 2374 589 2390 653
rect 2454 589 2470 653
rect 2534 589 2550 653
rect 2614 589 2630 653
rect 2694 589 2699 653
rect 2225 568 2699 589
rect 2225 504 2230 568
rect 2294 504 2310 568
rect 2374 504 2390 568
rect 2454 504 2470 568
rect 2534 504 2550 568
rect 2614 504 2630 568
rect 2694 504 2699 568
rect 14428 1486 15372 1487
rect 14428 1422 14438 1486
rect 14502 1422 14524 1486
rect 14588 1422 14610 1486
rect 14674 1422 14696 1486
rect 14760 1422 14782 1486
rect 14846 1422 14868 1486
rect 14932 1422 14954 1486
rect 15018 1422 15040 1486
rect 15104 1422 15126 1486
rect 15190 1422 15212 1486
rect 15276 1422 15298 1486
rect 15362 1422 15372 1486
rect 14428 1401 15372 1422
rect 14428 1337 14438 1401
rect 14502 1337 14524 1401
rect 14588 1337 14610 1401
rect 14674 1337 14696 1401
rect 14760 1337 14782 1401
rect 14846 1337 14868 1401
rect 14932 1337 14954 1401
rect 15018 1337 15040 1401
rect 15104 1337 15126 1401
rect 15190 1337 15212 1401
rect 15276 1337 15298 1401
rect 15362 1337 15372 1401
rect 14428 1316 15372 1337
rect 14428 1252 14438 1316
rect 14502 1252 14524 1316
rect 14588 1252 14610 1316
rect 14674 1252 14696 1316
rect 14760 1252 14782 1316
rect 14846 1252 14868 1316
rect 14932 1252 14954 1316
rect 15018 1252 15040 1316
rect 15104 1252 15126 1316
rect 15190 1252 15212 1316
rect 15276 1252 15298 1316
rect 15362 1252 15372 1316
rect 14428 1230 15372 1252
rect 14428 1166 14438 1230
rect 14502 1166 14524 1230
rect 14588 1166 14610 1230
rect 14674 1166 14696 1230
rect 14760 1166 14782 1230
rect 14846 1166 14868 1230
rect 14932 1166 14954 1230
rect 15018 1166 15040 1230
rect 15104 1166 15126 1230
rect 15190 1166 15212 1230
rect 15276 1166 15298 1230
rect 15362 1166 15372 1230
rect 14428 1144 15372 1166
rect 14428 1080 14438 1144
rect 14502 1080 14524 1144
rect 14588 1080 14610 1144
rect 14674 1080 14696 1144
rect 14760 1080 14782 1144
rect 14846 1080 14868 1144
rect 14932 1080 14954 1144
rect 15018 1080 15040 1144
rect 15104 1080 15126 1144
rect 15190 1080 15212 1144
rect 15276 1080 15298 1144
rect 15362 1080 15372 1144
rect 14428 1058 15372 1080
rect 14428 994 14438 1058
rect 14502 994 14524 1058
rect 14588 994 14610 1058
rect 14674 994 14696 1058
rect 14760 994 14782 1058
rect 14846 994 14868 1058
rect 14932 994 14954 1058
rect 15018 994 15040 1058
rect 15104 994 15126 1058
rect 15190 994 15212 1058
rect 15276 994 15298 1058
rect 15362 994 15372 1058
rect 14428 972 15372 994
rect 14428 908 14438 972
rect 14502 908 14524 972
rect 14588 908 14610 972
rect 14674 908 14696 972
rect 14760 908 14782 972
rect 14846 908 14868 972
rect 14932 908 14954 972
rect 15018 908 15040 972
rect 15104 908 15126 972
rect 15190 908 15212 972
rect 15276 908 15298 972
rect 15362 908 15372 972
rect 14428 886 15372 908
rect 14428 822 14438 886
rect 14502 822 14524 886
rect 14588 822 14610 886
rect 14674 822 14696 886
rect 14760 822 14782 886
rect 14846 822 14868 886
rect 14932 822 14954 886
rect 15018 822 15040 886
rect 15104 822 15126 886
rect 15190 822 15212 886
rect 15276 822 15298 886
rect 15362 822 15372 886
rect 14428 800 15372 822
rect 14428 736 14438 800
rect 14502 736 14524 800
rect 14588 736 14610 800
rect 14674 736 14696 800
rect 14760 736 14782 800
rect 14846 736 14868 800
rect 14932 736 14954 800
rect 15018 736 15040 800
rect 15104 736 15126 800
rect 15190 736 15212 800
rect 15276 736 15298 800
rect 15362 736 15372 800
rect 14428 714 15372 736
rect 14428 650 14438 714
rect 14502 650 14524 714
rect 14588 650 14610 714
rect 14674 650 14696 714
rect 14760 650 14782 714
rect 14846 650 14868 714
rect 14932 650 14954 714
rect 15018 650 15040 714
rect 15104 650 15126 714
rect 15190 650 15212 714
rect 15276 650 15298 714
rect 15362 650 15372 714
rect 14428 628 15372 650
rect 14428 564 14438 628
rect 14502 564 14524 628
rect 14588 564 14610 628
rect 14674 564 14696 628
rect 14760 564 14782 628
rect 14846 564 14868 628
rect 14932 564 14954 628
rect 15018 564 15040 628
rect 15104 564 15126 628
rect 15190 564 15212 628
rect 15276 564 15298 628
rect 15362 564 15372 628
rect 14428 563 15372 564
rect 2225 483 2699 504
rect 2225 419 2230 483
rect 2294 419 2310 483
rect 2374 419 2390 483
rect 2454 419 2470 483
rect 2534 419 2550 483
rect 2614 419 2630 483
rect 2694 419 2699 483
rect 2225 418 2699 419
rect 15746 407 16000 1497
rect 290 298 10488 299
rect 290 234 291 298
rect 355 234 371 298
rect 435 234 10343 298
rect 10407 234 10423 298
rect 10487 234 10488 298
rect 290 233 10488 234
rect 10713 298 11352 299
rect 10713 234 10714 298
rect 10778 234 10794 298
rect 10858 234 11207 298
rect 11271 234 11287 298
rect 11351 234 11352 298
rect 10713 233 11352 234
rect 13012 298 13463 299
rect 13012 234 13013 298
rect 13077 234 13093 298
rect 13157 234 13318 298
rect 13382 234 13398 298
rect 13462 234 13463 298
rect 13012 233 13463 234
rect 15029 298 15633 299
rect 15029 234 15030 298
rect 15094 234 15110 298
rect 15174 234 15488 298
rect 15552 234 15568 298
rect 15632 234 15633 298
rect 15029 233 15633 234
<< rmetal4 >>
rect 1460 21317 1467 23791
<< metal5 >>
rect 6423 25094 10731 29403
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1623348570
transform 1 0 13851 0 -1 792
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1623348570
transform 0 1 14463 1 0 884
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1623348570
transform 0 1 15482 1 0 884
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1623348570
transform 0 1 14982 1 0 884
box 0 0 882 404
use sky130_fd_io__gpio_opathv2  sky130_fd_io__gpio_opathv2_0
timestamp 1623348570
transform 1 0 815 0 1 3971
box -873 -2766 15315 31850
use sky130_fd_io__gpiov2_ctl  sky130_fd_io__gpiov2_ctl_0
timestamp 1623348570
transform 1 0 -3504 0 1 -3498
box 3421 3498 18546 11377
use sky130_fd_io__gpiov2_ipath  sky130_fd_io__gpiov2_ipath_0
timestamp 1623348570
transform 1 0 0 0 1 0
box 0 -136 16004 40000
use sky130_fd_io__gpiov2_amux  sky130_fd_io__gpiov2_amux_0
timestamp 1623348570
transform 1 0 1000 0 1 10260
box -1143 -10153 15134 9892
use sky130_fd_io__overlay_gpiov2_m4  sky130_fd_io__overlay_gpiov2_m4_0
timestamp 1623348570
transform 1 0 0 0 1 0
box 0 407 16000 40000
<< labels >>
flabel metal5 s 6423 25094 10731 29403 3 FreeSans 520 0 0 0 PAD
port 1 nsew signal bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 2 nsew ground bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 3 nsew signal bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 4 nsew signal bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 8 nsew ground bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 9 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 10 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 11 nsew power bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 13 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 400 21317 587 23791 3 FreeSans 520 0 0 0 PAD_A_NOESD_H
port 14 nsew signal bidirectional
flabel metal4 s 15746 7347 16000 8037 3 FreeSans 520 180 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 15746 8317 16000 9247 3 FreeSans 520 180 0 0 VSSD
port 2 nsew ground bidirectional
flabel metal4 s 15746 9673 16000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 3 nsew signal bidirectional
flabel metal4 s 15746 10625 16000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 4 nsew signal bidirectional
flabel metal4 s 15746 12817 16000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal4 s 15746 14007 16000 19000 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 15746 6377 16000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 15746 5167 16000 6097 3 FreeSans 520 180 0 0 VSSIO
port 8 nsew ground bidirectional
flabel metal4 s 15746 3957 16000 4887 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 15807 2987 16000 3677 3 FreeSans 520 180 0 0 VDDA
port 9 nsew power bidirectional
flabel metal4 s 15746 1777 16000 2707 3 FreeSans 520 180 0 0 VCCD
port 10 nsew power bidirectional
flabel metal4 s 15746 407 16000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 11 nsew power bidirectional
flabel metal4 s 15746 35157 16000 40000 3 FreeSans 520 180 0 0 VSSIO
port 8 nsew ground bidirectional
flabel metal4 s 15746 11281 16000 11347 3 FreeSans 520 180 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 15746 11647 16000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 13 nsew ground bidirectional
flabel metal4 s 15746 9547 16000 9613 3 FreeSans 520 180 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 15746 10329 16000 10565 3 FreeSans 520 180 0 0 VSSA
port 12 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 8 nsew ground bidirectional
flabel metal3 s 12564 0 12778 147 3 FreeSans 520 90 0 0 PAD_A_NOESD_H
port 14 nsew signal bidirectional
flabel metal3 s 9173 0 9239 52 3 FreeSans 520 90 0 0 ANALOG_POL
port 15 nsew signal input
flabel metal3 s 15716 0 15782 153 3 FreeSans 520 90 0 0 ENABLE_VDDIO
port 16 nsew signal input
flabel metal3 s 80 0 204 163 3 FreeSans 520 0 0 0 IN_H
port 17 nsew signal output
flabel metal3 s 15848 0 15914 163 3 FreeSans 520 0 0 0 IN
port 18 nsew signal output
flabel metal1 s 12486 0 12538 56 3 FreeSans 520 90 0 0 ANALOG_EN
port 19 nsew signal input
flabel metal2 s 4471 0 4523 67 0 FreeSans 400 0 0 0 OUT
port 20 nsew signal input
flabel metal2 s 15741 0 15781 44 3 FreeSans 520 90 0 0 TIE_HI_ESD
port 21 nsew signal output
flabel metal2 s 13655 0 13785 44 3 FreeSans 520 90 0 0 PAD_A_ESD_1_H
port 22 nsew signal bidirectional
flabel metal2 s 9971 0 10023 52 3 FreeSans 520 90 0 0 DM[0]
port 23 nsew signal input
flabel metal2 s 13367 0 13419 52 3 FreeSans 520 90 0 0 DM[1]
port 24 nsew signal input
flabel metal2 s 5698 0 5750 52 3 FreeSans 520 90 0 0 DM[2]
port 25 nsew signal input
flabel metal2 s 6363 0 6415 44 3 FreeSans 520 90 0 0 HLD_H_N
port 26 nsew signal input
flabel metal2 s 5320 0 5372 28 3 FreeSans 520 90 0 0 HLD_OVR
port 27 nsew signal input
flabel metal2 s 9049 0 9101 52 3 FreeSans 520 90 0 0 INP_DIS
port 28 nsew signal input
flabel metal2 s 2551 0 2603 44 3 FreeSans 520 90 0 0 ENABLE_VDDA_H
port 29 nsew signal input
flabel metal2 s 1226 0 1278 52 3 FreeSans 520 90 0 0 VTRIP_SEL
port 30 nsew signal input
flabel metal2 s 675 0 721 46 7 FreeSans 300 270 0 0 OE_N
port 31 nsew signal input
flabel metal2 s 15522 0 15574 44 3 FreeSans 520 90 0 0 SLOW
port 32 nsew signal input
flabel metal2 s 15943 0 15983 192 0 FreeSans 400 90 0 0 TIE_LO_ESD
port 33 nsew signal output
flabel metal2 s 15256 0 15384 44 3 FreeSans 520 90 0 0 PAD_A_ESD_0_H
port 34 nsew signal bidirectional
flabel metal2 s 6150 0 6202 56 3 FreeSans 520 90 0 0 ANALOG_SEL
port 35 nsew signal input
flabel metal2 s 7678 0 7730 89 3 FreeSans 520 90 0 0 ENABLE_INP_H
port 36 nsew signal input
flabel metal2 s 13683 22 13683 22 3 FreeSans 520 90 0 0 PAD_A_ESD_1_H
port 22 nsew
flabel metal2 s 15761 22 15761 22 3 FreeSans 520 90 0 0 TIE_HI_ESD
port 21 nsew
flabel metal2 s 7092 0 7144 56 3 FreeSans 520 90 0 0 ENABLE_H
port 37 nsew signal input
flabel metal2 s 1084 0 1130 79 3 FreeSans 520 90 0 0 IB_MODE_SEL
port 38 nsew signal input
flabel metal2 s 3262 0 3314 101 3 FreeSans 520 90 0 0 ENABLE_VSWITCH_H
port 39 nsew signal input
flabel comment s 13227 270 13227 270 0 FreeSans 200 0 0 0 ANTENNA FIX
flabel comment s 3335 37099 3335 37099 0 FreeSans 4000 0 0 0 VSSD
flabel comment s 1647 38266 1647 38266 0 FreeSans 4000 0 0 0 VDDIO_Q
flabel comment s 14714 37057 14714 37057 0 FreeSans 4000 0 0 0 VCCHIB
flabel comment s 5710 11509 5710 11509 0 FreeSans 200 0 0 0 ANTENNA FIX
flabel comment s 11003 274 11003 274 0 FreeSans 200 0 0 0 ANTENNA FIX
flabel comment s 15363 273 15363 273 0 FreeSans 200 0 0 0 ANTENNA FIX
rlabel metal2 s 13682 21 13684 23 1 PAD_A_ESD_1_H
port 22 nsew signal bidirectional
rlabel metal4 s 1503 23791 1714 24002 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1533 23791 2500 23821 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1563 23821 2500 23851 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1566 21242 1641 21317 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1570 21313 2500 21317 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1593 23851 2500 23881 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1600 21283 2500 21313 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1623 23881 2500 23911 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1641 21006 1877 21242 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1653 23911 2500 23941 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1660 21223 2500 21253 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1683 23941 2500 23971 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1690 21193 2500 21223 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1714 24002 1960 24248 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1720 21163 2500 21193 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1743 24001 2500 24031 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1750 21133 2500 21163 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1773 24031 2500 24061 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1780 21103 2500 21133 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1803 24061 2500 24091 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1810 21073 2500 21103 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1833 24091 2500 24121 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1840 21043 2500 21073 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1863 24121 2500 24151 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1877 20879 2004 21006 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1893 24151 2500 24181 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1900 20983 2500 21013 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1923 24181 2500 24211 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1930 20953 2500 20983 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1962 24241 2500 24250 1 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal2 s 15760 21 15762 23 1 TIE_HI_ESD
port 21 nsew signal output
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 16000 40000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string LEFsymmetry X Y R90
string GDS_END 8058748
string GDS_START 6287582
string MASKHINTS_HVI 1346 17198 5828 19224 13700 1890 15920 2360 24 17522 1778 20612
<< end >>
