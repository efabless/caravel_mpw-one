magic
tech sky130A
magscale 12 1
timestamp 1606780629
<< metal5 >>
rect 10 100 30 105
rect 5 95 30 100
rect 0 85 30 95
rect 0 20 15 85
rect 0 10 30 20
rect 5 5 30 10
rect 10 0 30 5
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
