magic
tech sky130A
magscale 1 2
timestamp 1625189325
<< fillblock >>
rect -262 -266 31304 2764
rect -140 -5140 35048 -1424
rect 26 -9464 13144 -6358
use font_20  font_20_4 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598785497
transform 1 0 12476 0 1 -9176
box 0 0 1 1
use font_47  font_47_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765398
transform 1 0 118 0 1 -4282
box 0 0 1080 2520
use font_6F  font_6F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777049
transform 1 0 1558 0 1 -4282
box 0 0 1080 1800
use font_6F  font_6F_1
timestamp 1598777049
transform 1 0 2998 0 1 -4282
box 0 0 1080 1800
use font_67  font_67_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776042
transform 1 0 4438 0 1 -4282
box 0 -720 1080 1800
use font_65  font_65_3 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775915
transform 1 0 6598 0 1 -4282
box 0 0 1080 1800
use font_6C  font_6C_2 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776550
transform 1 0 5878 0 1 -4282
box 0 0 360 2520
use font_53  font_53_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768855
transform 1 0 9838 0 1 -4282
box 0 0 1080 2520
use font_79  font_79_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777870
transform 1 0 12718 0 1 -4282
box 0 -720 1080 1800
use font_6B  font_6B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776472
transform 1 0 11278 0 1 -4282
box 0 0 1080 2520
use font_57  font_57_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769216
transform 1 0 14158 0 1 -4282
box 0 0 1800 2520
use font_74  font_74_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777367
transform 1 0 17758 0 1 -4282
box 0 0 1080 2160
use font_61  font_61_3 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775307
transform 1 0 16318 0 1 -4282
box 0 0 1080 1800
use font_65  font_65_4
timestamp 1598775915
transform 1 0 19198 0 1 -4282
box 0 0 1080 1800
use font_72  font_72_1 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777237
transform 1 0 20638 0 1 -4282
box 0 0 1080 1800
use font_20  font_20_2
timestamp 1598785497
transform 1 0 22078 0 1 -5002
box 0 0 1 1
use font_6F  font_6F_2
timestamp 1598777049
transform 1 0 23518 0 1 -4282
box 0 0 1080 1800
use font_65  font_65_5
timestamp 1598775915
transform 1 0 26398 0 1 -4282
box 0 0 1080 1800
use font_70  font_70_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777090
transform 1 0 24958 0 1 -4282
box 0 -720 1080 1800
use font_6E  font_6E_2 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776997
transform 1 0 27814 0 1 -4311
box 0 0 1080 1800
use font_20  font_20_3
timestamp 1598785497
transform 1 0 29278 0 1 -5362
box 0 0 1 1
use font_50  font_50_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 30718 0 1 -4282
box 0 0 1080 2520
use font_44  font_44_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763661
transform 1 0 32158 0 1 -4282
box 0 0 1080 2520
use font_4B  font_4B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766293
transform 1 0 33598 0 1 -4282
box 0 0 1080 2520
use font_2D  font_2D_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786817
transform 1 0 8038 0 1 -4642
box 0 1080 1440 1440
use font_61  font_61_0
timestamp 1598775307
transform 1 0 1440 0 1 0
box 0 0 1080 1800
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 0 0 1 0
box 0 0 1080 2520
use font_72  font_72_0
timestamp 1598777237
transform 1 0 2880 0 1 0
box 0 0 1080 1800
use font_61  font_61_1
timestamp 1598775307
transform 1 0 4320 0 1 0
box 0 0 1080 1800
use font_61  font_61_4
timestamp 1598775307
transform 1 0 7235 0 1 15
box 0 0 1080 1800
use font_76  font_76_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777472
transform 1 0 5760 0 1 0
box 0 0 1080 1800
use font_6E  font_6E_1
timestamp 1598776997
transform 1 0 8740 0 1 0
box 0 0 1080 1800
use font_20  font_20_0
timestamp 1598785497
transform 1 0 9360 0 1 0
box 0 0 1 1
use font_31  font_31_1 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787010
transform 1 0 12539 0 1 -1
box 0 0 1080 2520
use font_28  font_28_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1606780629
transform 1 0 15200 0 1 0
box 0 0 720 2520
use font_20  font_20_1
timestamp 1598785497
transform 1 0 14400 0 1 0
box 0 0 1 1
use font_29  font_29_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786350
transform 1 0 17720 0 1 0
box 0 0 720 2520
use font_43  font_43_1
timestamp 1598763351
transform 1 0 16280 0 1 0
box 0 0 1080 2520
use font_65  font_65_1
timestamp 1598775915
transform 1 0 20240 0 1 0
box 0 0 1080 1800
use font_61  font_61_2
timestamp 1598775307
transform 1 0 23120 0 1 0
box 0 0 1080 1800
use font_66  font_66_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775974
transform 1 0 21680 0 1 0
box 0 0 1080 2520
use font_6C  font_6C_1
timestamp 1598776550
transform 1 0 26000 0 1 0
box 0 0 360 2520
use font_62  font_62_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775406
transform 1 0 24560 0 1 0
box 0 0 1080 2520
use font_73  font_73_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777283
transform 1 0 28160 0 1 0
box 0 0 1080 1800
use font_65  font_65_2
timestamp 1598775915
transform 1 0 26720 0 1 0
box 0 0 1080 1800
use font_73  font_73_1
timestamp 1598777283
transform 1 0 29600 0 1 0
box 0 0 1080 1800
use font_56  font_56_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769117
transform 1 0 11128 0 1 15
box 0 0 1080 2520
use font_31  font_31_0
timestamp 1598787010
transform 1 0 11550 0 1 -9341
box 0 0 1080 2520
use font_32  font_32_1 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787041
transform 1 0 10116 0 1 -9321
box 0 0 1080 2520
use font_30  font_30_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786981
transform 1 0 8676 0 1 -9321
box 0 0 1080 2520
use font_32  font_32_0
timestamp 1598787041
transform 1 0 7236 0 1 -9321
box 0 0 1080 2520
use font_65  font_65_9
timestamp 1598775915
transform 1 0 4569 0 1 -9290
box 0 0 1080 1800
use font_6E  font_6E_0
timestamp 1598776997
transform 1 0 3142 0 1 -9290
box 0 0 1080 1800
use font_75  font_75_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777411
transform 1 0 1700 0 1 -9274
box 0 0 1080 1800
use font_4A  font_4A_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766195
transform 1 0 226 0 1 -9274
box 0 0 1080 2520
<< end >>
