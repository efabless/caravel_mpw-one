magic
tech sky130A
magscale 1 2
timestamp 1606790418
<< obsli1 >>
rect 1104 2159 428812 169983
<< metal1 >>
rect 1104 167504 428812 167600
rect 1104 166960 428812 167056
<< obsm1 >>
rect 566 167656 429350 169992
rect 566 167448 1048 167656
rect 428868 167448 429350 167656
rect 566 167112 429350 167448
rect 566 166904 1048 167112
rect 428868 166904 429350 167112
rect 566 620 429350 166904
<< metal2 >>
rect 570 169200 626 170000
rect 938 169200 994 170000
rect 1306 169200 1362 170000
rect 1674 169200 1730 170000
rect 2042 169200 2098 170000
rect 2410 169200 2466 170000
rect 2778 169200 2834 170000
rect 3146 169200 3202 170000
rect 3514 169200 3570 170000
rect 3882 169200 3938 170000
rect 4250 169200 4306 170000
rect 4618 169200 4674 170000
rect 4986 169200 5042 170000
rect 5354 169200 5410 170000
rect 5722 169200 5778 170000
rect 6090 169200 6146 170000
rect 6458 169200 6514 170000
rect 6826 169200 6882 170000
rect 7194 169200 7250 170000
rect 7562 169200 7618 170000
rect 7930 169200 7986 170000
rect 8298 169200 8354 170000
rect 8666 169200 8722 170000
rect 9034 169200 9090 170000
rect 9402 169200 9458 170000
rect 9770 169200 9826 170000
rect 10138 169200 10194 170000
rect 10506 169200 10562 170000
rect 10874 169200 10930 170000
rect 11242 169200 11298 170000
rect 37370 169200 37426 170000
rect 88890 169200 88946 170000
rect 114282 169200 114338 170000
rect 139306 169200 139362 170000
rect 140410 169200 140466 170000
rect 140778 169200 140834 170000
rect 141146 169200 141202 170000
rect 141514 169200 141570 170000
rect 141882 169200 141938 170000
rect 142250 169200 142306 170000
rect 142618 169200 142674 170000
rect 142986 169200 143042 170000
rect 143354 169200 143410 170000
rect 143722 169200 143778 170000
rect 144090 169200 144146 170000
rect 144458 169200 144514 170000
rect 144826 169200 144882 170000
rect 145194 169200 145250 170000
rect 145562 169200 145618 170000
rect 145930 169200 145986 170000
rect 146298 169200 146354 170000
rect 146666 169200 146722 170000
rect 147034 169200 147090 170000
rect 147402 169200 147458 170000
rect 147770 169200 147826 170000
rect 148138 169200 148194 170000
rect 148506 169200 148562 170000
rect 148874 169200 148930 170000
rect 149242 169200 149298 170000
rect 149610 169200 149666 170000
rect 149978 169200 150034 170000
rect 150346 169200 150402 170000
rect 150714 169200 150770 170000
rect 151082 169200 151138 170000
rect 151450 169200 151506 170000
rect 151818 169200 151874 170000
rect 152186 169200 152242 170000
rect 152554 169200 152610 170000
rect 152922 169200 152978 170000
rect 153290 169200 153346 170000
rect 153658 169200 153714 170000
rect 154026 169200 154082 170000
rect 154394 169200 154450 170000
rect 154762 169200 154818 170000
rect 155130 169200 155186 170000
rect 155498 169200 155554 170000
rect 155866 169200 155922 170000
rect 156234 169200 156290 170000
rect 156602 169200 156658 170000
rect 156970 169200 157026 170000
rect 157338 169200 157394 170000
rect 157706 169200 157762 170000
rect 158074 169200 158130 170000
rect 158442 169200 158498 170000
rect 158810 169200 158866 170000
rect 159178 169200 159234 170000
rect 159546 169200 159602 170000
rect 159914 169200 159970 170000
rect 160282 169200 160338 170000
rect 160650 169200 160706 170000
rect 161018 169200 161074 170000
rect 161386 169200 161442 170000
rect 161754 169200 161810 170000
rect 162122 169200 162178 170000
rect 162490 169200 162546 170000
rect 162858 169200 162914 170000
rect 163226 169200 163282 170000
rect 163594 169200 163650 170000
rect 163962 169200 164018 170000
rect 164330 169200 164386 170000
rect 164698 169200 164754 170000
rect 165066 169200 165122 170000
rect 165434 169200 165490 170000
rect 165802 169200 165858 170000
rect 166170 169200 166226 170000
rect 166538 169200 166594 170000
rect 166906 169200 166962 170000
rect 167274 169200 167330 170000
rect 167642 169200 167698 170000
rect 168010 169200 168066 170000
rect 168378 169200 168434 170000
rect 168746 169200 168802 170000
rect 169114 169200 169170 170000
rect 169482 169200 169538 170000
rect 169850 169200 169906 170000
rect 170218 169200 170274 170000
rect 170586 169200 170642 170000
rect 170954 169200 171010 170000
rect 171322 169200 171378 170000
rect 171690 169200 171746 170000
rect 172058 169200 172114 170000
rect 172426 169200 172482 170000
rect 172794 169200 172850 170000
rect 173162 169200 173218 170000
rect 173530 169200 173586 170000
rect 173898 169200 173954 170000
rect 174266 169200 174322 170000
rect 174634 169200 174690 170000
rect 175002 169200 175058 170000
rect 175370 169200 175426 170000
rect 175738 169200 175794 170000
rect 176106 169200 176162 170000
rect 176474 169200 176530 170000
rect 176842 169200 176898 170000
rect 177210 169200 177266 170000
rect 177578 169200 177634 170000
rect 177946 169200 178002 170000
rect 178314 169200 178370 170000
rect 178682 169200 178738 170000
rect 179050 169200 179106 170000
rect 179418 169200 179474 170000
rect 179786 169200 179842 170000
rect 180154 169200 180210 170000
rect 180522 169200 180578 170000
rect 180890 169200 180946 170000
rect 181258 169200 181314 170000
rect 181626 169200 181682 170000
rect 181994 169200 182050 170000
rect 182362 169200 182418 170000
rect 182730 169200 182786 170000
rect 183098 169200 183154 170000
rect 183466 169200 183522 170000
rect 183834 169200 183890 170000
rect 184202 169200 184258 170000
rect 184570 169200 184626 170000
rect 184938 169200 184994 170000
rect 185306 169200 185362 170000
rect 185674 169200 185730 170000
rect 186042 169200 186098 170000
rect 186410 169200 186466 170000
rect 186778 169200 186834 170000
rect 187146 169200 187202 170000
rect 187514 169200 187570 170000
rect 187882 169200 187938 170000
rect 188250 169200 188306 170000
rect 188618 169200 188674 170000
rect 188986 169200 189042 170000
rect 189354 169200 189410 170000
rect 189722 169200 189778 170000
rect 190090 169200 190146 170000
rect 190458 169200 190514 170000
rect 190826 169200 190882 170000
rect 191194 169200 191250 170000
rect 191562 169200 191618 170000
rect 191930 169200 191986 170000
rect 192298 169200 192354 170000
rect 192666 169200 192722 170000
rect 193034 169200 193090 170000
rect 193402 169200 193458 170000
rect 193770 169200 193826 170000
rect 194138 169200 194194 170000
rect 194506 169200 194562 170000
rect 194874 169200 194930 170000
rect 195242 169200 195298 170000
rect 195610 169200 195666 170000
rect 195978 169200 196034 170000
rect 196346 169200 196402 170000
rect 196714 169200 196770 170000
rect 197082 169200 197138 170000
rect 197450 169200 197506 170000
rect 197818 169200 197874 170000
rect 198186 169200 198242 170000
rect 198554 169200 198610 170000
rect 198922 169200 198978 170000
rect 199290 169200 199346 170000
rect 199658 169200 199714 170000
rect 200026 169200 200082 170000
rect 200394 169200 200450 170000
rect 200762 169200 200818 170000
rect 201130 169200 201186 170000
rect 201498 169200 201554 170000
rect 201866 169200 201922 170000
rect 202234 169200 202290 170000
rect 202602 169200 202658 170000
rect 202970 169200 203026 170000
rect 203338 169200 203394 170000
rect 203706 169200 203762 170000
rect 204074 169200 204130 170000
rect 204442 169200 204498 170000
rect 204810 169200 204866 170000
rect 205178 169200 205234 170000
rect 205546 169200 205602 170000
rect 205914 169200 205970 170000
rect 206282 169200 206338 170000
rect 206650 169200 206706 170000
rect 207018 169200 207074 170000
rect 207386 169200 207442 170000
rect 207754 169200 207810 170000
rect 208122 169200 208178 170000
rect 208490 169200 208546 170000
rect 208858 169200 208914 170000
rect 209226 169200 209282 170000
rect 209594 169200 209650 170000
rect 209962 169200 210018 170000
rect 210330 169200 210386 170000
rect 210698 169200 210754 170000
rect 211066 169200 211122 170000
rect 211434 169200 211490 170000
rect 211802 169200 211858 170000
rect 212170 169200 212226 170000
rect 212538 169200 212594 170000
rect 212906 169200 212962 170000
rect 213274 169200 213330 170000
rect 213642 169200 213698 170000
rect 214010 169200 214066 170000
rect 214378 169200 214434 170000
rect 214746 169200 214802 170000
rect 215114 169200 215170 170000
rect 215482 169200 215538 170000
rect 215850 169200 215906 170000
rect 216218 169200 216274 170000
rect 216586 169200 216642 170000
rect 216954 169200 217010 170000
rect 217322 169200 217378 170000
rect 217690 169200 217746 170000
rect 218058 169200 218114 170000
rect 218426 169200 218482 170000
rect 218794 169200 218850 170000
rect 219162 169200 219218 170000
rect 219530 169200 219586 170000
rect 219898 169200 219954 170000
rect 220266 169200 220322 170000
rect 220634 169200 220690 170000
rect 221002 169200 221058 170000
rect 221370 169200 221426 170000
rect 221738 169200 221794 170000
rect 222106 169200 222162 170000
rect 222474 169200 222530 170000
rect 222842 169200 222898 170000
rect 223210 169200 223266 170000
rect 223578 169200 223634 170000
rect 223946 169200 224002 170000
rect 224314 169200 224370 170000
rect 224682 169200 224738 170000
rect 225050 169200 225106 170000
rect 225418 169200 225474 170000
rect 225786 169200 225842 170000
rect 226154 169200 226210 170000
rect 226522 169200 226578 170000
rect 226890 169200 226946 170000
rect 227258 169200 227314 170000
rect 227626 169200 227682 170000
rect 227994 169200 228050 170000
rect 228362 169200 228418 170000
rect 228730 169200 228786 170000
rect 229098 169200 229154 170000
rect 229466 169200 229522 170000
rect 229834 169200 229890 170000
rect 230202 169200 230258 170000
rect 230570 169200 230626 170000
rect 230938 169200 230994 170000
rect 231306 169200 231362 170000
rect 231674 169200 231730 170000
rect 232042 169200 232098 170000
rect 232410 169200 232466 170000
rect 232778 169200 232834 170000
rect 233146 169200 233202 170000
rect 233514 169200 233570 170000
rect 233882 169200 233938 170000
rect 234250 169200 234306 170000
rect 234618 169200 234674 170000
rect 234986 169200 235042 170000
rect 235354 169200 235410 170000
rect 235722 169200 235778 170000
rect 236090 169200 236146 170000
rect 236458 169200 236514 170000
rect 236826 169200 236882 170000
rect 237194 169200 237250 170000
rect 237562 169200 237618 170000
rect 237930 169200 237986 170000
rect 238298 169200 238354 170000
rect 238666 169200 238722 170000
rect 239034 169200 239090 170000
rect 239402 169200 239458 170000
rect 239770 169200 239826 170000
rect 240138 169200 240194 170000
rect 240506 169200 240562 170000
rect 240874 169200 240930 170000
rect 241242 169200 241298 170000
rect 241610 169200 241666 170000
rect 241978 169200 242034 170000
rect 242346 169200 242402 170000
rect 242714 169200 242770 170000
rect 243082 169200 243138 170000
rect 243450 169200 243506 170000
rect 243818 169200 243874 170000
rect 244186 169200 244242 170000
rect 244554 169200 244610 170000
rect 244922 169200 244978 170000
rect 245290 169200 245346 170000
rect 245658 169200 245714 170000
rect 246026 169200 246082 170000
rect 246394 169200 246450 170000
rect 246762 169200 246818 170000
rect 247130 169200 247186 170000
rect 247498 169200 247554 170000
rect 247866 169200 247922 170000
rect 248234 169200 248290 170000
rect 248602 169200 248658 170000
rect 248970 169200 249026 170000
rect 249338 169200 249394 170000
rect 249706 169200 249762 170000
rect 250074 169200 250130 170000
rect 250442 169200 250498 170000
rect 250810 169200 250866 170000
rect 251178 169200 251234 170000
rect 251546 169200 251602 170000
rect 251914 169200 251970 170000
rect 252282 169200 252338 170000
rect 252650 169200 252706 170000
rect 253018 169200 253074 170000
rect 253386 169200 253442 170000
rect 253754 169200 253810 170000
rect 254122 169200 254178 170000
rect 254490 169200 254546 170000
rect 254858 169200 254914 170000
rect 255226 169200 255282 170000
rect 255594 169200 255650 170000
rect 255962 169200 256018 170000
rect 256330 169200 256386 170000
rect 256698 169200 256754 170000
rect 257066 169200 257122 170000
rect 257434 169200 257490 170000
rect 257802 169200 257858 170000
rect 258170 169200 258226 170000
rect 258538 169200 258594 170000
rect 258906 169200 258962 170000
rect 259274 169200 259330 170000
rect 259642 169200 259698 170000
rect 260010 169200 260066 170000
rect 260378 169200 260434 170000
rect 260746 169200 260802 170000
rect 261114 169200 261170 170000
rect 261482 169200 261538 170000
rect 261850 169200 261906 170000
rect 262218 169200 262274 170000
rect 262586 169200 262642 170000
rect 262954 169200 263010 170000
rect 263322 169200 263378 170000
rect 263690 169200 263746 170000
rect 264058 169200 264114 170000
rect 264426 169200 264482 170000
rect 264794 169200 264850 170000
rect 265162 169200 265218 170000
rect 265530 169200 265586 170000
rect 265898 169200 265954 170000
rect 266266 169200 266322 170000
rect 266634 169200 266690 170000
rect 267002 169200 267058 170000
rect 267370 169200 267426 170000
rect 267738 169200 267794 170000
rect 268106 169200 268162 170000
rect 268474 169200 268530 170000
rect 268842 169200 268898 170000
rect 269210 169200 269266 170000
rect 269578 169200 269634 170000
rect 269946 169200 270002 170000
rect 270314 169200 270370 170000
rect 270682 169200 270738 170000
rect 271050 169200 271106 170000
rect 271418 169200 271474 170000
rect 271786 169200 271842 170000
rect 272154 169200 272210 170000
rect 272522 169200 272578 170000
rect 272890 169200 272946 170000
rect 273258 169200 273314 170000
rect 273626 169200 273682 170000
rect 273994 169200 274050 170000
rect 274362 169200 274418 170000
rect 274730 169200 274786 170000
rect 275098 169200 275154 170000
rect 275466 169200 275522 170000
rect 275834 169200 275890 170000
rect 276202 169200 276258 170000
rect 276570 169200 276626 170000
rect 276938 169200 276994 170000
rect 277306 169200 277362 170000
rect 277674 169200 277730 170000
rect 278042 169200 278098 170000
rect 278410 169200 278466 170000
rect 278778 169200 278834 170000
rect 279146 169200 279202 170000
rect 279514 169200 279570 170000
rect 279882 169200 279938 170000
rect 280250 169200 280306 170000
rect 280618 169200 280674 170000
rect 280986 169200 281042 170000
rect 281354 169200 281410 170000
rect 281722 169200 281778 170000
rect 282090 169200 282146 170000
rect 282458 169200 282514 170000
rect 282826 169200 282882 170000
rect 283194 169200 283250 170000
rect 283562 169200 283618 170000
rect 283930 169200 283986 170000
rect 284298 169200 284354 170000
rect 284666 169200 284722 170000
rect 285034 169200 285090 170000
rect 285402 169200 285458 170000
rect 285770 169200 285826 170000
rect 286138 169200 286194 170000
rect 286506 169200 286562 170000
rect 286874 169200 286930 170000
rect 287242 169200 287298 170000
rect 287610 169200 287666 170000
rect 287978 169200 288034 170000
rect 288346 169200 288402 170000
rect 288714 169200 288770 170000
rect 289082 169200 289138 170000
rect 289450 169200 289506 170000
rect 289818 169200 289874 170000
rect 290186 169200 290242 170000
rect 290554 169200 290610 170000
rect 290922 169200 290978 170000
rect 291290 169200 291346 170000
rect 291658 169200 291714 170000
rect 292026 169200 292082 170000
rect 292394 169200 292450 170000
rect 292762 169200 292818 170000
rect 293130 169200 293186 170000
rect 293498 169200 293554 170000
rect 293866 169200 293922 170000
rect 294234 169200 294290 170000
rect 294602 169200 294658 170000
rect 294970 169200 295026 170000
rect 295338 169200 295394 170000
rect 295706 169200 295762 170000
rect 296074 169200 296130 170000
rect 296442 169200 296498 170000
rect 296810 169200 296866 170000
rect 297178 169200 297234 170000
rect 297546 169200 297602 170000
rect 297914 169200 297970 170000
rect 298282 169200 298338 170000
rect 298650 169200 298706 170000
rect 299018 169200 299074 170000
rect 299386 169200 299442 170000
rect 299754 169200 299810 170000
rect 300122 169200 300178 170000
rect 300490 169200 300546 170000
rect 300858 169200 300914 170000
rect 301226 169200 301282 170000
rect 301594 169200 301650 170000
rect 301962 169200 302018 170000
rect 302330 169200 302386 170000
rect 302698 169200 302754 170000
rect 303066 169200 303122 170000
rect 303434 169200 303490 170000
rect 303802 169200 303858 170000
rect 304170 169200 304226 170000
rect 304538 169200 304594 170000
rect 304906 169200 304962 170000
rect 305274 169200 305330 170000
rect 305642 169200 305698 170000
rect 306010 169200 306066 170000
rect 306378 169200 306434 170000
rect 306746 169200 306802 170000
rect 307114 169200 307170 170000
rect 307482 169200 307538 170000
rect 307850 169200 307906 170000
rect 308218 169200 308274 170000
rect 308586 169200 308642 170000
rect 308954 169200 309010 170000
rect 309322 169200 309378 170000
rect 309690 169200 309746 170000
rect 310058 169200 310114 170000
rect 310426 169200 310482 170000
rect 335082 169200 335138 170000
rect 426714 169200 426770 170000
rect 427082 169200 427138 170000
rect 427450 169200 427506 170000
rect 427818 169200 427874 170000
rect 428186 169200 428242 170000
rect 428554 169200 428610 170000
rect 428922 169200 428978 170000
rect 429290 169200 429346 170000
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 422298 0 422354 800
rect 422666 0 422722 800
rect 423034 0 423090 800
rect 423402 0 423458 800
rect 423770 0 423826 800
rect 424138 0 424194 800
rect 424506 0 424562 800
rect 424874 0 424930 800
rect 425242 0 425298 800
rect 425610 0 425666 800
rect 425978 0 426034 800
rect 426346 0 426402 800
rect 426714 0 426770 800
rect 427082 0 427138 800
rect 427450 0 427506 800
rect 427818 0 427874 800
rect 428186 0 428242 800
rect 428554 0 428610 800
rect 428922 0 428978 800
rect 429290 0 429346 800
<< obsm2 >>
rect 682 169144 882 169998
rect 1050 169144 1250 169998
rect 1418 169144 1618 169998
rect 1786 169144 1986 169998
rect 2154 169144 2354 169998
rect 2522 169144 2722 169998
rect 2890 169144 3090 169998
rect 3258 169144 3458 169998
rect 3626 169144 3826 169998
rect 3994 169144 4194 169998
rect 4362 169144 4562 169998
rect 4730 169144 4930 169998
rect 5098 169144 5298 169998
rect 5466 169144 5666 169998
rect 5834 169144 6034 169998
rect 6202 169144 6402 169998
rect 6570 169144 6770 169998
rect 6938 169144 7138 169998
rect 7306 169144 7506 169998
rect 7674 169144 7874 169998
rect 8042 169144 8242 169998
rect 8410 169144 8610 169998
rect 8778 169144 8978 169998
rect 9146 169144 9346 169998
rect 9514 169144 9714 169998
rect 9882 169144 10082 169998
rect 10250 169144 10450 169998
rect 10618 169144 10818 169998
rect 10986 169144 11186 169998
rect 11354 169144 37314 169998
rect 37482 169144 88834 169998
rect 89002 169144 114226 169998
rect 114394 169144 139250 169998
rect 139418 169144 140354 169998
rect 140522 169144 140722 169998
rect 140890 169144 141090 169998
rect 141258 169144 141458 169998
rect 141626 169144 141826 169998
rect 141994 169144 142194 169998
rect 142362 169144 142562 169998
rect 142730 169144 142930 169998
rect 143098 169144 143298 169998
rect 143466 169144 143666 169998
rect 143834 169144 144034 169998
rect 144202 169144 144402 169998
rect 144570 169144 144770 169998
rect 144938 169144 145138 169998
rect 145306 169144 145506 169998
rect 145674 169144 145874 169998
rect 146042 169144 146242 169998
rect 146410 169144 146610 169998
rect 146778 169144 146978 169998
rect 147146 169144 147346 169998
rect 147514 169144 147714 169998
rect 147882 169144 148082 169998
rect 148250 169144 148450 169998
rect 148618 169144 148818 169998
rect 148986 169144 149186 169998
rect 149354 169144 149554 169998
rect 149722 169144 149922 169998
rect 150090 169144 150290 169998
rect 150458 169144 150658 169998
rect 150826 169144 151026 169998
rect 151194 169144 151394 169998
rect 151562 169144 151762 169998
rect 151930 169144 152130 169998
rect 152298 169144 152498 169998
rect 152666 169144 152866 169998
rect 153034 169144 153234 169998
rect 153402 169144 153602 169998
rect 153770 169144 153970 169998
rect 154138 169144 154338 169998
rect 154506 169144 154706 169998
rect 154874 169144 155074 169998
rect 155242 169144 155442 169998
rect 155610 169144 155810 169998
rect 155978 169144 156178 169998
rect 156346 169144 156546 169998
rect 156714 169144 156914 169998
rect 157082 169144 157282 169998
rect 157450 169144 157650 169998
rect 157818 169144 158018 169998
rect 158186 169144 158386 169998
rect 158554 169144 158754 169998
rect 158922 169144 159122 169998
rect 159290 169144 159490 169998
rect 159658 169144 159858 169998
rect 160026 169144 160226 169998
rect 160394 169144 160594 169998
rect 160762 169144 160962 169998
rect 161130 169144 161330 169998
rect 161498 169144 161698 169998
rect 161866 169144 162066 169998
rect 162234 169144 162434 169998
rect 162602 169144 162802 169998
rect 162970 169144 163170 169998
rect 163338 169144 163538 169998
rect 163706 169144 163906 169998
rect 164074 169144 164274 169998
rect 164442 169144 164642 169998
rect 164810 169144 165010 169998
rect 165178 169144 165378 169998
rect 165546 169144 165746 169998
rect 165914 169144 166114 169998
rect 166282 169144 166482 169998
rect 166650 169144 166850 169998
rect 167018 169144 167218 169998
rect 167386 169144 167586 169998
rect 167754 169144 167954 169998
rect 168122 169144 168322 169998
rect 168490 169144 168690 169998
rect 168858 169144 169058 169998
rect 169226 169144 169426 169998
rect 169594 169144 169794 169998
rect 169962 169144 170162 169998
rect 170330 169144 170530 169998
rect 170698 169144 170898 169998
rect 171066 169144 171266 169998
rect 171434 169144 171634 169998
rect 171802 169144 172002 169998
rect 172170 169144 172370 169998
rect 172538 169144 172738 169998
rect 172906 169144 173106 169998
rect 173274 169144 173474 169998
rect 173642 169144 173842 169998
rect 174010 169144 174210 169998
rect 174378 169144 174578 169998
rect 174746 169144 174946 169998
rect 175114 169144 175314 169998
rect 175482 169144 175682 169998
rect 175850 169144 176050 169998
rect 176218 169144 176418 169998
rect 176586 169144 176786 169998
rect 176954 169144 177154 169998
rect 177322 169144 177522 169998
rect 177690 169144 177890 169998
rect 178058 169144 178258 169998
rect 178426 169144 178626 169998
rect 178794 169144 178994 169998
rect 179162 169144 179362 169998
rect 179530 169144 179730 169998
rect 179898 169144 180098 169998
rect 180266 169144 180466 169998
rect 180634 169144 180834 169998
rect 181002 169144 181202 169998
rect 181370 169144 181570 169998
rect 181738 169144 181938 169998
rect 182106 169144 182306 169998
rect 182474 169144 182674 169998
rect 182842 169144 183042 169998
rect 183210 169144 183410 169998
rect 183578 169144 183778 169998
rect 183946 169144 184146 169998
rect 184314 169144 184514 169998
rect 184682 169144 184882 169998
rect 185050 169144 185250 169998
rect 185418 169144 185618 169998
rect 185786 169144 185986 169998
rect 186154 169144 186354 169998
rect 186522 169144 186722 169998
rect 186890 169144 187090 169998
rect 187258 169144 187458 169998
rect 187626 169144 187826 169998
rect 187994 169144 188194 169998
rect 188362 169144 188562 169998
rect 188730 169144 188930 169998
rect 189098 169144 189298 169998
rect 189466 169144 189666 169998
rect 189834 169144 190034 169998
rect 190202 169144 190402 169998
rect 190570 169144 190770 169998
rect 190938 169144 191138 169998
rect 191306 169144 191506 169998
rect 191674 169144 191874 169998
rect 192042 169144 192242 169998
rect 192410 169144 192610 169998
rect 192778 169144 192978 169998
rect 193146 169144 193346 169998
rect 193514 169144 193714 169998
rect 193882 169144 194082 169998
rect 194250 169144 194450 169998
rect 194618 169144 194818 169998
rect 194986 169144 195186 169998
rect 195354 169144 195554 169998
rect 195722 169144 195922 169998
rect 196090 169144 196290 169998
rect 196458 169144 196658 169998
rect 196826 169144 197026 169998
rect 197194 169144 197394 169998
rect 197562 169144 197762 169998
rect 197930 169144 198130 169998
rect 198298 169144 198498 169998
rect 198666 169144 198866 169998
rect 199034 169144 199234 169998
rect 199402 169144 199602 169998
rect 199770 169144 199970 169998
rect 200138 169144 200338 169998
rect 200506 169144 200706 169998
rect 200874 169144 201074 169998
rect 201242 169144 201442 169998
rect 201610 169144 201810 169998
rect 201978 169144 202178 169998
rect 202346 169144 202546 169998
rect 202714 169144 202914 169998
rect 203082 169144 203282 169998
rect 203450 169144 203650 169998
rect 203818 169144 204018 169998
rect 204186 169144 204386 169998
rect 204554 169144 204754 169998
rect 204922 169144 205122 169998
rect 205290 169144 205490 169998
rect 205658 169144 205858 169998
rect 206026 169144 206226 169998
rect 206394 169144 206594 169998
rect 206762 169144 206962 169998
rect 207130 169144 207330 169998
rect 207498 169144 207698 169998
rect 207866 169144 208066 169998
rect 208234 169144 208434 169998
rect 208602 169144 208802 169998
rect 208970 169144 209170 169998
rect 209338 169144 209538 169998
rect 209706 169144 209906 169998
rect 210074 169144 210274 169998
rect 210442 169144 210642 169998
rect 210810 169144 211010 169998
rect 211178 169144 211378 169998
rect 211546 169144 211746 169998
rect 211914 169144 212114 169998
rect 212282 169144 212482 169998
rect 212650 169144 212850 169998
rect 213018 169144 213218 169998
rect 213386 169144 213586 169998
rect 213754 169144 213954 169998
rect 214122 169144 214322 169998
rect 214490 169144 214690 169998
rect 214858 169144 215058 169998
rect 215226 169144 215426 169998
rect 215594 169144 215794 169998
rect 215962 169144 216162 169998
rect 216330 169144 216530 169998
rect 216698 169144 216898 169998
rect 217066 169144 217266 169998
rect 217434 169144 217634 169998
rect 217802 169144 218002 169998
rect 218170 169144 218370 169998
rect 218538 169144 218738 169998
rect 218906 169144 219106 169998
rect 219274 169144 219474 169998
rect 219642 169144 219842 169998
rect 220010 169144 220210 169998
rect 220378 169144 220578 169998
rect 220746 169144 220946 169998
rect 221114 169144 221314 169998
rect 221482 169144 221682 169998
rect 221850 169144 222050 169998
rect 222218 169144 222418 169998
rect 222586 169144 222786 169998
rect 222954 169144 223154 169998
rect 223322 169144 223522 169998
rect 223690 169144 223890 169998
rect 224058 169144 224258 169998
rect 224426 169144 224626 169998
rect 224794 169144 224994 169998
rect 225162 169144 225362 169998
rect 225530 169144 225730 169998
rect 225898 169144 226098 169998
rect 226266 169144 226466 169998
rect 226634 169144 226834 169998
rect 227002 169144 227202 169998
rect 227370 169144 227570 169998
rect 227738 169144 227938 169998
rect 228106 169144 228306 169998
rect 228474 169144 228674 169998
rect 228842 169144 229042 169998
rect 229210 169144 229410 169998
rect 229578 169144 229778 169998
rect 229946 169144 230146 169998
rect 230314 169144 230514 169998
rect 230682 169144 230882 169998
rect 231050 169144 231250 169998
rect 231418 169144 231618 169998
rect 231786 169144 231986 169998
rect 232154 169144 232354 169998
rect 232522 169144 232722 169998
rect 232890 169144 233090 169998
rect 233258 169144 233458 169998
rect 233626 169144 233826 169998
rect 233994 169144 234194 169998
rect 234362 169144 234562 169998
rect 234730 169144 234930 169998
rect 235098 169144 235298 169998
rect 235466 169144 235666 169998
rect 235834 169144 236034 169998
rect 236202 169144 236402 169998
rect 236570 169144 236770 169998
rect 236938 169144 237138 169998
rect 237306 169144 237506 169998
rect 237674 169144 237874 169998
rect 238042 169144 238242 169998
rect 238410 169144 238610 169998
rect 238778 169144 238978 169998
rect 239146 169144 239346 169998
rect 239514 169144 239714 169998
rect 239882 169144 240082 169998
rect 240250 169144 240450 169998
rect 240618 169144 240818 169998
rect 240986 169144 241186 169998
rect 241354 169144 241554 169998
rect 241722 169144 241922 169998
rect 242090 169144 242290 169998
rect 242458 169144 242658 169998
rect 242826 169144 243026 169998
rect 243194 169144 243394 169998
rect 243562 169144 243762 169998
rect 243930 169144 244130 169998
rect 244298 169144 244498 169998
rect 244666 169144 244866 169998
rect 245034 169144 245234 169998
rect 245402 169144 245602 169998
rect 245770 169144 245970 169998
rect 246138 169144 246338 169998
rect 246506 169144 246706 169998
rect 246874 169144 247074 169998
rect 247242 169144 247442 169998
rect 247610 169144 247810 169998
rect 247978 169144 248178 169998
rect 248346 169144 248546 169998
rect 248714 169144 248914 169998
rect 249082 169144 249282 169998
rect 249450 169144 249650 169998
rect 249818 169144 250018 169998
rect 250186 169144 250386 169998
rect 250554 169144 250754 169998
rect 250922 169144 251122 169998
rect 251290 169144 251490 169998
rect 251658 169144 251858 169998
rect 252026 169144 252226 169998
rect 252394 169144 252594 169998
rect 252762 169144 252962 169998
rect 253130 169144 253330 169998
rect 253498 169144 253698 169998
rect 253866 169144 254066 169998
rect 254234 169144 254434 169998
rect 254602 169144 254802 169998
rect 254970 169144 255170 169998
rect 255338 169144 255538 169998
rect 255706 169144 255906 169998
rect 256074 169144 256274 169998
rect 256442 169144 256642 169998
rect 256810 169144 257010 169998
rect 257178 169144 257378 169998
rect 257546 169144 257746 169998
rect 257914 169144 258114 169998
rect 258282 169144 258482 169998
rect 258650 169144 258850 169998
rect 259018 169144 259218 169998
rect 259386 169144 259586 169998
rect 259754 169144 259954 169998
rect 260122 169144 260322 169998
rect 260490 169144 260690 169998
rect 260858 169144 261058 169998
rect 261226 169144 261426 169998
rect 261594 169144 261794 169998
rect 261962 169144 262162 169998
rect 262330 169144 262530 169998
rect 262698 169144 262898 169998
rect 263066 169144 263266 169998
rect 263434 169144 263634 169998
rect 263802 169144 264002 169998
rect 264170 169144 264370 169998
rect 264538 169144 264738 169998
rect 264906 169144 265106 169998
rect 265274 169144 265474 169998
rect 265642 169144 265842 169998
rect 266010 169144 266210 169998
rect 266378 169144 266578 169998
rect 266746 169144 266946 169998
rect 267114 169144 267314 169998
rect 267482 169144 267682 169998
rect 267850 169144 268050 169998
rect 268218 169144 268418 169998
rect 268586 169144 268786 169998
rect 268954 169144 269154 169998
rect 269322 169144 269522 169998
rect 269690 169144 269890 169998
rect 270058 169144 270258 169998
rect 270426 169144 270626 169998
rect 270794 169144 270994 169998
rect 271162 169144 271362 169998
rect 271530 169144 271730 169998
rect 271898 169144 272098 169998
rect 272266 169144 272466 169998
rect 272634 169144 272834 169998
rect 273002 169144 273202 169998
rect 273370 169144 273570 169998
rect 273738 169144 273938 169998
rect 274106 169144 274306 169998
rect 274474 169144 274674 169998
rect 274842 169144 275042 169998
rect 275210 169144 275410 169998
rect 275578 169144 275778 169998
rect 275946 169144 276146 169998
rect 276314 169144 276514 169998
rect 276682 169144 276882 169998
rect 277050 169144 277250 169998
rect 277418 169144 277618 169998
rect 277786 169144 277986 169998
rect 278154 169144 278354 169998
rect 278522 169144 278722 169998
rect 278890 169144 279090 169998
rect 279258 169144 279458 169998
rect 279626 169144 279826 169998
rect 279994 169144 280194 169998
rect 280362 169144 280562 169998
rect 280730 169144 280930 169998
rect 281098 169144 281298 169998
rect 281466 169144 281666 169998
rect 281834 169144 282034 169998
rect 282202 169144 282402 169998
rect 282570 169144 282770 169998
rect 282938 169144 283138 169998
rect 283306 169144 283506 169998
rect 283674 169144 283874 169998
rect 284042 169144 284242 169998
rect 284410 169144 284610 169998
rect 284778 169144 284978 169998
rect 285146 169144 285346 169998
rect 285514 169144 285714 169998
rect 285882 169144 286082 169998
rect 286250 169144 286450 169998
rect 286618 169144 286818 169998
rect 286986 169144 287186 169998
rect 287354 169144 287554 169998
rect 287722 169144 287922 169998
rect 288090 169144 288290 169998
rect 288458 169144 288658 169998
rect 288826 169144 289026 169998
rect 289194 169144 289394 169998
rect 289562 169144 289762 169998
rect 289930 169144 290130 169998
rect 290298 169144 290498 169998
rect 290666 169144 290866 169998
rect 291034 169144 291234 169998
rect 291402 169144 291602 169998
rect 291770 169144 291970 169998
rect 292138 169144 292338 169998
rect 292506 169144 292706 169998
rect 292874 169144 293074 169998
rect 293242 169144 293442 169998
rect 293610 169144 293810 169998
rect 293978 169144 294178 169998
rect 294346 169144 294546 169998
rect 294714 169144 294914 169998
rect 295082 169144 295282 169998
rect 295450 169144 295650 169998
rect 295818 169144 296018 169998
rect 296186 169144 296386 169998
rect 296554 169144 296754 169998
rect 296922 169144 297122 169998
rect 297290 169144 297490 169998
rect 297658 169144 297858 169998
rect 298026 169144 298226 169998
rect 298394 169144 298594 169998
rect 298762 169144 298962 169998
rect 299130 169144 299330 169998
rect 299498 169144 299698 169998
rect 299866 169144 300066 169998
rect 300234 169144 300434 169998
rect 300602 169144 300802 169998
rect 300970 169144 301170 169998
rect 301338 169144 301538 169998
rect 301706 169144 301906 169998
rect 302074 169144 302274 169998
rect 302442 169144 302642 169998
rect 302810 169144 303010 169998
rect 303178 169144 303378 169998
rect 303546 169144 303746 169998
rect 303914 169144 304114 169998
rect 304282 169144 304482 169998
rect 304650 169144 304850 169998
rect 305018 169144 305218 169998
rect 305386 169144 305586 169998
rect 305754 169144 305954 169998
rect 306122 169144 306322 169998
rect 306490 169144 306690 169998
rect 306858 169144 307058 169998
rect 307226 169144 307426 169998
rect 307594 169144 307794 169998
rect 307962 169144 308162 169998
rect 308330 169144 308530 169998
rect 308698 169144 308898 169998
rect 309066 169144 309266 169998
rect 309434 169144 309634 169998
rect 309802 169144 310002 169998
rect 310170 169144 310370 169998
rect 310538 169144 335026 169998
rect 335194 169144 426658 169998
rect 426826 169144 427026 169998
rect 427194 169144 427394 169998
rect 427562 169144 427762 169998
rect 427930 169144 428130 169998
rect 428298 169144 428498 169998
rect 428666 169144 428866 169998
rect 429034 169144 429234 169998
rect 570 856 429344 169144
rect 682 614 698 856
rect 866 614 882 856
rect 1050 614 1066 856
rect 1234 614 1250 856
rect 1418 614 1434 856
rect 1602 614 1618 856
rect 1786 614 1802 856
rect 1970 614 1986 856
rect 2154 614 2170 856
rect 2338 614 2354 856
rect 2522 614 2538 856
rect 2706 614 2722 856
rect 2890 614 2906 856
rect 3074 614 3090 856
rect 3258 614 3274 856
rect 3442 614 3458 856
rect 3626 614 3642 856
rect 3810 614 3826 856
rect 3994 614 4010 856
rect 4178 614 4194 856
rect 4362 614 4378 856
rect 4546 614 4562 856
rect 4730 614 4746 856
rect 4914 614 4930 856
rect 5098 614 5114 856
rect 5282 614 5298 856
rect 5466 614 5482 856
rect 5650 614 5666 856
rect 5834 614 5850 856
rect 6018 614 6034 856
rect 6202 614 6218 856
rect 6386 614 6402 856
rect 6570 614 6586 856
rect 6754 614 6770 856
rect 6938 614 6954 856
rect 7122 614 7138 856
rect 7306 614 7322 856
rect 7490 614 7506 856
rect 7674 614 7690 856
rect 7858 614 7874 856
rect 8042 614 8058 856
rect 8226 614 8242 856
rect 8410 614 8426 856
rect 8594 614 8610 856
rect 8778 614 8794 856
rect 8962 614 8978 856
rect 9146 614 9162 856
rect 9330 614 9346 856
rect 9514 614 9530 856
rect 9698 614 9714 856
rect 9882 614 9898 856
rect 10066 614 10082 856
rect 10250 614 10266 856
rect 10434 614 10450 856
rect 10618 614 10634 856
rect 10802 614 10818 856
rect 10986 614 11002 856
rect 11170 614 11186 856
rect 11354 614 11370 856
rect 11538 614 11554 856
rect 11722 614 11738 856
rect 11906 614 11922 856
rect 12090 614 12106 856
rect 12274 614 12290 856
rect 12458 614 12474 856
rect 12642 614 12658 856
rect 12826 614 12842 856
rect 13010 614 13026 856
rect 13194 614 13210 856
rect 13378 614 13394 856
rect 13562 614 13578 856
rect 13746 614 13762 856
rect 13930 614 13946 856
rect 14114 614 14130 856
rect 14298 614 14314 856
rect 14482 614 14498 856
rect 14666 614 14682 856
rect 14850 614 14866 856
rect 15034 614 15050 856
rect 15218 614 15234 856
rect 15402 614 15418 856
rect 15586 614 15602 856
rect 15770 614 15786 856
rect 15954 614 15970 856
rect 16138 614 16338 856
rect 16506 614 16706 856
rect 16874 614 17074 856
rect 17242 614 17442 856
rect 17610 614 17810 856
rect 17978 614 18178 856
rect 18346 614 18546 856
rect 18714 614 18914 856
rect 19082 614 19282 856
rect 19450 614 19650 856
rect 19818 614 20018 856
rect 20186 614 20386 856
rect 20554 614 20754 856
rect 20922 614 21122 856
rect 21290 614 21490 856
rect 21658 614 21858 856
rect 22026 614 22226 856
rect 22394 614 22594 856
rect 22762 614 22962 856
rect 23130 614 23330 856
rect 23498 614 23698 856
rect 23866 614 24066 856
rect 24234 614 24434 856
rect 24602 614 24802 856
rect 24970 614 25170 856
rect 25338 614 25538 856
rect 25706 614 25906 856
rect 26074 614 26274 856
rect 26442 614 26642 856
rect 26810 614 27010 856
rect 27178 614 27378 856
rect 27546 614 27746 856
rect 27914 614 28114 856
rect 28282 614 28482 856
rect 28650 614 28850 856
rect 29018 614 29218 856
rect 29386 614 29586 856
rect 29754 614 29954 856
rect 30122 614 30322 856
rect 30490 614 30690 856
rect 30858 614 31058 856
rect 31226 614 31426 856
rect 31594 614 31794 856
rect 31962 614 32162 856
rect 32330 614 32530 856
rect 32698 614 32898 856
rect 33066 614 33266 856
rect 33434 614 33634 856
rect 33802 614 34002 856
rect 34170 614 34370 856
rect 34538 614 34738 856
rect 34906 614 35106 856
rect 35274 614 35474 856
rect 35642 614 35842 856
rect 36010 614 36210 856
rect 36378 614 36578 856
rect 36746 614 36946 856
rect 37114 614 37314 856
rect 37482 614 37682 856
rect 37850 614 38050 856
rect 38218 614 38418 856
rect 38586 614 38786 856
rect 38954 614 39154 856
rect 39322 614 39522 856
rect 39690 614 422242 856
rect 422410 614 422610 856
rect 422778 614 422978 856
rect 423146 614 423346 856
rect 423514 614 423714 856
rect 423882 614 424082 856
rect 424250 614 424450 856
rect 424618 614 424818 856
rect 424986 614 425186 856
rect 425354 614 425554 856
rect 425722 614 425922 856
rect 426090 614 426290 856
rect 426458 614 426658 856
rect 426826 614 427026 856
rect 427194 614 427394 856
rect 427562 614 427762 856
rect 427930 614 428130 856
rect 428298 614 428498 856
rect 428666 614 428866 856
rect 429034 614 429234 856
<< metal3 >>
rect 0 168648 800 168768
rect 429200 168648 430000 168768
rect 0 168104 800 168224
rect 429200 168104 430000 168224
rect 0 167560 800 167680
rect 429200 167560 430000 167680
rect 0 167016 800 167136
rect 429200 167016 430000 167136
rect 0 166472 800 166592
rect 0 165928 800 166048
rect 0 165384 800 165504
rect 0 164840 800 164960
rect 0 164296 800 164416
rect 0 163752 800 163872
rect 0 163208 800 163328
rect 0 162664 800 162784
rect 0 162120 800 162240
rect 0 161576 800 161696
rect 0 161032 800 161152
rect 0 160488 800 160608
rect 0 159944 800 160064
rect 0 159400 800 159520
rect 0 158856 800 158976
rect 429200 157224 430000 157344
rect 0 149064 800 149184
rect 429200 113160 430000 113280
rect 429200 112616 430000 112736
rect 429200 112072 430000 112192
rect 429200 96296 430000 96416
rect 429200 89768 430000 89888
rect 429200 68008 430000 68128
rect 429200 67464 430000 67584
rect 429200 66920 430000 67040
rect 429200 66376 430000 66496
rect 0 39720 800 39840
rect 0 39176 800 39296
rect 0 38632 800 38752
rect 0 38088 800 38208
rect 0 37544 800 37664
rect 0 37000 800 37120
rect 0 36456 800 36576
rect 0 35912 800 36032
rect 0 35368 800 35488
rect 0 34824 800 34944
rect 0 34280 800 34400
rect 0 33736 800 33856
rect 0 33192 800 33312
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 0 31560 800 31680
rect 0 31016 800 31136
rect 0 30472 800 30592
rect 0 29928 800 30048
rect 0 29384 800 29504
rect 0 28840 800 28960
rect 0 28296 800 28416
rect 0 27752 800 27872
rect 0 27208 800 27328
rect 0 26664 800 26784
rect 0 26120 800 26240
rect 0 25576 800 25696
rect 0 25032 800 25152
rect 0 24488 800 24608
rect 0 23944 800 24064
rect 0 23400 800 23520
rect 0 22856 800 22976
rect 0 22312 800 22432
rect 0 21768 800 21888
rect 429200 21768 430000 21888
rect 0 21224 800 21344
rect 0 20680 800 20800
rect 0 20136 800 20256
rect 0 19592 800 19712
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 0 13608 800 13728
rect 0 13064 800 13184
rect 0 12520 800 12640
rect 0 11976 800 12096
rect 0 11432 800 11552
rect 0 10888 800 11008
rect 0 10344 800 10464
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8712 800 8832
rect 0 8168 800 8288
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 429200 7080 430000 7200
rect 0 6536 800 6656
rect 429200 6536 430000 6656
rect 0 5992 800 6112
rect 429200 5992 430000 6112
rect 0 5448 800 5568
rect 429200 5448 430000 5568
rect 0 4904 800 5024
rect 429200 4904 430000 5024
rect 0 4360 800 4480
rect 429200 4360 430000 4480
rect 0 3816 800 3936
rect 429200 3816 430000 3936
rect 0 3272 800 3392
rect 429200 3272 430000 3392
rect 0 2728 800 2848
rect 429200 2728 430000 2848
rect 0 2184 800 2304
rect 429200 2184 430000 2304
rect 0 1640 800 1760
rect 429200 1640 430000 1760
rect 0 1096 800 1216
rect 429200 1096 430000 1216
<< obsm3 >>
rect 880 168568 429120 168741
rect 565 168304 429210 168568
rect 880 168024 429120 168304
rect 565 167760 429210 168024
rect 880 167480 429120 167760
rect 565 167216 429210 167480
rect 880 166936 429120 167216
rect 565 166672 429210 166936
rect 880 166392 429210 166672
rect 565 166128 429210 166392
rect 880 165848 429210 166128
rect 565 165584 429210 165848
rect 880 165304 429210 165584
rect 565 165040 429210 165304
rect 880 164760 429210 165040
rect 565 164496 429210 164760
rect 880 164216 429210 164496
rect 565 163952 429210 164216
rect 880 163672 429210 163952
rect 565 163408 429210 163672
rect 880 163128 429210 163408
rect 565 162864 429210 163128
rect 880 162584 429210 162864
rect 565 162320 429210 162584
rect 880 162040 429210 162320
rect 565 161776 429210 162040
rect 880 161496 429210 161776
rect 565 161232 429210 161496
rect 880 160952 429210 161232
rect 565 160688 429210 160952
rect 880 160408 429210 160688
rect 565 160144 429210 160408
rect 880 159864 429210 160144
rect 565 159600 429210 159864
rect 880 159320 429210 159600
rect 565 159056 429210 159320
rect 880 158776 429210 159056
rect 565 157424 429210 158776
rect 565 157144 429120 157424
rect 565 149264 429210 157144
rect 880 148984 429210 149264
rect 565 113360 429210 148984
rect 565 113080 429120 113360
rect 565 112816 429210 113080
rect 565 112536 429120 112816
rect 565 112272 429210 112536
rect 565 111992 429120 112272
rect 565 96496 429210 111992
rect 565 96216 429120 96496
rect 565 89968 429210 96216
rect 565 89688 429120 89968
rect 565 68208 429210 89688
rect 565 67928 429120 68208
rect 565 67664 429210 67928
rect 565 67384 429120 67664
rect 565 67120 429210 67384
rect 565 66840 429120 67120
rect 565 66576 429210 66840
rect 565 66296 429120 66576
rect 565 39920 429210 66296
rect 880 39640 429210 39920
rect 565 39376 429210 39640
rect 880 39096 429210 39376
rect 565 38832 429210 39096
rect 880 38552 429210 38832
rect 565 38288 429210 38552
rect 880 38008 429210 38288
rect 565 37744 429210 38008
rect 880 37464 429210 37744
rect 565 37200 429210 37464
rect 880 36920 429210 37200
rect 565 36656 429210 36920
rect 880 36376 429210 36656
rect 565 36112 429210 36376
rect 880 35832 429210 36112
rect 565 35568 429210 35832
rect 880 35288 429210 35568
rect 565 35024 429210 35288
rect 880 34744 429210 35024
rect 565 34480 429210 34744
rect 880 34200 429210 34480
rect 565 33936 429210 34200
rect 880 33656 429210 33936
rect 565 33392 429210 33656
rect 880 33112 429210 33392
rect 565 32848 429210 33112
rect 880 32568 429210 32848
rect 565 32304 429210 32568
rect 880 32024 429210 32304
rect 565 31760 429210 32024
rect 880 31480 429210 31760
rect 565 31216 429210 31480
rect 880 30936 429210 31216
rect 565 30672 429210 30936
rect 880 30392 429210 30672
rect 565 30128 429210 30392
rect 880 29848 429210 30128
rect 565 29584 429210 29848
rect 880 29304 429210 29584
rect 565 29040 429210 29304
rect 880 28760 429210 29040
rect 565 28496 429210 28760
rect 880 28216 429210 28496
rect 565 27952 429210 28216
rect 880 27672 429210 27952
rect 565 27408 429210 27672
rect 880 27128 429210 27408
rect 565 26864 429210 27128
rect 880 26584 429210 26864
rect 565 26320 429210 26584
rect 880 26040 429210 26320
rect 565 25776 429210 26040
rect 880 25496 429210 25776
rect 565 25232 429210 25496
rect 880 24952 429210 25232
rect 565 24688 429210 24952
rect 880 24408 429210 24688
rect 565 24144 429210 24408
rect 880 23864 429210 24144
rect 565 23600 429210 23864
rect 880 23320 429210 23600
rect 565 23056 429210 23320
rect 880 22776 429210 23056
rect 565 22512 429210 22776
rect 880 22232 429210 22512
rect 565 21968 429210 22232
rect 880 21688 429120 21968
rect 565 21424 429210 21688
rect 880 21144 429210 21424
rect 565 20880 429210 21144
rect 880 20600 429210 20880
rect 565 20336 429210 20600
rect 880 20056 429210 20336
rect 565 19792 429210 20056
rect 880 19512 429210 19792
rect 565 19248 429210 19512
rect 880 18968 429210 19248
rect 565 18704 429210 18968
rect 880 18424 429210 18704
rect 565 18160 429210 18424
rect 880 17880 429210 18160
rect 565 17616 429210 17880
rect 880 17336 429210 17616
rect 565 17072 429210 17336
rect 880 16792 429210 17072
rect 565 16528 429210 16792
rect 880 16248 429210 16528
rect 565 15984 429210 16248
rect 880 15704 429210 15984
rect 565 15440 429210 15704
rect 880 15160 429210 15440
rect 565 14896 429210 15160
rect 880 14616 429210 14896
rect 565 14352 429210 14616
rect 880 14072 429210 14352
rect 565 13808 429210 14072
rect 880 13528 429210 13808
rect 565 13264 429210 13528
rect 880 12984 429210 13264
rect 565 12720 429210 12984
rect 880 12440 429210 12720
rect 565 12176 429210 12440
rect 880 11896 429210 12176
rect 565 11632 429210 11896
rect 880 11352 429210 11632
rect 565 11088 429210 11352
rect 880 10808 429210 11088
rect 565 10544 429210 10808
rect 880 10264 429210 10544
rect 565 10000 429210 10264
rect 880 9720 429210 10000
rect 565 9456 429210 9720
rect 880 9176 429210 9456
rect 565 8912 429210 9176
rect 880 8632 429210 8912
rect 565 8368 429210 8632
rect 880 8088 429210 8368
rect 565 7824 429210 8088
rect 880 7544 429210 7824
rect 565 7280 429210 7544
rect 880 7000 429120 7280
rect 565 6736 429210 7000
rect 880 6456 429120 6736
rect 565 6192 429210 6456
rect 880 5912 429120 6192
rect 565 5648 429210 5912
rect 880 5368 429120 5648
rect 565 5104 429210 5368
rect 880 4824 429120 5104
rect 565 4560 429210 4824
rect 880 4280 429120 4560
rect 565 4016 429210 4280
rect 880 3736 429120 4016
rect 565 3472 429210 3736
rect 880 3192 429120 3472
rect 565 2928 429210 3192
rect 880 2648 429120 2928
rect 565 2384 429210 2648
rect 880 2104 429120 2384
rect 565 1840 429210 2104
rect 880 1560 429120 1840
rect 565 1296 429210 1560
rect 880 1123 429120 1296
<< obsm4 >>
rect 3923 1259 427458 168333
<< obsm5 >>
rect 1104 5298 428812 167100
<< labels >>
rlabel metal2 s 570 0 626 800 6 clock
port 1 nsew
rlabel metal2 s 114282 169200 114338 170000 6 core_clk
port 2 nsew
rlabel metal2 s 225418 169200 225474 170000 6 core_rstn
port 3 nsew
rlabel metal2 s 938 0 994 800 6 flash_clk
port 4 nsew
rlabel metal3 s 0 1096 800 1216 6 flash_clk_ieb
port 5 nsew
rlabel metal2 s 1306 0 1362 800 6 flash_clk_oeb
port 6 nsew
rlabel metal3 s 0 1640 800 1760 6 flash_csb
port 7 nsew
rlabel metal2 s 1674 0 1730 800 6 flash_csb_ieb
port 8 nsew
rlabel metal2 s 2042 0 2098 800 6 flash_csb_oeb
port 9 nsew
rlabel metal3 s 0 2184 800 2304 6 flash_io0_di
port 10 nsew
rlabel metal2 s 2410 0 2466 800 6 flash_io0_do
port 11 nsew
rlabel metal3 s 0 2728 800 2848 6 flash_io0_ieb
port 12 nsew
rlabel metal2 s 2778 0 2834 800 6 flash_io0_oeb
port 13 nsew
rlabel metal2 s 3146 0 3202 800 6 flash_io1_di
port 14 nsew
rlabel metal3 s 0 3272 800 3392 6 flash_io1_do
port 15 nsew
rlabel metal2 s 3514 0 3570 800 6 flash_io1_ieb
port 16 nsew
rlabel metal3 s 0 3816 800 3936 6 flash_io1_oeb
port 17 nsew
rlabel metal2 s 3882 0 3938 800 6 gpio_in_pad
port 18 nsew
rlabel metal2 s 4250 0 4306 800 6 gpio_inenb_pad
port 19 nsew
rlabel metal3 s 0 4360 800 4480 6 gpio_mode0_pad
port 20 nsew
rlabel metal2 s 4618 0 4674 800 6 gpio_mode1_pad
port 21 nsew
rlabel metal3 s 0 4904 800 5024 6 gpio_out_pad
port 22 nsew
rlabel metal2 s 4986 0 5042 800 6 gpio_outenb_pad
port 23 nsew
rlabel metal3 s 429200 67464 430000 67584 6 jtag_out
port 24 nsew
rlabel metal3 s 429200 66920 430000 67040 6 jtag_outenb
port 25 nsew
rlabel metal2 s 225050 169200 225106 170000 6 la_input[0]
port 26 nsew
rlabel metal2 s 225786 169200 225842 170000 6 la_input[100]
port 27 nsew
rlabel metal2 s 224682 169200 224738 170000 6 la_input[101]
port 28 nsew
rlabel metal2 s 226154 169200 226210 170000 6 la_input[102]
port 29 nsew
rlabel metal2 s 224314 169200 224370 170000 6 la_input[103]
port 30 nsew
rlabel metal2 s 226522 169200 226578 170000 6 la_input[104]
port 31 nsew
rlabel metal2 s 223946 169200 224002 170000 6 la_input[105]
port 32 nsew
rlabel metal2 s 226890 169200 226946 170000 6 la_input[106]
port 33 nsew
rlabel metal2 s 223578 169200 223634 170000 6 la_input[107]
port 34 nsew
rlabel metal2 s 227258 169200 227314 170000 6 la_input[108]
port 35 nsew
rlabel metal2 s 223210 169200 223266 170000 6 la_input[109]
port 36 nsew
rlabel metal2 s 227626 169200 227682 170000 6 la_input[10]
port 37 nsew
rlabel metal2 s 222842 169200 222898 170000 6 la_input[110]
port 38 nsew
rlabel metal2 s 227994 169200 228050 170000 6 la_input[111]
port 39 nsew
rlabel metal2 s 222474 169200 222530 170000 6 la_input[112]
port 40 nsew
rlabel metal2 s 228362 169200 228418 170000 6 la_input[113]
port 41 nsew
rlabel metal2 s 222106 169200 222162 170000 6 la_input[114]
port 42 nsew
rlabel metal2 s 228730 169200 228786 170000 6 la_input[115]
port 43 nsew
rlabel metal2 s 221738 169200 221794 170000 6 la_input[116]
port 44 nsew
rlabel metal2 s 229098 169200 229154 170000 6 la_input[117]
port 45 nsew
rlabel metal2 s 221370 169200 221426 170000 6 la_input[118]
port 46 nsew
rlabel metal2 s 229466 169200 229522 170000 6 la_input[119]
port 47 nsew
rlabel metal2 s 221002 169200 221058 170000 6 la_input[11]
port 48 nsew
rlabel metal2 s 229834 169200 229890 170000 6 la_input[120]
port 49 nsew
rlabel metal2 s 220634 169200 220690 170000 6 la_input[121]
port 50 nsew
rlabel metal2 s 230202 169200 230258 170000 6 la_input[122]
port 51 nsew
rlabel metal2 s 220266 169200 220322 170000 6 la_input[123]
port 52 nsew
rlabel metal2 s 230570 169200 230626 170000 6 la_input[124]
port 53 nsew
rlabel metal2 s 219898 169200 219954 170000 6 la_input[125]
port 54 nsew
rlabel metal2 s 230938 169200 230994 170000 6 la_input[126]
port 55 nsew
rlabel metal2 s 219530 169200 219586 170000 6 la_input[127]
port 56 nsew
rlabel metal2 s 231306 169200 231362 170000 6 la_input[12]
port 57 nsew
rlabel metal2 s 219162 169200 219218 170000 6 la_input[13]
port 58 nsew
rlabel metal2 s 231674 169200 231730 170000 6 la_input[14]
port 59 nsew
rlabel metal2 s 218794 169200 218850 170000 6 la_input[15]
port 60 nsew
rlabel metal2 s 232042 169200 232098 170000 6 la_input[16]
port 61 nsew
rlabel metal2 s 218426 169200 218482 170000 6 la_input[17]
port 62 nsew
rlabel metal2 s 232410 169200 232466 170000 6 la_input[18]
port 63 nsew
rlabel metal2 s 218058 169200 218114 170000 6 la_input[19]
port 64 nsew
rlabel metal2 s 232778 169200 232834 170000 6 la_input[1]
port 65 nsew
rlabel metal2 s 217690 169200 217746 170000 6 la_input[20]
port 66 nsew
rlabel metal2 s 233146 169200 233202 170000 6 la_input[21]
port 67 nsew
rlabel metal2 s 217322 169200 217378 170000 6 la_input[22]
port 68 nsew
rlabel metal2 s 233514 169200 233570 170000 6 la_input[23]
port 69 nsew
rlabel metal2 s 216954 169200 217010 170000 6 la_input[24]
port 70 nsew
rlabel metal2 s 233882 169200 233938 170000 6 la_input[25]
port 71 nsew
rlabel metal2 s 216586 169200 216642 170000 6 la_input[26]
port 72 nsew
rlabel metal2 s 234250 169200 234306 170000 6 la_input[27]
port 73 nsew
rlabel metal2 s 216218 169200 216274 170000 6 la_input[28]
port 74 nsew
rlabel metal2 s 234618 169200 234674 170000 6 la_input[29]
port 75 nsew
rlabel metal2 s 215850 169200 215906 170000 6 la_input[2]
port 76 nsew
rlabel metal2 s 234986 169200 235042 170000 6 la_input[30]
port 77 nsew
rlabel metal2 s 215482 169200 215538 170000 6 la_input[31]
port 78 nsew
rlabel metal2 s 235354 169200 235410 170000 6 la_input[32]
port 79 nsew
rlabel metal2 s 215114 169200 215170 170000 6 la_input[33]
port 80 nsew
rlabel metal2 s 235722 169200 235778 170000 6 la_input[34]
port 81 nsew
rlabel metal2 s 214746 169200 214802 170000 6 la_input[35]
port 82 nsew
rlabel metal2 s 236090 169200 236146 170000 6 la_input[36]
port 83 nsew
rlabel metal2 s 214378 169200 214434 170000 6 la_input[37]
port 84 nsew
rlabel metal2 s 236458 169200 236514 170000 6 la_input[38]
port 85 nsew
rlabel metal2 s 214010 169200 214066 170000 6 la_input[39]
port 86 nsew
rlabel metal2 s 236826 169200 236882 170000 6 la_input[3]
port 87 nsew
rlabel metal2 s 213642 169200 213698 170000 6 la_input[40]
port 88 nsew
rlabel metal2 s 237194 169200 237250 170000 6 la_input[41]
port 89 nsew
rlabel metal2 s 213274 169200 213330 170000 6 la_input[42]
port 90 nsew
rlabel metal2 s 237562 169200 237618 170000 6 la_input[43]
port 91 nsew
rlabel metal2 s 212906 169200 212962 170000 6 la_input[44]
port 92 nsew
rlabel metal2 s 237930 169200 237986 170000 6 la_input[45]
port 93 nsew
rlabel metal2 s 212538 169200 212594 170000 6 la_input[46]
port 94 nsew
rlabel metal2 s 238298 169200 238354 170000 6 la_input[47]
port 95 nsew
rlabel metal2 s 212170 169200 212226 170000 6 la_input[48]
port 96 nsew
rlabel metal2 s 238666 169200 238722 170000 6 la_input[49]
port 97 nsew
rlabel metal2 s 211802 169200 211858 170000 6 la_input[4]
port 98 nsew
rlabel metal2 s 239034 169200 239090 170000 6 la_input[50]
port 99 nsew
rlabel metal2 s 211434 169200 211490 170000 6 la_input[51]
port 100 nsew
rlabel metal2 s 239402 169200 239458 170000 6 la_input[52]
port 101 nsew
rlabel metal2 s 211066 169200 211122 170000 6 la_input[53]
port 102 nsew
rlabel metal2 s 239770 169200 239826 170000 6 la_input[54]
port 103 nsew
rlabel metal2 s 210698 169200 210754 170000 6 la_input[55]
port 104 nsew
rlabel metal2 s 240138 169200 240194 170000 6 la_input[56]
port 105 nsew
rlabel metal2 s 210330 169200 210386 170000 6 la_input[57]
port 106 nsew
rlabel metal2 s 240506 169200 240562 170000 6 la_input[58]
port 107 nsew
rlabel metal2 s 209962 169200 210018 170000 6 la_input[59]
port 108 nsew
rlabel metal2 s 240874 169200 240930 170000 6 la_input[5]
port 109 nsew
rlabel metal2 s 209594 169200 209650 170000 6 la_input[60]
port 110 nsew
rlabel metal2 s 241242 169200 241298 170000 6 la_input[61]
port 111 nsew
rlabel metal2 s 209226 169200 209282 170000 6 la_input[62]
port 112 nsew
rlabel metal2 s 241610 169200 241666 170000 6 la_input[63]
port 113 nsew
rlabel metal2 s 208858 169200 208914 170000 6 la_input[64]
port 114 nsew
rlabel metal2 s 241978 169200 242034 170000 6 la_input[65]
port 115 nsew
rlabel metal2 s 208490 169200 208546 170000 6 la_input[66]
port 116 nsew
rlabel metal2 s 242346 169200 242402 170000 6 la_input[67]
port 117 nsew
rlabel metal2 s 208122 169200 208178 170000 6 la_input[68]
port 118 nsew
rlabel metal2 s 242714 169200 242770 170000 6 la_input[69]
port 119 nsew
rlabel metal2 s 207754 169200 207810 170000 6 la_input[6]
port 120 nsew
rlabel metal2 s 243082 169200 243138 170000 6 la_input[70]
port 121 nsew
rlabel metal2 s 207386 169200 207442 170000 6 la_input[71]
port 122 nsew
rlabel metal2 s 243450 169200 243506 170000 6 la_input[72]
port 123 nsew
rlabel metal2 s 207018 169200 207074 170000 6 la_input[73]
port 124 nsew
rlabel metal2 s 243818 169200 243874 170000 6 la_input[74]
port 125 nsew
rlabel metal2 s 206650 169200 206706 170000 6 la_input[75]
port 126 nsew
rlabel metal2 s 244186 169200 244242 170000 6 la_input[76]
port 127 nsew
rlabel metal2 s 206282 169200 206338 170000 6 la_input[77]
port 128 nsew
rlabel metal2 s 244554 169200 244610 170000 6 la_input[78]
port 129 nsew
rlabel metal2 s 205914 169200 205970 170000 6 la_input[79]
port 130 nsew
rlabel metal2 s 244922 169200 244978 170000 6 la_input[7]
port 131 nsew
rlabel metal2 s 205546 169200 205602 170000 6 la_input[80]
port 132 nsew
rlabel metal2 s 245290 169200 245346 170000 6 la_input[81]
port 133 nsew
rlabel metal2 s 205178 169200 205234 170000 6 la_input[82]
port 134 nsew
rlabel metal2 s 245658 169200 245714 170000 6 la_input[83]
port 135 nsew
rlabel metal2 s 204810 169200 204866 170000 6 la_input[84]
port 136 nsew
rlabel metal2 s 246026 169200 246082 170000 6 la_input[85]
port 137 nsew
rlabel metal2 s 204442 169200 204498 170000 6 la_input[86]
port 138 nsew
rlabel metal2 s 246394 169200 246450 170000 6 la_input[87]
port 139 nsew
rlabel metal2 s 204074 169200 204130 170000 6 la_input[88]
port 140 nsew
rlabel metal2 s 246762 169200 246818 170000 6 la_input[89]
port 141 nsew
rlabel metal2 s 203706 169200 203762 170000 6 la_input[8]
port 142 nsew
rlabel metal2 s 247130 169200 247186 170000 6 la_input[90]
port 143 nsew
rlabel metal2 s 203338 169200 203394 170000 6 la_input[91]
port 144 nsew
rlabel metal2 s 247498 169200 247554 170000 6 la_input[92]
port 145 nsew
rlabel metal2 s 202970 169200 203026 170000 6 la_input[93]
port 146 nsew
rlabel metal2 s 247866 169200 247922 170000 6 la_input[94]
port 147 nsew
rlabel metal2 s 202602 169200 202658 170000 6 la_input[95]
port 148 nsew
rlabel metal2 s 248234 169200 248290 170000 6 la_input[96]
port 149 nsew
rlabel metal2 s 202234 169200 202290 170000 6 la_input[97]
port 150 nsew
rlabel metal2 s 248602 169200 248658 170000 6 la_input[98]
port 151 nsew
rlabel metal2 s 201866 169200 201922 170000 6 la_input[99]
port 152 nsew
rlabel metal2 s 248970 169200 249026 170000 6 la_input[9]
port 153 nsew
rlabel metal2 s 201498 169200 201554 170000 6 la_oen[0]
port 154 nsew
rlabel metal2 s 249338 169200 249394 170000 6 la_oen[100]
port 155 nsew
rlabel metal2 s 201130 169200 201186 170000 6 la_oen[101]
port 156 nsew
rlabel metal2 s 249706 169200 249762 170000 6 la_oen[102]
port 157 nsew
rlabel metal2 s 200762 169200 200818 170000 6 la_oen[103]
port 158 nsew
rlabel metal2 s 250074 169200 250130 170000 6 la_oen[104]
port 159 nsew
rlabel metal2 s 200394 169200 200450 170000 6 la_oen[105]
port 160 nsew
rlabel metal2 s 250442 169200 250498 170000 6 la_oen[106]
port 161 nsew
rlabel metal2 s 200026 169200 200082 170000 6 la_oen[107]
port 162 nsew
rlabel metal2 s 250810 169200 250866 170000 6 la_oen[108]
port 163 nsew
rlabel metal2 s 199658 169200 199714 170000 6 la_oen[109]
port 164 nsew
rlabel metal2 s 251178 169200 251234 170000 6 la_oen[10]
port 165 nsew
rlabel metal2 s 199290 169200 199346 170000 6 la_oen[110]
port 166 nsew
rlabel metal2 s 251546 169200 251602 170000 6 la_oen[111]
port 167 nsew
rlabel metal2 s 198922 169200 198978 170000 6 la_oen[112]
port 168 nsew
rlabel metal2 s 251914 169200 251970 170000 6 la_oen[113]
port 169 nsew
rlabel metal2 s 198554 169200 198610 170000 6 la_oen[114]
port 170 nsew
rlabel metal2 s 252282 169200 252338 170000 6 la_oen[115]
port 171 nsew
rlabel metal2 s 198186 169200 198242 170000 6 la_oen[116]
port 172 nsew
rlabel metal2 s 252650 169200 252706 170000 6 la_oen[117]
port 173 nsew
rlabel metal2 s 197818 169200 197874 170000 6 la_oen[118]
port 174 nsew
rlabel metal2 s 253018 169200 253074 170000 6 la_oen[119]
port 175 nsew
rlabel metal2 s 197450 169200 197506 170000 6 la_oen[11]
port 176 nsew
rlabel metal2 s 253386 169200 253442 170000 6 la_oen[120]
port 177 nsew
rlabel metal2 s 197082 169200 197138 170000 6 la_oen[121]
port 178 nsew
rlabel metal2 s 253754 169200 253810 170000 6 la_oen[122]
port 179 nsew
rlabel metal2 s 196714 169200 196770 170000 6 la_oen[123]
port 180 nsew
rlabel metal2 s 254122 169200 254178 170000 6 la_oen[124]
port 181 nsew
rlabel metal2 s 196346 169200 196402 170000 6 la_oen[125]
port 182 nsew
rlabel metal2 s 254490 169200 254546 170000 6 la_oen[126]
port 183 nsew
rlabel metal2 s 195978 169200 196034 170000 6 la_oen[127]
port 184 nsew
rlabel metal2 s 254858 169200 254914 170000 6 la_oen[12]
port 185 nsew
rlabel metal2 s 195610 169200 195666 170000 6 la_oen[13]
port 186 nsew
rlabel metal2 s 255226 169200 255282 170000 6 la_oen[14]
port 187 nsew
rlabel metal2 s 195242 169200 195298 170000 6 la_oen[15]
port 188 nsew
rlabel metal2 s 255594 169200 255650 170000 6 la_oen[16]
port 189 nsew
rlabel metal2 s 194874 169200 194930 170000 6 la_oen[17]
port 190 nsew
rlabel metal2 s 255962 169200 256018 170000 6 la_oen[18]
port 191 nsew
rlabel metal2 s 194506 169200 194562 170000 6 la_oen[19]
port 192 nsew
rlabel metal2 s 256330 169200 256386 170000 6 la_oen[1]
port 193 nsew
rlabel metal2 s 194138 169200 194194 170000 6 la_oen[20]
port 194 nsew
rlabel metal2 s 256698 169200 256754 170000 6 la_oen[21]
port 195 nsew
rlabel metal2 s 193770 169200 193826 170000 6 la_oen[22]
port 196 nsew
rlabel metal2 s 257066 169200 257122 170000 6 la_oen[23]
port 197 nsew
rlabel metal2 s 193402 169200 193458 170000 6 la_oen[24]
port 198 nsew
rlabel metal2 s 257434 169200 257490 170000 6 la_oen[25]
port 199 nsew
rlabel metal2 s 193034 169200 193090 170000 6 la_oen[26]
port 200 nsew
rlabel metal2 s 257802 169200 257858 170000 6 la_oen[27]
port 201 nsew
rlabel metal2 s 192666 169200 192722 170000 6 la_oen[28]
port 202 nsew
rlabel metal2 s 258170 169200 258226 170000 6 la_oen[29]
port 203 nsew
rlabel metal2 s 192298 169200 192354 170000 6 la_oen[2]
port 204 nsew
rlabel metal2 s 258538 169200 258594 170000 6 la_oen[30]
port 205 nsew
rlabel metal2 s 191930 169200 191986 170000 6 la_oen[31]
port 206 nsew
rlabel metal2 s 258906 169200 258962 170000 6 la_oen[32]
port 207 nsew
rlabel metal2 s 191562 169200 191618 170000 6 la_oen[33]
port 208 nsew
rlabel metal2 s 259274 169200 259330 170000 6 la_oen[34]
port 209 nsew
rlabel metal2 s 191194 169200 191250 170000 6 la_oen[35]
port 210 nsew
rlabel metal2 s 259642 169200 259698 170000 6 la_oen[36]
port 211 nsew
rlabel metal2 s 190826 169200 190882 170000 6 la_oen[37]
port 212 nsew
rlabel metal2 s 260010 169200 260066 170000 6 la_oen[38]
port 213 nsew
rlabel metal2 s 190458 169200 190514 170000 6 la_oen[39]
port 214 nsew
rlabel metal2 s 260378 169200 260434 170000 6 la_oen[3]
port 215 nsew
rlabel metal2 s 190090 169200 190146 170000 6 la_oen[40]
port 216 nsew
rlabel metal2 s 260746 169200 260802 170000 6 la_oen[41]
port 217 nsew
rlabel metal2 s 189722 169200 189778 170000 6 la_oen[42]
port 218 nsew
rlabel metal2 s 261114 169200 261170 170000 6 la_oen[43]
port 219 nsew
rlabel metal2 s 189354 169200 189410 170000 6 la_oen[44]
port 220 nsew
rlabel metal2 s 261482 169200 261538 170000 6 la_oen[45]
port 221 nsew
rlabel metal2 s 188986 169200 189042 170000 6 la_oen[46]
port 222 nsew
rlabel metal2 s 261850 169200 261906 170000 6 la_oen[47]
port 223 nsew
rlabel metal2 s 188618 169200 188674 170000 6 la_oen[48]
port 224 nsew
rlabel metal2 s 262218 169200 262274 170000 6 la_oen[49]
port 225 nsew
rlabel metal2 s 188250 169200 188306 170000 6 la_oen[4]
port 226 nsew
rlabel metal2 s 262586 169200 262642 170000 6 la_oen[50]
port 227 nsew
rlabel metal2 s 187882 169200 187938 170000 6 la_oen[51]
port 228 nsew
rlabel metal2 s 262954 169200 263010 170000 6 la_oen[52]
port 229 nsew
rlabel metal2 s 187514 169200 187570 170000 6 la_oen[53]
port 230 nsew
rlabel metal2 s 263322 169200 263378 170000 6 la_oen[54]
port 231 nsew
rlabel metal2 s 187146 169200 187202 170000 6 la_oen[55]
port 232 nsew
rlabel metal2 s 263690 169200 263746 170000 6 la_oen[56]
port 233 nsew
rlabel metal2 s 186778 169200 186834 170000 6 la_oen[57]
port 234 nsew
rlabel metal2 s 264058 169200 264114 170000 6 la_oen[58]
port 235 nsew
rlabel metal2 s 186410 169200 186466 170000 6 la_oen[59]
port 236 nsew
rlabel metal2 s 264426 169200 264482 170000 6 la_oen[5]
port 237 nsew
rlabel metal2 s 186042 169200 186098 170000 6 la_oen[60]
port 238 nsew
rlabel metal2 s 264794 169200 264850 170000 6 la_oen[61]
port 239 nsew
rlabel metal2 s 185674 169200 185730 170000 6 la_oen[62]
port 240 nsew
rlabel metal2 s 265162 169200 265218 170000 6 la_oen[63]
port 241 nsew
rlabel metal2 s 185306 169200 185362 170000 6 la_oen[64]
port 242 nsew
rlabel metal2 s 265530 169200 265586 170000 6 la_oen[65]
port 243 nsew
rlabel metal2 s 184938 169200 184994 170000 6 la_oen[66]
port 244 nsew
rlabel metal2 s 265898 169200 265954 170000 6 la_oen[67]
port 245 nsew
rlabel metal2 s 184570 169200 184626 170000 6 la_oen[68]
port 246 nsew
rlabel metal2 s 266266 169200 266322 170000 6 la_oen[69]
port 247 nsew
rlabel metal2 s 184202 169200 184258 170000 6 la_oen[6]
port 248 nsew
rlabel metal2 s 266634 169200 266690 170000 6 la_oen[70]
port 249 nsew
rlabel metal2 s 183834 169200 183890 170000 6 la_oen[71]
port 250 nsew
rlabel metal2 s 267002 169200 267058 170000 6 la_oen[72]
port 251 nsew
rlabel metal2 s 183466 169200 183522 170000 6 la_oen[73]
port 252 nsew
rlabel metal2 s 267370 169200 267426 170000 6 la_oen[74]
port 253 nsew
rlabel metal2 s 183098 169200 183154 170000 6 la_oen[75]
port 254 nsew
rlabel metal2 s 267738 169200 267794 170000 6 la_oen[76]
port 255 nsew
rlabel metal2 s 182730 169200 182786 170000 6 la_oen[77]
port 256 nsew
rlabel metal2 s 268106 169200 268162 170000 6 la_oen[78]
port 257 nsew
rlabel metal2 s 182362 169200 182418 170000 6 la_oen[79]
port 258 nsew
rlabel metal2 s 268474 169200 268530 170000 6 la_oen[7]
port 259 nsew
rlabel metal2 s 181994 169200 182050 170000 6 la_oen[80]
port 260 nsew
rlabel metal2 s 268842 169200 268898 170000 6 la_oen[81]
port 261 nsew
rlabel metal2 s 181626 169200 181682 170000 6 la_oen[82]
port 262 nsew
rlabel metal2 s 269210 169200 269266 170000 6 la_oen[83]
port 263 nsew
rlabel metal2 s 181258 169200 181314 170000 6 la_oen[84]
port 264 nsew
rlabel metal2 s 269578 169200 269634 170000 6 la_oen[85]
port 265 nsew
rlabel metal2 s 180890 169200 180946 170000 6 la_oen[86]
port 266 nsew
rlabel metal2 s 269946 169200 270002 170000 6 la_oen[87]
port 267 nsew
rlabel metal2 s 180522 169200 180578 170000 6 la_oen[88]
port 268 nsew
rlabel metal2 s 270314 169200 270370 170000 6 la_oen[89]
port 269 nsew
rlabel metal2 s 180154 169200 180210 170000 6 la_oen[8]
port 270 nsew
rlabel metal2 s 270682 169200 270738 170000 6 la_oen[90]
port 271 nsew
rlabel metal2 s 179786 169200 179842 170000 6 la_oen[91]
port 272 nsew
rlabel metal2 s 271050 169200 271106 170000 6 la_oen[92]
port 273 nsew
rlabel metal2 s 179418 169200 179474 170000 6 la_oen[93]
port 274 nsew
rlabel metal2 s 271418 169200 271474 170000 6 la_oen[94]
port 275 nsew
rlabel metal2 s 179050 169200 179106 170000 6 la_oen[95]
port 276 nsew
rlabel metal2 s 271786 169200 271842 170000 6 la_oen[96]
port 277 nsew
rlabel metal2 s 178682 169200 178738 170000 6 la_oen[97]
port 278 nsew
rlabel metal2 s 272154 169200 272210 170000 6 la_oen[98]
port 279 nsew
rlabel metal2 s 178314 169200 178370 170000 6 la_oen[99]
port 280 nsew
rlabel metal2 s 272522 169200 272578 170000 6 la_oen[9]
port 281 nsew
rlabel metal2 s 177946 169200 178002 170000 6 la_output[0]
port 282 nsew
rlabel metal2 s 272890 169200 272946 170000 6 la_output[100]
port 283 nsew
rlabel metal2 s 177578 169200 177634 170000 6 la_output[101]
port 284 nsew
rlabel metal2 s 273258 169200 273314 170000 6 la_output[102]
port 285 nsew
rlabel metal2 s 177210 169200 177266 170000 6 la_output[103]
port 286 nsew
rlabel metal2 s 273626 169200 273682 170000 6 la_output[104]
port 287 nsew
rlabel metal2 s 176842 169200 176898 170000 6 la_output[105]
port 288 nsew
rlabel metal2 s 273994 169200 274050 170000 6 la_output[106]
port 289 nsew
rlabel metal2 s 176474 169200 176530 170000 6 la_output[107]
port 290 nsew
rlabel metal2 s 274362 169200 274418 170000 6 la_output[108]
port 291 nsew
rlabel metal2 s 176106 169200 176162 170000 6 la_output[109]
port 292 nsew
rlabel metal2 s 274730 169200 274786 170000 6 la_output[10]
port 293 nsew
rlabel metal2 s 175738 169200 175794 170000 6 la_output[110]
port 294 nsew
rlabel metal2 s 275098 169200 275154 170000 6 la_output[111]
port 295 nsew
rlabel metal2 s 175370 169200 175426 170000 6 la_output[112]
port 296 nsew
rlabel metal2 s 275466 169200 275522 170000 6 la_output[113]
port 297 nsew
rlabel metal2 s 175002 169200 175058 170000 6 la_output[114]
port 298 nsew
rlabel metal2 s 275834 169200 275890 170000 6 la_output[115]
port 299 nsew
rlabel metal2 s 174634 169200 174690 170000 6 la_output[116]
port 300 nsew
rlabel metal2 s 276202 169200 276258 170000 6 la_output[117]
port 301 nsew
rlabel metal2 s 174266 169200 174322 170000 6 la_output[118]
port 302 nsew
rlabel metal2 s 276570 169200 276626 170000 6 la_output[119]
port 303 nsew
rlabel metal2 s 173898 169200 173954 170000 6 la_output[11]
port 304 nsew
rlabel metal2 s 276938 169200 276994 170000 6 la_output[120]
port 305 nsew
rlabel metal2 s 173530 169200 173586 170000 6 la_output[121]
port 306 nsew
rlabel metal2 s 277306 169200 277362 170000 6 la_output[122]
port 307 nsew
rlabel metal2 s 173162 169200 173218 170000 6 la_output[123]
port 308 nsew
rlabel metal2 s 277674 169200 277730 170000 6 la_output[124]
port 309 nsew
rlabel metal2 s 172794 169200 172850 170000 6 la_output[125]
port 310 nsew
rlabel metal2 s 278042 169200 278098 170000 6 la_output[126]
port 311 nsew
rlabel metal2 s 172426 169200 172482 170000 6 la_output[127]
port 312 nsew
rlabel metal2 s 278410 169200 278466 170000 6 la_output[12]
port 313 nsew
rlabel metal2 s 172058 169200 172114 170000 6 la_output[13]
port 314 nsew
rlabel metal2 s 278778 169200 278834 170000 6 la_output[14]
port 315 nsew
rlabel metal2 s 171690 169200 171746 170000 6 la_output[15]
port 316 nsew
rlabel metal2 s 279146 169200 279202 170000 6 la_output[16]
port 317 nsew
rlabel metal2 s 171322 169200 171378 170000 6 la_output[17]
port 318 nsew
rlabel metal2 s 279514 169200 279570 170000 6 la_output[18]
port 319 nsew
rlabel metal2 s 170954 169200 171010 170000 6 la_output[19]
port 320 nsew
rlabel metal2 s 279882 169200 279938 170000 6 la_output[1]
port 321 nsew
rlabel metal2 s 170586 169200 170642 170000 6 la_output[20]
port 322 nsew
rlabel metal2 s 280250 169200 280306 170000 6 la_output[21]
port 323 nsew
rlabel metal2 s 170218 169200 170274 170000 6 la_output[22]
port 324 nsew
rlabel metal2 s 280618 169200 280674 170000 6 la_output[23]
port 325 nsew
rlabel metal2 s 169850 169200 169906 170000 6 la_output[24]
port 326 nsew
rlabel metal2 s 280986 169200 281042 170000 6 la_output[25]
port 327 nsew
rlabel metal2 s 169482 169200 169538 170000 6 la_output[26]
port 328 nsew
rlabel metal2 s 281354 169200 281410 170000 6 la_output[27]
port 329 nsew
rlabel metal2 s 169114 169200 169170 170000 6 la_output[28]
port 330 nsew
rlabel metal2 s 281722 169200 281778 170000 6 la_output[29]
port 331 nsew
rlabel metal2 s 168746 169200 168802 170000 6 la_output[2]
port 332 nsew
rlabel metal2 s 282090 169200 282146 170000 6 la_output[30]
port 333 nsew
rlabel metal2 s 168378 169200 168434 170000 6 la_output[31]
port 334 nsew
rlabel metal2 s 282458 169200 282514 170000 6 la_output[32]
port 335 nsew
rlabel metal2 s 168010 169200 168066 170000 6 la_output[33]
port 336 nsew
rlabel metal2 s 282826 169200 282882 170000 6 la_output[34]
port 337 nsew
rlabel metal2 s 167642 169200 167698 170000 6 la_output[35]
port 338 nsew
rlabel metal2 s 283194 169200 283250 170000 6 la_output[36]
port 339 nsew
rlabel metal2 s 167274 169200 167330 170000 6 la_output[37]
port 340 nsew
rlabel metal2 s 283562 169200 283618 170000 6 la_output[38]
port 341 nsew
rlabel metal2 s 166906 169200 166962 170000 6 la_output[39]
port 342 nsew
rlabel metal2 s 283930 169200 283986 170000 6 la_output[3]
port 343 nsew
rlabel metal2 s 166538 169200 166594 170000 6 la_output[40]
port 344 nsew
rlabel metal2 s 284298 169200 284354 170000 6 la_output[41]
port 345 nsew
rlabel metal2 s 166170 169200 166226 170000 6 la_output[42]
port 346 nsew
rlabel metal2 s 284666 169200 284722 170000 6 la_output[43]
port 347 nsew
rlabel metal2 s 165802 169200 165858 170000 6 la_output[44]
port 348 nsew
rlabel metal2 s 285034 169200 285090 170000 6 la_output[45]
port 349 nsew
rlabel metal2 s 165434 169200 165490 170000 6 la_output[46]
port 350 nsew
rlabel metal2 s 285402 169200 285458 170000 6 la_output[47]
port 351 nsew
rlabel metal2 s 165066 169200 165122 170000 6 la_output[48]
port 352 nsew
rlabel metal2 s 285770 169200 285826 170000 6 la_output[49]
port 353 nsew
rlabel metal2 s 164698 169200 164754 170000 6 la_output[4]
port 354 nsew
rlabel metal2 s 286138 169200 286194 170000 6 la_output[50]
port 355 nsew
rlabel metal2 s 164330 169200 164386 170000 6 la_output[51]
port 356 nsew
rlabel metal2 s 286506 169200 286562 170000 6 la_output[52]
port 357 nsew
rlabel metal2 s 163962 169200 164018 170000 6 la_output[53]
port 358 nsew
rlabel metal2 s 286874 169200 286930 170000 6 la_output[54]
port 359 nsew
rlabel metal2 s 163594 169200 163650 170000 6 la_output[55]
port 360 nsew
rlabel metal2 s 287242 169200 287298 170000 6 la_output[56]
port 361 nsew
rlabel metal2 s 163226 169200 163282 170000 6 la_output[57]
port 362 nsew
rlabel metal2 s 287610 169200 287666 170000 6 la_output[58]
port 363 nsew
rlabel metal2 s 162858 169200 162914 170000 6 la_output[59]
port 364 nsew
rlabel metal2 s 287978 169200 288034 170000 6 la_output[5]
port 365 nsew
rlabel metal2 s 162490 169200 162546 170000 6 la_output[60]
port 366 nsew
rlabel metal2 s 288346 169200 288402 170000 6 la_output[61]
port 367 nsew
rlabel metal2 s 162122 169200 162178 170000 6 la_output[62]
port 368 nsew
rlabel metal2 s 288714 169200 288770 170000 6 la_output[63]
port 369 nsew
rlabel metal2 s 161754 169200 161810 170000 6 la_output[64]
port 370 nsew
rlabel metal2 s 289082 169200 289138 170000 6 la_output[65]
port 371 nsew
rlabel metal2 s 161386 169200 161442 170000 6 la_output[66]
port 372 nsew
rlabel metal2 s 289450 169200 289506 170000 6 la_output[67]
port 373 nsew
rlabel metal2 s 161018 169200 161074 170000 6 la_output[68]
port 374 nsew
rlabel metal2 s 289818 169200 289874 170000 6 la_output[69]
port 375 nsew
rlabel metal2 s 160650 169200 160706 170000 6 la_output[6]
port 376 nsew
rlabel metal2 s 290186 169200 290242 170000 6 la_output[70]
port 377 nsew
rlabel metal2 s 160282 169200 160338 170000 6 la_output[71]
port 378 nsew
rlabel metal2 s 290554 169200 290610 170000 6 la_output[72]
port 379 nsew
rlabel metal2 s 159914 169200 159970 170000 6 la_output[73]
port 380 nsew
rlabel metal2 s 290922 169200 290978 170000 6 la_output[74]
port 381 nsew
rlabel metal2 s 159546 169200 159602 170000 6 la_output[75]
port 382 nsew
rlabel metal2 s 291290 169200 291346 170000 6 la_output[76]
port 383 nsew
rlabel metal2 s 159178 169200 159234 170000 6 la_output[77]
port 384 nsew
rlabel metal2 s 291658 169200 291714 170000 6 la_output[78]
port 385 nsew
rlabel metal2 s 158810 169200 158866 170000 6 la_output[79]
port 386 nsew
rlabel metal2 s 292026 169200 292082 170000 6 la_output[7]
port 387 nsew
rlabel metal2 s 158442 169200 158498 170000 6 la_output[80]
port 388 nsew
rlabel metal2 s 292394 169200 292450 170000 6 la_output[81]
port 389 nsew
rlabel metal2 s 158074 169200 158130 170000 6 la_output[82]
port 390 nsew
rlabel metal2 s 292762 169200 292818 170000 6 la_output[83]
port 391 nsew
rlabel metal2 s 157706 169200 157762 170000 6 la_output[84]
port 392 nsew
rlabel metal2 s 293130 169200 293186 170000 6 la_output[85]
port 393 nsew
rlabel metal2 s 157338 169200 157394 170000 6 la_output[86]
port 394 nsew
rlabel metal2 s 293498 169200 293554 170000 6 la_output[87]
port 395 nsew
rlabel metal2 s 156970 169200 157026 170000 6 la_output[88]
port 396 nsew
rlabel metal2 s 293866 169200 293922 170000 6 la_output[89]
port 397 nsew
rlabel metal2 s 156602 169200 156658 170000 6 la_output[8]
port 398 nsew
rlabel metal2 s 294234 169200 294290 170000 6 la_output[90]
port 399 nsew
rlabel metal2 s 156234 169200 156290 170000 6 la_output[91]
port 400 nsew
rlabel metal2 s 294602 169200 294658 170000 6 la_output[92]
port 401 nsew
rlabel metal2 s 155866 169200 155922 170000 6 la_output[93]
port 402 nsew
rlabel metal2 s 294970 169200 295026 170000 6 la_output[94]
port 403 nsew
rlabel metal2 s 155498 169200 155554 170000 6 la_output[95]
port 404 nsew
rlabel metal2 s 295338 169200 295394 170000 6 la_output[96]
port 405 nsew
rlabel metal2 s 155130 169200 155186 170000 6 la_output[97]
port 406 nsew
rlabel metal2 s 295706 169200 295762 170000 6 la_output[98]
port 407 nsew
rlabel metal2 s 154762 169200 154818 170000 6 la_output[99]
port 408 nsew
rlabel metal2 s 296074 169200 296130 170000 6 la_output[9]
port 409 nsew
rlabel metal2 s 429290 0 429346 800 6 mask_rev[0]
port 410 nsew
rlabel metal2 s 428922 0 428978 800 6 mask_rev[10]
port 411 nsew
rlabel metal3 s 429200 1096 430000 1216 6 mask_rev[11]
port 412 nsew
rlabel metal2 s 428554 0 428610 800 6 mask_rev[12]
port 413 nsew
rlabel metal3 s 429200 1640 430000 1760 6 mask_rev[13]
port 414 nsew
rlabel metal2 s 428186 0 428242 800 6 mask_rev[14]
port 415 nsew
rlabel metal2 s 427818 0 427874 800 6 mask_rev[15]
port 416 nsew
rlabel metal3 s 429200 2184 430000 2304 6 mask_rev[16]
port 417 nsew
rlabel metal2 s 427450 0 427506 800 6 mask_rev[17]
port 418 nsew
rlabel metal3 s 429200 2728 430000 2848 6 mask_rev[18]
port 419 nsew
rlabel metal2 s 427082 0 427138 800 6 mask_rev[19]
port 420 nsew
rlabel metal2 s 426714 0 426770 800 6 mask_rev[1]
port 421 nsew
rlabel metal3 s 429200 3272 430000 3392 6 mask_rev[20]
port 422 nsew
rlabel metal2 s 426346 0 426402 800 6 mask_rev[21]
port 423 nsew
rlabel metal3 s 429200 3816 430000 3936 6 mask_rev[22]
port 424 nsew
rlabel metal2 s 425978 0 426034 800 6 mask_rev[23]
port 425 nsew
rlabel metal2 s 425610 0 425666 800 6 mask_rev[24]
port 426 nsew
rlabel metal3 s 429200 4360 430000 4480 6 mask_rev[25]
port 427 nsew
rlabel metal2 s 425242 0 425298 800 6 mask_rev[26]
port 428 nsew
rlabel metal3 s 429200 4904 430000 5024 6 mask_rev[27]
port 429 nsew
rlabel metal2 s 424874 0 424930 800 6 mask_rev[28]
port 430 nsew
rlabel metal2 s 424506 0 424562 800 6 mask_rev[29]
port 431 nsew
rlabel metal3 s 429200 5448 430000 5568 6 mask_rev[2]
port 432 nsew
rlabel metal2 s 424138 0 424194 800 6 mask_rev[30]
port 433 nsew
rlabel metal3 s 429200 5992 430000 6112 6 mask_rev[31]
port 434 nsew
rlabel metal2 s 423770 0 423826 800 6 mask_rev[3]
port 435 nsew
rlabel metal2 s 423402 0 423458 800 6 mask_rev[4]
port 436 nsew
rlabel metal3 s 429200 6536 430000 6656 6 mask_rev[5]
port 437 nsew
rlabel metal2 s 423034 0 423090 800 6 mask_rev[6]
port 438 nsew
rlabel metal3 s 429200 7080 430000 7200 6 mask_rev[7]
port 439 nsew
rlabel metal2 s 422666 0 422722 800 6 mask_rev[8]
port 440 nsew
rlabel metal2 s 422298 0 422354 800 6 mask_rev[9]
port 441 nsew
rlabel metal2 s 5354 0 5410 800 6 mgmt_addr[0]
port 442 nsew
rlabel metal3 s 0 5448 800 5568 6 mgmt_addr[1]
port 443 nsew
rlabel metal2 s 5722 0 5778 800 6 mgmt_addr[2]
port 444 nsew
rlabel metal3 s 0 5992 800 6112 6 mgmt_addr[3]
port 445 nsew
rlabel metal2 s 6090 0 6146 800 6 mgmt_addr[4]
port 446 nsew
rlabel metal2 s 6458 0 6514 800 6 mgmt_addr[5]
port 447 nsew
rlabel metal3 s 0 6536 800 6656 6 mgmt_addr[6]
port 448 nsew
rlabel metal2 s 6826 0 6882 800 6 mgmt_addr[7]
port 449 nsew
rlabel metal3 s 0 7080 800 7200 6 mgmt_addr_ro[0]
port 450 nsew
rlabel metal2 s 7194 0 7250 800 6 mgmt_addr_ro[1]
port 451 nsew
rlabel metal2 s 7562 0 7618 800 6 mgmt_addr_ro[2]
port 452 nsew
rlabel metal3 s 0 7624 800 7744 6 mgmt_addr_ro[3]
port 453 nsew
rlabel metal2 s 7930 0 7986 800 6 mgmt_addr_ro[4]
port 454 nsew
rlabel metal3 s 0 8168 800 8288 6 mgmt_addr_ro[5]
port 455 nsew
rlabel metal2 s 8298 0 8354 800 6 mgmt_addr_ro[6]
port 456 nsew
rlabel metal2 s 8666 0 8722 800 6 mgmt_addr_ro[7]
port 457 nsew
rlabel metal3 s 0 8712 800 8832 6 mgmt_ena[0]
port 458 nsew
rlabel metal2 s 9034 0 9090 800 6 mgmt_ena[1]
port 459 nsew
rlabel metal3 s 0 9256 800 9376 6 mgmt_ena_ro
port 460 nsew
rlabel metal3 s 429200 68008 430000 68128 6 mgmt_in_data[0]
port 461 nsew
rlabel metal2 s 754 0 810 800 6 mgmt_in_data[10]
port 462 nsew
rlabel metal2 s 1122 0 1178 800 6 mgmt_in_data[11]
port 463 nsew
rlabel metal2 s 1490 0 1546 800 6 mgmt_in_data[12]
port 464 nsew
rlabel metal2 s 1858 0 1914 800 6 mgmt_in_data[13]
port 465 nsew
rlabel metal2 s 2226 0 2282 800 6 mgmt_in_data[14]
port 466 nsew
rlabel metal2 s 2594 0 2650 800 6 mgmt_in_data[15]
port 467 nsew
rlabel metal2 s 2962 0 3018 800 6 mgmt_in_data[16]
port 468 nsew
rlabel metal2 s 3330 0 3386 800 6 mgmt_in_data[17]
port 469 nsew
rlabel metal2 s 3698 0 3754 800 6 mgmt_in_data[18]
port 470 nsew
rlabel metal2 s 4066 0 4122 800 6 mgmt_in_data[19]
port 471 nsew
rlabel metal3 s 429200 112616 430000 112736 6 mgmt_in_data[1]
port 472 nsew
rlabel metal2 s 4434 0 4490 800 6 mgmt_in_data[20]
port 473 nsew
rlabel metal2 s 4802 0 4858 800 6 mgmt_in_data[21]
port 474 nsew
rlabel metal2 s 5170 0 5226 800 6 mgmt_in_data[22]
port 475 nsew
rlabel metal2 s 5538 0 5594 800 6 mgmt_in_data[23]
port 476 nsew
rlabel metal2 s 5906 0 5962 800 6 mgmt_in_data[24]
port 477 nsew
rlabel metal2 s 6274 0 6330 800 6 mgmt_in_data[25]
port 478 nsew
rlabel metal2 s 6642 0 6698 800 6 mgmt_in_data[26]
port 479 nsew
rlabel metal2 s 7010 0 7066 800 6 mgmt_in_data[27]
port 480 nsew
rlabel metal2 s 7378 0 7434 800 6 mgmt_in_data[28]
port 481 nsew
rlabel metal2 s 7746 0 7802 800 6 mgmt_in_data[29]
port 482 nsew
rlabel metal2 s 8114 0 8170 800 6 mgmt_in_data[2]
port 483 nsew
rlabel metal2 s 8482 0 8538 800 6 mgmt_in_data[30]
port 484 nsew
rlabel metal2 s 8850 0 8906 800 6 mgmt_in_data[31]
port 485 nsew
rlabel metal2 s 9218 0 9274 800 6 mgmt_in_data[32]
port 486 nsew
rlabel metal2 s 9586 0 9642 800 6 mgmt_in_data[33]
port 487 nsew
rlabel metal2 s 9954 0 10010 800 6 mgmt_in_data[34]
port 488 nsew
rlabel metal2 s 10322 0 10378 800 6 mgmt_in_data[35]
port 489 nsew
rlabel metal2 s 10690 0 10746 800 6 mgmt_in_data[36]
port 490 nsew
rlabel metal2 s 11058 0 11114 800 6 mgmt_in_data[37]
port 491 nsew
rlabel metal2 s 11426 0 11482 800 6 mgmt_in_data[3]
port 492 nsew
rlabel metal2 s 11794 0 11850 800 6 mgmt_in_data[4]
port 493 nsew
rlabel metal2 s 12162 0 12218 800 6 mgmt_in_data[5]
port 494 nsew
rlabel metal2 s 12530 0 12586 800 6 mgmt_in_data[6]
port 495 nsew
rlabel metal2 s 12898 0 12954 800 6 mgmt_in_data[7]
port 496 nsew
rlabel metal2 s 13266 0 13322 800 6 mgmt_in_data[8]
port 497 nsew
rlabel metal2 s 13634 0 13690 800 6 mgmt_in_data[9]
port 498 nsew
rlabel metal2 s 14002 0 14058 800 6 mgmt_out_data[0]
port 499 nsew
rlabel metal2 s 429290 169200 429346 170000 6 mgmt_out_data[10]
port 500 nsew
rlabel metal2 s 428922 169200 428978 170000 6 mgmt_out_data[11]
port 501 nsew
rlabel metal3 s 429200 168648 430000 168768 6 mgmt_out_data[12]
port 502 nsew
rlabel metal2 s 428554 169200 428610 170000 6 mgmt_out_data[13]
port 503 nsew
rlabel metal2 s 428186 169200 428242 170000 6 mgmt_out_data[14]
port 504 nsew
rlabel metal2 s 335082 169200 335138 170000 6 mgmt_out_data[15]
port 505 nsew
rlabel metal2 s 296442 169200 296498 170000 6 mgmt_out_data[16]
port 506 nsew
rlabel metal2 s 154394 169200 154450 170000 6 mgmt_out_data[17]
port 507 nsew
rlabel metal2 s 139306 169200 139362 170000 6 mgmt_out_data[18]
port 508 nsew
rlabel metal2 s 88890 169200 88946 170000 6 mgmt_out_data[19]
port 509 nsew
rlabel metal2 s 14370 0 14426 800 6 mgmt_out_data[1]
port 510 nsew
rlabel metal2 s 37370 169200 37426 170000 6 mgmt_out_data[20]
port 511 nsew
rlabel metal2 s 570 169200 626 170000 6 mgmt_out_data[21]
port 512 nsew
rlabel metal2 s 938 169200 994 170000 6 mgmt_out_data[22]
port 513 nsew
rlabel metal3 s 0 168648 800 168768 6 mgmt_out_data[23]
port 514 nsew
rlabel metal2 s 1306 169200 1362 170000 6 mgmt_out_data[24]
port 515 nsew
rlabel metal2 s 1674 169200 1730 170000 6 mgmt_out_data[25]
port 516 nsew
rlabel metal3 s 0 168104 800 168224 6 mgmt_out_data[26]
port 517 nsew
rlabel metal2 s 2042 169200 2098 170000 6 mgmt_out_data[27]
port 518 nsew
rlabel metal3 s 0 167560 800 167680 6 mgmt_out_data[28]
port 519 nsew
rlabel metal2 s 2410 169200 2466 170000 6 mgmt_out_data[29]
port 520 nsew
rlabel metal3 s 429200 157224 430000 157344 6 mgmt_out_data[2]
port 521 nsew
rlabel metal2 s 2778 169200 2834 170000 6 mgmt_out_data[30]
port 522 nsew
rlabel metal3 s 0 167016 800 167136 6 mgmt_out_data[31]
port 523 nsew
rlabel metal2 s 3146 169200 3202 170000 6 mgmt_out_data[32]
port 524 nsew
rlabel metal3 s 0 166472 800 166592 6 mgmt_out_data[33]
port 525 nsew
rlabel metal2 s 3514 169200 3570 170000 6 mgmt_out_data[34]
port 526 nsew
rlabel metal2 s 3882 169200 3938 170000 6 mgmt_out_data[35]
port 527 nsew
rlabel metal3 s 0 165928 800 166048 6 mgmt_out_data[36]
port 528 nsew
rlabel metal3 s 0 149064 800 149184 6 mgmt_out_data[37]
port 529 nsew
rlabel metal3 s 429200 168104 430000 168224 6 mgmt_out_data[3]
port 530 nsew
rlabel metal2 s 427818 169200 427874 170000 6 mgmt_out_data[4]
port 531 nsew
rlabel metal3 s 429200 167560 430000 167680 6 mgmt_out_data[5]
port 532 nsew
rlabel metal2 s 427450 169200 427506 170000 6 mgmt_out_data[6]
port 533 nsew
rlabel metal2 s 427082 169200 427138 170000 6 mgmt_out_data[7]
port 534 nsew
rlabel metal3 s 429200 167016 430000 167136 6 mgmt_out_data[8]
port 535 nsew
rlabel metal2 s 426714 169200 426770 170000 6 mgmt_out_data[9]
port 536 nsew
rlabel metal2 s 9402 0 9458 800 6 mgmt_rdata[0]
port 537 nsew
rlabel metal2 s 9770 0 9826 800 6 mgmt_rdata[10]
port 538 nsew
rlabel metal3 s 0 9800 800 9920 6 mgmt_rdata[11]
port 539 nsew
rlabel metal2 s 10138 0 10194 800 6 mgmt_rdata[12]
port 540 nsew
rlabel metal3 s 0 10344 800 10464 6 mgmt_rdata[13]
port 541 nsew
rlabel metal2 s 10506 0 10562 800 6 mgmt_rdata[14]
port 542 nsew
rlabel metal2 s 10874 0 10930 800 6 mgmt_rdata[15]
port 543 nsew
rlabel metal3 s 0 10888 800 11008 6 mgmt_rdata[16]
port 544 nsew
rlabel metal2 s 11242 0 11298 800 6 mgmt_rdata[17]
port 545 nsew
rlabel metal3 s 0 11432 800 11552 6 mgmt_rdata[18]
port 546 nsew
rlabel metal2 s 11610 0 11666 800 6 mgmt_rdata[19]
port 547 nsew
rlabel metal2 s 11978 0 12034 800 6 mgmt_rdata[1]
port 548 nsew
rlabel metal3 s 0 11976 800 12096 6 mgmt_rdata[20]
port 549 nsew
rlabel metal2 s 12346 0 12402 800 6 mgmt_rdata[21]
port 550 nsew
rlabel metal3 s 0 12520 800 12640 6 mgmt_rdata[22]
port 551 nsew
rlabel metal2 s 12714 0 12770 800 6 mgmt_rdata[23]
port 552 nsew
rlabel metal2 s 13082 0 13138 800 6 mgmt_rdata[24]
port 553 nsew
rlabel metal3 s 0 13064 800 13184 6 mgmt_rdata[25]
port 554 nsew
rlabel metal2 s 13450 0 13506 800 6 mgmt_rdata[26]
port 555 nsew
rlabel metal3 s 0 13608 800 13728 6 mgmt_rdata[27]
port 556 nsew
rlabel metal2 s 13818 0 13874 800 6 mgmt_rdata[28]
port 557 nsew
rlabel metal3 s 0 14152 800 14272 6 mgmt_rdata[29]
port 558 nsew
rlabel metal2 s 14186 0 14242 800 6 mgmt_rdata[2]
port 559 nsew
rlabel metal2 s 14554 0 14610 800 6 mgmt_rdata[30]
port 560 nsew
rlabel metal3 s 0 14696 800 14816 6 mgmt_rdata[31]
port 561 nsew
rlabel metal2 s 14922 0 14978 800 6 mgmt_rdata[32]
port 562 nsew
rlabel metal3 s 0 15240 800 15360 6 mgmt_rdata[33]
port 563 nsew
rlabel metal2 s 15290 0 15346 800 6 mgmt_rdata[34]
port 564 nsew
rlabel metal2 s 15658 0 15714 800 6 mgmt_rdata[35]
port 565 nsew
rlabel metal3 s 0 15784 800 15904 6 mgmt_rdata[36]
port 566 nsew
rlabel metal2 s 16026 0 16082 800 6 mgmt_rdata[37]
port 567 nsew
rlabel metal3 s 0 16328 800 16448 6 mgmt_rdata[38]
port 568 nsew
rlabel metal2 s 16394 0 16450 800 6 mgmt_rdata[39]
port 569 nsew
rlabel metal2 s 16762 0 16818 800 6 mgmt_rdata[3]
port 570 nsew
rlabel metal3 s 0 16872 800 16992 6 mgmt_rdata[40]
port 571 nsew
rlabel metal2 s 17130 0 17186 800 6 mgmt_rdata[41]
port 572 nsew
rlabel metal3 s 0 17416 800 17536 6 mgmt_rdata[42]
port 573 nsew
rlabel metal2 s 17498 0 17554 800 6 mgmt_rdata[43]
port 574 nsew
rlabel metal2 s 17866 0 17922 800 6 mgmt_rdata[44]
port 575 nsew
rlabel metal3 s 0 17960 800 18080 6 mgmt_rdata[45]
port 576 nsew
rlabel metal2 s 18234 0 18290 800 6 mgmt_rdata[46]
port 577 nsew
rlabel metal3 s 0 18504 800 18624 6 mgmt_rdata[47]
port 578 nsew
rlabel metal2 s 18602 0 18658 800 6 mgmt_rdata[48]
port 579 nsew
rlabel metal2 s 18970 0 19026 800 6 mgmt_rdata[49]
port 580 nsew
rlabel metal3 s 0 19048 800 19168 6 mgmt_rdata[4]
port 581 nsew
rlabel metal2 s 19338 0 19394 800 6 mgmt_rdata[50]
port 582 nsew
rlabel metal3 s 0 19592 800 19712 6 mgmt_rdata[51]
port 583 nsew
rlabel metal2 s 19706 0 19762 800 6 mgmt_rdata[52]
port 584 nsew
rlabel metal2 s 20074 0 20130 800 6 mgmt_rdata[53]
port 585 nsew
rlabel metal3 s 0 20136 800 20256 6 mgmt_rdata[54]
port 586 nsew
rlabel metal2 s 20442 0 20498 800 6 mgmt_rdata[55]
port 587 nsew
rlabel metal3 s 0 20680 800 20800 6 mgmt_rdata[56]
port 588 nsew
rlabel metal2 s 20810 0 20866 800 6 mgmt_rdata[57]
port 589 nsew
rlabel metal2 s 21178 0 21234 800 6 mgmt_rdata[58]
port 590 nsew
rlabel metal3 s 0 21224 800 21344 6 mgmt_rdata[59]
port 591 nsew
rlabel metal2 s 21546 0 21602 800 6 mgmt_rdata[5]
port 592 nsew
rlabel metal3 s 0 21768 800 21888 6 mgmt_rdata[60]
port 593 nsew
rlabel metal2 s 21914 0 21970 800 6 mgmt_rdata[61]
port 594 nsew
rlabel metal2 s 22282 0 22338 800 6 mgmt_rdata[62]
port 595 nsew
rlabel metal3 s 0 22312 800 22432 6 mgmt_rdata[63]
port 596 nsew
rlabel metal2 s 22650 0 22706 800 6 mgmt_rdata[6]
port 597 nsew
rlabel metal3 s 0 22856 800 22976 6 mgmt_rdata[7]
port 598 nsew
rlabel metal2 s 23018 0 23074 800 6 mgmt_rdata[8]
port 599 nsew
rlabel metal2 s 23386 0 23442 800 6 mgmt_rdata[9]
port 600 nsew
rlabel metal3 s 0 23400 800 23520 6 mgmt_rdata_ro[0]
port 601 nsew
rlabel metal2 s 23754 0 23810 800 6 mgmt_rdata_ro[10]
port 602 nsew
rlabel metal3 s 0 23944 800 24064 6 mgmt_rdata_ro[11]
port 603 nsew
rlabel metal2 s 24122 0 24178 800 6 mgmt_rdata_ro[12]
port 604 nsew
rlabel metal2 s 24490 0 24546 800 6 mgmt_rdata_ro[13]
port 605 nsew
rlabel metal3 s 0 24488 800 24608 6 mgmt_rdata_ro[14]
port 606 nsew
rlabel metal2 s 24858 0 24914 800 6 mgmt_rdata_ro[15]
port 607 nsew
rlabel metal3 s 0 25032 800 25152 6 mgmt_rdata_ro[16]
port 608 nsew
rlabel metal2 s 25226 0 25282 800 6 mgmt_rdata_ro[17]
port 609 nsew
rlabel metal2 s 25594 0 25650 800 6 mgmt_rdata_ro[18]
port 610 nsew
rlabel metal3 s 0 25576 800 25696 6 mgmt_rdata_ro[19]
port 611 nsew
rlabel metal2 s 25962 0 26018 800 6 mgmt_rdata_ro[1]
port 612 nsew
rlabel metal3 s 0 26120 800 26240 6 mgmt_rdata_ro[20]
port 613 nsew
rlabel metal2 s 26330 0 26386 800 6 mgmt_rdata_ro[21]
port 614 nsew
rlabel metal3 s 0 26664 800 26784 6 mgmt_rdata_ro[22]
port 615 nsew
rlabel metal2 s 26698 0 26754 800 6 mgmt_rdata_ro[23]
port 616 nsew
rlabel metal2 s 27066 0 27122 800 6 mgmt_rdata_ro[24]
port 617 nsew
rlabel metal3 s 0 27208 800 27328 6 mgmt_rdata_ro[25]
port 618 nsew
rlabel metal2 s 27434 0 27490 800 6 mgmt_rdata_ro[26]
port 619 nsew
rlabel metal3 s 0 27752 800 27872 6 mgmt_rdata_ro[27]
port 620 nsew
rlabel metal2 s 27802 0 27858 800 6 mgmt_rdata_ro[28]
port 621 nsew
rlabel metal2 s 28170 0 28226 800 6 mgmt_rdata_ro[29]
port 622 nsew
rlabel metal3 s 0 28296 800 28416 6 mgmt_rdata_ro[2]
port 623 nsew
rlabel metal2 s 28538 0 28594 800 6 mgmt_rdata_ro[30]
port 624 nsew
rlabel metal3 s 0 28840 800 28960 6 mgmt_rdata_ro[31]
port 625 nsew
rlabel metal2 s 28906 0 28962 800 6 mgmt_rdata_ro[3]
port 626 nsew
rlabel metal2 s 29274 0 29330 800 6 mgmt_rdata_ro[4]
port 627 nsew
rlabel metal3 s 0 29384 800 29504 6 mgmt_rdata_ro[5]
port 628 nsew
rlabel metal2 s 29642 0 29698 800 6 mgmt_rdata_ro[6]
port 629 nsew
rlabel metal3 s 0 29928 800 30048 6 mgmt_rdata_ro[7]
port 630 nsew
rlabel metal2 s 30010 0 30066 800 6 mgmt_rdata_ro[8]
port 631 nsew
rlabel metal2 s 30378 0 30434 800 6 mgmt_rdata_ro[9]
port 632 nsew
rlabel metal3 s 0 30472 800 30592 6 mgmt_wdata[0]
port 633 nsew
rlabel metal2 s 30746 0 30802 800 6 mgmt_wdata[10]
port 634 nsew
rlabel metal3 s 0 31016 800 31136 6 mgmt_wdata[11]
port 635 nsew
rlabel metal2 s 31114 0 31170 800 6 mgmt_wdata[12]
port 636 nsew
rlabel metal2 s 31482 0 31538 800 6 mgmt_wdata[13]
port 637 nsew
rlabel metal3 s 0 31560 800 31680 6 mgmt_wdata[14]
port 638 nsew
rlabel metal2 s 31850 0 31906 800 6 mgmt_wdata[15]
port 639 nsew
rlabel metal3 s 0 32104 800 32224 6 mgmt_wdata[16]
port 640 nsew
rlabel metal2 s 32218 0 32274 800 6 mgmt_wdata[17]
port 641 nsew
rlabel metal2 s 32586 0 32642 800 6 mgmt_wdata[18]
port 642 nsew
rlabel metal3 s 0 32648 800 32768 6 mgmt_wdata[19]
port 643 nsew
rlabel metal2 s 32954 0 33010 800 6 mgmt_wdata[1]
port 644 nsew
rlabel metal3 s 0 33192 800 33312 6 mgmt_wdata[20]
port 645 nsew
rlabel metal2 s 33322 0 33378 800 6 mgmt_wdata[21]
port 646 nsew
rlabel metal2 s 33690 0 33746 800 6 mgmt_wdata[22]
port 647 nsew
rlabel metal3 s 0 33736 800 33856 6 mgmt_wdata[23]
port 648 nsew
rlabel metal2 s 34058 0 34114 800 6 mgmt_wdata[24]
port 649 nsew
rlabel metal3 s 0 34280 800 34400 6 mgmt_wdata[25]
port 650 nsew
rlabel metal2 s 34426 0 34482 800 6 mgmt_wdata[26]
port 651 nsew
rlabel metal2 s 34794 0 34850 800 6 mgmt_wdata[27]
port 652 nsew
rlabel metal3 s 0 34824 800 34944 6 mgmt_wdata[28]
port 653 nsew
rlabel metal2 s 35162 0 35218 800 6 mgmt_wdata[29]
port 654 nsew
rlabel metal3 s 0 35368 800 35488 6 mgmt_wdata[2]
port 655 nsew
rlabel metal2 s 35530 0 35586 800 6 mgmt_wdata[30]
port 656 nsew
rlabel metal2 s 35898 0 35954 800 6 mgmt_wdata[31]
port 657 nsew
rlabel metal3 s 0 35912 800 36032 6 mgmt_wdata[3]
port 658 nsew
rlabel metal2 s 36266 0 36322 800 6 mgmt_wdata[4]
port 659 nsew
rlabel metal3 s 0 36456 800 36576 6 mgmt_wdata[5]
port 660 nsew
rlabel metal2 s 36634 0 36690 800 6 mgmt_wdata[6]
port 661 nsew
rlabel metal2 s 37002 0 37058 800 6 mgmt_wdata[7]
port 662 nsew
rlabel metal3 s 0 37000 800 37120 6 mgmt_wdata[8]
port 663 nsew
rlabel metal2 s 37370 0 37426 800 6 mgmt_wdata[9]
port 664 nsew
rlabel metal3 s 0 37544 800 37664 6 mgmt_wen[0]
port 665 nsew
rlabel metal2 s 37738 0 37794 800 6 mgmt_wen[1]
port 666 nsew
rlabel metal2 s 38106 0 38162 800 6 mgmt_wen_mask[0]
port 667 nsew
rlabel metal3 s 0 38088 800 38208 6 mgmt_wen_mask[1]
port 668 nsew
rlabel metal2 s 38474 0 38530 800 6 mgmt_wen_mask[2]
port 669 nsew
rlabel metal3 s 0 38632 800 38752 6 mgmt_wen_mask[3]
port 670 nsew
rlabel metal2 s 38842 0 38898 800 6 mgmt_wen_mask[4]
port 671 nsew
rlabel metal3 s 0 39176 800 39296 6 mgmt_wen_mask[5]
port 672 nsew
rlabel metal2 s 39210 0 39266 800 6 mgmt_wen_mask[6]
port 673 nsew
rlabel metal2 s 39578 0 39634 800 6 mgmt_wen_mask[7]
port 674 nsew
rlabel metal2 s 154026 169200 154082 170000 6 mprj2_vcc_pwrgood
port 675 nsew
rlabel metal2 s 296810 169200 296866 170000 6 mprj2_vdd_pwrgood
port 676 nsew
rlabel metal2 s 4250 169200 4306 170000 6 mprj_ack_i
port 677 nsew
rlabel metal2 s 153658 169200 153714 170000 6 mprj_adr_o[0]
port 678 nsew
rlabel metal2 s 297178 169200 297234 170000 6 mprj_adr_o[10]
port 679 nsew
rlabel metal2 s 153290 169200 153346 170000 6 mprj_adr_o[11]
port 680 nsew
rlabel metal2 s 297546 169200 297602 170000 6 mprj_adr_o[12]
port 681 nsew
rlabel metal2 s 152922 169200 152978 170000 6 mprj_adr_o[13]
port 682 nsew
rlabel metal2 s 297914 169200 297970 170000 6 mprj_adr_o[14]
port 683 nsew
rlabel metal2 s 152554 169200 152610 170000 6 mprj_adr_o[15]
port 684 nsew
rlabel metal2 s 298282 169200 298338 170000 6 mprj_adr_o[16]
port 685 nsew
rlabel metal2 s 152186 169200 152242 170000 6 mprj_adr_o[17]
port 686 nsew
rlabel metal2 s 298650 169200 298706 170000 6 mprj_adr_o[18]
port 687 nsew
rlabel metal2 s 151818 169200 151874 170000 6 mprj_adr_o[19]
port 688 nsew
rlabel metal2 s 299018 169200 299074 170000 6 mprj_adr_o[1]
port 689 nsew
rlabel metal2 s 151450 169200 151506 170000 6 mprj_adr_o[20]
port 690 nsew
rlabel metal2 s 299386 169200 299442 170000 6 mprj_adr_o[21]
port 691 nsew
rlabel metal2 s 151082 169200 151138 170000 6 mprj_adr_o[22]
port 692 nsew
rlabel metal2 s 299754 169200 299810 170000 6 mprj_adr_o[23]
port 693 nsew
rlabel metal2 s 150714 169200 150770 170000 6 mprj_adr_o[24]
port 694 nsew
rlabel metal2 s 300122 169200 300178 170000 6 mprj_adr_o[25]
port 695 nsew
rlabel metal2 s 150346 169200 150402 170000 6 mprj_adr_o[26]
port 696 nsew
rlabel metal2 s 300490 169200 300546 170000 6 mprj_adr_o[27]
port 697 nsew
rlabel metal2 s 149978 169200 150034 170000 6 mprj_adr_o[28]
port 698 nsew
rlabel metal2 s 300858 169200 300914 170000 6 mprj_adr_o[29]
port 699 nsew
rlabel metal2 s 149610 169200 149666 170000 6 mprj_adr_o[2]
port 700 nsew
rlabel metal2 s 301226 169200 301282 170000 6 mprj_adr_o[30]
port 701 nsew
rlabel metal2 s 149242 169200 149298 170000 6 mprj_adr_o[31]
port 702 nsew
rlabel metal2 s 301594 169200 301650 170000 6 mprj_adr_o[3]
port 703 nsew
rlabel metal2 s 148874 169200 148930 170000 6 mprj_adr_o[4]
port 704 nsew
rlabel metal2 s 301962 169200 302018 170000 6 mprj_adr_o[5]
port 705 nsew
rlabel metal2 s 148506 169200 148562 170000 6 mprj_adr_o[6]
port 706 nsew
rlabel metal2 s 302330 169200 302386 170000 6 mprj_adr_o[7]
port 707 nsew
rlabel metal2 s 148138 169200 148194 170000 6 mprj_adr_o[8]
port 708 nsew
rlabel metal2 s 302698 169200 302754 170000 6 mprj_adr_o[9]
port 709 nsew
rlabel metal2 s 147770 169200 147826 170000 6 mprj_cyc_o
port 710 nsew
rlabel metal3 s 0 165384 800 165504 6 mprj_dat_i[0]
port 711 nsew
rlabel metal2 s 4618 169200 4674 170000 6 mprj_dat_i[10]
port 712 nsew
rlabel metal2 s 4986 169200 5042 170000 6 mprj_dat_i[11]
port 713 nsew
rlabel metal3 s 0 164840 800 164960 6 mprj_dat_i[12]
port 714 nsew
rlabel metal2 s 5354 169200 5410 170000 6 mprj_dat_i[13]
port 715 nsew
rlabel metal3 s 0 164296 800 164416 6 mprj_dat_i[14]
port 716 nsew
rlabel metal2 s 5722 169200 5778 170000 6 mprj_dat_i[15]
port 717 nsew
rlabel metal2 s 6090 169200 6146 170000 6 mprj_dat_i[16]
port 718 nsew
rlabel metal3 s 0 163752 800 163872 6 mprj_dat_i[17]
port 719 nsew
rlabel metal2 s 6458 169200 6514 170000 6 mprj_dat_i[18]
port 720 nsew
rlabel metal3 s 0 163208 800 163328 6 mprj_dat_i[19]
port 721 nsew
rlabel metal2 s 6826 169200 6882 170000 6 mprj_dat_i[1]
port 722 nsew
rlabel metal2 s 7194 169200 7250 170000 6 mprj_dat_i[20]
port 723 nsew
rlabel metal3 s 0 162664 800 162784 6 mprj_dat_i[21]
port 724 nsew
rlabel metal2 s 7562 169200 7618 170000 6 mprj_dat_i[22]
port 725 nsew
rlabel metal3 s 0 162120 800 162240 6 mprj_dat_i[23]
port 726 nsew
rlabel metal2 s 7930 169200 7986 170000 6 mprj_dat_i[24]
port 727 nsew
rlabel metal2 s 8298 169200 8354 170000 6 mprj_dat_i[25]
port 728 nsew
rlabel metal3 s 0 161576 800 161696 6 mprj_dat_i[26]
port 729 nsew
rlabel metal2 s 8666 169200 8722 170000 6 mprj_dat_i[27]
port 730 nsew
rlabel metal3 s 0 161032 800 161152 6 mprj_dat_i[28]
port 731 nsew
rlabel metal2 s 9034 169200 9090 170000 6 mprj_dat_i[29]
port 732 nsew
rlabel metal2 s 9402 169200 9458 170000 6 mprj_dat_i[2]
port 733 nsew
rlabel metal3 s 0 160488 800 160608 6 mprj_dat_i[30]
port 734 nsew
rlabel metal2 s 9770 169200 9826 170000 6 mprj_dat_i[31]
port 735 nsew
rlabel metal3 s 0 159944 800 160064 6 mprj_dat_i[3]
port 736 nsew
rlabel metal2 s 10138 169200 10194 170000 6 mprj_dat_i[4]
port 737 nsew
rlabel metal2 s 10506 169200 10562 170000 6 mprj_dat_i[5]
port 738 nsew
rlabel metal3 s 0 159400 800 159520 6 mprj_dat_i[6]
port 739 nsew
rlabel metal2 s 10874 169200 10930 170000 6 mprj_dat_i[7]
port 740 nsew
rlabel metal3 s 0 158856 800 158976 6 mprj_dat_i[8]
port 741 nsew
rlabel metal2 s 11242 169200 11298 170000 6 mprj_dat_i[9]
port 742 nsew
rlabel metal2 s 303066 169200 303122 170000 6 mprj_dat_o[0]
port 743 nsew
rlabel metal2 s 147402 169200 147458 170000 6 mprj_dat_o[10]
port 744 nsew
rlabel metal2 s 303434 169200 303490 170000 6 mprj_dat_o[11]
port 745 nsew
rlabel metal2 s 147034 169200 147090 170000 6 mprj_dat_o[12]
port 746 nsew
rlabel metal2 s 303802 169200 303858 170000 6 mprj_dat_o[13]
port 747 nsew
rlabel metal2 s 146666 169200 146722 170000 6 mprj_dat_o[14]
port 748 nsew
rlabel metal2 s 304170 169200 304226 170000 6 mprj_dat_o[15]
port 749 nsew
rlabel metal2 s 146298 169200 146354 170000 6 mprj_dat_o[16]
port 750 nsew
rlabel metal2 s 304538 169200 304594 170000 6 mprj_dat_o[17]
port 751 nsew
rlabel metal2 s 145930 169200 145986 170000 6 mprj_dat_o[18]
port 752 nsew
rlabel metal2 s 304906 169200 304962 170000 6 mprj_dat_o[19]
port 753 nsew
rlabel metal2 s 145562 169200 145618 170000 6 mprj_dat_o[1]
port 754 nsew
rlabel metal2 s 305274 169200 305330 170000 6 mprj_dat_o[20]
port 755 nsew
rlabel metal2 s 145194 169200 145250 170000 6 mprj_dat_o[21]
port 756 nsew
rlabel metal2 s 305642 169200 305698 170000 6 mprj_dat_o[22]
port 757 nsew
rlabel metal2 s 144826 169200 144882 170000 6 mprj_dat_o[23]
port 758 nsew
rlabel metal2 s 306010 169200 306066 170000 6 mprj_dat_o[24]
port 759 nsew
rlabel metal2 s 144458 169200 144514 170000 6 mprj_dat_o[25]
port 760 nsew
rlabel metal2 s 306378 169200 306434 170000 6 mprj_dat_o[26]
port 761 nsew
rlabel metal2 s 144090 169200 144146 170000 6 mprj_dat_o[27]
port 762 nsew
rlabel metal2 s 306746 169200 306802 170000 6 mprj_dat_o[28]
port 763 nsew
rlabel metal2 s 143722 169200 143778 170000 6 mprj_dat_o[29]
port 764 nsew
rlabel metal2 s 307114 169200 307170 170000 6 mprj_dat_o[2]
port 765 nsew
rlabel metal2 s 143354 169200 143410 170000 6 mprj_dat_o[30]
port 766 nsew
rlabel metal2 s 307482 169200 307538 170000 6 mprj_dat_o[31]
port 767 nsew
rlabel metal2 s 142986 169200 143042 170000 6 mprj_dat_o[3]
port 768 nsew
rlabel metal2 s 307850 169200 307906 170000 6 mprj_dat_o[4]
port 769 nsew
rlabel metal2 s 142618 169200 142674 170000 6 mprj_dat_o[5]
port 770 nsew
rlabel metal2 s 308218 169200 308274 170000 6 mprj_dat_o[6]
port 771 nsew
rlabel metal2 s 142250 169200 142306 170000 6 mprj_dat_o[7]
port 772 nsew
rlabel metal2 s 308586 169200 308642 170000 6 mprj_dat_o[8]
port 773 nsew
rlabel metal2 s 141882 169200 141938 170000 6 mprj_dat_o[9]
port 774 nsew
rlabel metal3 s 429200 89768 430000 89888 6 mprj_io_loader_clock
port 775 nsew
rlabel metal3 s 429200 66376 430000 66496 6 mprj_io_loader_data
port 776 nsew
rlabel metal3 s 429200 96296 430000 96416 6 mprj_io_loader_resetn
port 777 nsew
rlabel metal2 s 308954 169200 309010 170000 6 mprj_sel_o[0]
port 778 nsew
rlabel metal2 s 141514 169200 141570 170000 6 mprj_sel_o[1]
port 779 nsew
rlabel metal2 s 309322 169200 309378 170000 6 mprj_sel_o[2]
port 780 nsew
rlabel metal2 s 141146 169200 141202 170000 6 mprj_sel_o[3]
port 781 nsew
rlabel metal2 s 309690 169200 309746 170000 6 mprj_stb_o
port 782 nsew
rlabel metal2 s 140778 169200 140834 170000 6 mprj_vcc_pwrgood
port 783 nsew
rlabel metal2 s 310058 169200 310114 170000 6 mprj_vdd_pwrgood
port 784 nsew
rlabel metal2 s 140410 169200 140466 170000 6 mprj_we_o
port 785 nsew
rlabel metal3 s 429200 21768 430000 21888 6 porb
port 786 nsew
rlabel metal2 s 14738 0 14794 800 6 pwr_ctrl_out[0]
port 787 nsew
rlabel metal2 s 15106 0 15162 800 6 pwr_ctrl_out[1]
port 788 nsew
rlabel metal2 s 15474 0 15530 800 6 pwr_ctrl_out[2]
port 789 nsew
rlabel metal2 s 15842 0 15898 800 6 pwr_ctrl_out[3]
port 790 nsew
rlabel metal3 s 0 39720 800 39840 6 resetb
port 791 nsew
rlabel metal3 s 429200 112072 430000 112192 6 sdo_out
port 792 nsew
rlabel metal3 s 429200 113160 430000 113280 6 sdo_outenb
port 793 nsew
rlabel metal2 s 310426 169200 310482 170000 6 user_clk
port 794 nsew
rlabel metal1 s 1104 167504 428812 167600 6 VPWR
port 795 nsew power default
rlabel metal1 s 1104 166960 428812 167056 6 VGND
port 796 nsew ground default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 430000 170000
string LEFview TRUE
string GDS_FILE mgmt_core.gds
string GDS_END 169521478
string GDS_START 2812312
<< end >>

