magic
tech sky130A
magscale 1 2
timestamp 1604412002
<< locali >>
rect 18573 17239 18607 17341
<< viali >>
rect 23633 34137 23667 34171
rect 25749 34137 25783 34171
rect 23449 33933 23483 33967
rect 25565 33933 25599 33967
rect 23357 33593 23391 33627
rect 24277 33593 24311 33627
rect 28969 33593 29003 33627
rect 19953 33525 19987 33559
rect 22437 33525 22471 33559
rect 23253 33525 23287 33559
rect 24185 33525 24219 33559
rect 24875 33525 24909 33559
rect 25013 33525 25047 33559
rect 25657 33525 25691 33559
rect 28049 33525 28083 33559
rect 28877 33525 28911 33559
rect 20597 33457 20631 33491
rect 20873 33457 20907 33491
rect 22529 33457 22563 33491
rect 26301 33457 26335 33491
rect 26577 33457 26611 33491
rect 28141 33457 28175 33491
rect 21333 33389 21367 33423
rect 21425 33389 21459 33423
rect 27037 33389 27071 33423
rect 27129 33389 27163 33423
rect 30993 33185 31027 33219
rect 25749 33117 25783 33151
rect 19677 33049 19711 33083
rect 20367 33049 20401 33083
rect 20505 33049 20539 33083
rect 21333 33049 21367 33083
rect 21790 33049 21824 33083
rect 23265 33049 23299 33083
rect 23817 33049 23851 33083
rect 26393 33049 26427 33083
rect 27865 33049 27899 33083
rect 28601 33049 28635 33083
rect 29061 33049 29095 33083
rect 30809 33049 30843 33083
rect 19769 32981 19803 33015
rect 24369 32981 24403 33015
rect 25197 32981 25231 33015
rect 23081 32913 23115 32947
rect 24277 32913 24311 32947
rect 25657 32913 25691 32947
rect 27681 32913 27715 32947
rect 21149 32845 21183 32879
rect 28417 32845 28451 32879
rect 29153 32845 29187 32879
rect 19493 32573 19527 32607
rect 21333 32573 21367 32607
rect 25657 32573 25691 32607
rect 19585 32505 19619 32539
rect 23817 32505 23851 32539
rect 27129 32505 27163 32539
rect 27221 32505 27255 32539
rect 19033 32437 19067 32471
rect 20045 32437 20079 32471
rect 21517 32437 21551 32471
rect 22897 32437 22931 32471
rect 23725 32437 23759 32471
rect 24369 32437 24403 32471
rect 25841 32437 25875 32471
rect 26669 32437 26703 32471
rect 27957 32437 27991 32471
rect 28693 32437 28727 32471
rect 22989 32369 23023 32403
rect 28877 32369 28911 32403
rect 21977 32097 22011 32131
rect 19769 32029 19803 32063
rect 21885 32029 21919 32063
rect 24369 32029 24403 32063
rect 25749 32029 25783 32063
rect 26301 32029 26335 32063
rect 26485 32029 26519 32063
rect 27865 32029 27899 32063
rect 27957 32029 27991 32063
rect 28785 32029 28819 32063
rect 20229 31961 20263 31995
rect 20413 31961 20447 31995
rect 20597 31961 20631 31995
rect 22805 31961 22839 31995
rect 23541 31961 23575 31995
rect 23725 31961 23759 31995
rect 24553 31961 24587 31995
rect 25197 31961 25231 31995
rect 25657 31961 25691 31995
rect 27405 31961 27439 31995
rect 28601 31961 28635 31995
rect 22437 31553 22471 31587
rect 20505 31485 20539 31519
rect 20045 31417 20079 31451
rect 20597 31417 20631 31451
rect 23541 31417 23575 31451
rect 21242 31349 21276 31383
rect 22989 31349 23023 31383
rect 24185 31349 24219 31383
rect 28325 31349 28359 31383
rect 29061 31349 29095 31383
rect 21057 31281 21091 31315
rect 22345 31281 22379 31315
rect 23449 31281 23483 31315
rect 24001 31281 24035 31315
rect 24553 31281 24587 31315
rect 28509 31281 28543 31315
rect 30165 31281 30199 31315
rect 21333 31213 21367 31247
rect 28969 31213 29003 31247
rect 30257 31213 30291 31247
rect 23357 31009 23391 31043
rect 22713 30941 22747 30975
rect 23909 30941 23943 30975
rect 20137 30873 20171 30907
rect 20321 30873 20355 30907
rect 22069 30873 22103 30907
rect 24093 30873 24127 30907
rect 26945 30873 26979 30907
rect 28233 30873 28267 30907
rect 29705 30873 29739 30907
rect 31269 30873 31303 30907
rect 20689 30805 20723 30839
rect 21241 30805 21275 30839
rect 21333 30805 21367 30839
rect 22161 30805 22195 30839
rect 23081 30805 23115 30839
rect 24369 30805 24403 30839
rect 26117 30805 26151 30839
rect 26209 30805 26243 30839
rect 27037 30805 27071 30839
rect 30809 30805 30843 30839
rect 31361 30805 31395 30839
rect 22989 30737 23023 30771
rect 29521 30737 29555 30771
rect 22878 30669 22912 30703
rect 32649 30465 32683 30499
rect 31361 30397 31395 30431
rect 20873 30329 20907 30363
rect 26025 30329 26059 30363
rect 28509 30329 28543 30363
rect 29061 30329 29095 30363
rect 17745 30261 17779 30295
rect 19125 30261 19159 30295
rect 19217 30261 19251 30295
rect 25105 30261 25139 30295
rect 25933 30261 25967 30295
rect 26761 30261 26795 30295
rect 26853 30261 26887 30295
rect 29889 30261 29923 30295
rect 31361 30261 31395 30295
rect 32097 30261 32131 30295
rect 20137 30193 20171 30227
rect 20497 30193 20531 30227
rect 22345 30193 22379 30227
rect 22713 30193 22747 30227
rect 23081 30193 23115 30227
rect 28969 30193 29003 30227
rect 17929 30125 17963 30159
rect 20321 30125 20355 30159
rect 20413 30125 20447 30159
rect 22529 30125 22563 30159
rect 22621 30125 22655 30159
rect 24737 30125 24771 30159
rect 31913 30125 31947 30159
rect 32557 30125 32591 30159
rect 24553 29921 24587 29955
rect 25473 29921 25507 29955
rect 20413 29853 20447 29887
rect 20597 29853 20631 29887
rect 20965 29853 20999 29887
rect 21425 29853 21459 29887
rect 21977 29853 22011 29887
rect 22713 29853 22747 29887
rect 22805 29853 22839 29887
rect 23173 29853 23207 29887
rect 23909 29853 23943 29887
rect 26761 29853 26795 29887
rect 28509 29853 28543 29887
rect 29705 29853 29739 29887
rect 30993 29853 31027 29887
rect 32925 29853 32959 29887
rect 16181 29785 16215 29819
rect 16825 29785 16859 29819
rect 20505 29785 20539 29819
rect 21609 29785 21643 29819
rect 22621 29785 22655 29819
rect 24056 29785 24090 29819
rect 25197 29785 25231 29819
rect 25381 29785 25415 29819
rect 26209 29785 26243 29819
rect 26393 29785 26427 29819
rect 27405 29785 27439 29819
rect 27865 29785 27899 29819
rect 27957 29785 27991 29819
rect 29061 29785 29095 29819
rect 29981 29785 30015 29819
rect 31729 29785 31763 29819
rect 31821 29785 31855 29819
rect 17101 29717 17135 29751
rect 18849 29717 18883 29751
rect 20229 29717 20263 29751
rect 22437 29717 22471 29751
rect 24277 29717 24311 29751
rect 27313 29717 27347 29751
rect 30901 29717 30935 29751
rect 32373 29717 32407 29751
rect 24185 29649 24219 29683
rect 32833 29649 32867 29683
rect 16365 29581 16399 29615
rect 24553 29377 24587 29411
rect 28233 29377 28267 29411
rect 29429 29309 29463 29343
rect 21333 29241 21367 29275
rect 25841 29241 25875 29275
rect 17009 29173 17043 29207
rect 17101 29173 17135 29207
rect 17285 29173 17319 29207
rect 18573 29173 18607 29207
rect 20781 29173 20815 29207
rect 23265 29173 23299 29207
rect 24461 29173 24495 29207
rect 25289 29173 25323 29207
rect 25474 29173 25508 29207
rect 26485 29173 26519 29207
rect 26853 29173 26887 29207
rect 28141 29173 28175 29207
rect 28969 29173 29003 29207
rect 30533 29173 30567 29207
rect 31269 29173 31303 29207
rect 19217 29105 19251 29139
rect 20597 29105 20631 29139
rect 20965 29105 20999 29139
rect 22989 29105 23023 29139
rect 23357 29105 23391 29139
rect 23725 29105 23759 29139
rect 24277 29105 24311 29139
rect 26301 29105 26335 29139
rect 27957 29105 27991 29139
rect 29521 29105 29555 29139
rect 31453 29105 31487 29139
rect 20873 29037 20907 29071
rect 23173 29037 23207 29071
rect 23081 28833 23115 28867
rect 25473 28833 25507 28867
rect 29153 28833 29187 28867
rect 31637 28833 31671 28867
rect 20597 28765 20631 28799
rect 21425 28765 21459 28799
rect 22897 28765 22931 28799
rect 23265 28765 23299 28799
rect 24093 28765 24127 28799
rect 27129 28765 27163 28799
rect 14433 28697 14467 28731
rect 15353 28697 15387 28731
rect 17837 28697 17871 28731
rect 18021 28697 18055 28731
rect 20505 28697 20539 28731
rect 21241 28697 21275 28731
rect 21333 28697 21367 28731
rect 23173 28697 23207 28731
rect 24277 28697 24311 28731
rect 25197 28697 25231 28731
rect 25381 28697 25415 28731
rect 27865 28697 27899 28731
rect 27957 28697 27991 28731
rect 29337 28697 29371 28731
rect 31545 28697 31579 28731
rect 15629 28629 15663 28663
rect 17377 28629 17411 28663
rect 18297 28629 18331 28663
rect 21057 28629 21091 28663
rect 21793 28629 21827 28663
rect 23633 28629 23667 28663
rect 27037 28629 27071 28663
rect 14617 28493 14651 28527
rect 24369 28493 24403 28527
rect 21517 28289 21551 28323
rect 26577 28289 26611 28323
rect 13789 28153 13823 28187
rect 16733 28153 16767 28187
rect 25197 28153 25231 28187
rect 29521 28153 29555 28187
rect 13513 28085 13547 28119
rect 17193 28085 17227 28119
rect 17469 28085 17503 28119
rect 17653 28085 17687 28119
rect 17837 28085 17871 28119
rect 18205 28085 18239 28119
rect 18849 28085 18883 28119
rect 20045 28085 20079 28119
rect 20689 28085 20723 28119
rect 21425 28085 21459 28119
rect 22345 28085 22379 28119
rect 22457 28085 22491 28119
rect 23541 28085 23575 28119
rect 25289 28085 25323 28119
rect 25657 28085 25691 28119
rect 25749 28085 25783 28119
rect 26485 28085 26519 28119
rect 28601 28085 28635 28119
rect 29429 28085 29463 28119
rect 15537 28017 15571 28051
rect 19493 28017 19527 28051
rect 21241 28017 21275 28051
rect 22897 28017 22931 28051
rect 23357 28017 23391 28051
rect 24645 28017 24679 28051
rect 26301 28017 26335 28051
rect 28693 28017 28727 28051
rect 23633 27949 23667 27983
rect 20229 27745 20263 27779
rect 27037 27745 27071 27779
rect 14065 27677 14099 27711
rect 16825 27677 16859 27711
rect 20413 27677 20447 27711
rect 21793 27677 21827 27711
rect 21885 27677 21919 27711
rect 22253 27677 22287 27711
rect 22897 27677 22931 27711
rect 23081 27677 23115 27711
rect 24093 27677 24127 27711
rect 24645 27677 24679 27711
rect 26393 27677 26427 27711
rect 29245 27677 29279 27711
rect 14525 27609 14559 27643
rect 14709 27609 14743 27643
rect 14985 27609 15019 27643
rect 17285 27609 17319 27643
rect 17561 27609 17595 27643
rect 17653 27609 17687 27643
rect 18113 27609 18147 27643
rect 20321 27609 20355 27643
rect 21701 27609 21735 27643
rect 22989 27609 23023 27643
rect 24277 27609 24311 27643
rect 25381 27609 25415 27643
rect 25565 27609 25599 27643
rect 28233 27609 28267 27643
rect 28417 27609 28451 27643
rect 28601 27609 28635 27643
rect 29429 27609 29463 27643
rect 15353 27541 15387 27575
rect 15445 27541 15479 27575
rect 18205 27541 18239 27575
rect 20045 27541 20079 27575
rect 20781 27541 20815 27575
rect 21517 27541 21551 27575
rect 22713 27541 22747 27575
rect 23449 27541 23483 27575
rect 25933 27541 25967 27575
rect 26761 27541 26795 27575
rect 29797 27541 29831 27575
rect 26669 27473 26703 27507
rect 28049 27473 28083 27507
rect 26531 27405 26565 27439
rect 26025 27201 26059 27235
rect 26393 27201 26427 27235
rect 18389 27133 18423 27167
rect 14617 27065 14651 27099
rect 16825 27065 16859 27099
rect 17377 27065 17411 27099
rect 17837 27065 17871 27099
rect 23173 27065 23207 27099
rect 24093 27065 24127 27099
rect 26117 27065 26151 27099
rect 30349 27065 30383 27099
rect 31269 27065 31303 27099
rect 14525 26997 14559 27031
rect 14985 26997 15019 27031
rect 16089 26997 16123 27031
rect 16181 26997 16215 27031
rect 17653 26997 17687 27031
rect 18297 26997 18331 27031
rect 18849 26997 18883 27031
rect 20965 26997 20999 27031
rect 21333 26997 21367 27031
rect 22713 26997 22747 27031
rect 24001 26997 24035 27031
rect 24277 26997 24311 27031
rect 24737 26997 24771 27031
rect 25896 26997 25930 27031
rect 28233 26997 28267 27031
rect 29705 26997 29739 27031
rect 31177 26997 31211 27031
rect 20781 26929 20815 26963
rect 22437 26929 22471 26963
rect 22805 26929 22839 26963
rect 25749 26929 25783 26963
rect 29797 26929 29831 26963
rect 30441 26929 30475 26963
rect 22621 26861 22655 26895
rect 17377 26657 17411 26691
rect 22621 26657 22655 26691
rect 28785 26657 28819 26691
rect 14617 26589 14651 26623
rect 22345 26589 22379 26623
rect 22713 26589 22747 26623
rect 23541 26589 23575 26623
rect 26117 26589 26151 26623
rect 26853 26589 26887 26623
rect 28509 26589 28543 26623
rect 29981 26589 30015 26623
rect 15261 26521 15295 26555
rect 15629 26521 15663 26555
rect 17745 26521 17779 26555
rect 18113 26521 18147 26555
rect 19585 26521 19619 26555
rect 20229 26521 20263 26555
rect 20413 26521 20447 26555
rect 20781 26521 20815 26555
rect 22529 26521 22563 26555
rect 27313 26521 27347 26555
rect 28693 26521 28727 26555
rect 29521 26521 29555 26555
rect 30993 26521 31027 26555
rect 31453 26521 31487 26555
rect 15353 26453 15387 26487
rect 15537 26453 15571 26487
rect 17653 26453 17687 26487
rect 18021 26453 18055 26487
rect 23081 26453 23115 26487
rect 23688 26453 23722 26487
rect 23909 26453 23943 26487
rect 24277 26453 24311 26487
rect 26264 26453 26298 26487
rect 26485 26453 26519 26487
rect 27681 26453 27715 26487
rect 30073 26453 30107 26487
rect 31545 26453 31579 26487
rect 20965 26385 20999 26419
rect 27451 26385 27485 26419
rect 27589 26385 27623 26419
rect 23817 26317 23851 26351
rect 26393 26317 26427 26351
rect 27957 26317 27991 26351
rect 30809 26317 30843 26351
rect 14709 26113 14743 26147
rect 22621 26113 22655 26147
rect 22989 26113 23023 26147
rect 25841 26113 25875 26147
rect 27037 26113 27071 26147
rect 25703 26045 25737 26079
rect 30165 26045 30199 26079
rect 16181 25977 16215 26011
rect 17837 25977 17871 26011
rect 22713 25977 22747 26011
rect 24461 25977 24495 26011
rect 25933 25977 25967 26011
rect 30257 25977 30291 26011
rect 13789 25909 13823 25943
rect 14433 25909 14467 25943
rect 14617 25909 14651 25943
rect 15813 25909 15847 25943
rect 17193 25909 17227 25943
rect 17377 25909 17411 25943
rect 17561 25909 17595 25943
rect 18205 25909 18239 25943
rect 19677 25909 19711 25943
rect 19861 25909 19895 25943
rect 20229 25909 20263 25943
rect 20965 25909 20999 25943
rect 21517 25909 21551 25943
rect 21701 25909 21735 25943
rect 22492 25909 22526 25943
rect 24185 25909 24219 25943
rect 25565 25909 25599 25943
rect 26761 25909 26795 25943
rect 26945 25909 26979 25943
rect 28325 25909 28359 25943
rect 29705 25909 29739 25943
rect 30809 25909 30843 25943
rect 31269 25909 31303 25943
rect 31821 25909 31855 25943
rect 15629 25841 15663 25875
rect 16733 25841 16767 25875
rect 20505 25841 20539 25875
rect 22345 25841 22379 25875
rect 24001 25841 24035 25875
rect 26301 25841 26335 25875
rect 29061 25841 29095 25875
rect 29245 25841 29279 25875
rect 31361 25841 31395 25875
rect 13973 25773 14007 25807
rect 31913 25773 31947 25807
rect 22989 25569 23023 25603
rect 29889 25569 29923 25603
rect 32189 25569 32223 25603
rect 17101 25501 17135 25535
rect 20689 25501 20723 25535
rect 25565 25501 25599 25535
rect 26761 25501 26795 25535
rect 28325 25501 28359 25535
rect 29797 25501 29831 25535
rect 31545 25501 31579 25535
rect 17745 25433 17779 25467
rect 18113 25433 18147 25467
rect 18297 25433 18331 25467
rect 19861 25433 19895 25467
rect 20045 25433 20079 25467
rect 20413 25433 20447 25467
rect 21425 25433 21459 25467
rect 21609 25433 21643 25467
rect 21885 25433 21919 25467
rect 22345 25433 22379 25467
rect 22492 25433 22526 25467
rect 23541 25433 23575 25467
rect 23725 25433 23759 25467
rect 25712 25433 25746 25467
rect 26945 25433 26979 25467
rect 28233 25433 28267 25467
rect 29061 25433 29095 25467
rect 29153 25433 29187 25467
rect 30809 25433 30843 25467
rect 31729 25433 31763 25467
rect 32373 25433 32407 25467
rect 13973 25365 14007 25399
rect 15997 25365 16031 25399
rect 17561 25365 17595 25399
rect 22713 25365 22747 25399
rect 24093 25365 24127 25399
rect 25933 25365 25967 25399
rect 27313 25365 27347 25399
rect 26209 25297 26243 25331
rect 14230 25229 14264 25263
rect 22621 25229 22655 25263
rect 25841 25229 25875 25263
rect 23725 25025 23759 25059
rect 28233 25025 28267 25059
rect 30717 24957 30751 24991
rect 32741 24957 32775 24991
rect 14157 24889 14191 24923
rect 15445 24889 15479 24923
rect 20689 24889 20723 24923
rect 25657 24889 25691 24923
rect 14709 24821 14743 24855
rect 14801 24821 14835 24855
rect 15077 24821 15111 24855
rect 15537 24821 15571 24855
rect 16917 24821 16951 24855
rect 19217 24821 19251 24855
rect 19401 24821 19435 24855
rect 19585 24821 19619 24855
rect 19861 24821 19895 24855
rect 20114 24821 20148 24855
rect 21241 24821 21275 24855
rect 21425 24821 21459 24855
rect 22345 24821 22379 24855
rect 22437 24821 22471 24855
rect 23449 24821 23483 24855
rect 23541 24821 23575 24855
rect 25381 24821 25415 24855
rect 26393 24821 26427 24855
rect 28141 24821 28175 24855
rect 29429 24821 29463 24855
rect 30349 24821 30383 24855
rect 31453 24821 31487 24855
rect 32373 24821 32407 24855
rect 17469 24753 17503 24787
rect 21793 24753 21827 24787
rect 22897 24753 22931 24787
rect 25197 24753 25231 24787
rect 26209 24753 26243 24787
rect 26761 24753 26795 24787
rect 27957 24753 27991 24787
rect 12869 24413 12903 24447
rect 13421 24413 13455 24447
rect 16549 24413 16583 24447
rect 25933 24413 25967 24447
rect 27129 24413 27163 24447
rect 31453 24413 31487 24447
rect 31545 24413 31579 24447
rect 32281 24413 32315 24447
rect 13053 24345 13087 24379
rect 14433 24345 14467 24379
rect 14801 24345 14835 24379
rect 15169 24345 15203 24379
rect 17009 24345 17043 24379
rect 17285 24345 17319 24379
rect 17469 24345 17503 24379
rect 17837 24345 17871 24379
rect 18021 24345 18055 24379
rect 18481 24345 18515 24379
rect 18665 24345 18699 24379
rect 19033 24345 19067 24379
rect 19677 24345 19711 24379
rect 22529 24345 22563 24379
rect 22897 24345 22931 24379
rect 23541 24345 23575 24379
rect 24369 24345 24403 24379
rect 24553 24345 24587 24379
rect 25197 24345 25231 24379
rect 25289 24345 25323 24379
rect 25473 24345 25507 24379
rect 27037 24345 27071 24379
rect 27865 24345 27899 24379
rect 28601 24345 28635 24379
rect 28693 24345 28727 24379
rect 29429 24345 29463 24379
rect 30257 24345 30291 24379
rect 32097 24345 32131 24379
rect 19585 24277 19619 24311
rect 22437 24277 22471 24311
rect 22989 24277 23023 24311
rect 24093 24277 24127 24311
rect 27957 24277 27991 24311
rect 29521 24277 29555 24311
rect 30993 24277 31027 24311
rect 19861 24141 19895 24175
rect 21977 24141 22011 24175
rect 30073 24141 30107 24175
rect 30717 23869 30751 23903
rect 14709 23801 14743 23835
rect 20597 23801 20631 23835
rect 23081 23801 23115 23835
rect 28325 23801 28359 23835
rect 30809 23801 30843 23835
rect 31821 23801 31855 23835
rect 15261 23733 15295 23767
rect 15537 23733 15571 23767
rect 15721 23733 15755 23767
rect 18205 23733 18239 23767
rect 19033 23733 19067 23767
rect 19309 23733 19343 23767
rect 19493 23733 19527 23767
rect 19769 23733 19803 23767
rect 19962 23733 19996 23767
rect 21057 23733 21091 23767
rect 21517 23733 21551 23767
rect 22897 23733 22931 23767
rect 23909 23733 23943 23767
rect 24093 23733 24127 23767
rect 24645 23733 24679 23767
rect 25013 23733 25047 23767
rect 26485 23733 26519 23767
rect 28877 23733 28911 23767
rect 30257 23733 30291 23767
rect 31269 23733 31303 23767
rect 18021 23665 18055 23699
rect 18573 23665 18607 23699
rect 21793 23665 21827 23699
rect 26301 23665 26335 23699
rect 26853 23665 26887 23699
rect 28233 23665 28267 23699
rect 29613 23665 29647 23699
rect 29797 23665 29831 23699
rect 31729 23665 31763 23699
rect 23725 23597 23759 23631
rect 16917 23393 16951 23427
rect 21057 23393 21091 23427
rect 22161 23393 22195 23427
rect 28233 23393 28267 23427
rect 30993 23393 31027 23427
rect 18481 23325 18515 23359
rect 19033 23325 19067 23359
rect 20321 23325 20355 23359
rect 22069 23325 22103 23359
rect 22253 23325 22287 23359
rect 22621 23325 22655 23359
rect 23081 23325 23115 23359
rect 23817 23325 23851 23359
rect 14709 23257 14743 23291
rect 14801 23257 14835 23291
rect 15077 23257 15111 23291
rect 15353 23257 15387 23291
rect 17469 23257 17503 23291
rect 17837 23257 17871 23291
rect 17929 23257 17963 23291
rect 18665 23257 18699 23291
rect 19677 23257 19711 23291
rect 20781 23257 20815 23291
rect 20965 23257 20999 23291
rect 23228 23257 23262 23291
rect 25197 23257 25231 23291
rect 25381 23257 25415 23291
rect 27313 23257 27347 23291
rect 28049 23257 28083 23291
rect 29245 23257 29279 23291
rect 30901 23257 30935 23291
rect 14157 23189 14191 23223
rect 15537 23189 15571 23223
rect 17561 23189 17595 23223
rect 21885 23189 21919 23223
rect 23449 23189 23483 23223
rect 26485 23189 26519 23223
rect 26577 23189 26611 23223
rect 27405 23189 27439 23223
rect 23357 23121 23391 23155
rect 25473 23053 25507 23087
rect 29613 23053 29647 23087
rect 15905 22849 15939 22883
rect 19861 22849 19895 22883
rect 18481 22781 18515 22815
rect 23909 22781 23943 22815
rect 13145 22713 13179 22747
rect 13421 22713 13455 22747
rect 15169 22713 15203 22747
rect 16825 22713 16859 22747
rect 21057 22713 21091 22747
rect 21793 22713 21827 22747
rect 22345 22713 22379 22747
rect 24001 22713 24035 22747
rect 25013 22713 25047 22747
rect 25933 22713 25967 22747
rect 30441 22713 30475 22747
rect 15629 22645 15663 22679
rect 15813 22645 15847 22679
rect 17469 22645 17503 22679
rect 18389 22645 18423 22679
rect 18665 22645 18699 22679
rect 19585 22645 19619 22679
rect 19769 22645 19803 22679
rect 21241 22645 21275 22679
rect 22529 22645 22563 22679
rect 23081 22645 23115 22679
rect 23633 22645 23667 22679
rect 23780 22645 23814 22679
rect 25105 22645 25139 22679
rect 25841 22645 25875 22679
rect 26669 22645 26703 22679
rect 28877 22645 28911 22679
rect 30257 22645 30291 22679
rect 21425 22577 21459 22611
rect 22621 22577 22655 22611
rect 22713 22577 22747 22611
rect 24369 22577 24403 22611
rect 26485 22577 26519 22611
rect 18849 22509 18883 22543
rect 21333 22509 21367 22543
rect 26761 22509 26795 22543
rect 18481 22305 18515 22339
rect 20045 22305 20079 22339
rect 21517 22305 21551 22339
rect 23817 22305 23851 22339
rect 25473 22305 25507 22339
rect 15169 22237 15203 22271
rect 19953 22237 19987 22271
rect 20137 22237 20171 22271
rect 21609 22237 21643 22271
rect 24001 22237 24035 22271
rect 25197 22237 25231 22271
rect 28877 22237 28911 22271
rect 31361 22237 31395 22271
rect 14249 22169 14283 22203
rect 14709 22169 14743 22203
rect 15813 22169 15847 22203
rect 16181 22169 16215 22203
rect 17837 22169 17871 22203
rect 21241 22169 21275 22203
rect 21425 22169 21459 22203
rect 22437 22169 22471 22203
rect 23633 22169 23667 22203
rect 23909 22169 23943 22203
rect 25381 22169 25415 22203
rect 26301 22169 26335 22203
rect 27773 22169 27807 22203
rect 28693 22169 28727 22203
rect 29337 22169 29371 22203
rect 29981 22169 30015 22203
rect 30257 22169 30291 22203
rect 30809 22169 30843 22203
rect 31269 22169 31303 22203
rect 14341 22101 14375 22135
rect 15629 22101 15663 22135
rect 16089 22101 16123 22135
rect 18205 22101 18239 22135
rect 19769 22101 19803 22135
rect 20505 22101 20539 22135
rect 21977 22101 22011 22135
rect 22584 22101 22618 22135
rect 22805 22101 22839 22135
rect 24369 22101 24403 22135
rect 27865 22101 27899 22135
rect 18113 22033 18147 22067
rect 23081 22033 23115 22067
rect 18002 21965 18036 21999
rect 22713 21965 22747 21999
rect 14341 21761 14375 21795
rect 15905 21693 15939 21727
rect 22989 21693 23023 21727
rect 27129 21693 27163 21727
rect 20781 21625 20815 21659
rect 23633 21625 23667 21659
rect 24185 21625 24219 21659
rect 25105 21625 25139 21659
rect 30533 21625 30567 21659
rect 30625 21625 30659 21659
rect 14157 21557 14191 21591
rect 15261 21557 15295 21591
rect 15445 21557 15479 21591
rect 15905 21557 15939 21591
rect 17469 21557 17503 21591
rect 18297 21557 18331 21591
rect 18481 21557 18515 21591
rect 18849 21557 18883 21591
rect 20413 21557 20447 21591
rect 21241 21557 21275 21591
rect 21425 21557 21459 21591
rect 22897 21557 22931 21591
rect 23173 21557 23207 21591
rect 24277 21557 24311 21591
rect 25013 21557 25047 21591
rect 26669 21557 26703 21591
rect 28141 21557 28175 21591
rect 28785 21557 28819 21591
rect 29705 21557 29739 21591
rect 29889 21557 29923 21591
rect 30073 21557 30107 21591
rect 31177 21557 31211 21591
rect 31637 21557 31671 21591
rect 32005 21557 32039 21591
rect 32097 21557 32131 21591
rect 21793 21489 21827 21523
rect 27221 21489 27255 21523
rect 29245 21489 29279 21523
rect 17285 21421 17319 21455
rect 19125 21421 19159 21455
rect 27957 21421 27991 21455
rect 28601 21421 28635 21455
rect 18297 21217 18331 21251
rect 21149 21217 21183 21251
rect 22805 21217 22839 21251
rect 28785 21217 28819 21251
rect 17561 21149 17595 21183
rect 18021 21149 18055 21183
rect 18389 21149 18423 21183
rect 19585 21149 19619 21183
rect 22529 21149 22563 21183
rect 27497 21149 27531 21183
rect 28049 21149 28083 21183
rect 30165 21149 30199 21183
rect 15813 21081 15847 21115
rect 16181 21081 16215 21115
rect 16365 21081 16399 21115
rect 16917 21081 16951 21115
rect 18205 21081 18239 21115
rect 19769 21081 19803 21115
rect 21517 21081 21551 21115
rect 21885 21081 21919 21115
rect 22069 21081 22103 21115
rect 22713 21081 22747 21115
rect 23817 21081 23851 21115
rect 26577 21081 26611 21115
rect 27313 21081 27347 21115
rect 28693 21081 28727 21115
rect 29613 21081 29647 21115
rect 30073 21081 30107 21115
rect 15905 21013 15939 21047
rect 18757 21013 18791 21047
rect 21609 21013 21643 21047
rect 25197 21013 25231 21047
rect 25749 21013 25783 21047
rect 25657 20945 25691 20979
rect 15445 20877 15479 20911
rect 19861 20877 19895 20911
rect 24001 20877 24035 20911
rect 28141 20877 28175 20911
rect 22345 20673 22379 20707
rect 27313 20605 27347 20639
rect 29889 20605 29923 20639
rect 15721 20537 15755 20571
rect 17469 20537 17503 20571
rect 24829 20537 24863 20571
rect 26853 20537 26887 20571
rect 27405 20537 27439 20571
rect 14985 20469 15019 20503
rect 15169 20469 15203 20503
rect 15353 20469 15387 20503
rect 15813 20469 15847 20503
rect 16825 20469 16859 20503
rect 18021 20469 18055 20503
rect 21149 20469 21183 20503
rect 21793 20469 21827 20503
rect 22621 20469 22655 20503
rect 24001 20469 24035 20503
rect 24185 20469 24219 20503
rect 24461 20469 24495 20503
rect 24921 20469 24955 20503
rect 25473 20469 25507 20503
rect 26393 20469 26427 20503
rect 14433 20401 14467 20435
rect 18297 20401 18331 20435
rect 20045 20401 20079 20435
rect 22529 20401 22563 20435
rect 23081 20401 23115 20435
rect 23541 20401 23575 20435
rect 26117 20401 26151 20435
rect 29705 20401 29739 20435
rect 16733 20129 16767 20163
rect 24461 20129 24495 20163
rect 28509 20129 28543 20163
rect 14249 20061 14283 20095
rect 15997 20061 16031 20095
rect 26853 20061 26887 20095
rect 13973 19993 14007 20027
rect 16457 19993 16491 20027
rect 16641 19993 16675 20027
rect 18021 19993 18055 20027
rect 18573 19993 18607 20027
rect 21425 19993 21459 20027
rect 22161 19993 22195 20027
rect 23633 19993 23667 20027
rect 24645 19993 24679 20027
rect 25289 19993 25323 20027
rect 26393 19993 26427 20027
rect 27313 19993 27347 20027
rect 27497 19993 27531 20027
rect 29613 19993 29647 20027
rect 17837 19925 17871 19959
rect 21793 19925 21827 19959
rect 28141 19925 28175 19959
rect 18481 19857 18515 19891
rect 27681 19857 27715 19891
rect 28509 19857 28543 19891
rect 23265 19789 23299 19823
rect 29705 19789 29739 19823
rect 14525 19585 14559 19619
rect 17929 19585 17963 19619
rect 19125 19585 19159 19619
rect 20045 19585 20079 19619
rect 29245 19517 29279 19551
rect 15537 19449 15571 19483
rect 25013 19449 25047 19483
rect 26117 19449 26151 19483
rect 14341 19381 14375 19415
rect 15353 19381 15387 19415
rect 15905 19381 15939 19415
rect 18297 19381 18331 19415
rect 19033 19381 19067 19415
rect 19861 19381 19895 19415
rect 22345 19381 22379 19415
rect 22529 19381 22563 19415
rect 23081 19381 23115 19415
rect 23265 19381 23299 19415
rect 25565 19381 25599 19415
rect 27957 19381 27991 19415
rect 28877 19381 28911 19415
rect 30073 19381 30107 19415
rect 18849 19313 18883 19347
rect 24921 19313 24955 19347
rect 26025 19313 26059 19347
rect 29981 19313 30015 19347
rect 23541 19245 23575 19279
rect 28785 19041 28819 19075
rect 19033 18973 19067 19007
rect 26669 18973 26703 19007
rect 27405 18973 27439 19007
rect 29429 18973 29463 19007
rect 18297 18905 18331 18939
rect 18573 18905 18607 18939
rect 19953 18905 19987 18939
rect 22437 18905 22471 18939
rect 23081 18905 23115 18939
rect 23173 18905 23207 18939
rect 23909 18905 23943 18939
rect 24369 18905 24403 18939
rect 26761 18905 26795 18939
rect 28141 18905 28175 18939
rect 20229 18837 20263 18871
rect 21977 18837 22011 18871
rect 26209 18837 26243 18871
rect 27313 18837 27347 18871
rect 28233 18837 28267 18871
rect 18389 18769 18423 18803
rect 22529 18701 22563 18735
rect 24553 18701 24587 18735
rect 29521 18701 29555 18735
rect 20873 18497 20907 18531
rect 21793 18429 21827 18463
rect 28417 18429 28451 18463
rect 17745 18361 17779 18395
rect 19769 18361 19803 18395
rect 23357 18361 23391 18395
rect 25105 18361 25139 18395
rect 27957 18361 27991 18395
rect 28509 18361 28543 18395
rect 14433 18293 14467 18327
rect 15813 18293 15847 18327
rect 20781 18293 20815 18327
rect 21609 18293 21643 18327
rect 23081 18293 23115 18327
rect 26485 18293 26519 18327
rect 27221 18293 27255 18327
rect 27405 18293 27439 18327
rect 18021 18225 18055 18259
rect 20597 18225 20631 18259
rect 14617 18157 14651 18191
rect 15629 18157 15663 18191
rect 21149 17953 21183 17987
rect 28141 17953 28175 17987
rect 15997 17885 16031 17919
rect 26761 17885 26795 17919
rect 13973 17817 14007 17851
rect 16457 17817 16491 17851
rect 16641 17817 16675 17851
rect 17193 17817 17227 17851
rect 17377 17817 17411 17851
rect 18389 17817 18423 17851
rect 19861 17817 19895 17851
rect 20965 17817 20999 17851
rect 22529 17817 22563 17851
rect 23081 17817 23115 17851
rect 23265 17817 23299 17851
rect 24461 17817 24495 17851
rect 26669 17817 26703 17851
rect 27497 17817 27531 17851
rect 28325 17817 28359 17851
rect 14249 17749 14283 17783
rect 18297 17749 18331 17783
rect 19769 17749 19803 17783
rect 22345 17749 22379 17783
rect 27589 17749 27623 17783
rect 17561 17681 17595 17715
rect 23541 17613 23575 17647
rect 24645 17613 24679 17647
rect 19953 17409 19987 17443
rect 15905 17341 15939 17375
rect 18573 17341 18607 17375
rect 11949 17273 11983 17307
rect 17009 17273 17043 17307
rect 23541 17273 23575 17307
rect 23817 17273 23851 17307
rect 25565 17273 25599 17307
rect 12041 17205 12075 17239
rect 14985 17205 15019 17239
rect 15077 17205 15111 17239
rect 15537 17205 15571 17239
rect 15721 17205 15755 17239
rect 17193 17205 17227 17239
rect 17377 17205 17411 17239
rect 17745 17205 17779 17239
rect 17929 17205 17963 17239
rect 18573 17205 18607 17239
rect 18665 17205 18699 17239
rect 18757 17205 18791 17239
rect 19861 17205 19895 17239
rect 12501 17137 12535 17171
rect 19217 17137 19251 17171
rect 19677 17137 19711 17171
rect 19861 16865 19895 16899
rect 16733 16797 16767 16831
rect 18297 16797 18331 16831
rect 18849 16797 18883 16831
rect 12133 16729 12167 16763
rect 12409 16729 12443 16763
rect 15445 16729 15479 16763
rect 15629 16729 15663 16763
rect 16181 16729 16215 16763
rect 16365 16729 16399 16763
rect 18205 16729 18239 16763
rect 18389 16729 18423 16763
rect 19585 16729 19619 16763
rect 19769 16729 19803 16763
rect 21057 16729 21091 16763
rect 21149 16729 21183 16763
rect 22253 16729 22287 16763
rect 22805 16729 22839 16763
rect 22989 16729 23023 16763
rect 24277 16729 24311 16763
rect 12593 16661 12627 16695
rect 22161 16661 22195 16695
rect 21333 16525 21367 16559
rect 23265 16525 23299 16559
rect 24461 16525 24495 16559
rect 12869 16185 12903 16219
rect 15353 16185 15387 16219
rect 17745 16185 17779 16219
rect 18941 16185 18975 16219
rect 21333 16185 21367 16219
rect 21517 16185 21551 16219
rect 23265 16185 23299 16219
rect 23541 16185 23575 16219
rect 25289 16185 25323 16219
rect 12409 16117 12443 16151
rect 12685 16117 12719 16151
rect 15629 16117 15663 16151
rect 15813 16117 15847 16151
rect 17377 16117 17411 16151
rect 18205 16117 18239 16151
rect 19033 16117 19067 16151
rect 19953 16117 19987 16151
rect 21241 16117 21275 16151
rect 21609 16117 21643 16151
rect 11857 16049 11891 16083
rect 14801 16049 14835 16083
rect 17193 16049 17227 16083
rect 19125 15981 19159 16015
rect 20137 15981 20171 16015
rect 20689 15981 20723 16015
rect 19033 15709 19067 15743
rect 12225 15641 12259 15675
rect 12777 15641 12811 15675
rect 12961 15641 12995 15675
rect 14341 15641 14375 15675
rect 16825 15641 16859 15675
rect 17193 15641 17227 15675
rect 17561 15641 17595 15675
rect 18481 15641 18515 15675
rect 18573 15641 18607 15675
rect 22161 15641 22195 15675
rect 22529 15641 22563 15675
rect 14617 15573 14651 15607
rect 16365 15573 16399 15607
rect 18297 15573 18331 15607
rect 19585 15573 19619 15607
rect 21609 15573 21643 15607
rect 12777 15505 12811 15539
rect 19842 15437 19876 15471
rect 24001 15437 24035 15471
rect 15997 15233 16031 15267
rect 20689 15233 20723 15267
rect 13881 15165 13915 15199
rect 12041 15097 12075 15131
rect 14893 15097 14927 15131
rect 19401 15097 19435 15131
rect 22345 15097 22379 15131
rect 11949 15029 11983 15063
rect 12777 15029 12811 15063
rect 13053 15029 13087 15063
rect 13421 15029 13455 15063
rect 13697 15029 13731 15063
rect 14985 15029 15019 15063
rect 15537 15029 15571 15063
rect 15721 15029 15755 15063
rect 17377 15029 17411 15063
rect 17929 15029 17963 15063
rect 18849 15029 18883 15063
rect 19033 15029 19067 15063
rect 20321 15029 20355 15063
rect 22437 15029 22471 15063
rect 24093 15029 24127 15063
rect 24369 15029 24403 15063
rect 17469 14961 17503 14995
rect 18113 14893 18147 14927
rect 23909 14893 23943 14927
rect 15721 14689 15755 14723
rect 21425 14689 21459 14723
rect 13053 14621 13087 14655
rect 23173 14621 23207 14655
rect 25197 14621 25231 14655
rect 12501 14553 12535 14587
rect 12777 14553 12811 14587
rect 13973 14553 14007 14587
rect 14801 14553 14835 14587
rect 15537 14553 15571 14587
rect 16733 14553 16767 14587
rect 18757 14553 18791 14587
rect 21333 14553 21367 14587
rect 21885 14553 21919 14587
rect 22161 14553 22195 14587
rect 23817 14553 23851 14587
rect 23909 14553 23943 14587
rect 24185 14553 24219 14587
rect 24277 14553 24311 14587
rect 25381 14553 25415 14587
rect 12041 14485 12075 14519
rect 14893 14485 14927 14519
rect 17009 14485 17043 14519
rect 14801 14417 14835 14451
rect 25473 14349 25507 14383
rect 12041 14145 12075 14179
rect 13053 14145 13087 14179
rect 17193 14145 17227 14179
rect 12777 14009 12811 14043
rect 14525 14009 14559 14043
rect 17653 14009 17687 14043
rect 19493 14009 19527 14043
rect 20045 14009 20079 14043
rect 20781 14009 20815 14043
rect 23725 14009 23759 14043
rect 11673 13941 11707 13975
rect 12869 13941 12903 13975
rect 14157 13941 14191 13975
rect 17745 13941 17779 13975
rect 18113 13941 18147 13975
rect 18297 13941 18331 13975
rect 18941 13941 18975 13975
rect 20689 13941 20723 13975
rect 21057 13941 21091 13975
rect 21149 13941 21183 13975
rect 23633 13941 23667 13975
rect 24461 13941 24495 13975
rect 24553 13941 24587 13975
rect 25565 13941 25599 13975
rect 26025 13941 26059 13975
rect 13973 13873 14007 13907
rect 18757 13873 18791 13907
rect 19125 13873 19159 13907
rect 19033 13805 19067 13839
rect 13421 13533 13455 13567
rect 15261 13533 15295 13567
rect 23265 13533 23299 13567
rect 27221 13533 27255 13567
rect 12961 13465 12995 13499
rect 14142 13465 14176 13499
rect 14617 13465 14651 13499
rect 14709 13465 14743 13499
rect 17561 13465 17595 13499
rect 17837 13465 17871 13499
rect 18573 13465 18607 13499
rect 19769 13465 19803 13499
rect 20873 13465 20907 13499
rect 20965 13465 20999 13499
rect 21425 13465 21459 13499
rect 21609 13465 21643 13499
rect 23817 13465 23851 13499
rect 24093 13465 24127 13499
rect 12869 13397 12903 13431
rect 13973 13397 14007 13431
rect 17009 13397 17043 13431
rect 18021 13397 18055 13431
rect 18481 13397 18515 13431
rect 19033 13397 19067 13431
rect 19677 13397 19711 13431
rect 20229 13397 20263 13431
rect 21977 13397 22011 13431
rect 24277 13397 24311 13431
rect 25197 13397 25231 13431
rect 25473 13397 25507 13431
rect 15353 13057 15387 13091
rect 25197 13057 25231 13091
rect 13513 12989 13547 13023
rect 18849 12989 18883 13023
rect 22621 12989 22655 13023
rect 12685 12921 12719 12955
rect 14249 12921 14283 12955
rect 18113 12921 18147 12955
rect 13145 12853 13179 12887
rect 13421 12853 13455 12887
rect 14341 12853 14375 12887
rect 14893 12853 14927 12887
rect 15077 12853 15111 12887
rect 18481 12853 18515 12887
rect 18757 12853 18791 12887
rect 20597 12853 20631 12887
rect 20689 12853 20723 12887
rect 21057 12853 21091 12887
rect 21149 12853 21183 12887
rect 22805 12853 22839 12887
rect 23173 12853 23207 12887
rect 23265 12853 23299 12887
rect 25013 12853 25047 12887
rect 25841 12853 25875 12887
rect 21701 12785 21735 12819
rect 25841 12717 25875 12751
rect 12501 12513 12535 12547
rect 16641 12445 16675 12479
rect 21701 12445 21735 12479
rect 23449 12445 23483 12479
rect 12869 12377 12903 12411
rect 13237 12377 13271 12411
rect 14525 12377 14559 12411
rect 14709 12377 14743 12411
rect 15261 12377 15295 12411
rect 15445 12377 15479 12411
rect 19585 12377 19619 12411
rect 20137 12377 20171 12411
rect 21425 12377 21459 12411
rect 25841 12377 25875 12411
rect 12961 12309 12995 12343
rect 13145 12309 13179 12343
rect 16365 12309 16399 12343
rect 18389 12309 18423 12343
rect 20413 12309 20447 12343
rect 19677 12241 19711 12275
rect 15721 12173 15755 12207
rect 25289 12173 25323 12207
rect 17653 11969 17687 12003
rect 21149 11969 21183 12003
rect 14433 11833 14467 11867
rect 16181 11833 16215 11867
rect 18389 11833 18423 11867
rect 18665 11833 18699 11867
rect 26853 11833 26887 11867
rect 14157 11765 14191 11799
rect 17837 11765 17871 11799
rect 20413 11765 20447 11799
rect 21517 11765 21551 11799
rect 22345 11765 22379 11799
rect 24829 11765 24863 11799
rect 22621 11697 22655 11731
rect 24369 11697 24403 11731
rect 25105 11697 25139 11731
rect 14985 11425 15019 11459
rect 16089 11425 16123 11459
rect 17469 11425 17503 11459
rect 19861 11425 19895 11459
rect 21333 11425 21367 11459
rect 23173 11425 23207 11459
rect 24737 11425 24771 11459
rect 25381 11357 25415 11391
rect 14801 11289 14835 11323
rect 15905 11289 15939 11323
rect 17285 11289 17319 11323
rect 19677 11289 19711 11323
rect 20965 11289 20999 11323
rect 22989 11289 23023 11323
rect 24553 11289 24587 11323
rect 26025 11289 26059 11323
<< metal1 >>
rect 11000 34418 34368 34440
rect 11000 34366 19142 34418
rect 19194 34366 19206 34418
rect 19258 34366 19270 34418
rect 19322 34366 19334 34418
rect 19386 34366 29142 34418
rect 29194 34366 29206 34418
rect 29258 34366 29270 34418
rect 29322 34366 29334 34418
rect 29386 34366 34368 34418
rect 11000 34344 34368 34366
rect 23618 34168 23624 34180
rect 23579 34140 23624 34168
rect 23618 34128 23624 34140
rect 23676 34128 23682 34180
rect 25737 34171 25795 34177
rect 25737 34137 25749 34171
rect 25783 34168 25795 34171
rect 26378 34168 26384 34180
rect 25783 34140 26384 34168
rect 25783 34137 25795 34140
rect 25737 34131 25795 34137
rect 26378 34128 26384 34140
rect 26436 34128 26442 34180
rect 23434 33964 23440 33976
rect 23395 33936 23440 33964
rect 23434 33924 23440 33936
rect 23492 33924 23498 33976
rect 25550 33964 25556 33976
rect 25511 33936 25556 33964
rect 25550 33924 25556 33936
rect 25608 33924 25614 33976
rect 11000 33874 34368 33896
rect 11000 33822 14142 33874
rect 14194 33822 14206 33874
rect 14258 33822 14270 33874
rect 14322 33822 14334 33874
rect 14386 33822 24142 33874
rect 24194 33822 24206 33874
rect 24258 33822 24270 33874
rect 24322 33822 24334 33874
rect 24386 33822 34368 33874
rect 11000 33800 34368 33822
rect 19864 33664 21732 33692
rect 19864 33488 19892 33664
rect 20122 33584 20128 33636
rect 20180 33624 20186 33636
rect 21704 33624 21732 33664
rect 23345 33627 23403 33633
rect 23345 33624 23357 33627
rect 20180 33596 21640 33624
rect 21704 33596 23357 33624
rect 20180 33584 20186 33596
rect 19941 33559 19999 33565
rect 19941 33525 19953 33559
rect 19987 33556 19999 33559
rect 20030 33556 20036 33568
rect 19987 33528 20036 33556
rect 19987 33525 19999 33528
rect 19941 33519 19999 33525
rect 20030 33516 20036 33528
rect 20088 33516 20094 33568
rect 15356 33460 19892 33488
rect 11014 33380 11020 33432
rect 11072 33420 11078 33432
rect 15356 33420 15384 33460
rect 20490 33448 20496 33500
rect 20548 33488 20554 33500
rect 20585 33491 20643 33497
rect 20585 33488 20597 33491
rect 20548 33460 20597 33488
rect 20548 33448 20554 33460
rect 20585 33457 20597 33460
rect 20631 33457 20643 33491
rect 20585 33451 20643 33457
rect 20861 33491 20919 33497
rect 20861 33457 20873 33491
rect 20907 33488 20919 33491
rect 21502 33488 21508 33500
rect 20907 33460 21508 33488
rect 20907 33457 20919 33460
rect 20861 33451 20919 33457
rect 11072 33392 15384 33420
rect 11072 33380 11078 33392
rect 15430 33380 15436 33432
rect 15488 33420 15494 33432
rect 16534 33420 16540 33432
rect 15488 33392 16540 33420
rect 15488 33380 15494 33392
rect 16534 33380 16540 33392
rect 16592 33380 16598 33432
rect 20600 33420 20628 33451
rect 21502 33448 21508 33460
rect 21560 33448 21566 33500
rect 21321 33423 21379 33429
rect 21321 33420 21333 33423
rect 20600 33392 21333 33420
rect 21321 33389 21333 33392
rect 21367 33389 21379 33423
rect 21321 33383 21379 33389
rect 21410 33380 21416 33432
rect 21468 33420 21474 33432
rect 21612 33420 21640 33596
rect 23345 33593 23357 33596
rect 23391 33593 23403 33627
rect 23345 33587 23403 33593
rect 24265 33627 24323 33633
rect 24265 33593 24277 33627
rect 24311 33624 24323 33627
rect 25090 33624 25096 33636
rect 24311 33596 25096 33624
rect 24311 33593 24323 33596
rect 24265 33587 24323 33593
rect 25090 33584 25096 33596
rect 25148 33624 25154 33636
rect 28957 33627 29015 33633
rect 25148 33596 25688 33624
rect 25148 33584 25154 33596
rect 22422 33556 22428 33568
rect 22383 33528 22428 33556
rect 22422 33516 22428 33528
rect 22480 33516 22486 33568
rect 23241 33559 23299 33565
rect 23241 33525 23253 33559
rect 23287 33556 23299 33559
rect 23526 33556 23532 33568
rect 23287 33528 23532 33556
rect 23287 33525 23299 33528
rect 23241 33519 23299 33525
rect 23526 33516 23532 33528
rect 23584 33516 23590 33568
rect 24170 33556 24176 33568
rect 24131 33528 24176 33556
rect 24170 33516 24176 33528
rect 24228 33516 24234 33568
rect 24863 33559 24921 33565
rect 24863 33556 24875 33559
rect 24464 33528 24875 33556
rect 22514 33488 22520 33500
rect 22475 33460 22520 33488
rect 22514 33448 22520 33460
rect 22572 33448 22578 33500
rect 24464 33420 24492 33528
rect 24863 33525 24875 33528
rect 24909 33525 24921 33559
rect 24863 33519 24921 33525
rect 24998 33516 25004 33568
rect 25056 33556 25062 33568
rect 25660 33565 25688 33596
rect 25752 33596 28816 33624
rect 25645 33559 25703 33565
rect 25056 33528 25504 33556
rect 25056 33516 25062 33528
rect 25476 33488 25504 33528
rect 25645 33525 25657 33559
rect 25691 33525 25703 33559
rect 25645 33519 25703 33525
rect 25752 33488 25780 33596
rect 28788 33568 28816 33596
rect 28957 33593 28969 33627
rect 29003 33624 29015 33627
rect 33646 33624 33652 33636
rect 29003 33596 33652 33624
rect 29003 33593 29015 33596
rect 28957 33587 29015 33593
rect 33646 33584 33652 33596
rect 33704 33584 33710 33636
rect 28034 33556 28040 33568
rect 27995 33528 28040 33556
rect 28034 33516 28040 33528
rect 28092 33516 28098 33568
rect 28770 33516 28776 33568
rect 28828 33556 28834 33568
rect 28865 33559 28923 33565
rect 28865 33556 28877 33559
rect 28828 33528 28877 33556
rect 28828 33516 28834 33528
rect 28865 33525 28877 33528
rect 28911 33525 28923 33559
rect 28865 33519 28923 33525
rect 25476 33460 25780 33488
rect 26194 33448 26200 33500
rect 26252 33488 26258 33500
rect 26289 33491 26347 33497
rect 26289 33488 26301 33491
rect 26252 33460 26301 33488
rect 26252 33448 26258 33460
rect 26289 33457 26301 33460
rect 26335 33457 26347 33491
rect 26289 33451 26347 33457
rect 21468 33392 21513 33420
rect 21612 33392 24492 33420
rect 26304 33420 26332 33451
rect 26470 33448 26476 33500
rect 26528 33488 26534 33500
rect 26565 33491 26623 33497
rect 26565 33488 26577 33491
rect 26528 33460 26577 33488
rect 26528 33448 26534 33460
rect 26565 33457 26577 33460
rect 26611 33457 26623 33491
rect 28126 33488 28132 33500
rect 28087 33460 28132 33488
rect 26565 33451 26623 33457
rect 28126 33448 28132 33460
rect 28184 33448 28190 33500
rect 27025 33423 27083 33429
rect 27025 33420 27037 33423
rect 26304 33392 27037 33420
rect 21468 33380 21474 33392
rect 27025 33389 27037 33392
rect 27071 33389 27083 33423
rect 27025 33383 27083 33389
rect 27114 33380 27120 33432
rect 27172 33420 27178 33432
rect 27172 33392 27217 33420
rect 27172 33380 27178 33392
rect 27390 33380 27396 33432
rect 27448 33420 27454 33432
rect 29506 33420 29512 33432
rect 27448 33392 29512 33420
rect 27448 33380 27454 33392
rect 29506 33380 29512 33392
rect 29564 33380 29570 33432
rect 11000 33330 34368 33352
rect 11000 33278 19142 33330
rect 19194 33278 19206 33330
rect 19258 33278 19270 33330
rect 19322 33278 19334 33330
rect 19386 33278 29142 33330
rect 29194 33278 29206 33330
rect 29258 33278 29270 33330
rect 29322 33278 29334 33330
rect 29386 33278 34368 33330
rect 11000 33256 34368 33278
rect 24446 33216 24452 33228
rect 19680 33188 24452 33216
rect 19680 33089 19708 33188
rect 24446 33176 24452 33188
rect 24504 33176 24510 33228
rect 30981 33219 31039 33225
rect 30981 33185 30993 33219
rect 31027 33216 31039 33219
rect 31438 33216 31444 33228
rect 31027 33188 31444 33216
rect 31027 33185 31039 33188
rect 30981 33179 31039 33185
rect 31438 33176 31444 33188
rect 31496 33176 31502 33228
rect 22514 33148 22520 33160
rect 21796 33120 22520 33148
rect 19665 33083 19723 33089
rect 19665 33049 19677 33083
rect 19711 33049 19723 33083
rect 20355 33083 20413 33089
rect 20355 33080 20367 33083
rect 19665 33043 19723 33049
rect 20140 33052 20367 33080
rect 19757 33015 19815 33021
rect 19757 32981 19769 33015
rect 19803 33012 19815 33015
rect 20030 33012 20036 33024
rect 19803 32984 20036 33012
rect 19803 32981 19815 32984
rect 19757 32975 19815 32981
rect 20030 32972 20036 32984
rect 20088 32972 20094 33024
rect 13958 32904 13964 32956
rect 14016 32944 14022 32956
rect 20140 32944 20168 33052
rect 20355 33049 20367 33052
rect 20401 33049 20413 33083
rect 20355 33043 20413 33049
rect 20493 33083 20551 33089
rect 20493 33049 20505 33083
rect 20539 33080 20551 33083
rect 20582 33080 20588 33092
rect 20539 33052 20588 33080
rect 20539 33049 20551 33052
rect 20493 33043 20551 33049
rect 20582 33040 20588 33052
rect 20640 33040 20646 33092
rect 21321 33083 21379 33089
rect 21321 33049 21333 33083
rect 21367 33080 21379 33083
rect 21502 33080 21508 33092
rect 21367 33052 21508 33080
rect 21367 33049 21379 33052
rect 21321 33043 21379 33049
rect 21502 33040 21508 33052
rect 21560 33040 21566 33092
rect 21796 33089 21824 33120
rect 22514 33108 22520 33120
rect 22572 33148 22578 33160
rect 25737 33151 25795 33157
rect 22572 33120 23848 33148
rect 22572 33108 22578 33120
rect 21778 33083 21836 33089
rect 21778 33049 21790 33083
rect 21824 33049 21836 33083
rect 21778 33043 21836 33049
rect 23253 33083 23311 33089
rect 23253 33049 23265 33083
rect 23299 33080 23311 33083
rect 23618 33080 23624 33092
rect 23299 33052 23624 33080
rect 23299 33049 23311 33052
rect 23253 33043 23311 33049
rect 23618 33040 23624 33052
rect 23676 33040 23682 33092
rect 23820 33089 23848 33120
rect 25737 33117 25749 33151
rect 25783 33148 25795 33151
rect 27114 33148 27120 33160
rect 25783 33120 27120 33148
rect 25783 33117 25795 33120
rect 25737 33111 25795 33117
rect 27114 33108 27120 33120
rect 27172 33108 27178 33160
rect 23805 33083 23863 33089
rect 23805 33049 23817 33083
rect 23851 33049 23863 33083
rect 23805 33043 23863 33049
rect 24170 33040 24176 33092
rect 24228 33080 24234 33092
rect 24906 33080 24912 33092
rect 24228 33052 24912 33080
rect 24228 33040 24234 33052
rect 24906 33040 24912 33052
rect 24964 33040 24970 33092
rect 26286 33040 26292 33092
rect 26344 33080 26350 33092
rect 26381 33083 26439 33089
rect 26381 33080 26393 33083
rect 26344 33052 26393 33080
rect 26344 33040 26350 33052
rect 26381 33049 26393 33052
rect 26427 33049 26439 33083
rect 26381 33043 26439 33049
rect 27853 33083 27911 33089
rect 27853 33049 27865 33083
rect 27899 33080 27911 33083
rect 28589 33083 28647 33089
rect 28589 33080 28601 33083
rect 27899 33052 28601 33080
rect 27899 33049 27911 33052
rect 27853 33043 27911 33049
rect 28589 33049 28601 33052
rect 28635 33080 28647 33083
rect 28862 33080 28868 33092
rect 28635 33052 28868 33080
rect 28635 33049 28647 33052
rect 28589 33043 28647 33049
rect 28862 33040 28868 33052
rect 28920 33040 28926 33092
rect 29046 33080 29052 33092
rect 29007 33052 29052 33080
rect 29046 33040 29052 33052
rect 29104 33040 29110 33092
rect 30610 33040 30616 33092
rect 30668 33080 30674 33092
rect 30797 33083 30855 33089
rect 30797 33080 30809 33083
rect 30668 33052 30809 33080
rect 30668 33040 30674 33052
rect 30797 33049 30809 33052
rect 30843 33049 30855 33083
rect 30797 33043 30855 33049
rect 23710 32972 23716 33024
rect 23768 33012 23774 33024
rect 24357 33015 24415 33021
rect 24357 33012 24369 33015
rect 23768 32984 24369 33012
rect 23768 32972 23774 32984
rect 24357 32981 24369 32984
rect 24403 32981 24415 33015
rect 25182 33012 25188 33024
rect 25143 32984 25188 33012
rect 24357 32975 24415 32981
rect 25182 32972 25188 32984
rect 25240 32972 25246 33024
rect 23066 32944 23072 32956
rect 14016 32916 20168 32944
rect 23027 32916 23072 32944
rect 14016 32904 14022 32916
rect 23066 32904 23072 32916
rect 23124 32944 23130 32956
rect 24265 32947 24323 32953
rect 24265 32944 24277 32947
rect 23124 32916 24277 32944
rect 23124 32904 23130 32916
rect 24265 32913 24277 32916
rect 24311 32913 24323 32947
rect 24265 32907 24323 32913
rect 25458 32904 25464 32956
rect 25516 32944 25522 32956
rect 25645 32947 25703 32953
rect 25645 32944 25657 32947
rect 25516 32916 25657 32944
rect 25516 32904 25522 32916
rect 25645 32913 25657 32916
rect 25691 32913 25703 32947
rect 25645 32907 25703 32913
rect 27114 32904 27120 32956
rect 27172 32944 27178 32956
rect 27669 32947 27727 32953
rect 27669 32944 27681 32947
rect 27172 32916 27681 32944
rect 27172 32904 27178 32916
rect 27669 32913 27681 32916
rect 27715 32913 27727 32947
rect 27669 32907 27727 32913
rect 21134 32876 21140 32888
rect 21095 32848 21140 32876
rect 21134 32836 21140 32848
rect 21192 32836 21198 32888
rect 28402 32876 28408 32888
rect 28363 32848 28408 32876
rect 28402 32836 28408 32848
rect 28460 32836 28466 32888
rect 29138 32876 29144 32888
rect 29099 32848 29144 32876
rect 29138 32836 29144 32848
rect 29196 32836 29202 32888
rect 11000 32786 34368 32808
rect 11000 32734 14142 32786
rect 14194 32734 14206 32786
rect 14258 32734 14270 32786
rect 14322 32734 14334 32786
rect 14386 32734 24142 32786
rect 24194 32734 24206 32786
rect 24258 32734 24270 32786
rect 24322 32734 24334 32786
rect 24386 32734 34368 32786
rect 11000 32712 34368 32734
rect 13222 32632 13228 32684
rect 13280 32672 13286 32684
rect 21686 32672 21692 32684
rect 13280 32644 21692 32672
rect 13280 32632 13286 32644
rect 21686 32632 21692 32644
rect 21744 32632 21750 32684
rect 19481 32607 19539 32613
rect 19481 32573 19493 32607
rect 19527 32604 19539 32607
rect 21318 32604 21324 32616
rect 19527 32576 21324 32604
rect 19527 32573 19539 32576
rect 19481 32567 19539 32573
rect 21318 32564 21324 32576
rect 21376 32564 21382 32616
rect 22238 32564 22244 32616
rect 22296 32604 22302 32616
rect 23526 32604 23532 32616
rect 22296 32576 23532 32604
rect 22296 32564 22302 32576
rect 23526 32564 23532 32576
rect 23584 32604 23590 32616
rect 24998 32604 25004 32616
rect 23584 32576 25004 32604
rect 23584 32564 23590 32576
rect 19573 32539 19631 32545
rect 19573 32505 19585 32539
rect 19619 32536 19631 32539
rect 21410 32536 21416 32548
rect 19619 32508 21416 32536
rect 19619 32505 19631 32508
rect 19573 32499 19631 32505
rect 21410 32496 21416 32508
rect 21468 32496 21474 32548
rect 19021 32471 19079 32477
rect 19021 32437 19033 32471
rect 19067 32468 19079 32471
rect 19754 32468 19760 32480
rect 19067 32440 19760 32468
rect 19067 32437 19079 32440
rect 19021 32431 19079 32437
rect 19754 32428 19760 32440
rect 19812 32468 19818 32480
rect 20033 32471 20091 32477
rect 20033 32468 20045 32471
rect 19812 32440 20045 32468
rect 19812 32428 19818 32440
rect 20033 32437 20045 32440
rect 20079 32437 20091 32471
rect 21502 32468 21508 32480
rect 21463 32440 21508 32468
rect 20033 32431 20091 32437
rect 21502 32428 21508 32440
rect 21560 32428 21566 32480
rect 22882 32468 22888 32480
rect 22843 32440 22888 32468
rect 22882 32428 22888 32440
rect 22940 32428 22946 32480
rect 23728 32477 23756 32576
rect 24998 32564 25004 32576
rect 25056 32564 25062 32616
rect 25458 32564 25464 32616
rect 25516 32604 25522 32616
rect 25645 32607 25703 32613
rect 25645 32604 25657 32607
rect 25516 32576 25657 32604
rect 25516 32564 25522 32576
rect 25645 32573 25657 32576
rect 25691 32573 25703 32607
rect 25645 32567 25703 32573
rect 23805 32539 23863 32545
rect 23805 32505 23817 32539
rect 23851 32536 23863 32539
rect 24630 32536 24636 32548
rect 23851 32508 24636 32536
rect 23851 32505 23863 32508
rect 23805 32499 23863 32505
rect 24630 32496 24636 32508
rect 24688 32496 24694 32548
rect 25918 32496 25924 32548
rect 25976 32536 25982 32548
rect 27114 32536 27120 32548
rect 25976 32508 27120 32536
rect 25976 32496 25982 32508
rect 27114 32496 27120 32508
rect 27172 32496 27178 32548
rect 27209 32539 27267 32545
rect 27209 32505 27221 32539
rect 27255 32536 27267 32539
rect 29138 32536 29144 32548
rect 27255 32508 29144 32536
rect 27255 32505 27267 32508
rect 27209 32499 27267 32505
rect 29138 32496 29144 32508
rect 29196 32496 29202 32548
rect 23713 32471 23771 32477
rect 23713 32437 23725 32471
rect 23759 32437 23771 32471
rect 23713 32431 23771 32437
rect 24357 32471 24415 32477
rect 24357 32437 24369 32471
rect 24403 32468 24415 32471
rect 25182 32468 25188 32480
rect 24403 32440 25188 32468
rect 24403 32437 24415 32440
rect 24357 32431 24415 32437
rect 22977 32403 23035 32409
rect 22977 32369 22989 32403
rect 23023 32400 23035 32403
rect 24372 32400 24400 32431
rect 25182 32428 25188 32440
rect 25240 32428 25246 32480
rect 25829 32471 25887 32477
rect 25829 32437 25841 32471
rect 25875 32437 25887 32471
rect 25829 32431 25887 32437
rect 23023 32372 24400 32400
rect 25844 32400 25872 32431
rect 26286 32428 26292 32480
rect 26344 32468 26350 32480
rect 26657 32471 26715 32477
rect 26657 32468 26669 32471
rect 26344 32440 26669 32468
rect 26344 32428 26350 32440
rect 26657 32437 26669 32440
rect 26703 32437 26715 32471
rect 26657 32431 26715 32437
rect 27945 32471 28003 32477
rect 27945 32437 27957 32471
rect 27991 32468 28003 32471
rect 28126 32468 28132 32480
rect 27991 32440 28132 32468
rect 27991 32437 28003 32440
rect 27945 32431 28003 32437
rect 28126 32428 28132 32440
rect 28184 32428 28190 32480
rect 28681 32471 28739 32477
rect 28681 32437 28693 32471
rect 28727 32468 28739 32471
rect 29046 32468 29052 32480
rect 28727 32440 29052 32468
rect 28727 32437 28739 32440
rect 28681 32431 28739 32437
rect 26470 32400 26476 32412
rect 25844 32372 26476 32400
rect 23023 32369 23035 32372
rect 22977 32363 23035 32369
rect 26470 32360 26476 32372
rect 26528 32360 26534 32412
rect 27850 32360 27856 32412
rect 27908 32400 27914 32412
rect 28696 32400 28724 32431
rect 29046 32428 29052 32440
rect 29104 32428 29110 32480
rect 28862 32400 28868 32412
rect 27908 32372 28724 32400
rect 28823 32372 28868 32400
rect 27908 32360 27914 32372
rect 28862 32360 28868 32372
rect 28920 32360 28926 32412
rect 11000 32242 34368 32264
rect 11000 32190 19142 32242
rect 19194 32190 19206 32242
rect 19258 32190 19270 32242
rect 19322 32190 19334 32242
rect 19386 32190 29142 32242
rect 29194 32190 29206 32242
rect 29258 32190 29270 32242
rect 29322 32190 29334 32242
rect 29386 32190 34368 32242
rect 11000 32168 34368 32190
rect 18190 32088 18196 32140
rect 18248 32128 18254 32140
rect 18248 32100 20352 32128
rect 18248 32088 18254 32100
rect 19754 32060 19760 32072
rect 19715 32032 19760 32060
rect 19754 32020 19760 32032
rect 19812 32020 19818 32072
rect 20217 31995 20275 32001
rect 20217 31961 20229 31995
rect 20263 31961 20275 31995
rect 20324 31992 20352 32100
rect 21502 32088 21508 32140
rect 21560 32128 21566 32140
rect 21965 32131 22023 32137
rect 21965 32128 21977 32131
rect 21560 32100 21977 32128
rect 21560 32088 21566 32100
rect 21965 32097 21977 32100
rect 22011 32097 22023 32131
rect 21965 32091 22023 32097
rect 21873 32063 21931 32069
rect 21873 32029 21885 32063
rect 21919 32060 21931 32063
rect 23066 32060 23072 32072
rect 21919 32032 23072 32060
rect 21919 32029 21931 32032
rect 21873 32023 21931 32029
rect 23066 32020 23072 32032
rect 23124 32020 23130 32072
rect 24357 32063 24415 32069
rect 24357 32029 24369 32063
rect 24403 32060 24415 32063
rect 25458 32060 25464 32072
rect 24403 32032 25464 32060
rect 24403 32029 24415 32032
rect 24357 32023 24415 32029
rect 25458 32020 25464 32032
rect 25516 32020 25522 32072
rect 25550 32020 25556 32072
rect 25608 32060 25614 32072
rect 25737 32063 25795 32069
rect 25737 32060 25749 32063
rect 25608 32032 25749 32060
rect 25608 32020 25614 32032
rect 25737 32029 25749 32032
rect 25783 32029 25795 32063
rect 25737 32023 25795 32029
rect 25918 32020 25924 32072
rect 25976 32060 25982 32072
rect 26289 32063 26347 32069
rect 26289 32060 26301 32063
rect 25976 32032 26301 32060
rect 25976 32020 25982 32032
rect 26289 32029 26301 32032
rect 26335 32029 26347 32063
rect 26470 32060 26476 32072
rect 26431 32032 26476 32060
rect 26289 32023 26347 32029
rect 26470 32020 26476 32032
rect 26528 32020 26534 32072
rect 27850 32060 27856 32072
rect 27811 32032 27856 32060
rect 27850 32020 27856 32032
rect 27908 32020 27914 32072
rect 27945 32063 28003 32069
rect 27945 32029 27957 32063
rect 27991 32060 28003 32063
rect 28402 32060 28408 32072
rect 27991 32032 28408 32060
rect 27991 32029 28003 32032
rect 27945 32023 28003 32029
rect 28402 32020 28408 32032
rect 28460 32020 28466 32072
rect 28773 32063 28831 32069
rect 28773 32029 28785 32063
rect 28819 32060 28831 32063
rect 28862 32060 28868 32072
rect 28819 32032 28868 32060
rect 28819 32029 28831 32032
rect 28773 32023 28831 32029
rect 28862 32020 28868 32032
rect 28920 32020 28926 32072
rect 20401 31995 20459 32001
rect 20401 31992 20413 31995
rect 20324 31964 20413 31992
rect 20217 31955 20275 31961
rect 20401 31961 20413 31964
rect 20447 31961 20459 31995
rect 20582 31992 20588 32004
rect 20495 31964 20588 31992
rect 20401 31955 20459 31961
rect 20232 31856 20260 31955
rect 20582 31952 20588 31964
rect 20640 31992 20646 32004
rect 22238 31992 22244 32004
rect 20640 31964 22244 31992
rect 20640 31952 20646 31964
rect 22238 31952 22244 31964
rect 22296 31952 22302 32004
rect 22793 31995 22851 32001
rect 22793 31961 22805 31995
rect 22839 31961 22851 31995
rect 23526 31992 23532 32004
rect 23487 31964 23532 31992
rect 22793 31955 22851 31961
rect 22808 31924 22836 31955
rect 23526 31952 23532 31964
rect 23584 31952 23590 32004
rect 23618 31952 23624 32004
rect 23676 31992 23682 32004
rect 23713 31995 23771 32001
rect 23713 31992 23725 31995
rect 23676 31964 23725 31992
rect 23676 31952 23682 31964
rect 23713 31961 23725 31964
rect 23759 31992 23771 31995
rect 24541 31995 24599 32001
rect 24541 31992 24553 31995
rect 23759 31964 24553 31992
rect 23759 31961 23771 31964
rect 23713 31955 23771 31961
rect 24541 31961 24553 31964
rect 24587 31961 24599 31995
rect 24541 31955 24599 31961
rect 25090 31952 25096 32004
rect 25148 31992 25154 32004
rect 25185 31995 25243 32001
rect 25185 31992 25197 31995
rect 25148 31964 25197 31992
rect 25148 31952 25154 31964
rect 25185 31961 25197 31964
rect 25231 31961 25243 31995
rect 25185 31955 25243 31961
rect 25645 31995 25703 32001
rect 25645 31961 25657 31995
rect 25691 31992 25703 31995
rect 26194 31992 26200 32004
rect 25691 31964 26200 31992
rect 25691 31961 25703 31964
rect 25645 31955 25703 31961
rect 26194 31952 26200 31964
rect 26252 31952 26258 32004
rect 27393 31995 27451 32001
rect 27393 31961 27405 31995
rect 27439 31992 27451 31995
rect 28126 31992 28132 32004
rect 27439 31964 28132 31992
rect 27439 31961 27451 31964
rect 27393 31955 27451 31961
rect 28126 31952 28132 31964
rect 28184 31952 28190 32004
rect 28586 31992 28592 32004
rect 28547 31964 28592 31992
rect 28586 31952 28592 31964
rect 28644 31952 28650 32004
rect 23802 31924 23808 31936
rect 22808 31896 23808 31924
rect 23802 31884 23808 31896
rect 23860 31884 23866 31936
rect 24722 31856 24728 31868
rect 20232 31828 24728 31856
rect 24722 31816 24728 31828
rect 24780 31816 24786 31868
rect 11000 31698 34368 31720
rect 11000 31646 14142 31698
rect 14194 31646 14206 31698
rect 14258 31646 14270 31698
rect 14322 31646 14334 31698
rect 14386 31646 24142 31698
rect 24194 31646 24206 31698
rect 24258 31646 24270 31698
rect 24322 31646 24334 31698
rect 24386 31646 34368 31698
rect 11000 31624 34368 31646
rect 22425 31587 22483 31593
rect 22425 31553 22437 31587
rect 22471 31584 22483 31587
rect 23710 31584 23716 31596
rect 22471 31556 23716 31584
rect 22471 31553 22483 31556
rect 22425 31547 22483 31553
rect 23710 31544 23716 31556
rect 23768 31544 23774 31596
rect 20490 31516 20496 31528
rect 20451 31488 20496 31516
rect 20490 31476 20496 31488
rect 20548 31476 20554 31528
rect 21318 31476 21324 31528
rect 21376 31516 21382 31528
rect 21376 31488 28356 31516
rect 21376 31476 21382 31488
rect 20030 31448 20036 31460
rect 19991 31420 20036 31448
rect 20030 31408 20036 31420
rect 20088 31408 20094 31460
rect 20585 31451 20643 31457
rect 20585 31417 20597 31451
rect 20631 31448 20643 31451
rect 21134 31448 21140 31460
rect 20631 31420 21140 31448
rect 20631 31417 20643 31420
rect 20585 31411 20643 31417
rect 21134 31408 21140 31420
rect 21192 31408 21198 31460
rect 23342 31448 23348 31460
rect 21244 31420 23348 31448
rect 21244 31389 21272 31420
rect 23342 31408 23348 31420
rect 23400 31408 23406 31460
rect 23434 31408 23440 31460
rect 23492 31448 23498 31460
rect 23529 31451 23587 31457
rect 23529 31448 23541 31451
rect 23492 31420 23541 31448
rect 23492 31408 23498 31420
rect 23529 31417 23541 31420
rect 23575 31417 23587 31451
rect 23529 31411 23587 31417
rect 21230 31383 21288 31389
rect 21230 31349 21242 31383
rect 21276 31349 21288 31383
rect 21230 31343 21288 31349
rect 22977 31383 23035 31389
rect 22977 31349 22989 31383
rect 23023 31380 23035 31383
rect 23802 31380 23808 31392
rect 23023 31352 23808 31380
rect 23023 31349 23035 31352
rect 22977 31343 23035 31349
rect 23802 31340 23808 31352
rect 23860 31340 23866 31392
rect 24173 31383 24231 31389
rect 24173 31349 24185 31383
rect 24219 31380 24231 31383
rect 25458 31380 25464 31392
rect 24219 31352 25464 31380
rect 24219 31349 24231 31352
rect 24173 31343 24231 31349
rect 25458 31340 25464 31352
rect 25516 31340 25522 31392
rect 28328 31389 28356 31488
rect 28313 31383 28371 31389
rect 28313 31349 28325 31383
rect 28359 31349 28371 31383
rect 28313 31343 28371 31349
rect 28954 31340 28960 31392
rect 29012 31380 29018 31392
rect 29049 31383 29107 31389
rect 29049 31380 29061 31383
rect 29012 31352 29061 31380
rect 29012 31340 29018 31352
rect 29049 31349 29061 31352
rect 29095 31349 29107 31383
rect 29049 31343 29107 31349
rect 20950 31272 20956 31324
rect 21008 31312 21014 31324
rect 21045 31315 21103 31321
rect 21045 31312 21057 31315
rect 21008 31284 21057 31312
rect 21008 31272 21014 31284
rect 21045 31281 21057 31284
rect 21091 31281 21103 31315
rect 21045 31275 21103 31281
rect 22333 31315 22391 31321
rect 22333 31281 22345 31315
rect 22379 31312 22391 31315
rect 23437 31315 23495 31321
rect 23437 31312 23449 31315
rect 22379 31284 23449 31312
rect 22379 31281 22391 31284
rect 22333 31275 22391 31281
rect 23437 31281 23449 31284
rect 23483 31312 23495 31315
rect 23526 31312 23532 31324
rect 23483 31284 23532 31312
rect 23483 31281 23495 31284
rect 23437 31275 23495 31281
rect 23526 31272 23532 31284
rect 23584 31272 23590 31324
rect 23989 31315 24047 31321
rect 23989 31281 24001 31315
rect 24035 31312 24047 31315
rect 24078 31312 24084 31324
rect 24035 31284 24084 31312
rect 24035 31281 24047 31284
rect 23989 31275 24047 31281
rect 24078 31272 24084 31284
rect 24136 31272 24142 31324
rect 24538 31312 24544 31324
rect 24499 31284 24544 31312
rect 24538 31272 24544 31284
rect 24596 31272 24602 31324
rect 28497 31315 28555 31321
rect 28497 31281 28509 31315
rect 28543 31312 28555 31315
rect 29782 31312 29788 31324
rect 28543 31284 29788 31312
rect 28543 31281 28555 31284
rect 28497 31275 28555 31281
rect 29782 31272 29788 31284
rect 29840 31272 29846 31324
rect 30153 31315 30211 31321
rect 30153 31281 30165 31315
rect 30199 31312 30211 31315
rect 31254 31312 31260 31324
rect 30199 31284 31260 31312
rect 30199 31281 30211 31284
rect 30153 31275 30211 31281
rect 31254 31272 31260 31284
rect 31312 31272 31318 31324
rect 21134 31204 21140 31256
rect 21192 31244 21198 31256
rect 21321 31247 21379 31253
rect 21321 31244 21333 31247
rect 21192 31216 21333 31244
rect 21192 31204 21198 31216
rect 21321 31213 21333 31216
rect 21367 31213 21379 31247
rect 21321 31207 21379 31213
rect 28957 31247 29015 31253
rect 28957 31213 28969 31247
rect 29003 31244 29015 31247
rect 29598 31244 29604 31256
rect 29003 31216 29604 31244
rect 29003 31213 29015 31216
rect 28957 31207 29015 31213
rect 29598 31204 29604 31216
rect 29656 31204 29662 31256
rect 29690 31204 29696 31256
rect 29748 31244 29754 31256
rect 30245 31247 30303 31253
rect 30245 31244 30257 31247
rect 29748 31216 30257 31244
rect 29748 31204 29754 31216
rect 30245 31213 30257 31216
rect 30291 31213 30303 31247
rect 30245 31207 30303 31213
rect 11000 31154 34368 31176
rect 11000 31102 19142 31154
rect 19194 31102 19206 31154
rect 19258 31102 19270 31154
rect 19322 31102 19334 31154
rect 19386 31102 29142 31154
rect 29194 31102 29206 31154
rect 29258 31102 29270 31154
rect 29322 31102 29334 31154
rect 29386 31102 34368 31154
rect 11000 31080 34368 31102
rect 22422 31000 22428 31052
rect 22480 31040 22486 31052
rect 23345 31043 23403 31049
rect 23345 31040 23357 31043
rect 22480 31012 23357 31040
rect 22480 31000 22486 31012
rect 23345 31009 23357 31012
rect 23391 31009 23403 31043
rect 23345 31003 23403 31009
rect 21134 30932 21140 30984
rect 21192 30972 21198 30984
rect 22701 30975 22759 30981
rect 22701 30972 22713 30975
rect 21192 30944 22713 30972
rect 21192 30932 21198 30944
rect 22701 30941 22713 30944
rect 22747 30941 22759 30975
rect 22882 30972 22888 30984
rect 22701 30935 22759 30941
rect 22808 30944 22888 30972
rect 20122 30904 20128 30916
rect 20083 30876 20128 30904
rect 20122 30864 20128 30876
rect 20180 30864 20186 30916
rect 20309 30907 20367 30913
rect 20309 30873 20321 30907
rect 20355 30873 20367 30907
rect 20309 30867 20367 30873
rect 22057 30907 22115 30913
rect 22057 30873 22069 30907
rect 22103 30904 22115 30907
rect 22238 30904 22244 30916
rect 22103 30876 22244 30904
rect 22103 30873 22115 30876
rect 22057 30867 22115 30873
rect 20324 30700 20352 30867
rect 22238 30864 22244 30876
rect 22296 30864 22302 30916
rect 22514 30864 22520 30916
rect 22572 30904 22578 30916
rect 22808 30904 22836 30944
rect 22882 30932 22888 30944
rect 22940 30972 22946 30984
rect 23897 30975 23955 30981
rect 23897 30972 23909 30975
rect 22940 30944 23909 30972
rect 22940 30932 22946 30944
rect 23897 30941 23909 30944
rect 23943 30941 23955 30975
rect 23897 30935 23955 30941
rect 22572 30876 22836 30904
rect 22572 30864 22578 30876
rect 23250 30864 23256 30916
rect 23308 30904 23314 30916
rect 24081 30907 24139 30913
rect 24081 30904 24093 30907
rect 23308 30876 24093 30904
rect 23308 30864 23314 30876
rect 24081 30873 24093 30876
rect 24127 30873 24139 30907
rect 24081 30867 24139 30873
rect 26746 30864 26752 30916
rect 26804 30904 26810 30916
rect 26933 30907 26991 30913
rect 26933 30904 26945 30907
rect 26804 30876 26945 30904
rect 26804 30864 26810 30876
rect 26933 30873 26945 30876
rect 26979 30873 26991 30907
rect 26933 30867 26991 30873
rect 28221 30907 28279 30913
rect 28221 30873 28233 30907
rect 28267 30904 28279 30907
rect 28494 30904 28500 30916
rect 28267 30876 28500 30904
rect 28267 30873 28279 30876
rect 28221 30867 28279 30873
rect 28494 30864 28500 30876
rect 28552 30864 28558 30916
rect 29690 30904 29696 30916
rect 29603 30876 29696 30904
rect 29690 30864 29696 30876
rect 29748 30904 29754 30916
rect 29966 30904 29972 30916
rect 29748 30876 29972 30904
rect 29748 30864 29754 30876
rect 29966 30864 29972 30876
rect 30024 30864 30030 30916
rect 31254 30904 31260 30916
rect 31215 30876 31260 30904
rect 31254 30864 31260 30876
rect 31312 30864 31318 30916
rect 20677 30839 20735 30845
rect 20677 30805 20689 30839
rect 20723 30805 20735 30839
rect 20677 30799 20735 30805
rect 20692 30768 20720 30799
rect 21134 30796 21140 30848
rect 21192 30836 21198 30848
rect 21229 30839 21287 30845
rect 21229 30836 21241 30839
rect 21192 30808 21241 30836
rect 21192 30796 21198 30808
rect 21229 30805 21241 30808
rect 21275 30805 21287 30839
rect 21229 30799 21287 30805
rect 21321 30839 21379 30845
rect 21321 30805 21333 30839
rect 21367 30836 21379 30839
rect 21594 30836 21600 30848
rect 21367 30808 21600 30836
rect 21367 30805 21379 30808
rect 21321 30799 21379 30805
rect 21594 30796 21600 30808
rect 21652 30796 21658 30848
rect 21686 30796 21692 30848
rect 21744 30836 21750 30848
rect 22149 30839 22207 30845
rect 22149 30836 22161 30839
rect 21744 30808 22161 30836
rect 21744 30796 21750 30808
rect 22149 30805 22161 30808
rect 22195 30805 22207 30839
rect 22149 30799 22207 30805
rect 22422 30796 22428 30848
rect 22480 30836 22486 30848
rect 23069 30839 23127 30845
rect 23069 30836 23081 30839
rect 22480 30808 23081 30836
rect 22480 30796 22486 30808
rect 23069 30805 23081 30808
rect 23115 30805 23127 30839
rect 23069 30799 23127 30805
rect 23342 30796 23348 30848
rect 23400 30836 23406 30848
rect 24357 30839 24415 30845
rect 24357 30836 24369 30839
rect 23400 30808 24369 30836
rect 23400 30796 23406 30808
rect 24357 30805 24369 30808
rect 24403 30836 24415 30839
rect 25366 30836 25372 30848
rect 24403 30808 25372 30836
rect 24403 30805 24415 30808
rect 24357 30799 24415 30805
rect 25366 30796 25372 30808
rect 25424 30836 25430 30848
rect 26105 30839 26163 30845
rect 26105 30836 26117 30839
rect 25424 30808 26117 30836
rect 25424 30796 25430 30808
rect 26105 30805 26117 30808
rect 26151 30805 26163 30839
rect 26105 30799 26163 30805
rect 26194 30796 26200 30848
rect 26252 30836 26258 30848
rect 26252 30808 26297 30836
rect 26252 30796 26258 30808
rect 26838 30796 26844 30848
rect 26896 30836 26902 30848
rect 27025 30839 27083 30845
rect 27025 30836 27037 30839
rect 26896 30808 27037 30836
rect 26896 30796 26902 30808
rect 27025 30805 27037 30808
rect 27071 30805 27083 30839
rect 30794 30836 30800 30848
rect 30755 30808 30800 30836
rect 27025 30799 27083 30805
rect 30794 30796 30800 30808
rect 30852 30796 30858 30848
rect 31349 30839 31407 30845
rect 31349 30805 31361 30839
rect 31395 30836 31407 30839
rect 32634 30836 32640 30848
rect 31395 30808 32640 30836
rect 31395 30805 31407 30808
rect 31349 30799 31407 30805
rect 32634 30796 32640 30808
rect 32692 30796 32698 30848
rect 22977 30771 23035 30777
rect 22977 30768 22989 30771
rect 20692 30740 22989 30768
rect 22977 30737 22989 30740
rect 23023 30737 23035 30771
rect 22977 30731 23035 30737
rect 24078 30728 24084 30780
rect 24136 30768 24142 30780
rect 26378 30768 26384 30780
rect 24136 30740 26384 30768
rect 24136 30728 24142 30740
rect 26378 30728 26384 30740
rect 26436 30728 26442 30780
rect 28586 30728 28592 30780
rect 28644 30768 28650 30780
rect 29046 30768 29052 30780
rect 28644 30740 29052 30768
rect 28644 30728 28650 30740
rect 29046 30728 29052 30740
rect 29104 30768 29110 30780
rect 29509 30771 29567 30777
rect 29509 30768 29521 30771
rect 29104 30740 29521 30768
rect 29104 30728 29110 30740
rect 29509 30737 29521 30740
rect 29555 30737 29567 30771
rect 29509 30731 29567 30737
rect 21226 30700 21232 30712
rect 20324 30672 21232 30700
rect 21226 30660 21232 30672
rect 21284 30660 21290 30712
rect 22866 30703 22924 30709
rect 22866 30669 22878 30703
rect 22912 30700 22924 30703
rect 23986 30700 23992 30712
rect 22912 30672 23992 30700
rect 22912 30669 22924 30672
rect 22866 30663 22924 30669
rect 23986 30660 23992 30672
rect 24044 30660 24050 30712
rect 11000 30610 34368 30632
rect 11000 30558 14142 30610
rect 14194 30558 14206 30610
rect 14258 30558 14270 30610
rect 14322 30558 14334 30610
rect 14386 30558 24142 30610
rect 24194 30558 24206 30610
rect 24258 30558 24270 30610
rect 24322 30558 24334 30610
rect 24386 30558 34368 30610
rect 11000 30536 34368 30558
rect 32634 30496 32640 30508
rect 32595 30468 32640 30496
rect 32634 30456 32640 30468
rect 32692 30456 32698 30508
rect 16810 30388 16816 30440
rect 16868 30428 16874 30440
rect 30610 30428 30616 30440
rect 16868 30400 30616 30428
rect 16868 30388 16874 30400
rect 30610 30388 30616 30400
rect 30668 30388 30674 30440
rect 31254 30388 31260 30440
rect 31312 30428 31318 30440
rect 31349 30431 31407 30437
rect 31349 30428 31361 30431
rect 31312 30400 31361 30428
rect 31312 30388 31318 30400
rect 31349 30397 31361 30400
rect 31395 30397 31407 30431
rect 31349 30391 31407 30397
rect 20122 30320 20128 30372
rect 20180 30360 20186 30372
rect 20861 30363 20919 30369
rect 20861 30360 20873 30363
rect 20180 30332 20873 30360
rect 20180 30320 20186 30332
rect 20861 30329 20873 30332
rect 20907 30329 20919 30363
rect 20861 30323 20919 30329
rect 26013 30363 26071 30369
rect 26013 30329 26025 30363
rect 26059 30360 26071 30363
rect 26286 30360 26292 30372
rect 26059 30332 26292 30360
rect 26059 30329 26071 30332
rect 26013 30323 26071 30329
rect 26286 30320 26292 30332
rect 26344 30320 26350 30372
rect 28494 30360 28500 30372
rect 28455 30332 28500 30360
rect 28494 30320 28500 30332
rect 28552 30320 28558 30372
rect 28954 30320 28960 30372
rect 29012 30360 29018 30372
rect 29049 30363 29107 30369
rect 29049 30360 29061 30363
rect 29012 30332 29061 30360
rect 29012 30320 29018 30332
rect 29049 30329 29061 30332
rect 29095 30329 29107 30363
rect 29049 30323 29107 30329
rect 16166 30252 16172 30304
rect 16224 30292 16230 30304
rect 17733 30295 17791 30301
rect 17733 30292 17745 30295
rect 16224 30264 17745 30292
rect 16224 30252 16230 30264
rect 17733 30261 17745 30264
rect 17779 30261 17791 30295
rect 17733 30255 17791 30261
rect 19113 30295 19171 30301
rect 19113 30261 19125 30295
rect 19159 30261 19171 30295
rect 19113 30255 19171 30261
rect 19205 30295 19263 30301
rect 19205 30261 19217 30295
rect 19251 30292 19263 30295
rect 20214 30292 20220 30304
rect 19251 30264 20220 30292
rect 19251 30261 19263 30264
rect 19205 30255 19263 30261
rect 17822 30116 17828 30168
rect 17880 30156 17886 30168
rect 17917 30159 17975 30165
rect 17917 30156 17929 30159
rect 17880 30128 17929 30156
rect 17880 30116 17886 30128
rect 17917 30125 17929 30128
rect 17963 30125 17975 30159
rect 17917 30119 17975 30125
rect 18466 30116 18472 30168
rect 18524 30156 18530 30168
rect 19128 30156 19156 30255
rect 20214 30252 20220 30264
rect 20272 30252 20278 30304
rect 20416 30264 20720 30292
rect 19938 30184 19944 30236
rect 19996 30224 20002 30236
rect 20125 30227 20183 30233
rect 20125 30224 20137 30227
rect 19996 30196 20137 30224
rect 19996 30184 20002 30196
rect 20125 30193 20137 30196
rect 20171 30224 20183 30227
rect 20416 30224 20444 30264
rect 20171 30196 20444 30224
rect 20485 30227 20543 30233
rect 20171 30193 20183 30196
rect 20125 30187 20183 30193
rect 20485 30193 20497 30227
rect 20531 30224 20543 30227
rect 20582 30224 20588 30236
rect 20531 30196 20588 30224
rect 20531 30193 20543 30196
rect 20485 30187 20543 30193
rect 20582 30184 20588 30196
rect 20640 30184 20646 30236
rect 20692 30224 20720 30264
rect 21594 30252 21600 30304
rect 21652 30292 21658 30304
rect 25090 30292 25096 30304
rect 21652 30264 24952 30292
rect 25051 30264 25096 30292
rect 21652 30252 21658 30264
rect 22330 30224 22336 30236
rect 20692 30196 22336 30224
rect 22330 30184 22336 30196
rect 22388 30224 22394 30236
rect 22701 30227 22759 30233
rect 22388 30196 22433 30224
rect 22388 30184 22394 30196
rect 22701 30193 22713 30227
rect 22747 30224 22759 30227
rect 23066 30224 23072 30236
rect 22747 30196 22928 30224
rect 23027 30196 23072 30224
rect 22747 30193 22759 30196
rect 22701 30187 22759 30193
rect 20309 30159 20367 30165
rect 20309 30156 20321 30159
rect 18524 30128 20321 30156
rect 18524 30116 18530 30128
rect 20309 30125 20321 30128
rect 20355 30125 20367 30159
rect 20309 30119 20367 30125
rect 20398 30116 20404 30168
rect 20456 30156 20462 30168
rect 20456 30128 20501 30156
rect 20456 30116 20462 30128
rect 22238 30116 22244 30168
rect 22296 30156 22302 30168
rect 22517 30159 22575 30165
rect 22517 30156 22529 30159
rect 22296 30128 22529 30156
rect 22296 30116 22302 30128
rect 22517 30125 22529 30128
rect 22563 30125 22575 30159
rect 22517 30119 22575 30125
rect 22606 30116 22612 30168
rect 22664 30156 22670 30168
rect 22900 30156 22928 30196
rect 23066 30184 23072 30196
rect 23124 30184 23130 30236
rect 24924 30224 24952 30264
rect 25090 30252 25096 30264
rect 25148 30252 25154 30304
rect 25826 30252 25832 30304
rect 25884 30292 25890 30304
rect 25921 30295 25979 30301
rect 25921 30292 25933 30295
rect 25884 30264 25933 30292
rect 25884 30252 25890 30264
rect 25921 30261 25933 30264
rect 25967 30261 25979 30295
rect 26746 30292 26752 30304
rect 26707 30264 26752 30292
rect 25921 30255 25979 30261
rect 26746 30252 26752 30264
rect 26804 30252 26810 30304
rect 26841 30295 26899 30301
rect 26841 30261 26853 30295
rect 26887 30292 26899 30295
rect 27114 30292 27120 30304
rect 26887 30264 27120 30292
rect 26887 30261 26899 30264
rect 26841 30255 26899 30261
rect 27114 30252 27120 30264
rect 27172 30252 27178 30304
rect 29877 30295 29935 30301
rect 29877 30292 29889 30295
rect 27684 30264 29889 30292
rect 27684 30224 27712 30264
rect 29877 30261 29889 30264
rect 29923 30292 29935 30295
rect 30794 30292 30800 30304
rect 29923 30264 30800 30292
rect 29923 30261 29935 30264
rect 29877 30255 29935 30261
rect 30794 30252 30800 30264
rect 30852 30252 30858 30304
rect 31349 30295 31407 30301
rect 31349 30261 31361 30295
rect 31395 30292 31407 30295
rect 31438 30292 31444 30304
rect 31395 30264 31444 30292
rect 31395 30261 31407 30264
rect 31349 30255 31407 30261
rect 31438 30252 31444 30264
rect 31496 30292 31502 30304
rect 32085 30295 32143 30301
rect 32085 30292 32097 30295
rect 31496 30264 32097 30292
rect 31496 30252 31502 30264
rect 32085 30261 32097 30264
rect 32131 30261 32143 30295
rect 32085 30255 32143 30261
rect 24924 30196 27712 30224
rect 28957 30227 29015 30233
rect 28957 30193 28969 30227
rect 29003 30224 29015 30227
rect 29046 30224 29052 30236
rect 29003 30196 29052 30224
rect 29003 30193 29015 30196
rect 28957 30187 29015 30193
rect 29046 30184 29052 30196
rect 29104 30184 29110 30236
rect 22974 30156 22980 30168
rect 22664 30128 22709 30156
rect 22900 30128 22980 30156
rect 22664 30116 22670 30128
rect 22974 30116 22980 30128
rect 23032 30116 23038 30168
rect 24722 30156 24728 30168
rect 24683 30128 24728 30156
rect 24722 30116 24728 30128
rect 24780 30116 24786 30168
rect 31898 30156 31904 30168
rect 31859 30128 31904 30156
rect 31898 30116 31904 30128
rect 31956 30116 31962 30168
rect 32545 30159 32603 30165
rect 32545 30125 32557 30159
rect 32591 30156 32603 30159
rect 32818 30156 32824 30168
rect 32591 30128 32824 30156
rect 32591 30125 32603 30128
rect 32545 30119 32603 30125
rect 32818 30116 32824 30128
rect 32876 30116 32882 30168
rect 11000 30066 34368 30088
rect 11000 30014 19142 30066
rect 19194 30014 19206 30066
rect 19258 30014 19270 30066
rect 19322 30014 19334 30066
rect 19386 30014 29142 30066
rect 29194 30014 29206 30066
rect 29258 30014 29270 30066
rect 29322 30014 29334 30066
rect 29386 30014 34368 30066
rect 11000 29992 34368 30014
rect 23066 29952 23072 29964
rect 21428 29924 23072 29952
rect 17822 29844 17828 29896
rect 17880 29844 17886 29896
rect 20214 29844 20220 29896
rect 20272 29884 20278 29896
rect 20401 29887 20459 29893
rect 20401 29884 20413 29887
rect 20272 29856 20413 29884
rect 20272 29844 20278 29856
rect 20401 29853 20413 29856
rect 20447 29853 20459 29887
rect 20401 29847 20459 29853
rect 20585 29887 20643 29893
rect 20585 29853 20597 29887
rect 20631 29884 20643 29887
rect 20950 29884 20956 29896
rect 20631 29856 20812 29884
rect 20911 29856 20956 29884
rect 20631 29853 20643 29856
rect 20585 29847 20643 29853
rect 14510 29776 14516 29828
rect 14568 29816 14574 29828
rect 16166 29816 16172 29828
rect 14568 29788 16172 29816
rect 14568 29776 14574 29788
rect 16166 29776 16172 29788
rect 16224 29776 16230 29828
rect 16810 29816 16816 29828
rect 16771 29788 16816 29816
rect 16810 29776 16816 29788
rect 16868 29776 16874 29828
rect 17086 29748 17092 29760
rect 17047 29720 17092 29748
rect 17086 29708 17092 29720
rect 17144 29708 17150 29760
rect 18466 29708 18472 29760
rect 18524 29748 18530 29760
rect 18837 29751 18895 29757
rect 18837 29748 18849 29751
rect 18524 29720 18849 29748
rect 18524 29708 18530 29720
rect 18837 29717 18849 29720
rect 18883 29717 18895 29751
rect 18837 29711 18895 29717
rect 19938 29708 19944 29760
rect 19996 29748 20002 29760
rect 20217 29751 20275 29757
rect 20217 29748 20229 29751
rect 19996 29720 20229 29748
rect 19996 29708 20002 29720
rect 20217 29717 20229 29720
rect 20263 29717 20275 29751
rect 20416 29748 20444 29847
rect 20493 29819 20551 29825
rect 20493 29785 20505 29819
rect 20539 29816 20551 29819
rect 20674 29816 20680 29828
rect 20539 29788 20680 29816
rect 20539 29785 20551 29788
rect 20493 29779 20551 29785
rect 20674 29776 20680 29788
rect 20732 29776 20738 29828
rect 20784 29816 20812 29856
rect 20950 29844 20956 29856
rect 21008 29844 21014 29896
rect 21428 29893 21456 29924
rect 23066 29912 23072 29924
rect 23124 29912 23130 29964
rect 24446 29912 24452 29964
rect 24504 29952 24510 29964
rect 24541 29955 24599 29961
rect 24541 29952 24553 29955
rect 24504 29924 24553 29952
rect 24504 29912 24510 29924
rect 24541 29921 24553 29924
rect 24587 29921 24599 29955
rect 24541 29915 24599 29921
rect 25090 29912 25096 29964
rect 25148 29952 25154 29964
rect 25461 29955 25519 29961
rect 25461 29952 25473 29955
rect 25148 29924 25473 29952
rect 25148 29912 25154 29924
rect 25461 29921 25473 29924
rect 25507 29921 25519 29955
rect 25461 29915 25519 29921
rect 26930 29912 26936 29964
rect 26988 29952 26994 29964
rect 26988 29924 27988 29952
rect 26988 29912 26994 29924
rect 21413 29887 21471 29893
rect 21413 29853 21425 29887
rect 21459 29853 21471 29887
rect 21965 29887 22023 29893
rect 21413 29847 21471 29853
rect 21520 29856 21732 29884
rect 20858 29816 20864 29828
rect 20784 29788 20864 29816
rect 20858 29776 20864 29788
rect 20916 29776 20922 29828
rect 21520 29748 21548 29856
rect 21597 29819 21655 29825
rect 21597 29785 21609 29819
rect 21643 29785 21655 29819
rect 21704 29816 21732 29856
rect 21965 29853 21977 29887
rect 22011 29884 22023 29887
rect 22514 29884 22520 29896
rect 22011 29856 22520 29884
rect 22011 29853 22023 29856
rect 21965 29847 22023 29853
rect 22514 29844 22520 29856
rect 22572 29844 22578 29896
rect 22698 29884 22704 29896
rect 22659 29856 22704 29884
rect 22698 29844 22704 29856
rect 22756 29844 22762 29896
rect 22793 29887 22851 29893
rect 22793 29853 22805 29887
rect 22839 29853 22851 29887
rect 22793 29847 22851 29853
rect 23161 29887 23219 29893
rect 23161 29853 23173 29887
rect 23207 29884 23219 29887
rect 23250 29884 23256 29896
rect 23207 29856 23256 29884
rect 23207 29853 23219 29856
rect 23161 29847 23219 29853
rect 22238 29816 22244 29828
rect 21704 29788 22244 29816
rect 21597 29779 21655 29785
rect 20416 29720 21548 29748
rect 21612 29748 21640 29779
rect 22238 29776 22244 29788
rect 22296 29816 22302 29828
rect 22609 29819 22667 29825
rect 22609 29816 22621 29819
rect 22296 29788 22621 29816
rect 22296 29776 22302 29788
rect 22609 29785 22621 29788
rect 22655 29785 22667 29819
rect 22808 29816 22836 29847
rect 23250 29844 23256 29856
rect 23308 29844 23314 29896
rect 23897 29887 23955 29893
rect 23897 29853 23909 29887
rect 23943 29884 23955 29887
rect 25274 29884 25280 29896
rect 23943 29856 25280 29884
rect 23943 29853 23955 29856
rect 23897 29847 23955 29853
rect 25274 29844 25280 29856
rect 25332 29844 25338 29896
rect 26749 29887 26807 29893
rect 26749 29853 26761 29887
rect 26795 29884 26807 29887
rect 26795 29856 27896 29884
rect 26795 29853 26807 29856
rect 26749 29847 26807 29853
rect 27868 29828 27896 29856
rect 23342 29816 23348 29828
rect 22808 29788 23348 29816
rect 22609 29779 22667 29785
rect 23342 29776 23348 29788
rect 23400 29776 23406 29828
rect 23986 29776 23992 29828
rect 24044 29825 24050 29828
rect 24044 29819 24102 29825
rect 24044 29785 24056 29819
rect 24090 29785 24102 29819
rect 25182 29816 25188 29828
rect 25143 29788 25188 29816
rect 24044 29779 24102 29785
rect 24044 29776 24050 29779
rect 25182 29776 25188 29788
rect 25240 29776 25246 29828
rect 25369 29819 25427 29825
rect 25369 29785 25381 29819
rect 25415 29816 25427 29819
rect 25458 29816 25464 29828
rect 25415 29788 25464 29816
rect 25415 29785 25427 29788
rect 25369 29779 25427 29785
rect 21612 29720 22284 29748
rect 20217 29711 20275 29717
rect 16350 29612 16356 29624
rect 16311 29584 16356 29612
rect 16350 29572 16356 29584
rect 16408 29572 16414 29624
rect 22256 29612 22284 29720
rect 22330 29708 22336 29760
rect 22388 29748 22394 29760
rect 22425 29751 22483 29757
rect 22425 29748 22437 29751
rect 22388 29720 22437 29748
rect 22388 29708 22394 29720
rect 22425 29717 22437 29720
rect 22471 29748 22483 29751
rect 22882 29748 22888 29760
rect 22471 29720 22888 29748
rect 22471 29717 22483 29720
rect 22425 29711 22483 29717
rect 22882 29708 22888 29720
rect 22940 29708 22946 29760
rect 24265 29751 24323 29757
rect 24265 29717 24277 29751
rect 24311 29748 24323 29751
rect 24630 29748 24636 29760
rect 24311 29720 24636 29748
rect 24311 29717 24323 29720
rect 24265 29711 24323 29717
rect 24630 29708 24636 29720
rect 24688 29708 24694 29760
rect 24173 29683 24231 29689
rect 24173 29649 24185 29683
rect 24219 29680 24231 29683
rect 24538 29680 24544 29692
rect 24219 29652 24544 29680
rect 24219 29649 24231 29652
rect 24173 29643 24231 29649
rect 24538 29640 24544 29652
rect 24596 29640 24602 29692
rect 25384 29612 25412 29779
rect 25458 29776 25464 29788
rect 25516 29776 25522 29828
rect 25826 29776 25832 29828
rect 25884 29816 25890 29828
rect 26197 29819 26255 29825
rect 26197 29816 26209 29819
rect 25884 29788 26209 29816
rect 25884 29776 25890 29788
rect 26197 29785 26209 29788
rect 26243 29785 26255 29819
rect 26378 29816 26384 29828
rect 26339 29788 26384 29816
rect 26197 29779 26255 29785
rect 26378 29776 26384 29788
rect 26436 29776 26442 29828
rect 27390 29816 27396 29828
rect 27351 29788 27396 29816
rect 27390 29776 27396 29788
rect 27448 29776 27454 29828
rect 27850 29816 27856 29828
rect 27763 29788 27856 29816
rect 27850 29776 27856 29788
rect 27908 29776 27914 29828
rect 27960 29825 27988 29924
rect 31806 29912 31812 29964
rect 31864 29912 31870 29964
rect 28494 29884 28500 29896
rect 28455 29856 28500 29884
rect 28494 29844 28500 29856
rect 28552 29844 28558 29896
rect 29598 29844 29604 29896
rect 29656 29884 29662 29896
rect 29693 29887 29751 29893
rect 29693 29884 29705 29887
rect 29656 29856 29705 29884
rect 29656 29844 29662 29856
rect 29693 29853 29705 29856
rect 29739 29853 29751 29887
rect 29693 29847 29751 29853
rect 30981 29887 31039 29893
rect 30981 29853 30993 29887
rect 31027 29884 31039 29887
rect 31162 29884 31168 29896
rect 31027 29856 31168 29884
rect 31027 29853 31039 29856
rect 30981 29847 31039 29853
rect 31162 29844 31168 29856
rect 31220 29844 31226 29896
rect 27945 29819 28003 29825
rect 27945 29785 27957 29819
rect 27991 29785 28003 29819
rect 27945 29779 28003 29785
rect 28954 29776 28960 29828
rect 29012 29816 29018 29828
rect 29049 29819 29107 29825
rect 29049 29816 29061 29819
rect 29012 29788 29061 29816
rect 29012 29776 29018 29788
rect 29049 29785 29061 29788
rect 29095 29785 29107 29819
rect 29966 29816 29972 29828
rect 29927 29788 29972 29816
rect 29049 29779 29107 29785
rect 29966 29776 29972 29788
rect 30024 29776 30030 29828
rect 31824 29825 31852 29912
rect 31898 29844 31904 29896
rect 31956 29884 31962 29896
rect 32913 29887 32971 29893
rect 32913 29884 32925 29887
rect 31956 29856 32925 29884
rect 31956 29844 31962 29856
rect 32913 29853 32925 29856
rect 32959 29853 32971 29887
rect 32913 29847 32971 29853
rect 31717 29819 31775 29825
rect 31717 29816 31729 29819
rect 30076 29788 31729 29816
rect 26746 29708 26752 29760
rect 26804 29748 26810 29760
rect 27301 29751 27359 29757
rect 27301 29748 27313 29751
rect 26804 29720 27313 29748
rect 26804 29708 26810 29720
rect 27301 29717 27313 29720
rect 27347 29717 27359 29751
rect 27301 29711 27359 29717
rect 27316 29680 27344 29711
rect 28862 29680 28868 29692
rect 27316 29652 28868 29680
rect 28862 29640 28868 29652
rect 28920 29680 28926 29692
rect 30076 29680 30104 29788
rect 31717 29785 31729 29788
rect 31763 29785 31775 29819
rect 31717 29779 31775 29785
rect 31809 29819 31867 29825
rect 31809 29785 31821 29819
rect 31855 29785 31867 29819
rect 31809 29779 31867 29785
rect 30886 29748 30892 29760
rect 30847 29720 30892 29748
rect 30886 29708 30892 29720
rect 30944 29708 30950 29760
rect 31162 29708 31168 29760
rect 31220 29748 31226 29760
rect 32361 29751 32419 29757
rect 32361 29748 32373 29751
rect 31220 29720 32373 29748
rect 31220 29708 31226 29720
rect 32361 29717 32373 29720
rect 32407 29717 32419 29751
rect 32361 29711 32419 29717
rect 32818 29680 32824 29692
rect 28920 29652 30104 29680
rect 32779 29652 32824 29680
rect 28920 29640 28926 29652
rect 32818 29640 32824 29652
rect 32876 29640 32882 29692
rect 26102 29612 26108 29624
rect 22256 29584 26108 29612
rect 26102 29572 26108 29584
rect 26160 29572 26166 29624
rect 11000 29522 34368 29544
rect 11000 29470 14142 29522
rect 14194 29470 14206 29522
rect 14258 29470 14270 29522
rect 14322 29470 14334 29522
rect 14386 29470 24142 29522
rect 24194 29470 24206 29522
rect 24258 29470 24270 29522
rect 24322 29470 24334 29522
rect 24386 29470 34368 29522
rect 11000 29448 34368 29470
rect 23986 29368 23992 29420
rect 24044 29408 24050 29420
rect 24541 29411 24599 29417
rect 24541 29408 24553 29411
rect 24044 29380 24553 29408
rect 24044 29368 24050 29380
rect 24541 29377 24553 29380
rect 24587 29377 24599 29411
rect 24541 29371 24599 29377
rect 28034 29368 28040 29420
rect 28092 29408 28098 29420
rect 28221 29411 28279 29417
rect 28221 29408 28233 29411
rect 28092 29380 28233 29408
rect 28092 29368 28098 29380
rect 28221 29377 28233 29380
rect 28267 29377 28279 29411
rect 28221 29371 28279 29377
rect 13958 29300 13964 29352
rect 14016 29340 14022 29352
rect 27942 29340 27948 29352
rect 14016 29312 27948 29340
rect 14016 29300 14022 29312
rect 27942 29300 27948 29312
rect 28000 29300 28006 29352
rect 29417 29343 29475 29349
rect 29417 29309 29429 29343
rect 29463 29340 29475 29343
rect 29598 29340 29604 29352
rect 29463 29312 29604 29340
rect 29463 29309 29475 29312
rect 29417 29303 29475 29309
rect 29598 29300 29604 29312
rect 29656 29300 29662 29352
rect 21226 29232 21232 29284
rect 21284 29272 21290 29284
rect 21321 29275 21379 29281
rect 21321 29272 21333 29275
rect 21284 29244 21333 29272
rect 21284 29232 21290 29244
rect 21321 29241 21333 29244
rect 21367 29272 21379 29275
rect 21870 29272 21876 29284
rect 21367 29244 21876 29272
rect 21367 29241 21379 29244
rect 21321 29235 21379 29241
rect 21870 29232 21876 29244
rect 21928 29232 21934 29284
rect 25826 29272 25832 29284
rect 25787 29244 25832 29272
rect 25826 29232 25832 29244
rect 25884 29232 25890 29284
rect 16994 29204 17000 29216
rect 16955 29176 17000 29204
rect 16994 29164 17000 29176
rect 17052 29164 17058 29216
rect 17089 29207 17147 29213
rect 17089 29173 17101 29207
rect 17135 29204 17147 29207
rect 17178 29204 17184 29216
rect 17135 29176 17184 29204
rect 17135 29173 17147 29176
rect 17089 29167 17147 29173
rect 17178 29164 17184 29176
rect 17236 29164 17242 29216
rect 17270 29164 17276 29216
rect 17328 29204 17334 29216
rect 17328 29176 17373 29204
rect 17328 29164 17334 29176
rect 17730 29164 17736 29216
rect 17788 29204 17794 29216
rect 18561 29207 18619 29213
rect 18561 29204 18573 29207
rect 17788 29176 18573 29204
rect 17788 29164 17794 29176
rect 18561 29173 18573 29176
rect 18607 29173 18619 29207
rect 18561 29167 18619 29173
rect 20769 29207 20827 29213
rect 20769 29173 20781 29207
rect 20815 29204 20827 29207
rect 21410 29204 21416 29216
rect 20815 29176 21416 29204
rect 20815 29173 20827 29176
rect 20769 29167 20827 29173
rect 21410 29164 21416 29176
rect 21468 29164 21474 29216
rect 22698 29164 22704 29216
rect 22756 29204 22762 29216
rect 23253 29207 23311 29213
rect 23253 29204 23265 29207
rect 22756 29176 23265 29204
rect 22756 29164 22762 29176
rect 23253 29173 23265 29176
rect 23299 29173 23311 29207
rect 24446 29204 24452 29216
rect 24407 29176 24452 29204
rect 23253 29167 23311 29173
rect 24446 29164 24452 29176
rect 24504 29164 24510 29216
rect 25090 29164 25096 29216
rect 25148 29204 25154 29216
rect 25277 29207 25335 29213
rect 25277 29204 25289 29207
rect 25148 29176 25289 29204
rect 25148 29164 25154 29176
rect 25277 29173 25289 29176
rect 25323 29173 25335 29207
rect 25277 29167 25335 29173
rect 25458 29164 25464 29216
rect 25516 29204 25522 29216
rect 26473 29207 26531 29213
rect 26473 29204 26485 29207
rect 25516 29176 25561 29204
rect 25660 29176 26485 29204
rect 25516 29164 25522 29176
rect 19205 29139 19263 29145
rect 19205 29105 19217 29139
rect 19251 29136 19263 29139
rect 19938 29136 19944 29148
rect 19251 29108 19944 29136
rect 19251 29105 19263 29108
rect 19205 29099 19263 29105
rect 19938 29096 19944 29108
rect 19996 29136 20002 29148
rect 20585 29139 20643 29145
rect 20585 29136 20597 29139
rect 19996 29108 20597 29136
rect 19996 29096 20002 29108
rect 20585 29105 20597 29108
rect 20631 29105 20643 29139
rect 20950 29136 20956 29148
rect 20911 29108 20956 29136
rect 20585 29099 20643 29105
rect 20950 29096 20956 29108
rect 21008 29096 21014 29148
rect 22882 29096 22888 29148
rect 22940 29136 22946 29148
rect 22977 29139 23035 29145
rect 22977 29136 22989 29139
rect 22940 29108 22989 29136
rect 22940 29096 22946 29108
rect 22977 29105 22989 29108
rect 23023 29105 23035 29139
rect 23342 29136 23348 29148
rect 23303 29108 23348 29136
rect 22977 29099 23035 29105
rect 23342 29096 23348 29108
rect 23400 29096 23406 29148
rect 23710 29136 23716 29148
rect 23671 29108 23716 29136
rect 23710 29096 23716 29108
rect 23768 29096 23774 29148
rect 23894 29096 23900 29148
rect 23952 29136 23958 29148
rect 24265 29139 24323 29145
rect 24265 29136 24277 29139
rect 23952 29108 24277 29136
rect 23952 29096 23958 29108
rect 24265 29105 24277 29108
rect 24311 29105 24323 29139
rect 24265 29099 24323 29105
rect 25550 29096 25556 29148
rect 25608 29136 25614 29148
rect 25660 29136 25688 29176
rect 26473 29173 26485 29176
rect 26519 29173 26531 29207
rect 26473 29167 26531 29173
rect 26562 29164 26568 29216
rect 26620 29204 26626 29216
rect 26841 29207 26899 29213
rect 26841 29204 26853 29207
rect 26620 29176 26853 29204
rect 26620 29164 26626 29176
rect 26841 29173 26853 29176
rect 26887 29204 26899 29207
rect 28129 29207 28187 29213
rect 28129 29204 28141 29207
rect 26887 29176 28141 29204
rect 26887 29173 26899 29176
rect 26841 29167 26899 29173
rect 28129 29173 28141 29176
rect 28175 29173 28187 29207
rect 28954 29204 28960 29216
rect 28915 29176 28960 29204
rect 28129 29167 28187 29173
rect 28954 29164 28960 29176
rect 29012 29164 29018 29216
rect 30521 29207 30579 29213
rect 30521 29173 30533 29207
rect 30567 29204 30579 29207
rect 31162 29204 31168 29216
rect 30567 29176 31168 29204
rect 30567 29173 30579 29176
rect 30521 29167 30579 29173
rect 31162 29164 31168 29176
rect 31220 29164 31226 29216
rect 31257 29207 31315 29213
rect 31257 29173 31269 29207
rect 31303 29204 31315 29207
rect 32818 29204 32824 29216
rect 31303 29176 32824 29204
rect 31303 29173 31315 29176
rect 31257 29167 31315 29173
rect 32818 29164 32824 29176
rect 32876 29164 32882 29216
rect 26286 29136 26292 29148
rect 25608 29108 25688 29136
rect 26247 29108 26292 29136
rect 25608 29096 25614 29108
rect 26286 29096 26292 29108
rect 26344 29096 26350 29148
rect 26654 29096 26660 29148
rect 26712 29136 26718 29148
rect 27945 29139 28003 29145
rect 27945 29136 27957 29139
rect 26712 29108 27957 29136
rect 26712 29096 26718 29108
rect 27945 29105 27957 29108
rect 27991 29105 28003 29139
rect 27945 29099 28003 29105
rect 29506 29096 29512 29148
rect 29564 29136 29570 29148
rect 31438 29136 31444 29148
rect 29564 29108 29609 29136
rect 31399 29108 31444 29136
rect 29564 29096 29570 29108
rect 31438 29096 31444 29108
rect 31496 29096 31502 29148
rect 20490 29028 20496 29080
rect 20548 29068 20554 29080
rect 20861 29071 20919 29077
rect 20861 29068 20873 29071
rect 20548 29040 20873 29068
rect 20548 29028 20554 29040
rect 20861 29037 20873 29040
rect 20907 29068 20919 29071
rect 22698 29068 22704 29080
rect 20907 29040 22704 29068
rect 20907 29037 20919 29040
rect 20861 29031 20919 29037
rect 22698 29028 22704 29040
rect 22756 29028 22762 29080
rect 23158 29068 23164 29080
rect 23119 29040 23164 29068
rect 23158 29028 23164 29040
rect 23216 29028 23222 29080
rect 25090 29028 25096 29080
rect 25148 29068 25154 29080
rect 26378 29068 26384 29080
rect 25148 29040 26384 29068
rect 25148 29028 25154 29040
rect 26378 29028 26384 29040
rect 26436 29028 26442 29080
rect 11000 28978 34368 29000
rect 11000 28926 19142 28978
rect 19194 28926 19206 28978
rect 19258 28926 19270 28978
rect 19322 28926 19334 28978
rect 19386 28926 29142 28978
rect 29194 28926 29206 28978
rect 29258 28926 29270 28978
rect 29322 28926 29334 28978
rect 29386 28926 34368 28978
rect 11000 28904 34368 28926
rect 16902 28864 16908 28876
rect 15356 28836 16908 28864
rect 15356 28740 15384 28836
rect 16902 28824 16908 28836
rect 16960 28824 16966 28876
rect 23069 28867 23127 28873
rect 23069 28864 23081 28867
rect 21704 28836 23081 28864
rect 21704 28808 21732 28836
rect 23069 28833 23081 28836
rect 23115 28864 23127 28867
rect 23158 28864 23164 28876
rect 23115 28836 23164 28864
rect 23115 28833 23127 28836
rect 23069 28827 23127 28833
rect 23158 28824 23164 28836
rect 23216 28824 23222 28876
rect 24446 28824 24452 28876
rect 24504 28864 24510 28876
rect 25458 28864 25464 28876
rect 24504 28836 25464 28864
rect 24504 28824 24510 28836
rect 25458 28824 25464 28836
rect 25516 28824 25522 28876
rect 29141 28867 29199 28873
rect 29141 28833 29153 28867
rect 29187 28864 29199 28867
rect 29506 28864 29512 28876
rect 29187 28836 29512 28864
rect 29187 28833 29199 28836
rect 29141 28827 29199 28833
rect 29506 28824 29512 28836
rect 29564 28824 29570 28876
rect 31438 28824 31444 28876
rect 31496 28864 31502 28876
rect 31625 28867 31683 28873
rect 31625 28864 31637 28867
rect 31496 28836 31637 28864
rect 31496 28824 31502 28836
rect 31625 28833 31637 28836
rect 31671 28833 31683 28867
rect 31625 28827 31683 28833
rect 16350 28756 16356 28808
rect 16408 28756 16414 28808
rect 17270 28756 17276 28808
rect 17328 28796 17334 28808
rect 20585 28799 20643 28805
rect 17328 28768 18052 28796
rect 17328 28756 17334 28768
rect 14421 28731 14479 28737
rect 14421 28697 14433 28731
rect 14467 28728 14479 28731
rect 14510 28728 14516 28740
rect 14467 28700 14516 28728
rect 14467 28697 14479 28700
rect 14421 28691 14479 28697
rect 14510 28688 14516 28700
rect 14568 28728 14574 28740
rect 14786 28728 14792 28740
rect 14568 28700 14792 28728
rect 14568 28688 14574 28700
rect 14786 28688 14792 28700
rect 14844 28688 14850 28740
rect 15338 28728 15344 28740
rect 15251 28700 15344 28728
rect 15338 28688 15344 28700
rect 15396 28688 15402 28740
rect 16994 28688 17000 28740
rect 17052 28728 17058 28740
rect 18024 28737 18052 28768
rect 20585 28765 20597 28799
rect 20631 28796 20643 28799
rect 20950 28796 20956 28808
rect 20631 28768 20956 28796
rect 20631 28765 20643 28768
rect 20585 28759 20643 28765
rect 20950 28756 20956 28768
rect 21008 28796 21014 28808
rect 21410 28796 21416 28808
rect 21008 28768 21272 28796
rect 21371 28768 21416 28796
rect 21008 28756 21014 28768
rect 21244 28737 21272 28768
rect 21410 28756 21416 28768
rect 21468 28796 21474 28808
rect 21686 28796 21692 28808
rect 21468 28768 21692 28796
rect 21468 28756 21474 28768
rect 21686 28756 21692 28768
rect 21744 28756 21750 28808
rect 22882 28796 22888 28808
rect 22843 28768 22888 28796
rect 22882 28756 22888 28768
rect 22940 28756 22946 28808
rect 22974 28756 22980 28808
rect 23032 28796 23038 28808
rect 23253 28799 23311 28805
rect 23253 28796 23265 28799
rect 23032 28768 23265 28796
rect 23032 28756 23038 28768
rect 23253 28765 23265 28768
rect 23299 28765 23311 28799
rect 23253 28759 23311 28765
rect 23710 28756 23716 28808
rect 23768 28796 23774 28808
rect 24081 28799 24139 28805
rect 24081 28796 24093 28799
rect 23768 28768 24093 28796
rect 23768 28756 23774 28768
rect 24081 28765 24093 28768
rect 24127 28796 24139 28799
rect 27117 28799 27175 28805
rect 24127 28768 25412 28796
rect 24127 28765 24139 28768
rect 24081 28759 24139 28765
rect 17825 28731 17883 28737
rect 17825 28728 17837 28731
rect 17052 28700 17837 28728
rect 17052 28688 17058 28700
rect 17825 28697 17837 28700
rect 17871 28697 17883 28731
rect 17825 28691 17883 28697
rect 18009 28731 18067 28737
rect 18009 28697 18021 28731
rect 18055 28697 18067 28731
rect 18009 28691 18067 28697
rect 20493 28731 20551 28737
rect 20493 28697 20505 28731
rect 20539 28728 20551 28731
rect 21229 28731 21287 28737
rect 20539 28700 21180 28728
rect 20539 28697 20551 28700
rect 20493 28691 20551 28697
rect 15617 28663 15675 28669
rect 15617 28629 15629 28663
rect 15663 28660 15675 28663
rect 16810 28660 16816 28672
rect 15663 28632 16816 28660
rect 15663 28629 15675 28632
rect 15617 28623 15675 28629
rect 16810 28620 16816 28632
rect 16868 28620 16874 28672
rect 17365 28663 17423 28669
rect 17365 28629 17377 28663
rect 17411 28660 17423 28663
rect 17730 28660 17736 28672
rect 17411 28632 17736 28660
rect 17411 28629 17423 28632
rect 17365 28623 17423 28629
rect 17730 28620 17736 28632
rect 17788 28620 17794 28672
rect 18282 28660 18288 28672
rect 18243 28632 18288 28660
rect 18282 28620 18288 28632
rect 18340 28620 18346 28672
rect 21045 28663 21103 28669
rect 21045 28629 21057 28663
rect 21091 28629 21103 28663
rect 21045 28623 21103 28629
rect 20490 28552 20496 28604
rect 20548 28592 20554 28604
rect 21060 28592 21088 28623
rect 20548 28564 21088 28592
rect 21152 28592 21180 28700
rect 21229 28697 21241 28731
rect 21275 28697 21287 28731
rect 21229 28691 21287 28697
rect 21321 28731 21379 28737
rect 21321 28697 21333 28731
rect 21367 28728 21379 28731
rect 21502 28728 21508 28740
rect 21367 28700 21508 28728
rect 21367 28697 21379 28700
rect 21321 28691 21379 28697
rect 21244 28660 21272 28691
rect 21502 28688 21508 28700
rect 21560 28688 21566 28740
rect 22606 28728 22612 28740
rect 21612 28700 22612 28728
rect 21612 28660 21640 28700
rect 22606 28688 22612 28700
rect 22664 28688 22670 28740
rect 22698 28688 22704 28740
rect 22756 28728 22762 28740
rect 23161 28731 23219 28737
rect 23161 28728 23173 28731
rect 22756 28700 23173 28728
rect 22756 28688 22762 28700
rect 23161 28697 23173 28700
rect 23207 28697 23219 28731
rect 24265 28731 24323 28737
rect 24265 28728 24277 28731
rect 23161 28691 23219 28697
rect 23544 28700 24277 28728
rect 21778 28660 21784 28672
rect 21244 28632 21640 28660
rect 21739 28632 21784 28660
rect 21778 28620 21784 28632
rect 21836 28620 21842 28672
rect 21870 28620 21876 28672
rect 21928 28660 21934 28672
rect 23544 28660 23572 28700
rect 24265 28697 24277 28700
rect 24311 28728 24323 28731
rect 25090 28728 25096 28740
rect 24311 28700 25096 28728
rect 24311 28697 24323 28700
rect 24265 28691 24323 28697
rect 25090 28688 25096 28700
rect 25148 28688 25154 28740
rect 25384 28737 25412 28768
rect 27117 28765 27129 28799
rect 27163 28796 27175 28799
rect 28954 28796 28960 28808
rect 27163 28768 28960 28796
rect 27163 28765 27175 28768
rect 27117 28759 27175 28765
rect 28954 28756 28960 28768
rect 29012 28756 29018 28808
rect 25185 28731 25243 28737
rect 25185 28697 25197 28731
rect 25231 28697 25243 28731
rect 25185 28691 25243 28697
rect 25369 28731 25427 28737
rect 25369 28697 25381 28731
rect 25415 28697 25427 28731
rect 25369 28691 25427 28697
rect 27853 28731 27911 28737
rect 27853 28697 27865 28731
rect 27899 28697 27911 28731
rect 27853 28691 27911 28697
rect 21928 28632 23572 28660
rect 23621 28663 23679 28669
rect 21928 28620 21934 28632
rect 23621 28629 23633 28663
rect 23667 28660 23679 28663
rect 24446 28660 24452 28672
rect 23667 28632 24452 28660
rect 23667 28629 23679 28632
rect 23621 28623 23679 28629
rect 24446 28620 24452 28632
rect 24504 28660 24510 28672
rect 25200 28660 25228 28691
rect 27022 28660 27028 28672
rect 24504 28632 25228 28660
rect 26983 28632 27028 28660
rect 24504 28620 24510 28632
rect 27022 28620 27028 28632
rect 27080 28620 27086 28672
rect 27868 28660 27896 28691
rect 27942 28688 27948 28740
rect 28000 28728 28006 28740
rect 29325 28731 29383 28737
rect 28000 28700 28045 28728
rect 28000 28688 28006 28700
rect 29325 28697 29337 28731
rect 29371 28728 29383 28731
rect 29966 28728 29972 28740
rect 29371 28700 29972 28728
rect 29371 28697 29383 28700
rect 29325 28691 29383 28697
rect 29966 28688 29972 28700
rect 30024 28688 30030 28740
rect 31346 28688 31352 28740
rect 31404 28728 31410 28740
rect 31533 28731 31591 28737
rect 31533 28728 31545 28731
rect 31404 28700 31545 28728
rect 31404 28688 31410 28700
rect 31533 28697 31545 28700
rect 31579 28697 31591 28731
rect 31533 28691 31591 28697
rect 28954 28660 28960 28672
rect 27868 28632 28960 28660
rect 28954 28620 28960 28632
rect 29012 28620 29018 28672
rect 23066 28592 23072 28604
rect 21152 28564 23072 28592
rect 20548 28552 20554 28564
rect 23066 28552 23072 28564
rect 23124 28552 23130 28604
rect 14510 28484 14516 28536
rect 14568 28524 14574 28536
rect 14605 28527 14663 28533
rect 14605 28524 14617 28527
rect 14568 28496 14617 28524
rect 14568 28484 14574 28496
rect 14605 28493 14617 28496
rect 14651 28493 14663 28527
rect 14605 28487 14663 28493
rect 24357 28527 24415 28533
rect 24357 28493 24369 28527
rect 24403 28524 24415 28527
rect 26746 28524 26752 28536
rect 24403 28496 26752 28524
rect 24403 28493 24415 28496
rect 24357 28487 24415 28493
rect 26746 28484 26752 28496
rect 26804 28484 26810 28536
rect 11000 28434 34368 28456
rect 11000 28382 14142 28434
rect 14194 28382 14206 28434
rect 14258 28382 14270 28434
rect 14322 28382 14334 28434
rect 14386 28382 24142 28434
rect 24194 28382 24206 28434
rect 24258 28382 24270 28434
rect 24322 28382 24334 28434
rect 24386 28382 34368 28434
rect 11000 28360 34368 28382
rect 21505 28323 21563 28329
rect 21505 28289 21517 28323
rect 21551 28320 21563 28323
rect 22422 28320 22428 28332
rect 21551 28292 22428 28320
rect 21551 28289 21563 28292
rect 21505 28283 21563 28289
rect 22422 28280 22428 28292
rect 22480 28280 22486 28332
rect 25826 28280 25832 28332
rect 25884 28320 25890 28332
rect 26565 28323 26623 28329
rect 26565 28320 26577 28323
rect 25884 28292 26577 28320
rect 25884 28280 25890 28292
rect 26565 28289 26577 28292
rect 26611 28289 26623 28323
rect 26565 28283 26623 28289
rect 23342 28252 23348 28264
rect 22348 28224 23348 28252
rect 13777 28187 13835 28193
rect 13777 28153 13789 28187
rect 13823 28184 13835 28187
rect 14142 28184 14148 28196
rect 13823 28156 14148 28184
rect 13823 28153 13835 28156
rect 13777 28147 13835 28153
rect 14142 28144 14148 28156
rect 14200 28144 14206 28196
rect 16721 28187 16779 28193
rect 16721 28153 16733 28187
rect 16767 28184 16779 28187
rect 16810 28184 16816 28196
rect 16767 28156 16816 28184
rect 16767 28153 16779 28156
rect 16721 28147 16779 28153
rect 16810 28144 16816 28156
rect 16868 28144 16874 28196
rect 22348 28184 22376 28224
rect 23342 28212 23348 28224
rect 23400 28252 23406 28264
rect 27114 28252 27120 28264
rect 23400 28224 23664 28252
rect 23400 28212 23406 28224
rect 22606 28184 22612 28196
rect 21336 28156 21548 28184
rect 13501 28119 13559 28125
rect 13501 28085 13513 28119
rect 13547 28085 13559 28119
rect 17178 28116 17184 28128
rect 17139 28088 17184 28116
rect 13501 28079 13559 28085
rect 13516 27980 13544 28079
rect 17178 28076 17184 28088
rect 17236 28076 17242 28128
rect 17457 28119 17515 28125
rect 17457 28085 17469 28119
rect 17503 28085 17515 28119
rect 17638 28116 17644 28128
rect 17599 28088 17644 28116
rect 17457 28079 17515 28085
rect 14510 28008 14516 28060
rect 14568 28008 14574 28060
rect 15430 28008 15436 28060
rect 15488 28048 15494 28060
rect 15525 28051 15583 28057
rect 15525 28048 15537 28051
rect 15488 28020 15537 28048
rect 15488 28008 15494 28020
rect 15525 28017 15537 28020
rect 15571 28017 15583 28051
rect 17472 28048 17500 28079
rect 17638 28076 17644 28088
rect 17696 28076 17702 28128
rect 17730 28076 17736 28128
rect 17788 28116 17794 28128
rect 17825 28119 17883 28125
rect 17825 28116 17837 28119
rect 17788 28088 17837 28116
rect 17788 28076 17794 28088
rect 17825 28085 17837 28088
rect 17871 28085 17883 28119
rect 18190 28116 18196 28128
rect 18151 28088 18196 28116
rect 17825 28079 17883 28085
rect 18190 28076 18196 28088
rect 18248 28076 18254 28128
rect 18837 28119 18895 28125
rect 18837 28116 18849 28119
rect 18760 28088 18849 28116
rect 18282 28048 18288 28060
rect 17472 28020 18288 28048
rect 15525 28011 15583 28017
rect 13774 27980 13780 27992
rect 13516 27952 13780 27980
rect 13774 27940 13780 27952
rect 13832 27980 13838 27992
rect 15338 27980 15344 27992
rect 13832 27952 15344 27980
rect 13832 27940 13838 27952
rect 15338 27940 15344 27952
rect 15396 27940 15402 27992
rect 15540 27980 15568 28011
rect 18282 28008 18288 28020
rect 18340 28008 18346 28060
rect 18760 27980 18788 28088
rect 18837 28085 18849 28088
rect 18883 28085 18895 28119
rect 20030 28116 20036 28128
rect 19991 28088 20036 28116
rect 18837 28079 18895 28085
rect 20030 28076 20036 28088
rect 20088 28076 20094 28128
rect 20677 28119 20735 28125
rect 20677 28085 20689 28119
rect 20723 28116 20735 28119
rect 21336 28116 21364 28156
rect 20723 28088 21364 28116
rect 21413 28119 21471 28125
rect 20723 28085 20735 28088
rect 20677 28079 20735 28085
rect 21413 28085 21425 28119
rect 21459 28085 21471 28119
rect 21520 28116 21548 28156
rect 22164 28156 22376 28184
rect 22440 28156 22612 28184
rect 22164 28116 22192 28156
rect 22330 28116 22336 28128
rect 21520 28088 22192 28116
rect 22291 28088 22336 28116
rect 21413 28079 21471 28085
rect 19481 28051 19539 28057
rect 19481 28017 19493 28051
rect 19527 28048 19539 28051
rect 20490 28048 20496 28060
rect 19527 28020 20496 28048
rect 19527 28017 19539 28020
rect 19481 28011 19539 28017
rect 20490 28008 20496 28020
rect 20548 28008 20554 28060
rect 21229 28051 21287 28057
rect 21229 28017 21241 28051
rect 21275 28017 21287 28051
rect 21428 28048 21456 28079
rect 22330 28076 22336 28088
rect 22388 28076 22394 28128
rect 22440 28125 22468 28156
rect 22606 28144 22612 28156
rect 22664 28144 22670 28196
rect 22440 28119 22503 28125
rect 22440 28088 22457 28119
rect 22445 28085 22457 28088
rect 22491 28085 22503 28119
rect 23529 28119 23587 28125
rect 23529 28116 23541 28119
rect 22445 28079 22503 28085
rect 22716 28088 23541 28116
rect 22606 28048 22612 28060
rect 21428 28020 22612 28048
rect 21229 28011 21287 28017
rect 20398 27980 20404 27992
rect 15540 27952 20404 27980
rect 20398 27940 20404 27952
rect 20456 27940 20462 27992
rect 21244 27980 21272 28011
rect 22606 28008 22612 28020
rect 22664 28048 22670 28060
rect 22716 28048 22744 28088
rect 23529 28085 23541 28088
rect 23575 28085 23587 28119
rect 23636 28116 23664 28224
rect 26856 28224 27120 28252
rect 26856 28196 26884 28224
rect 27114 28212 27120 28224
rect 27172 28212 27178 28264
rect 25090 28144 25096 28196
rect 25148 28184 25154 28196
rect 25185 28187 25243 28193
rect 25185 28184 25197 28187
rect 25148 28156 25197 28184
rect 25148 28144 25154 28156
rect 25185 28153 25197 28156
rect 25231 28153 25243 28187
rect 25185 28147 25243 28153
rect 25476 28156 25872 28184
rect 25476 28128 25504 28156
rect 25277 28119 25335 28125
rect 23636 28088 24768 28116
rect 23529 28079 23587 28085
rect 22882 28048 22888 28060
rect 22664 28020 22744 28048
rect 22843 28020 22888 28048
rect 22664 28008 22670 28020
rect 22882 28008 22888 28020
rect 22940 28008 22946 28060
rect 23342 28048 23348 28060
rect 23303 28020 23348 28048
rect 23342 28008 23348 28020
rect 23400 28008 23406 28060
rect 24633 28051 24691 28057
rect 24633 28017 24645 28051
rect 24679 28017 24691 28051
rect 24740 28048 24768 28088
rect 25277 28085 25289 28119
rect 25323 28116 25335 28119
rect 25458 28116 25464 28128
rect 25323 28088 25464 28116
rect 25323 28085 25335 28088
rect 25277 28079 25335 28085
rect 25458 28076 25464 28088
rect 25516 28076 25522 28128
rect 25645 28119 25703 28125
rect 25645 28085 25657 28119
rect 25691 28085 25703 28119
rect 25645 28079 25703 28085
rect 25737 28119 25795 28125
rect 25737 28085 25749 28119
rect 25783 28085 25795 28119
rect 25844 28116 25872 28156
rect 26838 28144 26844 28196
rect 26896 28144 26902 28196
rect 29509 28187 29567 28193
rect 29509 28153 29521 28187
rect 29555 28184 29567 28187
rect 31070 28184 31076 28196
rect 29555 28156 31076 28184
rect 29555 28153 29567 28156
rect 29509 28147 29567 28153
rect 31070 28144 31076 28156
rect 31128 28144 31134 28196
rect 26473 28119 26531 28125
rect 26473 28116 26485 28119
rect 25844 28088 26485 28116
rect 25737 28079 25795 28085
rect 26473 28085 26485 28088
rect 26519 28085 26531 28119
rect 28586 28116 28592 28128
rect 28547 28088 28592 28116
rect 26473 28079 26531 28085
rect 25660 28048 25688 28079
rect 24740 28020 25688 28048
rect 25752 28048 25780 28079
rect 28586 28076 28592 28088
rect 28644 28076 28650 28128
rect 28954 28076 28960 28128
rect 29012 28116 29018 28128
rect 29417 28119 29475 28125
rect 29417 28116 29429 28119
rect 29012 28088 29429 28116
rect 29012 28076 29018 28088
rect 29417 28085 29429 28088
rect 29463 28085 29475 28119
rect 29417 28079 29475 28085
rect 25918 28048 25924 28060
rect 25752 28020 25924 28048
rect 24633 28011 24691 28017
rect 22900 27980 22928 28008
rect 23618 27980 23624 27992
rect 21244 27952 22928 27980
rect 23579 27952 23624 27980
rect 23618 27940 23624 27952
rect 23676 27940 23682 27992
rect 24648 27980 24676 28011
rect 25918 28008 25924 28020
rect 25976 28008 25982 28060
rect 26286 28048 26292 28060
rect 26199 28020 26292 28048
rect 26286 28008 26292 28020
rect 26344 28008 26350 28060
rect 28681 28051 28739 28057
rect 28681 28017 28693 28051
rect 28727 28017 28739 28051
rect 28681 28011 28739 28017
rect 24998 27980 25004 27992
rect 24648 27952 25004 27980
rect 24998 27940 25004 27952
rect 25056 27940 25062 27992
rect 25642 27940 25648 27992
rect 25700 27980 25706 27992
rect 26304 27980 26332 28008
rect 25700 27952 26332 27980
rect 28696 27980 28724 28011
rect 29506 27980 29512 27992
rect 28696 27952 29512 27980
rect 25700 27940 25706 27952
rect 29506 27940 29512 27952
rect 29564 27940 29570 27992
rect 11000 27890 34368 27912
rect 11000 27838 19142 27890
rect 19194 27838 19206 27890
rect 19258 27838 19270 27890
rect 19322 27838 19334 27890
rect 19386 27838 29142 27890
rect 29194 27838 29206 27890
rect 29258 27838 29270 27890
rect 29322 27838 29334 27890
rect 29386 27838 34368 27890
rect 11000 27816 34368 27838
rect 20214 27776 20220 27788
rect 20175 27748 20220 27776
rect 20214 27736 20220 27748
rect 20272 27736 20278 27788
rect 20582 27736 20588 27788
rect 20640 27776 20646 27788
rect 24814 27776 24820 27788
rect 20640 27748 24820 27776
rect 20640 27736 20646 27748
rect 14053 27711 14111 27717
rect 14053 27677 14065 27711
rect 14099 27708 14111 27711
rect 14142 27708 14148 27720
rect 14099 27680 14148 27708
rect 14099 27677 14111 27680
rect 14053 27671 14111 27677
rect 14142 27668 14148 27680
rect 14200 27668 14206 27720
rect 16813 27711 16871 27717
rect 16813 27677 16825 27711
rect 16859 27708 16871 27711
rect 17086 27708 17092 27720
rect 16859 27680 17092 27708
rect 16859 27677 16871 27680
rect 16813 27671 16871 27677
rect 17086 27668 17092 27680
rect 17144 27668 17150 27720
rect 20398 27708 20404 27720
rect 20359 27680 20404 27708
rect 20398 27668 20404 27680
rect 20456 27668 20462 27720
rect 20490 27668 20496 27720
rect 20548 27708 20554 27720
rect 21410 27708 21416 27720
rect 20548 27680 21416 27708
rect 20548 27668 20554 27680
rect 21410 27668 21416 27680
rect 21468 27708 21474 27720
rect 21888 27717 21916 27748
rect 24814 27736 24820 27748
rect 24872 27776 24878 27788
rect 27025 27779 27083 27785
rect 24872 27748 26884 27776
rect 24872 27736 24878 27748
rect 21781 27711 21839 27717
rect 21781 27708 21793 27711
rect 21468 27680 21793 27708
rect 21468 27668 21474 27680
rect 21781 27677 21793 27680
rect 21827 27677 21839 27711
rect 21781 27671 21839 27677
rect 21873 27711 21931 27717
rect 21873 27677 21885 27711
rect 21919 27677 21931 27711
rect 21873 27671 21931 27677
rect 22241 27711 22299 27717
rect 22241 27677 22253 27711
rect 22287 27708 22299 27711
rect 22606 27708 22612 27720
rect 22287 27680 22612 27708
rect 22287 27677 22299 27680
rect 22241 27671 22299 27677
rect 14513 27643 14571 27649
rect 14513 27609 14525 27643
rect 14559 27609 14571 27643
rect 14694 27640 14700 27652
rect 14655 27612 14700 27640
rect 14513 27603 14571 27609
rect 14528 27572 14556 27603
rect 14694 27600 14700 27612
rect 14752 27600 14758 27652
rect 14973 27643 15031 27649
rect 14973 27609 14985 27643
rect 15019 27640 15031 27643
rect 15062 27640 15068 27652
rect 15019 27612 15068 27640
rect 15019 27609 15031 27612
rect 14973 27603 15031 27609
rect 15062 27600 15068 27612
rect 15120 27640 15126 27652
rect 15120 27612 16856 27640
rect 15120 27600 15126 27612
rect 14602 27572 14608 27584
rect 14528 27544 14608 27572
rect 14602 27532 14608 27544
rect 14660 27532 14666 27584
rect 15338 27572 15344 27584
rect 15299 27544 15344 27572
rect 15338 27532 15344 27544
rect 15396 27532 15402 27584
rect 15433 27575 15491 27581
rect 15433 27541 15445 27575
rect 15479 27572 15491 27575
rect 15522 27572 15528 27584
rect 15479 27544 15528 27572
rect 15479 27541 15491 27544
rect 15433 27535 15491 27541
rect 15522 27532 15528 27544
rect 15580 27532 15586 27584
rect 16828 27572 16856 27612
rect 16902 27600 16908 27652
rect 16960 27640 16966 27652
rect 17273 27643 17331 27649
rect 17273 27640 17285 27643
rect 16960 27612 17285 27640
rect 16960 27600 16966 27612
rect 17273 27609 17285 27612
rect 17319 27609 17331 27643
rect 17546 27640 17552 27652
rect 17507 27612 17552 27640
rect 17273 27603 17331 27609
rect 17546 27600 17552 27612
rect 17604 27600 17610 27652
rect 17638 27600 17644 27652
rect 17696 27640 17702 27652
rect 18098 27640 18104 27652
rect 17696 27612 17789 27640
rect 18059 27612 18104 27640
rect 17696 27600 17702 27612
rect 18098 27600 18104 27612
rect 18156 27640 18162 27652
rect 18466 27640 18472 27652
rect 18156 27612 18472 27640
rect 18156 27600 18162 27612
rect 18466 27600 18472 27612
rect 18524 27600 18530 27652
rect 20306 27600 20312 27652
rect 20364 27640 20370 27652
rect 20582 27640 20588 27652
rect 20364 27612 20588 27640
rect 20364 27600 20370 27612
rect 20582 27600 20588 27612
rect 20640 27600 20646 27652
rect 21686 27640 21692 27652
rect 21647 27612 21692 27640
rect 21686 27600 21692 27612
rect 21744 27600 21750 27652
rect 21796 27640 21824 27671
rect 22606 27668 22612 27680
rect 22664 27668 22670 27720
rect 22790 27668 22796 27720
rect 22848 27708 22854 27720
rect 22885 27711 22943 27717
rect 22885 27708 22897 27711
rect 22848 27680 22897 27708
rect 22848 27668 22854 27680
rect 22885 27677 22897 27680
rect 22931 27677 22943 27711
rect 23066 27708 23072 27720
rect 23027 27680 23072 27708
rect 22885 27671 22943 27677
rect 23066 27668 23072 27680
rect 23124 27668 23130 27720
rect 24081 27711 24139 27717
rect 24081 27677 24093 27711
rect 24127 27708 24139 27711
rect 24538 27708 24544 27720
rect 24127 27680 24544 27708
rect 24127 27677 24139 27680
rect 24081 27671 24139 27677
rect 24538 27668 24544 27680
rect 24596 27668 24602 27720
rect 24633 27711 24691 27717
rect 24633 27677 24645 27711
rect 24679 27708 24691 27711
rect 26381 27711 26439 27717
rect 24679 27680 25596 27708
rect 24679 27677 24691 27680
rect 24633 27671 24691 27677
rect 25568 27652 25596 27680
rect 26381 27677 26393 27711
rect 26427 27708 26439 27711
rect 26562 27708 26568 27720
rect 26427 27680 26568 27708
rect 26427 27677 26439 27680
rect 26381 27671 26439 27677
rect 26562 27668 26568 27680
rect 26620 27668 26626 27720
rect 22977 27643 23035 27649
rect 22977 27640 22989 27643
rect 21796 27612 22989 27640
rect 22977 27609 22989 27612
rect 23023 27609 23035 27643
rect 22977 27603 23035 27609
rect 24265 27643 24323 27649
rect 24265 27609 24277 27643
rect 24311 27640 24323 27643
rect 24446 27640 24452 27652
rect 24311 27612 24452 27640
rect 24311 27609 24323 27612
rect 24265 27603 24323 27609
rect 24446 27600 24452 27612
rect 24504 27600 24510 27652
rect 25366 27640 25372 27652
rect 25327 27612 25372 27640
rect 25366 27600 25372 27612
rect 25424 27600 25430 27652
rect 25550 27640 25556 27652
rect 25511 27612 25556 27640
rect 25550 27600 25556 27612
rect 25608 27600 25614 27652
rect 17656 27572 17684 27600
rect 18190 27572 18196 27584
rect 16828 27544 17684 27572
rect 18103 27544 18196 27572
rect 18190 27532 18196 27544
rect 18248 27532 18254 27584
rect 19938 27532 19944 27584
rect 19996 27572 20002 27584
rect 20033 27575 20091 27581
rect 20033 27572 20045 27575
rect 19996 27544 20045 27572
rect 19996 27532 20002 27544
rect 20033 27541 20045 27544
rect 20079 27541 20091 27575
rect 20033 27535 20091 27541
rect 20769 27575 20827 27581
rect 20769 27541 20781 27575
rect 20815 27572 20827 27575
rect 20950 27572 20956 27584
rect 20815 27544 20956 27572
rect 20815 27541 20827 27544
rect 20769 27535 20827 27541
rect 20950 27532 20956 27544
rect 21008 27532 21014 27584
rect 21502 27572 21508 27584
rect 21463 27544 21508 27572
rect 21502 27532 21508 27544
rect 21560 27572 21566 27584
rect 22701 27575 22759 27581
rect 22701 27572 22713 27575
rect 21560 27544 22713 27572
rect 21560 27532 21566 27544
rect 22701 27541 22713 27544
rect 22747 27541 22759 27575
rect 22701 27535 22759 27541
rect 23437 27575 23495 27581
rect 23437 27541 23449 27575
rect 23483 27572 23495 27575
rect 23526 27572 23532 27584
rect 23483 27544 23532 27572
rect 23483 27541 23495 27544
rect 23437 27535 23495 27541
rect 23526 27532 23532 27544
rect 23584 27572 23590 27584
rect 25642 27572 25648 27584
rect 23584 27544 25648 27572
rect 23584 27532 23590 27544
rect 25642 27532 25648 27544
rect 25700 27532 25706 27584
rect 25921 27575 25979 27581
rect 25921 27541 25933 27575
rect 25967 27572 25979 27575
rect 26286 27572 26292 27584
rect 25967 27544 26292 27572
rect 25967 27541 25979 27544
rect 25921 27535 25979 27541
rect 26286 27532 26292 27544
rect 26344 27532 26350 27584
rect 26470 27532 26476 27584
rect 26528 27572 26534 27584
rect 26749 27575 26807 27581
rect 26749 27572 26761 27575
rect 26528 27544 26761 27572
rect 26528 27532 26534 27544
rect 26749 27541 26761 27544
rect 26795 27541 26807 27575
rect 26856 27572 26884 27748
rect 27025 27745 27037 27779
rect 27071 27776 27083 27779
rect 30886 27776 30892 27788
rect 27071 27748 30892 27776
rect 27071 27745 27083 27748
rect 27025 27739 27083 27745
rect 30886 27736 30892 27748
rect 30944 27736 30950 27788
rect 29233 27711 29291 27717
rect 29233 27708 29245 27711
rect 28236 27680 29245 27708
rect 27850 27600 27856 27652
rect 27908 27640 27914 27652
rect 28236 27649 28264 27680
rect 29233 27677 29245 27680
rect 29279 27677 29291 27711
rect 29233 27671 29291 27677
rect 28221 27643 28279 27649
rect 28221 27640 28233 27643
rect 27908 27612 28233 27640
rect 27908 27600 27914 27612
rect 28221 27609 28233 27612
rect 28267 27609 28279 27643
rect 28221 27603 28279 27609
rect 28405 27643 28463 27649
rect 28405 27609 28417 27643
rect 28451 27640 28463 27643
rect 28494 27640 28500 27652
rect 28451 27612 28500 27640
rect 28451 27609 28463 27612
rect 28405 27603 28463 27609
rect 28494 27600 28500 27612
rect 28552 27600 28558 27652
rect 28589 27643 28647 27649
rect 28589 27609 28601 27643
rect 28635 27609 28647 27643
rect 28589 27603 28647 27609
rect 29417 27643 29475 27649
rect 29417 27609 29429 27643
rect 29463 27609 29475 27643
rect 29417 27603 29475 27609
rect 28604 27572 28632 27603
rect 26856 27544 28632 27572
rect 26749 27535 26807 27541
rect 15540 27504 15568 27532
rect 18208 27504 18236 27532
rect 15540 27476 18236 27504
rect 26657 27507 26715 27513
rect 26657 27473 26669 27507
rect 26703 27504 26715 27507
rect 27850 27504 27856 27516
rect 26703 27476 27856 27504
rect 26703 27473 26715 27476
rect 26657 27467 26715 27473
rect 27850 27464 27856 27476
rect 27908 27464 27914 27516
rect 28037 27507 28095 27513
rect 28037 27473 28049 27507
rect 28083 27504 28095 27507
rect 28586 27504 28592 27516
rect 28083 27476 28592 27504
rect 28083 27473 28095 27476
rect 28037 27467 28095 27473
rect 28586 27464 28592 27476
rect 28644 27464 28650 27516
rect 21686 27396 21692 27448
rect 21744 27436 21750 27448
rect 22790 27436 22796 27448
rect 21744 27408 22796 27436
rect 21744 27396 21750 27408
rect 22790 27396 22796 27408
rect 22848 27396 22854 27448
rect 25366 27396 25372 27448
rect 25424 27436 25430 27448
rect 26519 27439 26577 27445
rect 26519 27436 26531 27439
rect 25424 27408 26531 27436
rect 25424 27396 25430 27408
rect 26519 27405 26531 27408
rect 26565 27436 26577 27439
rect 27298 27436 27304 27448
rect 26565 27408 27304 27436
rect 26565 27405 26577 27408
rect 26519 27399 26577 27405
rect 27298 27396 27304 27408
rect 27356 27396 27362 27448
rect 28494 27396 28500 27448
rect 28552 27436 28558 27448
rect 29432 27436 29460 27603
rect 29785 27575 29843 27581
rect 29785 27541 29797 27575
rect 29831 27572 29843 27575
rect 30334 27572 30340 27584
rect 29831 27544 30340 27572
rect 29831 27541 29843 27544
rect 29785 27535 29843 27541
rect 30334 27532 30340 27544
rect 30392 27532 30398 27584
rect 28552 27408 29460 27436
rect 28552 27396 28558 27408
rect 11000 27346 34368 27368
rect 11000 27294 14142 27346
rect 14194 27294 14206 27346
rect 14258 27294 14270 27346
rect 14322 27294 14334 27346
rect 14386 27294 24142 27346
rect 24194 27294 24206 27346
rect 24258 27294 24270 27346
rect 24322 27294 24334 27346
rect 24386 27294 34368 27346
rect 11000 27272 34368 27294
rect 22422 27192 22428 27244
rect 22480 27232 22486 27244
rect 23434 27232 23440 27244
rect 22480 27204 23440 27232
rect 22480 27192 22486 27204
rect 23434 27192 23440 27204
rect 23492 27192 23498 27244
rect 25458 27192 25464 27244
rect 25516 27232 25522 27244
rect 26013 27235 26071 27241
rect 26013 27232 26025 27235
rect 25516 27204 26025 27232
rect 25516 27192 25522 27204
rect 26013 27201 26025 27204
rect 26059 27201 26071 27235
rect 26013 27195 26071 27201
rect 26381 27235 26439 27241
rect 26381 27201 26393 27235
rect 26427 27232 26439 27235
rect 26654 27232 26660 27244
rect 26427 27204 26660 27232
rect 26427 27201 26439 27204
rect 26381 27195 26439 27201
rect 26654 27192 26660 27204
rect 26712 27192 26718 27244
rect 17546 27164 17552 27176
rect 17380 27136 17552 27164
rect 14605 27099 14663 27105
rect 14605 27065 14617 27099
rect 14651 27096 14663 27099
rect 14694 27096 14700 27108
rect 14651 27068 14700 27096
rect 14651 27065 14663 27068
rect 14605 27059 14663 27065
rect 14694 27056 14700 27068
rect 14752 27056 14758 27108
rect 16813 27099 16871 27105
rect 16813 27065 16825 27099
rect 16859 27096 16871 27099
rect 16994 27096 17000 27108
rect 16859 27068 17000 27096
rect 16859 27065 16871 27068
rect 16813 27059 16871 27065
rect 16994 27056 17000 27068
rect 17052 27056 17058 27108
rect 17380 27105 17408 27136
rect 17546 27124 17552 27136
rect 17604 27164 17610 27176
rect 18377 27167 18435 27173
rect 18377 27164 18389 27167
rect 17604 27136 18389 27164
rect 17604 27124 17610 27136
rect 18377 27133 18389 27136
rect 18423 27133 18435 27167
rect 18377 27127 18435 27133
rect 17365 27099 17423 27105
rect 17365 27065 17377 27099
rect 17411 27065 17423 27099
rect 17365 27059 17423 27065
rect 17825 27099 17883 27105
rect 17825 27065 17837 27099
rect 17871 27096 17883 27099
rect 18006 27096 18012 27108
rect 17871 27068 18012 27096
rect 17871 27065 17883 27068
rect 17825 27059 17883 27065
rect 18006 27056 18012 27068
rect 18064 27056 18070 27108
rect 21226 27056 21232 27108
rect 21284 27096 21290 27108
rect 23161 27099 23219 27105
rect 23161 27096 23173 27099
rect 21284 27068 23173 27096
rect 21284 27056 21290 27068
rect 23161 27065 23173 27068
rect 23207 27065 23219 27099
rect 23161 27059 23219 27065
rect 14510 27028 14516 27040
rect 14471 27000 14516 27028
rect 14510 26988 14516 27000
rect 14568 26988 14574 27040
rect 14970 27028 14976 27040
rect 14931 27000 14976 27028
rect 14970 26988 14976 27000
rect 15028 26988 15034 27040
rect 16077 27031 16135 27037
rect 16077 26997 16089 27031
rect 16123 26997 16135 27031
rect 16077 26991 16135 26997
rect 16169 27031 16227 27037
rect 16169 26997 16181 27031
rect 16215 27028 16227 27031
rect 17270 27028 17276 27040
rect 16215 27000 17276 27028
rect 16215 26997 16227 27000
rect 16169 26991 16227 26997
rect 16092 26892 16120 26991
rect 17270 26988 17276 27000
rect 17328 26988 17334 27040
rect 17638 27028 17644 27040
rect 17599 27000 17644 27028
rect 17638 26988 17644 27000
rect 17696 26988 17702 27040
rect 17914 26988 17920 27040
rect 17972 27028 17978 27040
rect 18285 27031 18343 27037
rect 18285 27028 18297 27031
rect 17972 27000 18297 27028
rect 17972 26988 17978 27000
rect 18285 26997 18297 27000
rect 18331 26997 18343 27031
rect 18285 26991 18343 26997
rect 18837 27031 18895 27037
rect 18837 26997 18849 27031
rect 18883 26997 18895 27031
rect 20950 27028 20956 27040
rect 20911 27000 20956 27028
rect 18837 26991 18895 26997
rect 16626 26920 16632 26972
rect 16684 26960 16690 26972
rect 18852 26960 18880 26991
rect 20950 26988 20956 27000
rect 21008 26988 21014 27040
rect 21318 27028 21324 27040
rect 21279 27000 21324 27028
rect 21318 26988 21324 27000
rect 21376 26988 21382 27040
rect 22606 26988 22612 27040
rect 22664 27028 22670 27040
rect 22701 27031 22759 27037
rect 22701 27028 22713 27031
rect 22664 27000 22713 27028
rect 22664 26988 22670 27000
rect 22701 26997 22713 27000
rect 22747 26997 22759 27031
rect 23176 27028 23204 27059
rect 23802 27056 23808 27108
rect 23860 27096 23866 27108
rect 24081 27099 24139 27105
rect 24081 27096 24093 27099
rect 23860 27068 24093 27096
rect 23860 27056 23866 27068
rect 24081 27065 24093 27068
rect 24127 27065 24139 27099
rect 26102 27096 26108 27108
rect 26063 27068 26108 27096
rect 24081 27059 24139 27065
rect 26102 27056 26108 27068
rect 26160 27056 26166 27108
rect 29782 27096 29788 27108
rect 29708 27068 29788 27096
rect 23250 27028 23256 27040
rect 23163 27000 23256 27028
rect 22701 26991 22759 26997
rect 23250 26988 23256 27000
rect 23308 27028 23314 27040
rect 23989 27031 24047 27037
rect 23989 27028 24001 27031
rect 23308 27000 24001 27028
rect 23308 26988 23314 27000
rect 23989 26997 24001 27000
rect 24035 26997 24047 27031
rect 23989 26991 24047 26997
rect 24265 27031 24323 27037
rect 24265 26997 24277 27031
rect 24311 26997 24323 27031
rect 24265 26991 24323 26997
rect 24725 27031 24783 27037
rect 24725 26997 24737 27031
rect 24771 27028 24783 27031
rect 25884 27031 25942 27037
rect 25884 27028 25896 27031
rect 24771 27000 25896 27028
rect 24771 26997 24783 27000
rect 24725 26991 24783 26997
rect 25884 26997 25896 27000
rect 25930 26997 25942 27031
rect 25884 26991 25942 26997
rect 28221 27031 28279 27037
rect 28221 26997 28233 27031
rect 28267 26997 28279 27031
rect 28221 26991 28279 26997
rect 16684 26932 18880 26960
rect 20769 26963 20827 26969
rect 16684 26920 16690 26932
rect 20769 26929 20781 26963
rect 20815 26960 20827 26963
rect 21778 26960 21784 26972
rect 20815 26932 21784 26960
rect 20815 26929 20827 26932
rect 20769 26923 20827 26929
rect 21778 26920 21784 26932
rect 21836 26920 21842 26972
rect 22422 26960 22428 26972
rect 22383 26932 22428 26960
rect 22422 26920 22428 26932
rect 22480 26920 22486 26972
rect 22793 26963 22851 26969
rect 22793 26929 22805 26963
rect 22839 26960 22851 26963
rect 22974 26960 22980 26972
rect 22839 26932 22980 26960
rect 22839 26929 22851 26932
rect 22793 26923 22851 26929
rect 22974 26920 22980 26932
rect 23032 26920 23038 26972
rect 23434 26920 23440 26972
rect 23492 26960 23498 26972
rect 24280 26960 24308 26991
rect 23492 26932 24308 26960
rect 23492 26920 23498 26932
rect 17086 26892 17092 26904
rect 16092 26864 17092 26892
rect 17086 26852 17092 26864
rect 17144 26852 17150 26904
rect 20214 26852 20220 26904
rect 20272 26892 20278 26904
rect 21962 26892 21968 26904
rect 20272 26864 21968 26892
rect 20272 26852 20278 26864
rect 21962 26852 21968 26864
rect 22020 26892 22026 26904
rect 22609 26895 22667 26901
rect 22609 26892 22621 26895
rect 22020 26864 22621 26892
rect 22020 26852 22026 26864
rect 22609 26861 22621 26864
rect 22655 26861 22667 26895
rect 24280 26892 24308 26932
rect 25642 26920 25648 26972
rect 25700 26960 25706 26972
rect 25737 26963 25795 26969
rect 25737 26960 25749 26963
rect 25700 26932 25749 26960
rect 25700 26920 25706 26932
rect 25737 26929 25749 26932
rect 25783 26929 25795 26963
rect 28236 26960 28264 26991
rect 29598 26988 29604 27040
rect 29656 27028 29662 27040
rect 29708 27037 29736 27068
rect 29782 27056 29788 27068
rect 29840 27056 29846 27108
rect 30334 27096 30340 27108
rect 30295 27068 30340 27096
rect 30334 27056 30340 27068
rect 30392 27056 30398 27108
rect 31254 27096 31260 27108
rect 31215 27068 31260 27096
rect 31254 27056 31260 27068
rect 31312 27056 31318 27108
rect 29693 27031 29751 27037
rect 29693 27028 29705 27031
rect 29656 27000 29705 27028
rect 29656 26988 29662 27000
rect 29693 26997 29705 27000
rect 29739 26997 29751 27031
rect 29693 26991 29751 26997
rect 31165 27031 31223 27037
rect 31165 26997 31177 27031
rect 31211 26997 31223 27031
rect 31165 26991 31223 26997
rect 29506 26960 29512 26972
rect 28236 26932 29512 26960
rect 25737 26923 25795 26929
rect 29506 26920 29512 26932
rect 29564 26920 29570 26972
rect 29782 26960 29788 26972
rect 29743 26932 29788 26960
rect 29782 26920 29788 26932
rect 29840 26920 29846 26972
rect 29874 26920 29880 26972
rect 29932 26960 29938 26972
rect 30429 26963 30487 26969
rect 30429 26960 30441 26963
rect 29932 26932 30441 26960
rect 29932 26920 29938 26932
rect 30429 26929 30441 26932
rect 30475 26929 30487 26963
rect 30429 26923 30487 26929
rect 25918 26892 25924 26904
rect 24280 26864 25924 26892
rect 22609 26855 22667 26861
rect 25918 26852 25924 26864
rect 25976 26852 25982 26904
rect 28954 26852 28960 26904
rect 29012 26892 29018 26904
rect 31180 26892 31208 26991
rect 29012 26864 31208 26892
rect 29012 26852 29018 26864
rect 11000 26802 34368 26824
rect 11000 26750 19142 26802
rect 19194 26750 19206 26802
rect 19258 26750 19270 26802
rect 19322 26750 19334 26802
rect 19386 26750 29142 26802
rect 29194 26750 29206 26802
rect 29258 26750 29270 26802
rect 29322 26750 29334 26802
rect 29386 26750 34368 26802
rect 11000 26728 34368 26750
rect 17365 26691 17423 26697
rect 17365 26657 17377 26691
rect 17411 26688 17423 26691
rect 17546 26688 17552 26700
rect 17411 26660 17552 26688
rect 17411 26657 17423 26660
rect 17365 26651 17423 26657
rect 17546 26648 17552 26660
rect 17604 26688 17610 26700
rect 17914 26688 17920 26700
rect 17604 26660 17920 26688
rect 17604 26648 17610 26660
rect 17914 26648 17920 26660
rect 17972 26648 17978 26700
rect 20398 26648 20404 26700
rect 20456 26688 20462 26700
rect 22606 26688 22612 26700
rect 20456 26660 22612 26688
rect 20456 26648 20462 26660
rect 22606 26648 22612 26660
rect 22664 26648 22670 26700
rect 24998 26648 25004 26700
rect 25056 26688 25062 26700
rect 27574 26688 27580 26700
rect 25056 26660 27580 26688
rect 25056 26648 25062 26660
rect 27574 26648 27580 26660
rect 27632 26648 27638 26700
rect 27850 26648 27856 26700
rect 27908 26688 27914 26700
rect 28773 26691 28831 26697
rect 28773 26688 28785 26691
rect 27908 26660 28785 26688
rect 27908 26648 27914 26660
rect 28773 26657 28785 26660
rect 28819 26657 28831 26691
rect 28773 26651 28831 26657
rect 14510 26580 14516 26632
rect 14568 26620 14574 26632
rect 14605 26623 14663 26629
rect 14605 26620 14617 26623
rect 14568 26592 14617 26620
rect 14568 26580 14574 26592
rect 14605 26589 14617 26592
rect 14651 26589 14663 26623
rect 17638 26620 17644 26632
rect 14605 26583 14663 26589
rect 15264 26592 17644 26620
rect 15264 26561 15292 26592
rect 17638 26580 17644 26592
rect 17696 26620 17702 26632
rect 19938 26620 19944 26632
rect 17696 26592 18144 26620
rect 17696 26580 17702 26592
rect 15249 26555 15307 26561
rect 15249 26521 15261 26555
rect 15295 26521 15307 26555
rect 15249 26515 15307 26521
rect 15617 26555 15675 26561
rect 15617 26521 15629 26555
rect 15663 26552 15675 26555
rect 17733 26555 17791 26561
rect 17733 26552 17745 26555
rect 15663 26524 17745 26552
rect 15663 26521 15675 26524
rect 15617 26515 15675 26521
rect 17733 26521 17745 26524
rect 17779 26552 17791 26555
rect 17822 26552 17828 26564
rect 17779 26524 17828 26552
rect 17779 26521 17791 26524
rect 17733 26515 17791 26521
rect 17822 26512 17828 26524
rect 17880 26512 17886 26564
rect 18116 26561 18144 26592
rect 19588 26592 19944 26620
rect 19588 26564 19616 26592
rect 19938 26580 19944 26592
rect 19996 26620 20002 26632
rect 22333 26623 22391 26629
rect 22333 26620 22345 26623
rect 19996 26592 22345 26620
rect 19996 26580 20002 26592
rect 22333 26589 22345 26592
rect 22379 26620 22391 26623
rect 22422 26620 22428 26632
rect 22379 26592 22428 26620
rect 22379 26589 22391 26592
rect 22333 26583 22391 26589
rect 22422 26580 22428 26592
rect 22480 26580 22486 26632
rect 22701 26623 22759 26629
rect 22701 26589 22713 26623
rect 22747 26620 22759 26623
rect 23066 26620 23072 26632
rect 22747 26592 23072 26620
rect 22747 26589 22759 26592
rect 22701 26583 22759 26589
rect 23066 26580 23072 26592
rect 23124 26580 23130 26632
rect 23529 26623 23587 26629
rect 23529 26589 23541 26623
rect 23575 26620 23587 26623
rect 23618 26620 23624 26632
rect 23575 26592 23624 26620
rect 23575 26589 23587 26592
rect 23529 26583 23587 26589
rect 23618 26580 23624 26592
rect 23676 26580 23682 26632
rect 26105 26623 26163 26629
rect 26105 26589 26117 26623
rect 26151 26620 26163 26623
rect 26286 26620 26292 26632
rect 26151 26592 26292 26620
rect 26151 26589 26163 26592
rect 26105 26583 26163 26589
rect 26286 26580 26292 26592
rect 26344 26580 26350 26632
rect 26841 26623 26899 26629
rect 26841 26589 26853 26623
rect 26887 26620 26899 26623
rect 27022 26620 27028 26632
rect 26887 26592 27028 26620
rect 26887 26589 26899 26592
rect 26841 26583 26899 26589
rect 27022 26580 27028 26592
rect 27080 26580 27086 26632
rect 28497 26623 28555 26629
rect 28497 26620 28509 26623
rect 27132 26592 28509 26620
rect 18101 26555 18159 26561
rect 18101 26521 18113 26555
rect 18147 26521 18159 26555
rect 19570 26552 19576 26564
rect 19531 26524 19576 26552
rect 18101 26515 18159 26521
rect 19570 26512 19576 26524
rect 19628 26512 19634 26564
rect 20214 26552 20220 26564
rect 20175 26524 20220 26552
rect 20214 26512 20220 26524
rect 20272 26512 20278 26564
rect 20398 26552 20404 26564
rect 20359 26524 20404 26552
rect 20398 26512 20404 26524
rect 20456 26512 20462 26564
rect 20490 26512 20496 26564
rect 20548 26552 20554 26564
rect 20769 26555 20827 26561
rect 20769 26552 20781 26555
rect 20548 26524 20781 26552
rect 20548 26512 20554 26524
rect 20769 26521 20781 26524
rect 20815 26521 20827 26555
rect 20769 26515 20827 26521
rect 21686 26512 21692 26564
rect 21744 26552 21750 26564
rect 22238 26552 22244 26564
rect 21744 26524 22244 26552
rect 21744 26512 21750 26524
rect 22238 26512 22244 26524
rect 22296 26552 22302 26564
rect 22517 26555 22575 26561
rect 22517 26552 22529 26555
rect 22296 26524 22529 26552
rect 22296 26512 22302 26524
rect 22517 26521 22529 26524
rect 22563 26521 22575 26555
rect 22517 26515 22575 26521
rect 23342 26512 23348 26564
rect 23400 26552 23406 26564
rect 27132 26552 27160 26592
rect 28497 26589 28509 26592
rect 28543 26589 28555 26623
rect 28497 26583 28555 26589
rect 29782 26580 29788 26632
rect 29840 26620 29846 26632
rect 29969 26623 30027 26629
rect 29969 26620 29981 26623
rect 29840 26592 29981 26620
rect 29840 26580 29846 26592
rect 29969 26589 29981 26592
rect 30015 26589 30027 26623
rect 29969 26583 30027 26589
rect 27298 26552 27304 26564
rect 23400 26524 27160 26552
rect 27259 26524 27304 26552
rect 23400 26512 23406 26524
rect 27298 26512 27304 26524
rect 27356 26512 27362 26564
rect 28681 26555 28739 26561
rect 28681 26552 28693 26555
rect 27776 26524 28693 26552
rect 15341 26487 15399 26493
rect 15341 26453 15353 26487
rect 15387 26453 15399 26487
rect 15341 26447 15399 26453
rect 15356 26416 15384 26447
rect 15430 26444 15436 26496
rect 15488 26484 15494 26496
rect 15525 26487 15583 26493
rect 15525 26484 15537 26487
rect 15488 26456 15537 26484
rect 15488 26444 15494 26456
rect 15525 26453 15537 26456
rect 15571 26453 15583 26487
rect 15525 26447 15583 26453
rect 17641 26487 17699 26493
rect 17641 26453 17653 26487
rect 17687 26453 17699 26487
rect 18006 26484 18012 26496
rect 17919 26456 18012 26484
rect 17641 26447 17699 26453
rect 17656 26416 17684 26447
rect 18006 26444 18012 26456
rect 18064 26484 18070 26496
rect 19662 26484 19668 26496
rect 18064 26456 19668 26484
rect 18064 26444 18070 26456
rect 19662 26444 19668 26456
rect 19720 26484 19726 26496
rect 20232 26484 20260 26512
rect 19720 26456 20260 26484
rect 23069 26487 23127 26493
rect 19720 26444 19726 26456
rect 23069 26453 23081 26487
rect 23115 26484 23127 26487
rect 23676 26487 23734 26493
rect 23676 26484 23688 26487
rect 23115 26456 23688 26484
rect 23115 26453 23127 26456
rect 23069 26447 23127 26453
rect 23676 26453 23688 26456
rect 23722 26453 23734 26487
rect 23676 26447 23734 26453
rect 23897 26487 23955 26493
rect 23897 26453 23909 26487
rect 23943 26453 23955 26487
rect 23897 26447 23955 26453
rect 24265 26487 24323 26493
rect 24265 26453 24277 26487
rect 24311 26484 24323 26487
rect 26252 26487 26310 26493
rect 26252 26484 26264 26487
rect 24311 26456 26264 26484
rect 24311 26453 24323 26456
rect 24265 26447 24323 26453
rect 26252 26453 26264 26456
rect 26298 26453 26310 26487
rect 26470 26484 26476 26496
rect 26431 26456 26476 26484
rect 26252 26447 26310 26453
rect 18098 26416 18104 26428
rect 15356 26388 15476 26416
rect 17656 26388 18104 26416
rect 15448 26348 15476 26388
rect 18098 26376 18104 26388
rect 18156 26416 18162 26428
rect 18466 26416 18472 26428
rect 18156 26388 18472 26416
rect 18156 26376 18162 26388
rect 18466 26376 18472 26388
rect 18524 26376 18530 26428
rect 20953 26419 21011 26425
rect 20953 26385 20965 26419
rect 20999 26416 21011 26419
rect 22606 26416 22612 26428
rect 20999 26388 22612 26416
rect 20999 26385 21011 26388
rect 20953 26379 21011 26385
rect 22606 26376 22612 26388
rect 22664 26416 22670 26428
rect 23912 26416 23940 26447
rect 26470 26444 26476 26456
rect 26528 26484 26534 26496
rect 27669 26487 27727 26493
rect 27669 26484 27681 26487
rect 26528 26456 27681 26484
rect 26528 26444 26534 26456
rect 27669 26453 27681 26456
rect 27715 26453 27727 26487
rect 27669 26447 27727 26453
rect 22664 26388 23940 26416
rect 22664 26376 22670 26388
rect 23986 26376 23992 26428
rect 24044 26416 24050 26428
rect 27439 26419 27497 26425
rect 27439 26416 27451 26419
rect 24044 26388 27451 26416
rect 24044 26376 24050 26388
rect 27439 26385 27451 26388
rect 27485 26385 27497 26419
rect 27574 26416 27580 26428
rect 27535 26388 27580 26416
rect 27439 26379 27497 26385
rect 27574 26376 27580 26388
rect 27632 26376 27638 26428
rect 19846 26348 19852 26360
rect 15448 26320 19852 26348
rect 19846 26308 19852 26320
rect 19904 26308 19910 26360
rect 23250 26308 23256 26360
rect 23308 26348 23314 26360
rect 23805 26351 23863 26357
rect 23805 26348 23817 26351
rect 23308 26320 23817 26348
rect 23308 26308 23314 26320
rect 23805 26317 23817 26320
rect 23851 26317 23863 26351
rect 23805 26311 23863 26317
rect 25642 26308 25648 26360
rect 25700 26348 25706 26360
rect 26381 26351 26439 26357
rect 26381 26348 26393 26351
rect 25700 26320 26393 26348
rect 25700 26308 25706 26320
rect 26381 26317 26393 26320
rect 26427 26317 26439 26351
rect 26381 26311 26439 26317
rect 26746 26308 26752 26360
rect 26804 26348 26810 26360
rect 27776 26348 27804 26524
rect 28681 26521 28693 26524
rect 28727 26521 28739 26555
rect 29506 26552 29512 26564
rect 29467 26524 29512 26552
rect 28681 26515 28739 26521
rect 29506 26512 29512 26524
rect 29564 26512 29570 26564
rect 29598 26512 29604 26564
rect 29656 26552 29662 26564
rect 30981 26555 31039 26561
rect 30981 26552 30993 26555
rect 29656 26524 30993 26552
rect 29656 26512 29662 26524
rect 30981 26521 30993 26524
rect 31027 26521 31039 26555
rect 31438 26552 31444 26564
rect 31399 26524 31444 26552
rect 30981 26515 31039 26521
rect 31438 26512 31444 26524
rect 31496 26512 31502 26564
rect 30061 26487 30119 26493
rect 30061 26453 30073 26487
rect 30107 26484 30119 26487
rect 31533 26487 31591 26493
rect 31533 26484 31545 26487
rect 30107 26456 31545 26484
rect 30107 26453 30119 26456
rect 30061 26447 30119 26453
rect 31533 26453 31545 26456
rect 31579 26453 31591 26487
rect 31533 26447 31591 26453
rect 26804 26320 27804 26348
rect 27945 26351 28003 26357
rect 26804 26308 26810 26320
rect 27945 26317 27957 26351
rect 27991 26348 28003 26351
rect 28402 26348 28408 26360
rect 27991 26320 28408 26348
rect 27991 26317 28003 26320
rect 27945 26311 28003 26317
rect 28402 26308 28408 26320
rect 28460 26308 28466 26360
rect 30242 26308 30248 26360
rect 30300 26348 30306 26360
rect 30797 26351 30855 26357
rect 30797 26348 30809 26351
rect 30300 26320 30809 26348
rect 30300 26308 30306 26320
rect 30797 26317 30809 26320
rect 30843 26317 30855 26351
rect 30797 26311 30855 26317
rect 11000 26258 34368 26280
rect 11000 26206 14142 26258
rect 14194 26206 14206 26258
rect 14258 26206 14270 26258
rect 14322 26206 14334 26258
rect 14386 26206 24142 26258
rect 24194 26206 24206 26258
rect 24258 26206 24270 26258
rect 24322 26206 24334 26258
rect 24386 26206 34368 26258
rect 11000 26184 34368 26206
rect 14602 26104 14608 26156
rect 14660 26144 14666 26156
rect 14697 26147 14755 26153
rect 14697 26144 14709 26147
rect 14660 26116 14709 26144
rect 14660 26104 14666 26116
rect 14697 26113 14709 26116
rect 14743 26113 14755 26147
rect 22606 26144 22612 26156
rect 22567 26116 22612 26144
rect 14697 26107 14755 26113
rect 22606 26104 22612 26116
rect 22664 26104 22670 26156
rect 22977 26147 23035 26153
rect 22977 26113 22989 26147
rect 23023 26144 23035 26147
rect 23986 26144 23992 26156
rect 23023 26116 23992 26144
rect 23023 26113 23035 26116
rect 22977 26107 23035 26113
rect 23986 26104 23992 26116
rect 24044 26104 24050 26156
rect 25458 26144 25464 26156
rect 24556 26116 25464 26144
rect 21318 26036 21324 26088
rect 21376 26076 21382 26088
rect 24556 26076 24584 26116
rect 25458 26104 25464 26116
rect 25516 26144 25522 26156
rect 25829 26147 25887 26153
rect 25829 26144 25841 26147
rect 25516 26116 25841 26144
rect 25516 26104 25522 26116
rect 25829 26113 25841 26116
rect 25875 26113 25887 26147
rect 25829 26107 25887 26113
rect 21376 26048 24584 26076
rect 21376 26036 21382 26048
rect 25550 26036 25556 26088
rect 25608 26076 25614 26088
rect 25691 26079 25749 26085
rect 25691 26076 25703 26079
rect 25608 26048 25703 26076
rect 25608 26036 25614 26048
rect 25691 26045 25703 26048
rect 25737 26045 25749 26079
rect 25844 26076 25872 26107
rect 26470 26104 26476 26156
rect 26528 26144 26534 26156
rect 27025 26147 27083 26153
rect 27025 26144 27037 26147
rect 26528 26116 27037 26144
rect 26528 26104 26534 26116
rect 27025 26113 27037 26116
rect 27071 26113 27083 26147
rect 27025 26107 27083 26113
rect 30153 26079 30211 26085
rect 30153 26076 30165 26079
rect 25844 26048 26792 26076
rect 25691 26039 25749 26045
rect 14786 26008 14792 26020
rect 13792 25980 14792 26008
rect 13792 25949 13820 25980
rect 14786 25968 14792 25980
rect 14844 25968 14850 26020
rect 16169 26011 16227 26017
rect 16169 25977 16181 26011
rect 16215 26008 16227 26011
rect 16902 26008 16908 26020
rect 16215 25980 16908 26008
rect 16215 25977 16227 25980
rect 16169 25971 16227 25977
rect 16902 25968 16908 25980
rect 16960 25968 16966 26020
rect 17822 26008 17828 26020
rect 17783 25980 17828 26008
rect 17822 25968 17828 25980
rect 17880 25968 17886 26020
rect 19478 26008 19484 26020
rect 18208 25980 19484 26008
rect 13777 25943 13835 25949
rect 13777 25909 13789 25943
rect 13823 25909 13835 25943
rect 13777 25903 13835 25909
rect 14421 25943 14479 25949
rect 14421 25909 14433 25943
rect 14467 25940 14479 25943
rect 14510 25940 14516 25952
rect 14467 25912 14516 25940
rect 14467 25909 14479 25912
rect 14421 25903 14479 25909
rect 14510 25900 14516 25912
rect 14568 25900 14574 25952
rect 14605 25943 14663 25949
rect 14605 25909 14617 25943
rect 14651 25940 14663 25943
rect 14970 25940 14976 25952
rect 14651 25912 14976 25940
rect 14651 25909 14663 25912
rect 14605 25903 14663 25909
rect 14970 25900 14976 25912
rect 15028 25940 15034 25952
rect 15801 25943 15859 25949
rect 15028 25912 15752 25940
rect 15028 25900 15034 25912
rect 15617 25875 15675 25881
rect 15617 25841 15629 25875
rect 15663 25841 15675 25875
rect 15724 25872 15752 25912
rect 15801 25909 15813 25943
rect 15847 25940 15859 25943
rect 16626 25940 16632 25952
rect 15847 25912 16632 25940
rect 15847 25909 15859 25912
rect 15801 25903 15859 25909
rect 16626 25900 16632 25912
rect 16684 25940 16690 25952
rect 17181 25943 17239 25949
rect 17181 25940 17193 25943
rect 16684 25912 17193 25940
rect 16684 25900 16690 25912
rect 17181 25909 17193 25912
rect 17227 25909 17239 25943
rect 17181 25903 17239 25909
rect 17270 25900 17276 25952
rect 17328 25940 17334 25952
rect 17365 25943 17423 25949
rect 17365 25940 17377 25943
rect 17328 25912 17377 25940
rect 17328 25900 17334 25912
rect 17365 25909 17377 25912
rect 17411 25909 17423 25943
rect 17546 25940 17552 25952
rect 17507 25912 17552 25940
rect 17365 25903 17423 25909
rect 17546 25900 17552 25912
rect 17604 25900 17610 25952
rect 18208 25949 18236 25980
rect 19478 25968 19484 25980
rect 19536 26008 19542 26020
rect 19536 25980 19892 26008
rect 19536 25968 19542 25980
rect 19864 25949 19892 25980
rect 20306 25968 20312 26020
rect 20364 26008 20370 26020
rect 22698 26008 22704 26020
rect 20364 25980 20996 26008
rect 22659 25980 22704 26008
rect 20364 25968 20370 25980
rect 20968 25952 20996 25980
rect 22698 25968 22704 25980
rect 22756 25968 22762 26020
rect 24449 26011 24507 26017
rect 24449 25977 24461 26011
rect 24495 26008 24507 26011
rect 25182 26008 25188 26020
rect 24495 25980 25188 26008
rect 24495 25977 24507 25980
rect 24449 25971 24507 25977
rect 25182 25968 25188 25980
rect 25240 26008 25246 26020
rect 25568 26008 25596 26036
rect 25240 25980 25596 26008
rect 25921 26011 25979 26017
rect 25240 25968 25246 25980
rect 25921 25977 25933 26011
rect 25967 26008 25979 26011
rect 26102 26008 26108 26020
rect 25967 25980 26108 26008
rect 25967 25977 25979 25980
rect 25921 25971 25979 25977
rect 26102 25968 26108 25980
rect 26160 25968 26166 26020
rect 18193 25943 18251 25949
rect 18193 25909 18205 25943
rect 18239 25909 18251 25943
rect 18193 25903 18251 25909
rect 19665 25943 19723 25949
rect 19665 25909 19677 25943
rect 19711 25909 19723 25943
rect 19665 25903 19723 25909
rect 19849 25943 19907 25949
rect 19849 25909 19861 25943
rect 19895 25909 19907 25943
rect 19849 25903 19907 25909
rect 20217 25943 20275 25949
rect 20217 25909 20229 25943
rect 20263 25940 20275 25943
rect 20398 25940 20404 25952
rect 20263 25912 20404 25940
rect 20263 25909 20275 25912
rect 20217 25903 20275 25909
rect 16721 25875 16779 25881
rect 16721 25872 16733 25875
rect 15724 25844 16733 25872
rect 15617 25835 15675 25841
rect 16721 25841 16733 25844
rect 16767 25841 16779 25875
rect 16721 25835 16779 25841
rect 13958 25804 13964 25816
rect 13919 25776 13964 25804
rect 13958 25764 13964 25776
rect 14016 25764 14022 25816
rect 15632 25804 15660 25835
rect 17564 25804 17592 25900
rect 19680 25872 19708 25903
rect 20398 25900 20404 25912
rect 20456 25900 20462 25952
rect 20950 25940 20956 25952
rect 20863 25912 20956 25940
rect 20950 25900 20956 25912
rect 21008 25900 21014 25952
rect 21505 25943 21563 25949
rect 21505 25909 21517 25943
rect 21551 25940 21563 25943
rect 21594 25940 21600 25952
rect 21551 25912 21600 25940
rect 21551 25909 21563 25912
rect 21505 25903 21563 25909
rect 21594 25900 21600 25912
rect 21652 25900 21658 25952
rect 21689 25943 21747 25949
rect 21689 25909 21701 25943
rect 21735 25940 21747 25943
rect 22480 25943 22538 25949
rect 22480 25940 22492 25943
rect 21735 25912 22492 25940
rect 21735 25909 21747 25912
rect 21689 25903 21747 25909
rect 22480 25909 22492 25912
rect 22526 25940 22538 25943
rect 24173 25943 24231 25949
rect 24173 25940 24185 25943
rect 22526 25912 24185 25940
rect 22526 25909 22538 25912
rect 22480 25903 22538 25909
rect 24173 25909 24185 25912
rect 24219 25940 24231 25943
rect 24538 25940 24544 25952
rect 24219 25912 24544 25940
rect 24219 25909 24231 25912
rect 24173 25903 24231 25909
rect 24538 25900 24544 25912
rect 24596 25900 24602 25952
rect 25553 25943 25611 25949
rect 25553 25909 25565 25943
rect 25599 25940 25611 25943
rect 25826 25940 25832 25952
rect 25599 25912 25832 25940
rect 25599 25909 25611 25912
rect 25553 25903 25611 25909
rect 25826 25900 25832 25912
rect 25884 25900 25890 25952
rect 26764 25949 26792 26048
rect 30076 26048 30165 26076
rect 26749 25943 26807 25949
rect 25936 25912 26516 25940
rect 20306 25872 20312 25884
rect 19680 25844 20312 25872
rect 20306 25832 20312 25844
rect 20364 25832 20370 25884
rect 20493 25875 20551 25881
rect 20493 25841 20505 25875
rect 20539 25872 20551 25875
rect 20539 25844 21180 25872
rect 20539 25841 20551 25844
rect 20493 25835 20551 25841
rect 15632 25776 17592 25804
rect 21152 25804 21180 25844
rect 22330 25832 22336 25884
rect 22388 25872 22394 25884
rect 23989 25875 24047 25881
rect 22388 25844 22433 25872
rect 22388 25832 22394 25844
rect 23989 25841 24001 25875
rect 24035 25841 24047 25875
rect 23989 25835 24047 25841
rect 23802 25804 23808 25816
rect 21152 25776 23808 25804
rect 23802 25764 23808 25776
rect 23860 25804 23866 25816
rect 24004 25804 24032 25835
rect 24078 25832 24084 25884
rect 24136 25872 24142 25884
rect 25936 25872 25964 25912
rect 24136 25844 25964 25872
rect 26289 25875 26347 25881
rect 24136 25832 24142 25844
rect 26289 25841 26301 25875
rect 26335 25872 26347 25875
rect 26378 25872 26384 25884
rect 26335 25844 26384 25872
rect 26335 25841 26347 25844
rect 26289 25835 26347 25841
rect 26378 25832 26384 25844
rect 26436 25832 26442 25884
rect 26488 25872 26516 25912
rect 26749 25909 26761 25943
rect 26795 25909 26807 25943
rect 26930 25940 26936 25952
rect 26891 25912 26936 25940
rect 26749 25903 26807 25909
rect 26930 25900 26936 25912
rect 26988 25900 26994 25952
rect 28310 25940 28316 25952
rect 28223 25912 28316 25940
rect 28310 25900 28316 25912
rect 28368 25940 28374 25952
rect 29693 25943 29751 25949
rect 29693 25940 29705 25943
rect 28368 25912 29705 25940
rect 28368 25900 28374 25912
rect 29693 25909 29705 25912
rect 29739 25909 29751 25943
rect 29693 25903 29751 25909
rect 26948 25872 26976 25900
rect 26488 25844 26976 25872
rect 29049 25875 29107 25881
rect 29049 25841 29061 25875
rect 29095 25841 29107 25875
rect 29049 25835 29107 25841
rect 29233 25875 29291 25881
rect 29233 25841 29245 25875
rect 29279 25872 29291 25875
rect 29598 25872 29604 25884
rect 29279 25844 29604 25872
rect 29279 25841 29291 25844
rect 29233 25835 29291 25841
rect 23860 25776 24032 25804
rect 23860 25764 23866 25776
rect 25274 25764 25280 25816
rect 25332 25804 25338 25816
rect 28218 25804 28224 25816
rect 25332 25776 28224 25804
rect 25332 25764 25338 25776
rect 28218 25764 28224 25776
rect 28276 25764 28282 25816
rect 29064 25804 29092 25835
rect 29598 25832 29604 25844
rect 29656 25832 29662 25884
rect 30076 25804 30104 26048
rect 30153 26045 30165 26048
rect 30199 26076 30211 26079
rect 31438 26076 31444 26088
rect 30199 26048 31444 26076
rect 30199 26045 30211 26048
rect 30153 26039 30211 26045
rect 31438 26036 31444 26048
rect 31496 26036 31502 26088
rect 30242 26008 30248 26020
rect 30203 25980 30248 26008
rect 30242 25968 30248 25980
rect 30300 25968 30306 26020
rect 30518 25900 30524 25952
rect 30576 25940 30582 25952
rect 30797 25943 30855 25949
rect 30797 25940 30809 25943
rect 30576 25912 30809 25940
rect 30576 25900 30582 25912
rect 30797 25909 30809 25912
rect 30843 25909 30855 25943
rect 30797 25903 30855 25909
rect 31257 25943 31315 25949
rect 31257 25909 31269 25943
rect 31303 25940 31315 25943
rect 31530 25940 31536 25952
rect 31303 25912 31536 25940
rect 31303 25909 31315 25912
rect 31257 25903 31315 25909
rect 31530 25900 31536 25912
rect 31588 25940 31594 25952
rect 31809 25943 31867 25949
rect 31809 25940 31821 25943
rect 31588 25912 31821 25940
rect 31588 25900 31594 25912
rect 31809 25909 31821 25912
rect 31855 25909 31867 25943
rect 31809 25903 31867 25909
rect 31349 25875 31407 25881
rect 31349 25841 31361 25875
rect 31395 25872 31407 25875
rect 32174 25872 32180 25884
rect 31395 25844 32180 25872
rect 31395 25841 31407 25844
rect 31349 25835 31407 25841
rect 32174 25832 32180 25844
rect 32232 25832 32238 25884
rect 31898 25804 31904 25816
rect 29064 25776 30104 25804
rect 31859 25776 31904 25804
rect 31898 25764 31904 25776
rect 31956 25764 31962 25816
rect 11000 25714 34368 25736
rect 11000 25662 19142 25714
rect 19194 25662 19206 25714
rect 19258 25662 19270 25714
rect 19322 25662 19334 25714
rect 19386 25662 29142 25714
rect 29194 25662 29206 25714
rect 29258 25662 29270 25714
rect 29322 25662 29334 25714
rect 29386 25662 34368 25714
rect 11000 25640 34368 25662
rect 22977 25603 23035 25609
rect 22977 25569 22989 25603
rect 23023 25600 23035 25603
rect 23023 25572 26792 25600
rect 23023 25569 23035 25572
rect 22977 25563 23035 25569
rect 13958 25492 13964 25544
rect 14016 25532 14022 25544
rect 17086 25532 17092 25544
rect 14016 25504 14726 25532
rect 17047 25504 17092 25532
rect 14016 25492 14022 25504
rect 17086 25492 17092 25504
rect 17144 25492 17150 25544
rect 19478 25492 19484 25544
rect 19536 25532 19542 25544
rect 20677 25535 20735 25541
rect 19536 25504 20076 25532
rect 19536 25492 19542 25504
rect 13774 25424 13780 25476
rect 13832 25464 13838 25476
rect 13832 25436 14004 25464
rect 13832 25424 13838 25436
rect 13976 25405 14004 25436
rect 16718 25424 16724 25476
rect 16776 25464 16782 25476
rect 17638 25464 17644 25476
rect 16776 25436 17644 25464
rect 16776 25424 16782 25436
rect 17638 25424 17644 25436
rect 17696 25464 17702 25476
rect 17733 25467 17791 25473
rect 17733 25464 17745 25467
rect 17696 25436 17745 25464
rect 17696 25424 17702 25436
rect 17733 25433 17745 25436
rect 17779 25433 17791 25467
rect 17733 25427 17791 25433
rect 17822 25424 17828 25476
rect 17880 25464 17886 25476
rect 18101 25467 18159 25473
rect 18101 25464 18113 25467
rect 17880 25436 18113 25464
rect 17880 25424 17886 25436
rect 18101 25433 18113 25436
rect 18147 25433 18159 25467
rect 18101 25427 18159 25433
rect 18285 25467 18343 25473
rect 18285 25433 18297 25467
rect 18331 25464 18343 25467
rect 19018 25464 19024 25476
rect 18331 25436 19024 25464
rect 18331 25433 18343 25436
rect 18285 25427 18343 25433
rect 19018 25424 19024 25436
rect 19076 25464 19082 25476
rect 19570 25464 19576 25476
rect 19076 25436 19576 25464
rect 19076 25424 19082 25436
rect 19570 25424 19576 25436
rect 19628 25424 19634 25476
rect 19846 25464 19852 25476
rect 19759 25436 19852 25464
rect 19846 25424 19852 25436
rect 19904 25464 19910 25476
rect 20048 25473 20076 25504
rect 20677 25501 20689 25535
rect 20723 25532 20735 25535
rect 22698 25532 22704 25544
rect 20723 25504 22704 25532
rect 20723 25501 20735 25504
rect 20677 25495 20735 25501
rect 20033 25467 20091 25473
rect 19904 25436 19984 25464
rect 19904 25424 19910 25436
rect 13961 25399 14019 25405
rect 13961 25365 13973 25399
rect 14007 25365 14019 25399
rect 15982 25396 15988 25408
rect 15943 25368 15988 25396
rect 13961 25359 14019 25365
rect 15982 25356 15988 25368
rect 16040 25356 16046 25408
rect 17549 25399 17607 25405
rect 17549 25365 17561 25399
rect 17595 25365 17607 25399
rect 19956 25396 19984 25436
rect 20033 25433 20045 25467
rect 20079 25433 20091 25467
rect 20398 25464 20404 25476
rect 20359 25436 20404 25464
rect 20033 25427 20091 25433
rect 20398 25424 20404 25436
rect 20456 25424 20462 25476
rect 21410 25464 21416 25476
rect 20508 25436 21416 25464
rect 20508 25396 20536 25436
rect 21410 25424 21416 25436
rect 21468 25424 21474 25476
rect 21594 25464 21600 25476
rect 21555 25436 21600 25464
rect 21594 25424 21600 25436
rect 21652 25424 21658 25476
rect 22532 25473 22560 25504
rect 22698 25492 22704 25504
rect 22756 25492 22762 25544
rect 22882 25492 22888 25544
rect 22940 25532 22946 25544
rect 22940 25504 23756 25532
rect 22940 25492 22946 25504
rect 21873 25467 21931 25473
rect 21873 25433 21885 25467
rect 21919 25464 21931 25467
rect 22333 25467 22391 25473
rect 22333 25464 22345 25467
rect 21919 25436 22345 25464
rect 21919 25433 21931 25436
rect 21873 25427 21931 25433
rect 22333 25433 22345 25436
rect 22379 25433 22391 25467
rect 22333 25427 22391 25433
rect 22480 25467 22560 25473
rect 22480 25433 22492 25467
rect 22526 25436 22560 25467
rect 23526 25464 23532 25476
rect 23487 25436 23532 25464
rect 22526 25433 22538 25436
rect 22480 25427 22538 25433
rect 23526 25424 23532 25436
rect 23584 25424 23590 25476
rect 23728 25473 23756 25504
rect 25274 25492 25280 25544
rect 25332 25532 25338 25544
rect 26764 25541 26792 25572
rect 29506 25560 29512 25612
rect 29564 25600 29570 25612
rect 29877 25603 29935 25609
rect 29877 25600 29889 25603
rect 29564 25572 29889 25600
rect 29564 25560 29570 25572
rect 29877 25569 29889 25572
rect 29923 25569 29935 25603
rect 32174 25600 32180 25612
rect 32135 25572 32180 25600
rect 29877 25563 29935 25569
rect 32174 25560 32180 25572
rect 32232 25560 32238 25612
rect 25553 25535 25611 25541
rect 25553 25532 25565 25535
rect 25332 25504 25565 25532
rect 25332 25492 25338 25504
rect 25553 25501 25565 25504
rect 25599 25501 25611 25535
rect 25553 25495 25611 25501
rect 26749 25535 26807 25541
rect 26749 25501 26761 25535
rect 26795 25501 26807 25535
rect 28310 25532 28316 25544
rect 28271 25504 28316 25532
rect 26749 25495 26807 25501
rect 28310 25492 28316 25504
rect 28368 25492 28374 25544
rect 29782 25532 29788 25544
rect 29743 25504 29788 25532
rect 29782 25492 29788 25504
rect 29840 25492 29846 25544
rect 30518 25492 30524 25544
rect 30576 25532 30582 25544
rect 31530 25532 31536 25544
rect 30576 25504 30840 25532
rect 31491 25504 31536 25532
rect 30576 25492 30582 25504
rect 23713 25467 23771 25473
rect 23713 25433 23725 25467
rect 23759 25433 23771 25467
rect 23713 25427 23771 25433
rect 25700 25467 25758 25473
rect 25700 25433 25712 25467
rect 25746 25464 25758 25467
rect 25826 25464 25832 25476
rect 25746 25436 25832 25464
rect 25746 25433 25758 25436
rect 25700 25427 25758 25433
rect 25826 25424 25832 25436
rect 25884 25424 25890 25476
rect 26102 25464 26108 25476
rect 25936 25436 26108 25464
rect 22698 25396 22704 25408
rect 19956 25368 20536 25396
rect 22659 25368 22704 25396
rect 17549 25359 17607 25365
rect 17564 25328 17592 25359
rect 22698 25356 22704 25368
rect 22756 25356 22762 25408
rect 24081 25399 24139 25405
rect 24081 25365 24093 25399
rect 24127 25396 24139 25399
rect 24630 25396 24636 25408
rect 24127 25368 24636 25396
rect 24127 25365 24139 25368
rect 24081 25359 24139 25365
rect 24630 25356 24636 25368
rect 24688 25356 24694 25408
rect 25936 25405 25964 25436
rect 26102 25424 26108 25436
rect 26160 25424 26166 25476
rect 26378 25424 26384 25476
rect 26436 25464 26442 25476
rect 26933 25467 26991 25473
rect 26933 25464 26945 25467
rect 26436 25436 26700 25464
rect 26436 25424 26442 25436
rect 25921 25399 25979 25405
rect 25921 25365 25933 25399
rect 25967 25365 25979 25399
rect 26672 25396 26700 25436
rect 26856 25436 26945 25464
rect 26856 25396 26884 25436
rect 26933 25433 26945 25436
rect 26979 25433 26991 25467
rect 28221 25467 28279 25473
rect 28221 25464 28233 25467
rect 26933 25427 26991 25433
rect 27040 25436 28233 25464
rect 26672 25368 26884 25396
rect 25921 25359 25979 25365
rect 17730 25328 17736 25340
rect 17564 25300 17736 25328
rect 17730 25288 17736 25300
rect 17788 25328 17794 25340
rect 18650 25328 18656 25340
rect 17788 25300 18656 25328
rect 17788 25288 17794 25300
rect 18650 25288 18656 25300
rect 18708 25288 18714 25340
rect 26197 25331 26255 25337
rect 26197 25297 26209 25331
rect 26243 25328 26255 25331
rect 27040 25328 27068 25436
rect 28221 25433 28233 25436
rect 28267 25433 28279 25467
rect 28221 25427 28279 25433
rect 28954 25424 28960 25476
rect 29012 25464 29018 25476
rect 29049 25467 29107 25473
rect 29049 25464 29061 25467
rect 29012 25436 29061 25464
rect 29012 25424 29018 25436
rect 29049 25433 29061 25436
rect 29095 25433 29107 25467
rect 29049 25427 29107 25433
rect 29141 25467 29199 25473
rect 29141 25433 29153 25467
rect 29187 25464 29199 25467
rect 30610 25464 30616 25476
rect 29187 25436 30616 25464
rect 29187 25433 29199 25436
rect 29141 25427 29199 25433
rect 30610 25424 30616 25436
rect 30668 25424 30674 25476
rect 30812 25473 30840 25504
rect 31530 25492 31536 25504
rect 31588 25492 31594 25544
rect 30797 25467 30855 25473
rect 30797 25433 30809 25467
rect 30843 25433 30855 25467
rect 30797 25427 30855 25433
rect 31717 25467 31775 25473
rect 31717 25433 31729 25467
rect 31763 25464 31775 25467
rect 32358 25464 32364 25476
rect 31763 25436 32364 25464
rect 31763 25433 31775 25436
rect 31717 25427 31775 25433
rect 32358 25424 32364 25436
rect 32416 25424 32422 25476
rect 27301 25399 27359 25405
rect 27301 25365 27313 25399
rect 27347 25396 27359 25399
rect 28586 25396 28592 25408
rect 27347 25368 28592 25396
rect 27347 25365 27359 25368
rect 27301 25359 27359 25365
rect 28586 25356 28592 25368
rect 28644 25356 28650 25408
rect 26243 25300 27068 25328
rect 26243 25297 26255 25300
rect 26197 25291 26255 25297
rect 13958 25220 13964 25272
rect 14016 25260 14022 25272
rect 14218 25263 14276 25269
rect 14218 25260 14230 25263
rect 14016 25232 14230 25260
rect 14016 25220 14022 25232
rect 14218 25229 14230 25232
rect 14264 25229 14276 25263
rect 22606 25260 22612 25272
rect 22567 25232 22612 25260
rect 14218 25223 14276 25229
rect 22606 25220 22612 25232
rect 22664 25220 22670 25272
rect 25829 25263 25887 25269
rect 25829 25229 25841 25263
rect 25875 25260 25887 25263
rect 25918 25260 25924 25272
rect 25875 25232 25924 25260
rect 25875 25229 25887 25232
rect 25829 25223 25887 25229
rect 25918 25220 25924 25232
rect 25976 25220 25982 25272
rect 11000 25170 34368 25192
rect 11000 25118 14142 25170
rect 14194 25118 14206 25170
rect 14258 25118 14270 25170
rect 14322 25118 14334 25170
rect 14386 25118 24142 25170
rect 24194 25118 24206 25170
rect 24258 25118 24270 25170
rect 24322 25118 24334 25170
rect 24386 25118 34368 25170
rect 11000 25096 34368 25118
rect 21042 25056 21048 25068
rect 20600 25028 21048 25056
rect 13958 24880 13964 24932
rect 14016 24920 14022 24932
rect 14145 24923 14203 24929
rect 14145 24920 14157 24923
rect 14016 24892 14157 24920
rect 14016 24880 14022 24892
rect 14145 24889 14157 24892
rect 14191 24889 14203 24923
rect 14145 24883 14203 24889
rect 15433 24923 15491 24929
rect 15433 24889 15445 24923
rect 15479 24920 15491 24923
rect 15982 24920 15988 24932
rect 15479 24892 15988 24920
rect 15479 24889 15491 24892
rect 15433 24883 15491 24889
rect 15982 24880 15988 24892
rect 16040 24880 16046 24932
rect 19478 24880 19484 24932
rect 19536 24920 19542 24932
rect 19536 24892 19892 24920
rect 19536 24880 19542 24892
rect 14694 24852 14700 24864
rect 14655 24824 14700 24852
rect 14694 24812 14700 24824
rect 14752 24812 14758 24864
rect 14789 24855 14847 24861
rect 14789 24821 14801 24855
rect 14835 24821 14847 24855
rect 15062 24852 15068 24864
rect 15023 24824 15068 24852
rect 14789 24815 14847 24821
rect 13406 24744 13412 24796
rect 13464 24784 13470 24796
rect 14804 24784 14832 24815
rect 15062 24812 15068 24824
rect 15120 24812 15126 24864
rect 15522 24852 15528 24864
rect 15483 24824 15528 24852
rect 15522 24812 15528 24824
rect 15580 24812 15586 24864
rect 16902 24852 16908 24864
rect 16863 24824 16908 24852
rect 16902 24812 16908 24824
rect 16960 24812 16966 24864
rect 19205 24855 19263 24861
rect 19205 24821 19217 24855
rect 19251 24821 19263 24855
rect 19205 24815 19263 24821
rect 19389 24855 19447 24861
rect 19389 24821 19401 24855
rect 19435 24821 19447 24855
rect 19570 24852 19576 24864
rect 19531 24824 19576 24852
rect 19389 24815 19447 24821
rect 17454 24784 17460 24796
rect 13464 24756 14832 24784
rect 17415 24756 17460 24784
rect 13464 24744 13470 24756
rect 17454 24744 17460 24756
rect 17512 24744 17518 24796
rect 19220 24784 19248 24815
rect 19404 24784 19432 24815
rect 19570 24812 19576 24824
rect 19628 24812 19634 24864
rect 19864 24861 19892 24892
rect 19849 24855 19907 24861
rect 19849 24821 19861 24855
rect 19895 24821 19907 24855
rect 19849 24815 19907 24821
rect 20102 24855 20160 24861
rect 20102 24821 20114 24855
rect 20148 24852 20160 24855
rect 20600 24852 20628 25028
rect 21042 25016 21048 25028
rect 21100 25056 21106 25068
rect 23066 25056 23072 25068
rect 21100 25028 23072 25056
rect 21100 25016 21106 25028
rect 23066 25016 23072 25028
rect 23124 25016 23130 25068
rect 23713 25059 23771 25065
rect 23713 25025 23725 25059
rect 23759 25056 23771 25059
rect 23894 25056 23900 25068
rect 23759 25028 23900 25056
rect 23759 25025 23771 25028
rect 23713 25019 23771 25025
rect 23894 25016 23900 25028
rect 23952 25016 23958 25068
rect 25550 25016 25556 25068
rect 25608 25056 25614 25068
rect 25608 25028 28172 25056
rect 25608 25016 25614 25028
rect 22698 24988 22704 25000
rect 22440 24960 22704 24988
rect 20677 24923 20735 24929
rect 20677 24889 20689 24923
rect 20723 24920 20735 24923
rect 21594 24920 21600 24932
rect 20723 24892 21600 24920
rect 20723 24889 20735 24892
rect 20677 24883 20735 24889
rect 21594 24880 21600 24892
rect 21652 24880 21658 24932
rect 21226 24852 21232 24864
rect 20148 24824 20628 24852
rect 21187 24824 21232 24852
rect 20148 24821 20160 24824
rect 20102 24815 20160 24821
rect 21226 24812 21232 24824
rect 21284 24812 21290 24864
rect 21318 24812 21324 24864
rect 21376 24852 21382 24864
rect 21413 24855 21471 24861
rect 21413 24852 21425 24855
rect 21376 24824 21425 24852
rect 21376 24812 21382 24824
rect 21413 24821 21425 24824
rect 21459 24821 21471 24855
rect 22330 24852 22336 24864
rect 22291 24824 22336 24852
rect 21413 24815 21471 24821
rect 22330 24812 22336 24824
rect 22388 24812 22394 24864
rect 22440 24861 22468 24960
rect 22698 24948 22704 24960
rect 22756 24988 22762 25000
rect 23434 24988 23440 25000
rect 22756 24960 23440 24988
rect 22756 24948 22762 24960
rect 23434 24948 23440 24960
rect 23492 24948 23498 25000
rect 23066 24880 23072 24932
rect 23124 24920 23130 24932
rect 25642 24920 25648 24932
rect 23124 24892 23572 24920
rect 25603 24892 25648 24920
rect 23124 24880 23130 24892
rect 22425 24855 22483 24861
rect 22425 24821 22437 24855
rect 22471 24821 22483 24855
rect 23434 24852 23440 24864
rect 23395 24824 23440 24852
rect 22425 24815 22483 24821
rect 23434 24812 23440 24824
rect 23492 24812 23498 24864
rect 23544 24861 23572 24892
rect 25642 24880 25648 24892
rect 25700 24880 25706 24932
rect 26746 24920 26752 24932
rect 26212 24892 26752 24920
rect 23529 24855 23587 24861
rect 23529 24821 23541 24855
rect 23575 24821 23587 24855
rect 23529 24815 23587 24821
rect 25369 24855 25427 24861
rect 25369 24821 25381 24855
rect 25415 24852 25427 24855
rect 26212 24852 26240 24892
rect 26746 24880 26752 24892
rect 26804 24880 26810 24932
rect 26378 24852 26384 24864
rect 25415 24824 26240 24852
rect 26339 24824 26384 24852
rect 25415 24821 25427 24824
rect 25369 24815 25427 24821
rect 26378 24812 26384 24824
rect 26436 24812 26442 24864
rect 28144 24861 28172 25028
rect 28218 25016 28224 25068
rect 28276 25056 28282 25068
rect 28276 25028 28321 25056
rect 28276 25016 28282 25028
rect 30702 24988 30708 25000
rect 30663 24960 30708 24988
rect 30702 24948 30708 24960
rect 30760 24948 30766 25000
rect 31346 24948 31352 25000
rect 31404 24988 31410 25000
rect 32729 24991 32787 24997
rect 32729 24988 32741 24991
rect 31404 24960 32741 24988
rect 31404 24948 31410 24960
rect 32729 24957 32741 24960
rect 32775 24957 32787 24991
rect 32729 24951 32787 24957
rect 28129 24855 28187 24861
rect 28129 24821 28141 24855
rect 28175 24821 28187 24855
rect 28129 24815 28187 24821
rect 29417 24855 29475 24861
rect 29417 24821 29429 24855
rect 29463 24852 29475 24855
rect 29874 24852 29880 24864
rect 29463 24824 29880 24852
rect 29463 24821 29475 24824
rect 29417 24815 29475 24821
rect 29874 24812 29880 24824
rect 29932 24812 29938 24864
rect 30334 24852 30340 24864
rect 30295 24824 30340 24852
rect 30334 24812 30340 24824
rect 30392 24812 30398 24864
rect 31162 24812 31168 24864
rect 31220 24852 31226 24864
rect 31441 24855 31499 24861
rect 31441 24852 31453 24855
rect 31220 24824 31453 24852
rect 31220 24812 31226 24824
rect 31441 24821 31453 24824
rect 31487 24821 31499 24855
rect 32358 24852 32364 24864
rect 32319 24824 32364 24852
rect 31441 24815 31499 24821
rect 32358 24812 32364 24824
rect 32416 24812 32422 24864
rect 19662 24784 19668 24796
rect 19220 24756 19340 24784
rect 19404 24756 19668 24784
rect 18650 24676 18656 24728
rect 18708 24716 18714 24728
rect 19312 24716 19340 24756
rect 19662 24744 19668 24756
rect 19720 24744 19726 24796
rect 21781 24787 21839 24793
rect 21781 24753 21793 24787
rect 21827 24753 21839 24787
rect 21781 24747 21839 24753
rect 22885 24787 22943 24793
rect 22885 24753 22897 24787
rect 22931 24784 22943 24787
rect 23250 24784 23256 24796
rect 22931 24756 23256 24784
rect 22931 24753 22943 24756
rect 22885 24747 22943 24753
rect 21502 24716 21508 24728
rect 18708 24688 21508 24716
rect 18708 24676 18714 24688
rect 21502 24676 21508 24688
rect 21560 24676 21566 24728
rect 21796 24716 21824 24747
rect 23250 24744 23256 24756
rect 23308 24744 23314 24796
rect 23342 24744 23348 24796
rect 23400 24784 23406 24796
rect 25185 24787 25243 24793
rect 25185 24784 25197 24787
rect 23400 24756 25197 24784
rect 23400 24744 23406 24756
rect 25185 24753 25197 24756
rect 25231 24753 25243 24787
rect 25185 24747 25243 24753
rect 25274 24744 25280 24796
rect 25332 24784 25338 24796
rect 26197 24787 26255 24793
rect 26197 24784 26209 24787
rect 25332 24756 26209 24784
rect 25332 24744 25338 24756
rect 26197 24753 26209 24756
rect 26243 24753 26255 24787
rect 26197 24747 26255 24753
rect 26749 24787 26807 24793
rect 26749 24753 26761 24787
rect 26795 24784 26807 24787
rect 27022 24784 27028 24796
rect 26795 24756 27028 24784
rect 26795 24753 26807 24756
rect 26749 24747 26807 24753
rect 27022 24744 27028 24756
rect 27080 24744 27086 24796
rect 27942 24784 27948 24796
rect 27903 24756 27948 24784
rect 27942 24744 27948 24756
rect 28000 24744 28006 24796
rect 29892 24784 29920 24812
rect 30242 24784 30248 24796
rect 29892 24756 30248 24784
rect 30242 24744 30248 24756
rect 30300 24744 30306 24796
rect 22514 24716 22520 24728
rect 21796 24688 22520 24716
rect 22514 24676 22520 24688
rect 22572 24676 22578 24728
rect 22974 24676 22980 24728
rect 23032 24716 23038 24728
rect 24354 24716 24360 24728
rect 23032 24688 24360 24716
rect 23032 24676 23038 24688
rect 24354 24676 24360 24688
rect 24412 24676 24418 24728
rect 11000 24626 34368 24648
rect 11000 24574 19142 24626
rect 19194 24574 19206 24626
rect 19258 24574 19270 24626
rect 19322 24574 19334 24626
rect 19386 24574 29142 24626
rect 29194 24574 29206 24626
rect 29258 24574 29270 24626
rect 29322 24574 29334 24626
rect 29386 24574 34368 24626
rect 11000 24552 34368 24574
rect 22606 24472 22612 24524
rect 22664 24512 22670 24524
rect 25090 24512 25096 24524
rect 22664 24484 25096 24512
rect 22664 24472 22670 24484
rect 25090 24472 25096 24484
rect 25148 24512 25154 24524
rect 25148 24484 25320 24512
rect 25148 24472 25154 24484
rect 12857 24447 12915 24453
rect 12857 24413 12869 24447
rect 12903 24444 12915 24447
rect 13406 24444 13412 24456
rect 12903 24416 13268 24444
rect 13367 24416 13412 24444
rect 12903 24413 12915 24416
rect 12857 24407 12915 24413
rect 13041 24379 13099 24385
rect 13041 24345 13053 24379
rect 13087 24345 13099 24379
rect 13240 24376 13268 24416
rect 13406 24404 13412 24416
rect 13464 24404 13470 24456
rect 16537 24447 16595 24453
rect 16537 24413 16549 24447
rect 16583 24444 16595 24447
rect 16626 24444 16632 24456
rect 16583 24416 16632 24444
rect 16583 24413 16595 24416
rect 16537 24407 16595 24413
rect 16626 24404 16632 24416
rect 16684 24404 16690 24456
rect 19570 24444 19576 24456
rect 18024 24416 19576 24444
rect 14421 24379 14479 24385
rect 14421 24376 14433 24379
rect 13240 24348 14433 24376
rect 13041 24339 13099 24345
rect 14421 24345 14433 24348
rect 14467 24376 14479 24379
rect 14602 24376 14608 24388
rect 14467 24348 14608 24376
rect 14467 24345 14479 24348
rect 14421 24339 14479 24345
rect 13056 24308 13084 24339
rect 14602 24336 14608 24348
rect 14660 24336 14666 24388
rect 14694 24336 14700 24388
rect 14752 24376 14758 24388
rect 14789 24379 14847 24385
rect 14789 24376 14801 24379
rect 14752 24348 14801 24376
rect 14752 24336 14758 24348
rect 14789 24345 14801 24348
rect 14835 24345 14847 24379
rect 14789 24339 14847 24345
rect 15157 24379 15215 24385
rect 15157 24345 15169 24379
rect 15203 24376 15215 24379
rect 16902 24376 16908 24388
rect 15203 24348 16908 24376
rect 15203 24345 15215 24348
rect 15157 24339 15215 24345
rect 15172 24308 15200 24339
rect 16902 24336 16908 24348
rect 16960 24336 16966 24388
rect 16997 24379 17055 24385
rect 16997 24345 17009 24379
rect 17043 24345 17055 24379
rect 16997 24339 17055 24345
rect 17273 24379 17331 24385
rect 17273 24345 17285 24379
rect 17319 24345 17331 24379
rect 17454 24376 17460 24388
rect 17415 24348 17460 24376
rect 17273 24339 17331 24345
rect 13056 24280 15200 24308
rect 16626 24268 16632 24320
rect 16684 24308 16690 24320
rect 17012 24308 17040 24339
rect 16684 24280 17040 24308
rect 16684 24268 16690 24280
rect 17288 24172 17316 24339
rect 17454 24336 17460 24348
rect 17512 24336 17518 24388
rect 17822 24376 17828 24388
rect 17783 24348 17828 24376
rect 17822 24336 17828 24348
rect 17880 24336 17886 24388
rect 18024 24385 18052 24416
rect 19570 24404 19576 24416
rect 19628 24404 19634 24456
rect 22716 24416 25228 24444
rect 18009 24379 18067 24385
rect 18009 24345 18021 24379
rect 18055 24345 18067 24379
rect 18466 24376 18472 24388
rect 18379 24348 18472 24376
rect 18009 24339 18067 24345
rect 18466 24336 18472 24348
rect 18524 24336 18530 24388
rect 18650 24376 18656 24388
rect 18611 24348 18656 24376
rect 18650 24336 18656 24348
rect 18708 24336 18714 24388
rect 19021 24379 19079 24385
rect 19021 24345 19033 24379
rect 19067 24376 19079 24379
rect 19202 24376 19208 24388
rect 19067 24348 19208 24376
rect 19067 24345 19079 24348
rect 19021 24339 19079 24345
rect 19202 24336 19208 24348
rect 19260 24376 19266 24388
rect 19478 24376 19484 24388
rect 19260 24348 19484 24376
rect 19260 24336 19266 24348
rect 19478 24336 19484 24348
rect 19536 24336 19542 24388
rect 19662 24376 19668 24388
rect 19575 24348 19668 24376
rect 19662 24336 19668 24348
rect 19720 24376 19726 24388
rect 20030 24376 20036 24388
rect 19720 24348 20036 24376
rect 19720 24336 19726 24348
rect 20030 24336 20036 24348
rect 20088 24336 20094 24388
rect 22514 24376 22520 24388
rect 22475 24348 22520 24376
rect 22514 24336 22520 24348
rect 22572 24336 22578 24388
rect 18484 24308 18512 24336
rect 18926 24308 18932 24320
rect 18484 24280 18932 24308
rect 18926 24268 18932 24280
rect 18984 24268 18990 24320
rect 19573 24311 19631 24317
rect 19573 24277 19585 24311
rect 19619 24308 19631 24311
rect 19846 24308 19852 24320
rect 19619 24280 19852 24308
rect 19619 24277 19631 24280
rect 19573 24271 19631 24277
rect 19846 24268 19852 24280
rect 19904 24268 19910 24320
rect 22422 24308 22428 24320
rect 22383 24280 22428 24308
rect 22422 24268 22428 24280
rect 22480 24308 22486 24320
rect 22716 24308 22744 24416
rect 22882 24376 22888 24388
rect 22843 24348 22888 24376
rect 22882 24336 22888 24348
rect 22940 24336 22946 24388
rect 23529 24379 23587 24385
rect 23529 24345 23541 24379
rect 23575 24376 23587 24379
rect 23802 24376 23808 24388
rect 23575 24348 23808 24376
rect 23575 24345 23587 24348
rect 23529 24339 23587 24345
rect 23802 24336 23808 24348
rect 23860 24376 23866 24388
rect 23986 24376 23992 24388
rect 23860 24348 23992 24376
rect 23860 24336 23866 24348
rect 23986 24336 23992 24348
rect 24044 24336 24050 24388
rect 24354 24376 24360 24388
rect 24315 24348 24360 24376
rect 24354 24336 24360 24348
rect 24412 24336 24418 24388
rect 24541 24379 24599 24385
rect 24541 24345 24553 24379
rect 24587 24376 24599 24379
rect 24814 24376 24820 24388
rect 24587 24348 24820 24376
rect 24587 24345 24599 24348
rect 24541 24339 24599 24345
rect 24814 24336 24820 24348
rect 24872 24336 24878 24388
rect 25200 24385 25228 24416
rect 25292 24385 25320 24484
rect 25918 24444 25924 24456
rect 25879 24416 25924 24444
rect 25918 24404 25924 24416
rect 25976 24404 25982 24456
rect 27117 24447 27175 24453
rect 27117 24413 27129 24447
rect 27163 24444 27175 24447
rect 28862 24444 28868 24456
rect 27163 24416 28868 24444
rect 27163 24413 27175 24416
rect 27117 24407 27175 24413
rect 28862 24404 28868 24416
rect 28920 24404 28926 24456
rect 30518 24444 30524 24456
rect 29340 24416 30524 24444
rect 25185 24379 25243 24385
rect 25185 24345 25197 24379
rect 25231 24345 25243 24379
rect 25185 24339 25243 24345
rect 25277 24379 25335 24385
rect 25277 24345 25289 24379
rect 25323 24345 25335 24379
rect 25458 24376 25464 24388
rect 25419 24348 25464 24376
rect 25277 24339 25335 24345
rect 22480 24280 22744 24308
rect 22977 24311 23035 24317
rect 22480 24268 22486 24280
rect 22977 24277 22989 24311
rect 23023 24308 23035 24311
rect 23434 24308 23440 24320
rect 23023 24280 23440 24308
rect 23023 24277 23035 24280
rect 22977 24271 23035 24277
rect 23434 24268 23440 24280
rect 23492 24308 23498 24320
rect 24081 24311 24139 24317
rect 24081 24308 24093 24311
rect 23492 24280 24093 24308
rect 23492 24268 23498 24280
rect 24081 24277 24093 24280
rect 24127 24277 24139 24311
rect 25200 24308 25228 24339
rect 25458 24336 25464 24348
rect 25516 24336 25522 24388
rect 27022 24376 27028 24388
rect 26983 24348 27028 24376
rect 27022 24336 27028 24348
rect 27080 24336 27086 24388
rect 27850 24376 27856 24388
rect 27811 24348 27856 24376
rect 27850 24336 27856 24348
rect 27908 24376 27914 24388
rect 28586 24376 28592 24388
rect 27908 24348 28448 24376
rect 28547 24348 28592 24376
rect 27908 24336 27914 24348
rect 26378 24308 26384 24320
rect 25200 24280 26384 24308
rect 24081 24271 24139 24277
rect 24096 24240 24124 24271
rect 26378 24268 26384 24280
rect 26436 24268 26442 24320
rect 27942 24308 27948 24320
rect 27903 24280 27948 24308
rect 27942 24268 27948 24280
rect 28000 24268 28006 24320
rect 28420 24308 28448 24348
rect 28586 24336 28592 24348
rect 28644 24336 28650 24388
rect 28681 24379 28739 24385
rect 28681 24345 28693 24379
rect 28727 24376 28739 24379
rect 29340 24376 29368 24416
rect 30518 24404 30524 24416
rect 30576 24404 30582 24456
rect 31346 24404 31352 24456
rect 31404 24444 31410 24456
rect 31441 24447 31499 24453
rect 31441 24444 31453 24447
rect 31404 24416 31453 24444
rect 31404 24404 31410 24416
rect 31441 24413 31453 24416
rect 31487 24413 31499 24447
rect 31441 24407 31499 24413
rect 31533 24447 31591 24453
rect 31533 24413 31545 24447
rect 31579 24444 31591 24447
rect 31898 24444 31904 24456
rect 31579 24416 31904 24444
rect 31579 24413 31591 24416
rect 31533 24407 31591 24413
rect 31898 24404 31904 24416
rect 31956 24404 31962 24456
rect 32269 24447 32327 24453
rect 32269 24413 32281 24447
rect 32315 24444 32327 24447
rect 32358 24444 32364 24456
rect 32315 24416 32364 24444
rect 32315 24413 32327 24416
rect 32269 24407 32327 24413
rect 32358 24404 32364 24416
rect 32416 24404 32422 24456
rect 28727 24348 29368 24376
rect 29417 24379 29475 24385
rect 28727 24345 28739 24348
rect 28681 24339 28739 24345
rect 29417 24345 29429 24379
rect 29463 24345 29475 24379
rect 29417 24339 29475 24345
rect 28954 24308 28960 24320
rect 28420 24280 28960 24308
rect 28954 24268 28960 24280
rect 29012 24308 29018 24320
rect 29432 24308 29460 24339
rect 29782 24336 29788 24388
rect 29840 24376 29846 24388
rect 30245 24379 30303 24385
rect 30245 24376 30257 24379
rect 29840 24348 30257 24376
rect 29840 24336 29846 24348
rect 30245 24345 30257 24348
rect 30291 24376 30303 24379
rect 30334 24376 30340 24388
rect 30291 24348 30340 24376
rect 30291 24345 30303 24348
rect 30245 24339 30303 24345
rect 30334 24336 30340 24348
rect 30392 24336 30398 24388
rect 30702 24336 30708 24388
rect 30760 24376 30766 24388
rect 32085 24379 32143 24385
rect 32085 24376 32097 24379
rect 30760 24348 32097 24376
rect 30760 24336 30766 24348
rect 32085 24345 32097 24348
rect 32131 24345 32143 24379
rect 32085 24339 32143 24345
rect 29012 24280 29460 24308
rect 29509 24311 29567 24317
rect 29012 24268 29018 24280
rect 29509 24277 29521 24311
rect 29555 24308 29567 24311
rect 29966 24308 29972 24320
rect 29555 24280 29972 24308
rect 29555 24277 29567 24280
rect 29509 24271 29567 24277
rect 29966 24268 29972 24280
rect 30024 24268 30030 24320
rect 30981 24311 31039 24317
rect 30981 24277 30993 24311
rect 31027 24308 31039 24311
rect 31162 24308 31168 24320
rect 31027 24280 31168 24308
rect 31027 24277 31039 24280
rect 30981 24271 31039 24277
rect 31162 24268 31168 24280
rect 31220 24268 31226 24320
rect 25458 24240 25464 24252
rect 24096 24212 25464 24240
rect 25458 24200 25464 24212
rect 25516 24200 25522 24252
rect 19849 24175 19907 24181
rect 19849 24172 19861 24175
rect 17288 24144 19861 24172
rect 19849 24141 19861 24144
rect 19895 24172 19907 24175
rect 20398 24172 20404 24184
rect 19895 24144 20404 24172
rect 19895 24141 19907 24144
rect 19849 24135 19907 24141
rect 20398 24132 20404 24144
rect 20456 24132 20462 24184
rect 21965 24175 22023 24181
rect 21965 24141 21977 24175
rect 22011 24172 22023 24175
rect 23066 24172 23072 24184
rect 22011 24144 23072 24172
rect 22011 24141 22023 24144
rect 21965 24135 22023 24141
rect 23066 24132 23072 24144
rect 23124 24132 23130 24184
rect 30061 24175 30119 24181
rect 30061 24141 30073 24175
rect 30107 24172 30119 24175
rect 31806 24172 31812 24184
rect 30107 24144 31812 24172
rect 30107 24141 30119 24144
rect 30061 24135 30119 24141
rect 31806 24132 31812 24144
rect 31864 24132 31870 24184
rect 11000 24082 34368 24104
rect 11000 24030 14142 24082
rect 14194 24030 14206 24082
rect 14258 24030 14270 24082
rect 14322 24030 14334 24082
rect 14386 24030 24142 24082
rect 24194 24030 24206 24082
rect 24258 24030 24270 24082
rect 24322 24030 24334 24082
rect 24386 24030 34368 24082
rect 11000 24008 34368 24030
rect 13130 23928 13136 23980
rect 13188 23968 13194 23980
rect 27942 23968 27948 23980
rect 13188 23940 27948 23968
rect 13188 23928 13194 23940
rect 27942 23928 27948 23940
rect 28000 23928 28006 23980
rect 16534 23860 16540 23912
rect 16592 23900 16598 23912
rect 27298 23900 27304 23912
rect 16592 23872 27304 23900
rect 16592 23860 16598 23872
rect 27298 23860 27304 23872
rect 27356 23860 27362 23912
rect 30702 23900 30708 23912
rect 30663 23872 30708 23900
rect 30702 23860 30708 23872
rect 30760 23860 30766 23912
rect 14602 23792 14608 23844
rect 14660 23832 14666 23844
rect 14697 23835 14755 23841
rect 14697 23832 14709 23835
rect 14660 23804 14709 23832
rect 14660 23792 14666 23804
rect 14697 23801 14709 23804
rect 14743 23801 14755 23835
rect 16718 23832 16724 23844
rect 14697 23795 14755 23801
rect 15540 23804 16724 23832
rect 14786 23724 14792 23776
rect 14844 23764 14850 23776
rect 15540 23773 15568 23804
rect 16718 23792 16724 23804
rect 16776 23792 16782 23844
rect 18926 23792 18932 23844
rect 18984 23832 18990 23844
rect 18984 23804 19156 23832
rect 18984 23792 18990 23804
rect 15249 23767 15307 23773
rect 15249 23764 15261 23767
rect 14844 23736 15261 23764
rect 14844 23724 14850 23736
rect 15249 23733 15261 23736
rect 15295 23733 15307 23767
rect 15249 23727 15307 23733
rect 15525 23767 15583 23773
rect 15525 23733 15537 23767
rect 15571 23733 15583 23767
rect 15525 23727 15583 23733
rect 15709 23767 15767 23773
rect 15709 23733 15721 23767
rect 15755 23764 15767 23767
rect 16074 23764 16080 23776
rect 15755 23736 16080 23764
rect 15755 23733 15767 23736
rect 15709 23727 15767 23733
rect 16074 23724 16080 23736
rect 16132 23724 16138 23776
rect 18193 23767 18251 23773
rect 18193 23733 18205 23767
rect 18239 23764 18251 23767
rect 18374 23764 18380 23776
rect 18239 23736 18380 23764
rect 18239 23733 18251 23736
rect 18193 23727 18251 23733
rect 18374 23724 18380 23736
rect 18432 23724 18438 23776
rect 19018 23764 19024 23776
rect 18979 23736 19024 23764
rect 19018 23724 19024 23736
rect 19076 23724 19082 23776
rect 19128 23764 19156 23804
rect 19202 23792 19208 23844
rect 19260 23832 19266 23844
rect 20585 23835 20643 23841
rect 19260 23804 19800 23832
rect 19260 23792 19266 23804
rect 19297 23767 19355 23773
rect 19297 23764 19309 23767
rect 19128 23736 19309 23764
rect 19297 23733 19309 23736
rect 19343 23733 19355 23767
rect 19297 23727 19355 23733
rect 19481 23767 19539 23773
rect 19481 23733 19493 23767
rect 19527 23764 19539 23767
rect 19570 23764 19576 23776
rect 19527 23736 19576 23764
rect 19527 23733 19539 23736
rect 19481 23727 19539 23733
rect 19570 23724 19576 23736
rect 19628 23724 19634 23776
rect 19772 23773 19800 23804
rect 20585 23801 20597 23835
rect 20631 23832 20643 23835
rect 20631 23804 21548 23832
rect 20631 23801 20643 23804
rect 20585 23795 20643 23801
rect 19757 23767 19815 23773
rect 19757 23733 19769 23767
rect 19803 23733 19815 23767
rect 19757 23727 19815 23733
rect 19846 23724 19852 23776
rect 19904 23764 19910 23776
rect 19950 23767 20008 23773
rect 19950 23764 19962 23767
rect 19904 23736 19962 23764
rect 19904 23724 19910 23736
rect 19950 23733 19962 23736
rect 19996 23733 20008 23767
rect 19950 23727 20008 23733
rect 18006 23696 18012 23708
rect 17967 23668 18012 23696
rect 18006 23656 18012 23668
rect 18064 23656 18070 23708
rect 18561 23699 18619 23705
rect 18561 23665 18573 23699
rect 18607 23696 18619 23699
rect 19662 23696 19668 23708
rect 18607 23668 19668 23696
rect 18607 23665 18619 23668
rect 18561 23659 18619 23665
rect 19662 23656 19668 23668
rect 19720 23656 19726 23708
rect 19956 23696 19984 23727
rect 20122 23724 20128 23776
rect 20180 23764 20186 23776
rect 21045 23767 21103 23773
rect 21045 23764 21057 23767
rect 20180 23736 21057 23764
rect 20180 23724 20186 23736
rect 21045 23733 21057 23736
rect 21091 23764 21103 23767
rect 21410 23764 21416 23776
rect 21091 23736 21416 23764
rect 21091 23733 21103 23736
rect 21045 23727 21103 23733
rect 21410 23724 21416 23736
rect 21468 23724 21474 23776
rect 21520 23773 21548 23804
rect 22974 23792 22980 23844
rect 23032 23832 23038 23844
rect 23069 23835 23127 23841
rect 23069 23832 23081 23835
rect 23032 23804 23081 23832
rect 23032 23792 23038 23804
rect 23069 23801 23081 23804
rect 23115 23801 23127 23835
rect 23069 23795 23127 23801
rect 23802 23792 23808 23844
rect 23860 23792 23866 23844
rect 28313 23835 28371 23841
rect 28313 23801 28325 23835
rect 28359 23832 28371 23835
rect 30797 23835 30855 23841
rect 30797 23832 30809 23835
rect 28359 23804 30809 23832
rect 28359 23801 28371 23804
rect 28313 23795 28371 23801
rect 30797 23801 30809 23804
rect 30843 23801 30855 23835
rect 31806 23832 31812 23844
rect 31767 23804 31812 23832
rect 30797 23795 30855 23801
rect 31806 23792 31812 23804
rect 31864 23792 31870 23844
rect 21505 23767 21563 23773
rect 21505 23733 21517 23767
rect 21551 23733 21563 23767
rect 22882 23764 22888 23776
rect 21505 23727 21563 23733
rect 21612 23736 22888 23764
rect 21612 23696 21640 23736
rect 22882 23724 22888 23736
rect 22940 23724 22946 23776
rect 23820 23764 23848 23792
rect 23897 23767 23955 23773
rect 23897 23764 23909 23767
rect 23820 23736 23909 23764
rect 23897 23733 23909 23736
rect 23943 23733 23955 23767
rect 23897 23727 23955 23733
rect 23986 23724 23992 23776
rect 24044 23764 24050 23776
rect 24081 23767 24139 23773
rect 24081 23764 24093 23767
rect 24044 23736 24093 23764
rect 24044 23724 24050 23736
rect 24081 23733 24093 23736
rect 24127 23733 24139 23767
rect 24630 23764 24636 23776
rect 24591 23736 24636 23764
rect 24081 23727 24139 23733
rect 24630 23724 24636 23736
rect 24688 23724 24694 23776
rect 24998 23764 25004 23776
rect 24959 23736 25004 23764
rect 24998 23724 25004 23736
rect 25056 23724 25062 23776
rect 26473 23767 26531 23773
rect 26473 23733 26485 23767
rect 26519 23764 26531 23767
rect 26746 23764 26752 23776
rect 26519 23736 26752 23764
rect 26519 23733 26531 23736
rect 26473 23727 26531 23733
rect 26746 23724 26752 23736
rect 26804 23724 26810 23776
rect 28862 23764 28868 23776
rect 28823 23736 28868 23764
rect 28862 23724 28868 23736
rect 28920 23764 28926 23776
rect 28920 23736 30196 23764
rect 28920 23724 28926 23736
rect 19956 23668 21640 23696
rect 21781 23699 21839 23705
rect 21781 23665 21793 23699
rect 21827 23696 21839 23699
rect 23158 23696 23164 23708
rect 21827 23668 23164 23696
rect 21827 23665 21839 23668
rect 21781 23659 21839 23665
rect 23158 23656 23164 23668
rect 23216 23656 23222 23708
rect 26286 23696 26292 23708
rect 26247 23668 26292 23696
rect 26286 23656 26292 23668
rect 26344 23656 26350 23708
rect 26841 23699 26899 23705
rect 26841 23665 26853 23699
rect 26887 23696 26899 23699
rect 28126 23696 28132 23708
rect 26887 23668 28132 23696
rect 26887 23665 26899 23668
rect 26841 23659 26899 23665
rect 28126 23656 28132 23668
rect 28184 23656 28190 23708
rect 28221 23699 28279 23705
rect 28221 23665 28233 23699
rect 28267 23696 28279 23699
rect 29601 23699 29659 23705
rect 29601 23696 29613 23699
rect 28267 23668 29613 23696
rect 28267 23665 28279 23668
rect 28221 23659 28279 23665
rect 29601 23665 29613 23668
rect 29647 23665 29659 23699
rect 29782 23696 29788 23708
rect 29743 23668 29788 23696
rect 29601 23659 29659 23665
rect 23710 23628 23716 23640
rect 23671 23600 23716 23628
rect 23710 23588 23716 23600
rect 23768 23588 23774 23640
rect 29616 23628 29644 23659
rect 29782 23656 29788 23668
rect 29840 23656 29846 23708
rect 30168 23696 30196 23736
rect 30242 23724 30248 23776
rect 30300 23764 30306 23776
rect 31257 23767 31315 23773
rect 30300 23736 30345 23764
rect 30300 23724 30306 23736
rect 31257 23733 31269 23767
rect 31303 23733 31315 23767
rect 31257 23727 31315 23733
rect 31272 23696 31300 23727
rect 30168 23668 31300 23696
rect 31717 23699 31775 23705
rect 31717 23665 31729 23699
rect 31763 23665 31775 23699
rect 31717 23659 31775 23665
rect 31732 23628 31760 23659
rect 29616 23600 31760 23628
rect 11000 23538 34368 23560
rect 11000 23486 19142 23538
rect 19194 23486 19206 23538
rect 19258 23486 19270 23538
rect 19322 23486 19334 23538
rect 19386 23486 29142 23538
rect 29194 23486 29206 23538
rect 29258 23486 29270 23538
rect 29322 23486 29334 23538
rect 29386 23486 34368 23538
rect 11000 23464 34368 23486
rect 16902 23424 16908 23436
rect 16863 23396 16908 23424
rect 16902 23384 16908 23396
rect 16960 23384 16966 23436
rect 21042 23424 21048 23436
rect 21003 23396 21048 23424
rect 21042 23384 21048 23396
rect 21100 23384 21106 23436
rect 21410 23384 21416 23436
rect 21468 23424 21474 23436
rect 22149 23427 22207 23433
rect 22149 23424 22161 23427
rect 21468 23396 22161 23424
rect 21468 23384 21474 23396
rect 22149 23393 22161 23396
rect 22195 23393 22207 23427
rect 22974 23424 22980 23436
rect 22149 23387 22207 23393
rect 22256 23396 22980 23424
rect 15430 23356 15436 23368
rect 15343 23328 15436 23356
rect 14694 23288 14700 23300
rect 14655 23260 14700 23288
rect 14694 23248 14700 23260
rect 14752 23248 14758 23300
rect 14786 23248 14792 23300
rect 14844 23288 14850 23300
rect 15062 23288 15068 23300
rect 14844 23260 14889 23288
rect 14975 23260 15068 23288
rect 14844 23248 14850 23260
rect 15062 23248 15068 23260
rect 15120 23288 15126 23300
rect 15246 23288 15252 23300
rect 15120 23260 15252 23288
rect 15120 23248 15126 23260
rect 15246 23248 15252 23260
rect 15304 23248 15310 23300
rect 15356 23297 15384 23328
rect 15430 23316 15436 23328
rect 15488 23356 15494 23368
rect 18006 23356 18012 23368
rect 15488 23328 18012 23356
rect 15488 23316 15494 23328
rect 18006 23316 18012 23328
rect 18064 23356 18070 23368
rect 18469 23359 18527 23365
rect 18469 23356 18481 23359
rect 18064 23328 18481 23356
rect 18064 23316 18070 23328
rect 18469 23325 18481 23328
rect 18515 23325 18527 23359
rect 18469 23319 18527 23325
rect 19021 23359 19079 23365
rect 19021 23325 19033 23359
rect 19067 23356 19079 23359
rect 19067 23328 19340 23356
rect 19067 23325 19079 23328
rect 19021 23319 19079 23325
rect 15341 23291 15399 23297
rect 15341 23257 15353 23291
rect 15387 23257 15399 23291
rect 15341 23251 15399 23257
rect 16718 23248 16724 23300
rect 16776 23288 16782 23300
rect 17457 23291 17515 23297
rect 17457 23288 17469 23291
rect 16776 23260 17469 23288
rect 16776 23248 16782 23260
rect 17457 23257 17469 23260
rect 17503 23257 17515 23291
rect 17822 23288 17828 23300
rect 17783 23260 17828 23288
rect 17457 23251 17515 23257
rect 17822 23248 17828 23260
rect 17880 23248 17886 23300
rect 17917 23291 17975 23297
rect 17917 23257 17929 23291
rect 17963 23288 17975 23291
rect 18374 23288 18380 23300
rect 17963 23260 18380 23288
rect 17963 23257 17975 23260
rect 17917 23251 17975 23257
rect 18374 23248 18380 23260
rect 18432 23248 18438 23300
rect 18653 23291 18711 23297
rect 18653 23257 18665 23291
rect 18699 23288 18711 23291
rect 19202 23288 19208 23300
rect 18699 23260 19208 23288
rect 18699 23257 18711 23260
rect 18653 23251 18711 23257
rect 13406 23180 13412 23232
rect 13464 23220 13470 23232
rect 14145 23223 14203 23229
rect 14145 23220 14157 23223
rect 13464 23192 14157 23220
rect 13464 23180 13470 23192
rect 14145 23189 14157 23192
rect 14191 23189 14203 23223
rect 15522 23220 15528 23232
rect 15483 23192 15528 23220
rect 14145 23183 14203 23189
rect 15522 23180 15528 23192
rect 15580 23180 15586 23232
rect 15982 23180 15988 23232
rect 16040 23220 16046 23232
rect 17549 23223 17607 23229
rect 17549 23220 17561 23223
rect 16040 23192 17561 23220
rect 16040 23180 16046 23192
rect 17549 23189 17561 23192
rect 17595 23220 17607 23223
rect 18668 23220 18696 23251
rect 19202 23248 19208 23260
rect 19260 23248 19266 23300
rect 19312 23288 19340 23328
rect 19478 23316 19484 23368
rect 19536 23356 19542 23368
rect 19754 23356 19760 23368
rect 19536 23328 19760 23356
rect 19536 23316 19542 23328
rect 19754 23316 19760 23328
rect 19812 23316 19818 23368
rect 20309 23359 20367 23365
rect 20309 23325 20321 23359
rect 20355 23356 20367 23359
rect 20582 23356 20588 23368
rect 20355 23328 20588 23356
rect 20355 23325 20367 23328
rect 20309 23319 20367 23325
rect 20582 23316 20588 23328
rect 20640 23316 20646 23368
rect 21962 23316 21968 23368
rect 22020 23356 22026 23368
rect 22256 23365 22284 23396
rect 22974 23384 22980 23396
rect 23032 23384 23038 23436
rect 25458 23384 25464 23436
rect 25516 23424 25522 23436
rect 28221 23427 28279 23433
rect 28221 23424 28233 23427
rect 25516 23396 28233 23424
rect 25516 23384 25522 23396
rect 28221 23393 28233 23396
rect 28267 23424 28279 23427
rect 28494 23424 28500 23436
rect 28267 23396 28500 23424
rect 28267 23393 28279 23396
rect 28221 23387 28279 23393
rect 28494 23384 28500 23396
rect 28552 23384 28558 23436
rect 29782 23384 29788 23436
rect 29840 23424 29846 23436
rect 30981 23427 31039 23433
rect 30981 23424 30993 23427
rect 29840 23396 30993 23424
rect 29840 23384 29846 23396
rect 30981 23393 30993 23396
rect 31027 23393 31039 23427
rect 30981 23387 31039 23393
rect 22057 23359 22115 23365
rect 22057 23356 22069 23359
rect 22020 23328 22069 23356
rect 22020 23316 22026 23328
rect 22057 23325 22069 23328
rect 22103 23325 22115 23359
rect 22057 23319 22115 23325
rect 22241 23359 22299 23365
rect 22241 23325 22253 23359
rect 22287 23325 22299 23359
rect 22241 23319 22299 23325
rect 22514 23316 22520 23368
rect 22572 23356 22578 23368
rect 22609 23359 22667 23365
rect 22609 23356 22621 23359
rect 22572 23328 22621 23356
rect 22572 23316 22578 23328
rect 22609 23325 22621 23328
rect 22655 23325 22667 23359
rect 23066 23356 23072 23368
rect 23027 23328 23072 23356
rect 22609 23319 22667 23325
rect 23066 23316 23072 23328
rect 23124 23316 23130 23368
rect 23805 23359 23863 23365
rect 23805 23325 23817 23359
rect 23851 23356 23863 23359
rect 25274 23356 25280 23368
rect 23851 23328 25280 23356
rect 23851 23325 23863 23328
rect 23805 23319 23863 23325
rect 25274 23316 25280 23328
rect 25332 23316 25338 23368
rect 25384 23328 28172 23356
rect 19570 23288 19576 23300
rect 19312 23260 19576 23288
rect 19570 23248 19576 23260
rect 19628 23288 19634 23300
rect 19665 23291 19723 23297
rect 19665 23288 19677 23291
rect 19628 23260 19677 23288
rect 19628 23248 19634 23260
rect 19665 23257 19677 23260
rect 19711 23257 19723 23291
rect 20766 23288 20772 23300
rect 20727 23260 20772 23288
rect 19665 23251 19723 23257
rect 20766 23248 20772 23260
rect 20824 23248 20830 23300
rect 20953 23291 21011 23297
rect 20953 23257 20965 23291
rect 20999 23257 21011 23291
rect 20953 23251 21011 23257
rect 17595 23192 18696 23220
rect 17595 23189 17607 23192
rect 17549 23183 17607 23189
rect 19478 23180 19484 23232
rect 19536 23220 19542 23232
rect 20968 23220 20996 23251
rect 23158 23248 23164 23300
rect 23216 23297 23222 23300
rect 23216 23291 23274 23297
rect 23216 23257 23228 23291
rect 23262 23257 23274 23291
rect 23216 23251 23274 23257
rect 23216 23248 23222 23251
rect 23894 23248 23900 23300
rect 23952 23288 23958 23300
rect 25384 23297 25412 23328
rect 28144 23300 28172 23328
rect 25185 23291 25243 23297
rect 25185 23288 25197 23291
rect 23952 23260 25197 23288
rect 23952 23248 23958 23260
rect 25185 23257 25197 23260
rect 25231 23257 25243 23291
rect 25185 23251 25243 23257
rect 25369 23291 25427 23297
rect 25369 23257 25381 23291
rect 25415 23257 25427 23291
rect 27298 23288 27304 23300
rect 27259 23260 27304 23288
rect 25369 23251 25427 23257
rect 27298 23248 27304 23260
rect 27356 23248 27362 23300
rect 28034 23288 28040 23300
rect 27995 23260 28040 23288
rect 28034 23248 28040 23260
rect 28092 23248 28098 23300
rect 28126 23248 28132 23300
rect 28184 23288 28190 23300
rect 29233 23291 29291 23297
rect 29233 23288 29245 23291
rect 28184 23260 29245 23288
rect 28184 23248 28190 23260
rect 29233 23257 29245 23260
rect 29279 23257 29291 23291
rect 30886 23288 30892 23300
rect 30847 23260 30892 23288
rect 29233 23251 29291 23257
rect 30886 23248 30892 23260
rect 30944 23248 30950 23300
rect 21410 23220 21416 23232
rect 19536 23192 21416 23220
rect 19536 23180 19542 23192
rect 21410 23180 21416 23192
rect 21468 23180 21474 23232
rect 21502 23180 21508 23232
rect 21560 23220 21566 23232
rect 21873 23223 21931 23229
rect 21873 23220 21885 23223
rect 21560 23192 21885 23220
rect 21560 23180 21566 23192
rect 21873 23189 21885 23192
rect 21919 23189 21931 23223
rect 21873 23183 21931 23189
rect 22606 23180 22612 23232
rect 22664 23220 22670 23232
rect 23437 23223 23495 23229
rect 23437 23220 23449 23223
rect 22664 23192 23449 23220
rect 22664 23180 22670 23192
rect 23437 23189 23449 23192
rect 23483 23189 23495 23223
rect 23437 23183 23495 23189
rect 26102 23180 26108 23232
rect 26160 23220 26166 23232
rect 26473 23223 26531 23229
rect 26473 23220 26485 23223
rect 26160 23192 26485 23220
rect 26160 23180 26166 23192
rect 26473 23189 26485 23192
rect 26519 23189 26531 23223
rect 26473 23183 26531 23189
rect 26565 23223 26623 23229
rect 26565 23189 26577 23223
rect 26611 23220 26623 23223
rect 27206 23220 27212 23232
rect 26611 23192 27212 23220
rect 26611 23189 26623 23192
rect 26565 23183 26623 23189
rect 27206 23180 27212 23192
rect 27264 23180 27270 23232
rect 27390 23220 27396 23232
rect 27351 23192 27396 23220
rect 27390 23180 27396 23192
rect 27448 23220 27454 23232
rect 27850 23220 27856 23232
rect 27448 23192 27856 23220
rect 27448 23180 27454 23192
rect 27850 23180 27856 23192
rect 27908 23180 27914 23232
rect 11934 23112 11940 23164
rect 11992 23152 11998 23164
rect 19570 23152 19576 23164
rect 11992 23124 19576 23152
rect 11992 23112 11998 23124
rect 19570 23112 19576 23124
rect 19628 23112 19634 23164
rect 23345 23155 23403 23161
rect 23345 23121 23357 23155
rect 23391 23152 23403 23155
rect 23986 23152 23992 23164
rect 23391 23124 23992 23152
rect 23391 23121 23403 23124
rect 23345 23115 23403 23121
rect 23986 23112 23992 23124
rect 24044 23112 24050 23164
rect 18926 23044 18932 23096
rect 18984 23084 18990 23096
rect 19478 23084 19484 23096
rect 18984 23056 19484 23084
rect 18984 23044 18990 23056
rect 19478 23044 19484 23056
rect 19536 23044 19542 23096
rect 23618 23044 23624 23096
rect 23676 23084 23682 23096
rect 24906 23084 24912 23096
rect 23676 23056 24912 23084
rect 23676 23044 23682 23056
rect 24906 23044 24912 23056
rect 24964 23044 24970 23096
rect 25458 23084 25464 23096
rect 25419 23056 25464 23084
rect 25458 23044 25464 23056
rect 25516 23044 25522 23096
rect 29598 23084 29604 23096
rect 29559 23056 29604 23084
rect 29598 23044 29604 23056
rect 29656 23044 29662 23096
rect 11000 22994 34368 23016
rect 11000 22942 14142 22994
rect 14194 22942 14206 22994
rect 14258 22942 14270 22994
rect 14322 22942 14334 22994
rect 14386 22942 24142 22994
rect 24194 22942 24206 22994
rect 24258 22942 24270 22994
rect 24322 22942 24334 22994
rect 24386 22942 34368 22994
rect 11000 22920 34368 22942
rect 13774 22880 13780 22892
rect 13148 22852 13780 22880
rect 13148 22753 13176 22852
rect 13774 22840 13780 22852
rect 13832 22840 13838 22892
rect 14694 22840 14700 22892
rect 14752 22880 14758 22892
rect 15893 22883 15951 22889
rect 15893 22880 15905 22883
rect 14752 22852 15905 22880
rect 14752 22840 14758 22852
rect 15893 22849 15905 22852
rect 15939 22849 15951 22883
rect 19846 22880 19852 22892
rect 19807 22852 19852 22880
rect 15893 22843 15951 22849
rect 19846 22840 19852 22852
rect 19904 22840 19910 22892
rect 22330 22840 22336 22892
rect 22388 22880 22394 22892
rect 22698 22880 22704 22892
rect 22388 22852 22704 22880
rect 22388 22840 22394 22852
rect 22698 22840 22704 22852
rect 22756 22840 22762 22892
rect 18466 22812 18472 22824
rect 18427 22784 18472 22812
rect 18466 22772 18472 22784
rect 18524 22772 18530 22824
rect 23897 22815 23955 22821
rect 23897 22812 23909 22815
rect 21796 22784 23909 22812
rect 13133 22747 13191 22753
rect 13133 22713 13145 22747
rect 13179 22713 13191 22747
rect 13406 22744 13412 22756
rect 13367 22716 13412 22744
rect 13133 22707 13191 22713
rect 13406 22704 13412 22716
rect 13464 22704 13470 22756
rect 15157 22747 15215 22753
rect 15157 22713 15169 22747
rect 15203 22744 15215 22747
rect 15430 22744 15436 22756
rect 15203 22716 15436 22744
rect 15203 22713 15215 22716
rect 15157 22707 15215 22713
rect 15430 22704 15436 22716
rect 15488 22704 15494 22756
rect 16074 22704 16080 22756
rect 16132 22744 16138 22756
rect 16813 22747 16871 22753
rect 16813 22744 16825 22747
rect 16132 22716 16825 22744
rect 16132 22704 16138 22716
rect 16813 22713 16825 22716
rect 16859 22744 16871 22747
rect 20766 22744 20772 22756
rect 16859 22716 20772 22744
rect 16859 22713 16871 22716
rect 16813 22707 16871 22713
rect 15614 22676 15620 22688
rect 15575 22648 15620 22676
rect 15614 22636 15620 22648
rect 15672 22636 15678 22688
rect 15801 22679 15859 22685
rect 15801 22645 15813 22679
rect 15847 22676 15859 22679
rect 15890 22676 15896 22688
rect 15847 22648 15896 22676
rect 15847 22645 15859 22648
rect 15801 22639 15859 22645
rect 15890 22636 15896 22648
rect 15948 22676 15954 22688
rect 16626 22676 16632 22688
rect 15948 22648 16632 22676
rect 15948 22636 15954 22648
rect 16626 22636 16632 22648
rect 16684 22636 16690 22688
rect 17457 22679 17515 22685
rect 17457 22645 17469 22679
rect 17503 22676 17515 22679
rect 18006 22676 18012 22688
rect 17503 22648 18012 22676
rect 17503 22645 17515 22648
rect 17457 22639 17515 22645
rect 18006 22636 18012 22648
rect 18064 22636 18070 22688
rect 18374 22676 18380 22688
rect 18335 22648 18380 22676
rect 18374 22636 18380 22648
rect 18432 22636 18438 22688
rect 19588 22685 19616 22716
rect 20766 22704 20772 22716
rect 20824 22704 20830 22756
rect 21045 22747 21103 22753
rect 21045 22713 21057 22747
rect 21091 22744 21103 22747
rect 21502 22744 21508 22756
rect 21091 22716 21508 22744
rect 21091 22713 21103 22716
rect 21045 22707 21103 22713
rect 21502 22704 21508 22716
rect 21560 22704 21566 22756
rect 21796 22753 21824 22784
rect 23897 22781 23909 22784
rect 23943 22781 23955 22815
rect 23897 22775 23955 22781
rect 21781 22747 21839 22753
rect 21781 22713 21793 22747
rect 21827 22713 21839 22747
rect 21781 22707 21839 22713
rect 22333 22747 22391 22753
rect 22333 22713 22345 22747
rect 22379 22744 22391 22747
rect 23158 22744 23164 22756
rect 22379 22716 23164 22744
rect 22379 22713 22391 22716
rect 22333 22707 22391 22713
rect 23158 22704 23164 22716
rect 23216 22704 23222 22756
rect 23986 22704 23992 22756
rect 24044 22744 24050 22756
rect 25001 22747 25059 22753
rect 24044 22716 24089 22744
rect 24044 22704 24050 22716
rect 25001 22713 25013 22747
rect 25047 22744 25059 22747
rect 25458 22744 25464 22756
rect 25047 22716 25464 22744
rect 25047 22713 25059 22716
rect 25001 22707 25059 22713
rect 25458 22704 25464 22716
rect 25516 22704 25522 22756
rect 25918 22744 25924 22756
rect 25879 22716 25924 22744
rect 25918 22704 25924 22716
rect 25976 22704 25982 22756
rect 27390 22744 27396 22756
rect 26304 22716 27396 22744
rect 18653 22679 18711 22685
rect 18653 22645 18665 22679
rect 18699 22676 18711 22679
rect 19573 22679 19631 22685
rect 18699 22648 19432 22676
rect 18699 22645 18711 22648
rect 18653 22639 18711 22645
rect 14694 22608 14700 22620
rect 14634 22580 14700 22608
rect 14694 22568 14700 22580
rect 14752 22568 14758 22620
rect 18834 22540 18840 22552
rect 18795 22512 18840 22540
rect 18834 22500 18840 22512
rect 18892 22500 18898 22552
rect 19404 22540 19432 22648
rect 19573 22645 19585 22679
rect 19619 22645 19631 22679
rect 19754 22676 19760 22688
rect 19715 22648 19760 22676
rect 19573 22639 19631 22645
rect 19754 22636 19760 22648
rect 19812 22636 19818 22688
rect 19938 22636 19944 22688
rect 19996 22676 20002 22688
rect 21229 22679 21287 22685
rect 21229 22676 21241 22679
rect 19996 22648 21241 22676
rect 19996 22636 20002 22648
rect 21229 22645 21241 22648
rect 21275 22676 21287 22679
rect 21962 22676 21968 22688
rect 21275 22648 21968 22676
rect 21275 22645 21287 22648
rect 21229 22639 21287 22645
rect 21962 22636 21968 22648
rect 22020 22676 22026 22688
rect 22517 22679 22575 22685
rect 22517 22676 22529 22679
rect 22020 22648 22529 22676
rect 22020 22636 22026 22648
rect 22517 22645 22529 22648
rect 22563 22645 22575 22679
rect 22882 22676 22888 22688
rect 22517 22639 22575 22645
rect 22624 22648 22888 22676
rect 19478 22568 19484 22620
rect 19536 22608 19542 22620
rect 21134 22608 21140 22620
rect 19536 22580 21140 22608
rect 19536 22568 19542 22580
rect 21134 22568 21140 22580
rect 21192 22568 21198 22620
rect 21410 22608 21416 22620
rect 21371 22580 21416 22608
rect 21410 22568 21416 22580
rect 21468 22568 21474 22620
rect 22624 22617 22652 22648
rect 22882 22636 22888 22648
rect 22940 22636 22946 22688
rect 23069 22679 23127 22685
rect 23069 22645 23081 22679
rect 23115 22676 23127 22679
rect 23342 22676 23348 22688
rect 23115 22648 23348 22676
rect 23115 22645 23127 22648
rect 23069 22639 23127 22645
rect 23342 22636 23348 22648
rect 23400 22636 23406 22688
rect 23618 22676 23624 22688
rect 23579 22648 23624 22676
rect 23618 22636 23624 22648
rect 23676 22636 23682 22688
rect 23768 22679 23826 22685
rect 23768 22645 23780 22679
rect 23814 22645 23826 22679
rect 23768 22639 23826 22645
rect 22609 22611 22667 22617
rect 22609 22608 22621 22611
rect 21612 22580 22621 22608
rect 20122 22540 20128 22552
rect 19404 22512 20128 22540
rect 20122 22500 20128 22512
rect 20180 22500 20186 22552
rect 20950 22500 20956 22552
rect 21008 22540 21014 22552
rect 21321 22543 21379 22549
rect 21321 22540 21333 22543
rect 21008 22512 21333 22540
rect 21008 22500 21014 22512
rect 21321 22509 21333 22512
rect 21367 22540 21379 22543
rect 21502 22540 21508 22552
rect 21367 22512 21508 22540
rect 21367 22509 21379 22512
rect 21321 22503 21379 22509
rect 21502 22500 21508 22512
rect 21560 22540 21566 22552
rect 21612 22540 21640 22580
rect 22609 22577 22621 22580
rect 22655 22577 22667 22611
rect 22609 22571 22667 22577
rect 22698 22568 22704 22620
rect 22756 22608 22762 22620
rect 22756 22580 22801 22608
rect 22756 22568 22762 22580
rect 23783 22552 23811 22639
rect 25090 22636 25096 22688
rect 25148 22676 25154 22688
rect 25829 22679 25887 22685
rect 25829 22676 25841 22679
rect 25148 22648 25193 22676
rect 25292 22648 25841 22676
rect 25148 22636 25154 22648
rect 24357 22611 24415 22617
rect 24357 22577 24369 22611
rect 24403 22608 24415 22611
rect 24446 22608 24452 22620
rect 24403 22580 24452 22608
rect 24403 22577 24415 22580
rect 24357 22571 24415 22577
rect 24446 22568 24452 22580
rect 24504 22568 24510 22620
rect 24998 22568 25004 22620
rect 25056 22608 25062 22620
rect 25292 22608 25320 22648
rect 25829 22645 25841 22648
rect 25875 22676 25887 22679
rect 26304 22676 26332 22716
rect 27390 22704 27396 22716
rect 27448 22744 27454 22756
rect 28770 22744 28776 22756
rect 27448 22716 28776 22744
rect 27448 22704 27454 22716
rect 28770 22704 28776 22716
rect 28828 22704 28834 22756
rect 30429 22747 30487 22753
rect 28880 22716 30380 22744
rect 25875 22648 26332 22676
rect 25875 22645 25887 22648
rect 25829 22639 25887 22645
rect 26378 22636 26384 22688
rect 26436 22676 26442 22688
rect 26657 22679 26715 22685
rect 26657 22676 26669 22679
rect 26436 22648 26669 22676
rect 26436 22636 26442 22648
rect 26657 22645 26669 22648
rect 26703 22645 26715 22679
rect 26657 22639 26715 22645
rect 27206 22636 27212 22688
rect 27264 22676 27270 22688
rect 28880 22685 28908 22716
rect 28865 22679 28923 22685
rect 28865 22676 28877 22679
rect 27264 22648 28877 22676
rect 27264 22636 27270 22648
rect 28865 22645 28877 22648
rect 28911 22645 28923 22679
rect 30242 22676 30248 22688
rect 30203 22648 30248 22676
rect 28865 22639 28923 22645
rect 30242 22636 30248 22648
rect 30300 22636 30306 22688
rect 30352 22676 30380 22716
rect 30429 22713 30441 22747
rect 30475 22744 30487 22747
rect 30886 22744 30892 22756
rect 30475 22716 30892 22744
rect 30475 22713 30487 22716
rect 30429 22707 30487 22713
rect 30886 22704 30892 22716
rect 30944 22744 30950 22756
rect 31254 22744 31260 22756
rect 30944 22716 31260 22744
rect 30944 22704 30950 22716
rect 31254 22704 31260 22716
rect 31312 22704 31318 22756
rect 30794 22676 30800 22688
rect 30352 22648 30800 22676
rect 30794 22636 30800 22648
rect 30852 22636 30858 22688
rect 26470 22608 26476 22620
rect 25056 22580 25320 22608
rect 26431 22580 26476 22608
rect 25056 22568 25062 22580
rect 26470 22568 26476 22580
rect 26528 22568 26534 22620
rect 23783 22540 23808 22552
rect 21560 22512 21640 22540
rect 23715 22512 23808 22540
rect 21560 22500 21566 22512
rect 23802 22500 23808 22512
rect 23860 22540 23866 22552
rect 26749 22543 26807 22549
rect 26749 22540 26761 22543
rect 23860 22512 26761 22540
rect 23860 22500 23866 22512
rect 26749 22509 26761 22512
rect 26795 22509 26807 22543
rect 26749 22503 26807 22509
rect 11000 22450 34368 22472
rect 11000 22398 19142 22450
rect 19194 22398 19206 22450
rect 19258 22398 19270 22450
rect 19322 22398 19334 22450
rect 19386 22398 29142 22450
rect 29194 22398 29206 22450
rect 29258 22398 29270 22450
rect 29322 22398 29334 22450
rect 29386 22398 34368 22450
rect 11000 22376 34368 22398
rect 17822 22296 17828 22348
rect 17880 22296 17886 22348
rect 18374 22296 18380 22348
rect 18432 22336 18438 22348
rect 18469 22339 18527 22345
rect 18469 22336 18481 22339
rect 18432 22308 18481 22336
rect 18432 22296 18438 22308
rect 18469 22305 18481 22308
rect 18515 22305 18527 22339
rect 18469 22299 18527 22305
rect 20033 22339 20091 22345
rect 20033 22305 20045 22339
rect 20079 22336 20091 22339
rect 20582 22336 20588 22348
rect 20079 22308 20588 22336
rect 20079 22305 20091 22308
rect 20033 22299 20091 22305
rect 20582 22296 20588 22308
rect 20640 22296 20646 22348
rect 21410 22296 21416 22348
rect 21468 22296 21474 22348
rect 21502 22296 21508 22348
rect 21560 22336 21566 22348
rect 21560 22308 21605 22336
rect 21560 22296 21566 22308
rect 22698 22296 22704 22348
rect 22756 22336 22762 22348
rect 23805 22339 23863 22345
rect 23805 22336 23817 22339
rect 22756 22308 23817 22336
rect 22756 22296 22762 22308
rect 23805 22305 23817 22308
rect 23851 22305 23863 22339
rect 23805 22299 23863 22305
rect 25274 22296 25280 22348
rect 25332 22336 25338 22348
rect 25461 22339 25519 22345
rect 25461 22336 25473 22339
rect 25332 22308 25473 22336
rect 25332 22296 25338 22308
rect 25461 22305 25473 22308
rect 25507 22305 25519 22339
rect 29506 22336 29512 22348
rect 25461 22299 25519 22305
rect 28236 22308 29512 22336
rect 15157 22271 15215 22277
rect 15157 22268 15169 22271
rect 14252 22240 15169 22268
rect 14252 22209 14280 22240
rect 15157 22237 15169 22240
rect 15203 22268 15215 22271
rect 15614 22268 15620 22280
rect 15203 22240 15620 22268
rect 15203 22237 15215 22240
rect 15157 22231 15215 22237
rect 15614 22228 15620 22240
rect 15672 22228 15678 22280
rect 17840 22268 17868 22296
rect 19938 22268 19944 22280
rect 15816 22240 17868 22268
rect 19899 22240 19944 22268
rect 15816 22209 15844 22240
rect 19938 22228 19944 22240
rect 19996 22228 20002 22280
rect 20122 22268 20128 22280
rect 20083 22240 20128 22268
rect 20122 22228 20128 22240
rect 20180 22228 20186 22280
rect 21134 22228 21140 22280
rect 21192 22268 21198 22280
rect 21428 22268 21456 22296
rect 21597 22271 21655 22277
rect 21597 22268 21609 22271
rect 21192 22240 21364 22268
rect 21428 22240 21609 22268
rect 21192 22228 21198 22240
rect 14237 22203 14295 22209
rect 14237 22169 14249 22203
rect 14283 22169 14295 22203
rect 14237 22163 14295 22169
rect 14697 22203 14755 22209
rect 14697 22169 14709 22203
rect 14743 22200 14755 22203
rect 15801 22203 15859 22209
rect 14743 22172 15752 22200
rect 14743 22169 14755 22172
rect 14697 22163 14755 22169
rect 14329 22135 14387 22141
rect 14329 22101 14341 22135
rect 14375 22132 14387 22135
rect 14786 22132 14792 22144
rect 14375 22104 14792 22132
rect 14375 22101 14387 22104
rect 14329 22095 14387 22101
rect 14786 22092 14792 22104
rect 14844 22092 14850 22144
rect 15430 22092 15436 22144
rect 15488 22132 15494 22144
rect 15617 22135 15675 22141
rect 15617 22132 15629 22135
rect 15488 22104 15629 22132
rect 15488 22092 15494 22104
rect 15617 22101 15629 22104
rect 15663 22101 15675 22135
rect 15724 22132 15752 22172
rect 15801 22169 15813 22203
rect 15847 22169 15859 22203
rect 16166 22200 16172 22212
rect 16079 22172 16172 22200
rect 15801 22163 15859 22169
rect 16166 22160 16172 22172
rect 16224 22200 16230 22212
rect 16718 22200 16724 22212
rect 16224 22172 16724 22200
rect 16224 22160 16230 22172
rect 16718 22160 16724 22172
rect 16776 22160 16782 22212
rect 17825 22203 17883 22209
rect 17825 22169 17837 22203
rect 17871 22200 17883 22203
rect 17914 22200 17920 22212
rect 17871 22172 17920 22200
rect 17871 22169 17883 22172
rect 17825 22163 17883 22169
rect 17914 22160 17920 22172
rect 17972 22160 17978 22212
rect 19956 22200 19984 22228
rect 21229 22203 21287 22209
rect 21229 22200 21241 22203
rect 18208 22172 19984 22200
rect 20140 22172 21241 22200
rect 15890 22132 15896 22144
rect 15724 22104 15896 22132
rect 15617 22095 15675 22101
rect 15890 22092 15896 22104
rect 15948 22092 15954 22144
rect 16074 22132 16080 22144
rect 16035 22104 16080 22132
rect 16074 22092 16080 22104
rect 16132 22092 16138 22144
rect 18208 22141 18236 22172
rect 18193 22135 18251 22141
rect 18193 22101 18205 22135
rect 18239 22101 18251 22135
rect 18193 22095 18251 22101
rect 18282 22092 18288 22144
rect 18340 22132 18346 22144
rect 19018 22132 19024 22144
rect 18340 22104 19024 22132
rect 18340 22092 18346 22104
rect 19018 22092 19024 22104
rect 19076 22132 19082 22144
rect 19757 22135 19815 22141
rect 19757 22132 19769 22135
rect 19076 22104 19769 22132
rect 19076 22092 19082 22104
rect 19757 22101 19769 22104
rect 19803 22132 19815 22135
rect 20140 22132 20168 22172
rect 21229 22169 21241 22172
rect 21275 22169 21287 22203
rect 21336 22200 21364 22240
rect 21597 22237 21609 22240
rect 21643 22237 21655 22271
rect 21597 22231 21655 22237
rect 22974 22228 22980 22280
rect 23032 22268 23038 22280
rect 23989 22271 24047 22277
rect 23989 22268 24001 22271
rect 23032 22240 24001 22268
rect 23032 22228 23038 22240
rect 23989 22237 24001 22240
rect 24035 22237 24047 22271
rect 23989 22231 24047 22237
rect 24630 22228 24636 22280
rect 24688 22268 24694 22280
rect 25185 22271 25243 22277
rect 25185 22268 25197 22271
rect 24688 22240 25197 22268
rect 24688 22228 24694 22240
rect 25185 22237 25197 22240
rect 25231 22237 25243 22271
rect 25185 22231 25243 22237
rect 21413 22203 21471 22209
rect 21413 22200 21425 22203
rect 21336 22172 21425 22200
rect 21229 22163 21287 22169
rect 21413 22169 21425 22172
rect 21459 22200 21471 22203
rect 22238 22200 22244 22212
rect 21459 22172 22244 22200
rect 21459 22169 21471 22172
rect 21413 22163 21471 22169
rect 20490 22132 20496 22144
rect 19803 22104 20168 22132
rect 20451 22104 20496 22132
rect 19803 22101 19815 22104
rect 19757 22095 19815 22101
rect 20490 22092 20496 22104
rect 20548 22092 20554 22144
rect 16092 22064 16120 22092
rect 18101 22067 18159 22073
rect 18101 22064 18113 22067
rect 16092 22036 18113 22064
rect 18101 22033 18113 22036
rect 18147 22033 18159 22067
rect 21244 22064 21272 22163
rect 22238 22160 22244 22172
rect 22296 22160 22302 22212
rect 22330 22160 22336 22212
rect 22388 22200 22394 22212
rect 22425 22203 22483 22209
rect 22425 22200 22437 22203
rect 22388 22172 22437 22200
rect 22388 22160 22394 22172
rect 22425 22169 22437 22172
rect 22471 22169 22483 22203
rect 22882 22200 22888 22212
rect 22425 22163 22483 22169
rect 22587 22172 22888 22200
rect 22587 22141 22615 22172
rect 22882 22160 22888 22172
rect 22940 22200 22946 22212
rect 23621 22203 23679 22209
rect 23621 22200 23633 22203
rect 22940 22172 23633 22200
rect 22940 22160 22946 22172
rect 23621 22169 23633 22172
rect 23667 22169 23679 22203
rect 23621 22163 23679 22169
rect 23897 22203 23955 22209
rect 23897 22169 23909 22203
rect 23943 22169 23955 22203
rect 23897 22163 23955 22169
rect 25369 22203 25427 22209
rect 25369 22169 25381 22203
rect 25415 22200 25427 22203
rect 25458 22200 25464 22212
rect 25415 22172 25464 22200
rect 25415 22169 25427 22172
rect 25369 22163 25427 22169
rect 21965 22135 22023 22141
rect 21965 22101 21977 22135
rect 22011 22132 22023 22135
rect 22572 22135 22630 22141
rect 22011 22104 22468 22132
rect 22011 22101 22023 22104
rect 21965 22095 22023 22101
rect 22440 22076 22468 22104
rect 22572 22101 22584 22135
rect 22618 22101 22630 22135
rect 22572 22095 22630 22101
rect 22793 22135 22851 22141
rect 22793 22101 22805 22135
rect 22839 22132 22851 22135
rect 23158 22132 23164 22144
rect 22839 22104 23164 22132
rect 22839 22101 22851 22104
rect 22793 22095 22851 22101
rect 23158 22092 23164 22104
rect 23216 22132 23222 22144
rect 23912 22132 23940 22163
rect 25458 22160 25464 22172
rect 25516 22160 25522 22212
rect 26194 22160 26200 22212
rect 26252 22200 26258 22212
rect 26289 22203 26347 22209
rect 26289 22200 26301 22203
rect 26252 22172 26301 22200
rect 26252 22160 26258 22172
rect 26289 22169 26301 22172
rect 26335 22169 26347 22203
rect 27758 22200 27764 22212
rect 27671 22172 27764 22200
rect 26289 22163 26347 22169
rect 27758 22160 27764 22172
rect 27816 22200 27822 22212
rect 28236 22200 28264 22308
rect 29506 22296 29512 22308
rect 29564 22296 29570 22348
rect 28865 22271 28923 22277
rect 28865 22237 28877 22271
rect 28911 22268 28923 22271
rect 31349 22271 31407 22277
rect 31349 22268 31361 22271
rect 28911 22240 31361 22268
rect 28911 22237 28923 22240
rect 28865 22231 28923 22237
rect 31349 22237 31361 22240
rect 31395 22237 31407 22271
rect 31349 22231 31407 22237
rect 27816 22172 28264 22200
rect 28681 22203 28739 22209
rect 27816 22160 27822 22172
rect 28681 22169 28693 22203
rect 28727 22169 28739 22203
rect 28681 22163 28739 22169
rect 29325 22203 29383 22209
rect 29325 22169 29337 22203
rect 29371 22200 29383 22203
rect 29506 22200 29512 22212
rect 29371 22172 29512 22200
rect 29371 22169 29383 22172
rect 29325 22163 29383 22169
rect 23216 22104 23940 22132
rect 23216 22092 23222 22104
rect 23986 22092 23992 22144
rect 24044 22132 24050 22144
rect 24357 22135 24415 22141
rect 24357 22132 24369 22135
rect 24044 22104 24369 22132
rect 24044 22092 24050 22104
rect 24357 22101 24369 22104
rect 24403 22101 24415 22135
rect 27850 22132 27856 22144
rect 27811 22104 27856 22132
rect 24357 22095 24415 22101
rect 27850 22092 27856 22104
rect 27908 22092 27914 22144
rect 28696 22132 28724 22163
rect 29506 22160 29512 22172
rect 29564 22160 29570 22212
rect 29969 22203 30027 22209
rect 29969 22169 29981 22203
rect 30015 22169 30027 22203
rect 30242 22200 30248 22212
rect 30203 22172 30248 22200
rect 29969 22163 30027 22169
rect 29984 22132 30012 22163
rect 30242 22160 30248 22172
rect 30300 22160 30306 22212
rect 30794 22200 30800 22212
rect 30755 22172 30800 22200
rect 30794 22160 30800 22172
rect 30852 22160 30858 22212
rect 31254 22200 31260 22212
rect 31215 22172 31260 22200
rect 31254 22160 31260 22172
rect 31312 22160 31318 22212
rect 30058 22132 30064 22144
rect 28696 22104 30064 22132
rect 30058 22092 30064 22104
rect 30116 22092 30122 22144
rect 22330 22064 22336 22076
rect 21244 22036 22336 22064
rect 18101 22027 18159 22033
rect 22330 22024 22336 22036
rect 22388 22024 22394 22076
rect 22422 22024 22428 22076
rect 22480 22024 22486 22076
rect 23069 22067 23127 22073
rect 23069 22033 23081 22067
rect 23115 22064 23127 22067
rect 29874 22064 29880 22076
rect 23115 22036 29880 22064
rect 23115 22033 23127 22036
rect 23069 22027 23127 22033
rect 29874 22024 29880 22036
rect 29932 22024 29938 22076
rect 18006 22005 18012 22008
rect 17990 21999 18012 22005
rect 17990 21965 18002 21999
rect 17990 21959 18012 21965
rect 18006 21956 18012 21959
rect 18064 21956 18070 22008
rect 21962 21956 21968 22008
rect 22020 21996 22026 22008
rect 22701 21999 22759 22005
rect 22701 21996 22713 21999
rect 22020 21968 22713 21996
rect 22020 21956 22026 21968
rect 22701 21965 22713 21968
rect 22747 21965 22759 21999
rect 22701 21959 22759 21965
rect 29322 21956 29328 22008
rect 29380 21996 29386 22008
rect 30242 21996 30248 22008
rect 29380 21968 30248 21996
rect 29380 21956 29386 21968
rect 30242 21956 30248 21968
rect 30300 21956 30306 22008
rect 11000 21906 34368 21928
rect 11000 21854 14142 21906
rect 14194 21854 14206 21906
rect 14258 21854 14270 21906
rect 14322 21854 14334 21906
rect 14386 21854 24142 21906
rect 24194 21854 24206 21906
rect 24258 21854 24270 21906
rect 24322 21854 24334 21906
rect 24386 21854 34368 21906
rect 11000 21832 34368 21854
rect 14329 21795 14387 21801
rect 14329 21761 14341 21795
rect 14375 21792 14387 21795
rect 14694 21792 14700 21804
rect 14375 21764 14700 21792
rect 14375 21761 14387 21764
rect 14329 21755 14387 21761
rect 14694 21752 14700 21764
rect 14752 21752 14758 21804
rect 22698 21792 22704 21804
rect 20692 21764 22704 21792
rect 15890 21724 15896 21736
rect 15851 21696 15896 21724
rect 15890 21684 15896 21696
rect 15948 21684 15954 21736
rect 16166 21656 16172 21668
rect 15448 21628 16172 21656
rect 14145 21591 14203 21597
rect 14145 21557 14157 21591
rect 14191 21588 14203 21591
rect 14602 21588 14608 21600
rect 14191 21560 14608 21588
rect 14191 21557 14203 21560
rect 14145 21551 14203 21557
rect 14602 21548 14608 21560
rect 14660 21588 14666 21600
rect 14878 21588 14884 21600
rect 14660 21560 14884 21588
rect 14660 21548 14666 21560
rect 14878 21548 14884 21560
rect 14936 21548 14942 21600
rect 15448 21597 15476 21628
rect 16166 21616 16172 21628
rect 16224 21616 16230 21668
rect 19754 21616 19760 21668
rect 19812 21656 19818 21668
rect 20692 21656 20720 21764
rect 22698 21752 22704 21764
rect 22756 21752 22762 21804
rect 28034 21792 28040 21804
rect 23636 21764 28040 21792
rect 21410 21724 21416 21736
rect 20784 21696 21416 21724
rect 20784 21665 20812 21696
rect 21410 21684 21416 21696
rect 21468 21684 21474 21736
rect 22238 21684 22244 21736
rect 22296 21724 22302 21736
rect 22974 21724 22980 21736
rect 22296 21696 22980 21724
rect 22296 21684 22302 21696
rect 22974 21684 22980 21696
rect 23032 21684 23038 21736
rect 19812 21628 20720 21656
rect 20769 21659 20827 21665
rect 19812 21616 19818 21628
rect 15249 21591 15307 21597
rect 15249 21557 15261 21591
rect 15295 21557 15307 21591
rect 15249 21551 15307 21557
rect 15433 21591 15491 21597
rect 15433 21557 15445 21591
rect 15479 21557 15491 21591
rect 15433 21551 15491 21557
rect 15264 21520 15292 21551
rect 15522 21548 15528 21600
rect 15580 21588 15586 21600
rect 15893 21591 15951 21597
rect 15893 21588 15905 21591
rect 15580 21560 15905 21588
rect 15580 21548 15586 21560
rect 15893 21557 15905 21560
rect 15939 21557 15951 21591
rect 17454 21588 17460 21600
rect 17415 21560 17460 21588
rect 15893 21551 15951 21557
rect 17454 21548 17460 21560
rect 17512 21548 17518 21600
rect 17822 21548 17828 21600
rect 17880 21588 17886 21600
rect 18098 21588 18104 21600
rect 17880 21560 18104 21588
rect 17880 21548 17886 21560
rect 18098 21548 18104 21560
rect 18156 21548 18162 21600
rect 18282 21588 18288 21600
rect 18243 21560 18288 21588
rect 18282 21548 18288 21560
rect 18340 21548 18346 21600
rect 18469 21591 18527 21597
rect 18469 21557 18481 21591
rect 18515 21557 18527 21591
rect 18834 21588 18840 21600
rect 18795 21560 18840 21588
rect 18469 21551 18527 21557
rect 16074 21520 16080 21532
rect 15264 21492 16080 21520
rect 16074 21480 16080 21492
rect 16132 21480 16138 21532
rect 18116 21520 18144 21548
rect 18484 21520 18512 21551
rect 18834 21548 18840 21560
rect 18892 21548 18898 21600
rect 20416 21597 20444 21628
rect 20769 21625 20781 21659
rect 20815 21625 20827 21659
rect 20769 21619 20827 21625
rect 22330 21616 22336 21668
rect 22388 21656 22394 21668
rect 23636 21665 23664 21764
rect 28034 21752 28040 21764
rect 28092 21752 28098 21804
rect 28862 21752 28868 21804
rect 28920 21792 28926 21804
rect 28920 21764 30564 21792
rect 28920 21752 28926 21764
rect 27117 21727 27175 21733
rect 27117 21693 27129 21727
rect 27163 21724 27175 21727
rect 27850 21724 27856 21736
rect 27163 21696 27856 21724
rect 27163 21693 27175 21696
rect 27117 21687 27175 21693
rect 27850 21684 27856 21696
rect 27908 21684 27914 21736
rect 28052 21724 28080 21752
rect 30536 21724 30564 21764
rect 31990 21724 31996 21736
rect 28052 21696 30104 21724
rect 23621 21659 23679 21665
rect 22388 21628 23204 21656
rect 22388 21616 22394 21628
rect 23176 21600 23204 21628
rect 23621 21625 23633 21659
rect 23667 21625 23679 21659
rect 23621 21619 23679 21625
rect 24173 21659 24231 21665
rect 24173 21625 24185 21659
rect 24219 21656 24231 21659
rect 24446 21656 24452 21668
rect 24219 21628 24452 21656
rect 24219 21625 24231 21628
rect 24173 21619 24231 21625
rect 24446 21616 24452 21628
rect 24504 21616 24510 21668
rect 25093 21659 25151 21665
rect 25093 21625 25105 21659
rect 25139 21656 25151 21659
rect 28310 21656 28316 21668
rect 25139 21628 28316 21656
rect 25139 21625 25151 21628
rect 25093 21619 25151 21625
rect 28310 21616 28316 21628
rect 28368 21616 28374 21668
rect 20401 21591 20459 21597
rect 20401 21557 20413 21591
rect 20447 21557 20459 21591
rect 20401 21551 20459 21557
rect 20490 21548 20496 21600
rect 20548 21588 20554 21600
rect 21229 21591 21287 21597
rect 21229 21588 21241 21591
rect 20548 21560 21241 21588
rect 20548 21548 20554 21560
rect 21229 21557 21241 21560
rect 21275 21557 21287 21591
rect 21410 21588 21416 21600
rect 21371 21560 21416 21588
rect 21229 21551 21287 21557
rect 21410 21548 21416 21560
rect 21468 21548 21474 21600
rect 22146 21548 22152 21600
rect 22204 21588 22210 21600
rect 22882 21588 22888 21600
rect 22204 21560 22888 21588
rect 22204 21548 22210 21560
rect 22882 21548 22888 21560
rect 22940 21548 22946 21600
rect 23158 21588 23164 21600
rect 23119 21560 23164 21588
rect 23158 21548 23164 21560
rect 23216 21548 23222 21600
rect 23894 21548 23900 21600
rect 23952 21588 23958 21600
rect 24265 21591 24323 21597
rect 24265 21588 24277 21591
rect 23952 21560 24277 21588
rect 23952 21548 23958 21560
rect 24265 21557 24277 21560
rect 24311 21557 24323 21591
rect 24265 21551 24323 21557
rect 24630 21548 24636 21600
rect 24688 21588 24694 21600
rect 24998 21588 25004 21600
rect 24688 21560 25004 21588
rect 24688 21548 24694 21560
rect 24998 21548 25004 21560
rect 25056 21548 25062 21600
rect 26194 21548 26200 21600
rect 26252 21588 26258 21600
rect 26657 21591 26715 21597
rect 26657 21588 26669 21591
rect 26252 21560 26669 21588
rect 26252 21548 26258 21560
rect 26657 21557 26669 21560
rect 26703 21557 26715 21591
rect 26657 21551 26715 21557
rect 27758 21548 27764 21600
rect 27816 21588 27822 21600
rect 28129 21591 28187 21597
rect 28129 21588 28141 21591
rect 27816 21560 28141 21588
rect 27816 21548 27822 21560
rect 28129 21557 28141 21560
rect 28175 21557 28187 21591
rect 28129 21551 28187 21557
rect 28773 21591 28831 21597
rect 28773 21557 28785 21591
rect 28819 21588 28831 21591
rect 29322 21588 29328 21600
rect 28819 21560 29328 21588
rect 28819 21557 28831 21560
rect 28773 21551 28831 21557
rect 29322 21548 29328 21560
rect 29380 21548 29386 21600
rect 29598 21548 29604 21600
rect 29656 21588 29662 21600
rect 29693 21591 29751 21597
rect 29693 21588 29705 21591
rect 29656 21560 29705 21588
rect 29656 21548 29662 21560
rect 29693 21557 29705 21560
rect 29739 21557 29751 21591
rect 29874 21588 29880 21600
rect 29835 21560 29880 21588
rect 29693 21551 29751 21557
rect 18116 21492 18512 21520
rect 21781 21523 21839 21529
rect 21781 21489 21793 21523
rect 21827 21520 21839 21523
rect 26102 21520 26108 21532
rect 21827 21492 26108 21520
rect 21827 21489 21839 21492
rect 21781 21483 21839 21489
rect 26102 21480 26108 21492
rect 26160 21480 26166 21532
rect 27209 21523 27267 21529
rect 27209 21489 27221 21523
rect 27255 21520 27267 21523
rect 28494 21520 28500 21532
rect 27255 21492 28500 21520
rect 27255 21489 27267 21492
rect 27209 21483 27267 21489
rect 28494 21480 28500 21492
rect 28552 21480 28558 21532
rect 29233 21523 29291 21529
rect 29233 21489 29245 21523
rect 29279 21520 29291 21523
rect 29506 21520 29512 21532
rect 29279 21492 29512 21520
rect 29279 21489 29291 21492
rect 29233 21483 29291 21489
rect 29506 21480 29512 21492
rect 29564 21480 29570 21532
rect 29708 21520 29736 21551
rect 29874 21548 29880 21560
rect 29932 21548 29938 21600
rect 30076 21597 30104 21696
rect 30536 21696 31996 21724
rect 30536 21665 30564 21696
rect 31990 21684 31996 21696
rect 32048 21684 32054 21736
rect 30521 21659 30579 21665
rect 30521 21625 30533 21659
rect 30567 21625 30579 21659
rect 30521 21619 30579 21625
rect 30613 21659 30671 21665
rect 30613 21625 30625 21659
rect 30659 21656 30671 21659
rect 32174 21656 32180 21668
rect 30659 21628 32180 21656
rect 30659 21625 30671 21628
rect 30613 21619 30671 21625
rect 32174 21616 32180 21628
rect 32232 21616 32238 21668
rect 30061 21591 30119 21597
rect 30061 21557 30073 21591
rect 30107 21557 30119 21591
rect 31162 21588 31168 21600
rect 30061 21551 30119 21557
rect 30260 21560 31024 21588
rect 31123 21560 31168 21588
rect 30260 21520 30288 21560
rect 29708 21492 30288 21520
rect 30996 21520 31024 21560
rect 31162 21548 31168 21560
rect 31220 21548 31226 21600
rect 31625 21591 31683 21597
rect 31625 21557 31637 21591
rect 31671 21557 31683 21591
rect 31990 21588 31996 21600
rect 31951 21560 31996 21588
rect 31625 21551 31683 21557
rect 31640 21520 31668 21551
rect 31990 21548 31996 21560
rect 32048 21548 32054 21600
rect 32082 21548 32088 21600
rect 32140 21588 32146 21600
rect 32140 21560 32185 21588
rect 32140 21548 32146 21560
rect 30996 21492 31668 21520
rect 17270 21452 17276 21464
rect 17231 21424 17276 21452
rect 17270 21412 17276 21424
rect 17328 21412 17334 21464
rect 19113 21455 19171 21461
rect 19113 21421 19125 21455
rect 19159 21452 19171 21455
rect 19570 21452 19576 21464
rect 19159 21424 19576 21452
rect 19159 21421 19171 21424
rect 19113 21415 19171 21421
rect 19570 21412 19576 21424
rect 19628 21412 19634 21464
rect 21410 21412 21416 21464
rect 21468 21452 21474 21464
rect 24630 21452 24636 21464
rect 21468 21424 24636 21452
rect 21468 21412 21474 21424
rect 24630 21412 24636 21424
rect 24688 21412 24694 21464
rect 27942 21452 27948 21464
rect 27903 21424 27948 21452
rect 27942 21412 27948 21424
rect 28000 21412 28006 21464
rect 28589 21455 28647 21461
rect 28589 21421 28601 21455
rect 28635 21452 28647 21455
rect 30150 21452 30156 21464
rect 28635 21424 30156 21452
rect 28635 21421 28647 21424
rect 28589 21415 28647 21421
rect 30150 21412 30156 21424
rect 30208 21412 30214 21464
rect 11000 21362 34368 21384
rect 11000 21310 19142 21362
rect 19194 21310 19206 21362
rect 19258 21310 19270 21362
rect 19322 21310 19334 21362
rect 19386 21310 29142 21362
rect 29194 21310 29206 21362
rect 29258 21310 29270 21362
rect 29322 21310 29334 21362
rect 29386 21310 34368 21362
rect 11000 21288 34368 21310
rect 18285 21251 18343 21257
rect 18285 21217 18297 21251
rect 18331 21248 18343 21251
rect 20490 21248 20496 21260
rect 18331 21220 20496 21248
rect 18331 21217 18343 21220
rect 18285 21211 18343 21217
rect 20490 21208 20496 21220
rect 20548 21208 20554 21260
rect 21137 21251 21195 21257
rect 21137 21217 21149 21251
rect 21183 21217 21195 21251
rect 21137 21211 21195 21217
rect 17549 21183 17607 21189
rect 17549 21180 17561 21183
rect 15816 21152 17561 21180
rect 15816 21121 15844 21152
rect 17549 21149 17561 21152
rect 17595 21180 17607 21183
rect 17822 21180 17828 21192
rect 17595 21152 17828 21180
rect 17595 21149 17607 21152
rect 17549 21143 17607 21149
rect 17822 21140 17828 21152
rect 17880 21140 17886 21192
rect 18006 21180 18012 21192
rect 17967 21152 18012 21180
rect 18006 21140 18012 21152
rect 18064 21140 18070 21192
rect 18098 21140 18104 21192
rect 18156 21180 18162 21192
rect 18377 21183 18435 21189
rect 18377 21180 18389 21183
rect 18156 21152 18389 21180
rect 18156 21140 18162 21152
rect 18377 21149 18389 21152
rect 18423 21149 18435 21183
rect 19570 21180 19576 21192
rect 19531 21152 19576 21180
rect 18377 21143 18435 21149
rect 19570 21140 19576 21152
rect 19628 21140 19634 21192
rect 21152 21180 21180 21211
rect 22606 21208 22612 21260
rect 22664 21248 22670 21260
rect 22793 21251 22851 21257
rect 22793 21248 22805 21251
rect 22664 21220 22805 21248
rect 22664 21208 22670 21220
rect 22793 21217 22805 21220
rect 22839 21217 22851 21251
rect 22793 21211 22851 21217
rect 28494 21208 28500 21260
rect 28552 21248 28558 21260
rect 28773 21251 28831 21257
rect 28773 21248 28785 21251
rect 28552 21220 28785 21248
rect 28552 21208 28558 21220
rect 28773 21217 28785 21220
rect 28819 21217 28831 21251
rect 28773 21211 28831 21217
rect 21152 21152 22376 21180
rect 15801 21115 15859 21121
rect 15801 21081 15813 21115
rect 15847 21081 15859 21115
rect 16166 21112 16172 21124
rect 16127 21084 16172 21112
rect 15801 21075 15859 21081
rect 16166 21072 16172 21084
rect 16224 21072 16230 21124
rect 16353 21115 16411 21121
rect 16353 21081 16365 21115
rect 16399 21081 16411 21115
rect 16353 21075 16411 21081
rect 15893 21047 15951 21053
rect 15893 21013 15905 21047
rect 15939 21044 15951 21047
rect 15982 21044 15988 21056
rect 15939 21016 15988 21044
rect 15939 21013 15951 21016
rect 15893 21007 15951 21013
rect 15982 21004 15988 21016
rect 16040 21004 16046 21056
rect 16074 21004 16080 21056
rect 16132 21044 16138 21056
rect 16368 21044 16396 21075
rect 16442 21072 16448 21124
rect 16500 21112 16506 21124
rect 16905 21115 16963 21121
rect 16905 21112 16917 21115
rect 16500 21084 16917 21112
rect 16500 21072 16506 21084
rect 16905 21081 16917 21084
rect 16951 21081 16963 21115
rect 16905 21075 16963 21081
rect 17914 21072 17920 21124
rect 17972 21112 17978 21124
rect 18193 21115 18251 21121
rect 18193 21112 18205 21115
rect 17972 21084 18205 21112
rect 17972 21072 17978 21084
rect 18193 21081 18205 21084
rect 18239 21081 18251 21115
rect 19754 21112 19760 21124
rect 19715 21084 19760 21112
rect 18193 21075 18251 21081
rect 19754 21072 19760 21084
rect 19812 21072 19818 21124
rect 21042 21072 21048 21124
rect 21100 21112 21106 21124
rect 21505 21115 21563 21121
rect 21505 21112 21517 21115
rect 21100 21084 21517 21112
rect 21100 21072 21106 21084
rect 21505 21081 21517 21084
rect 21551 21081 21563 21115
rect 21873 21115 21931 21121
rect 21873 21112 21885 21115
rect 21505 21075 21563 21081
rect 21704 21084 21885 21112
rect 18006 21044 18012 21056
rect 16132 21016 18012 21044
rect 16132 21004 16138 21016
rect 18006 21004 18012 21016
rect 18064 21004 18070 21056
rect 18374 21004 18380 21056
rect 18432 21044 18438 21056
rect 18745 21047 18803 21053
rect 18745 21044 18757 21047
rect 18432 21016 18757 21044
rect 18432 21004 18438 21016
rect 18745 21013 18757 21016
rect 18791 21013 18803 21047
rect 21594 21044 21600 21056
rect 21555 21016 21600 21044
rect 18745 21007 18803 21013
rect 21594 21004 21600 21016
rect 21652 21004 21658 21056
rect 21410 20936 21416 20988
rect 21468 20976 21474 20988
rect 21704 20976 21732 21084
rect 21873 21081 21885 21084
rect 21919 21081 21931 21115
rect 21873 21075 21931 21081
rect 22057 21115 22115 21121
rect 22057 21081 22069 21115
rect 22103 21112 22115 21115
rect 22146 21112 22152 21124
rect 22103 21084 22152 21112
rect 22103 21081 22115 21084
rect 22057 21075 22115 21081
rect 22146 21072 22152 21084
rect 22204 21072 22210 21124
rect 22348 21044 22376 21152
rect 22422 21140 22428 21192
rect 22480 21180 22486 21192
rect 22517 21183 22575 21189
rect 22517 21180 22529 21183
rect 22480 21152 22529 21180
rect 22480 21140 22486 21152
rect 22517 21149 22529 21152
rect 22563 21149 22575 21183
rect 22517 21143 22575 21149
rect 27485 21183 27543 21189
rect 27485 21149 27497 21183
rect 27531 21180 27543 21183
rect 27758 21180 27764 21192
rect 27531 21152 27764 21180
rect 27531 21149 27543 21152
rect 27485 21143 27543 21149
rect 27758 21140 27764 21152
rect 27816 21140 27822 21192
rect 27850 21140 27856 21192
rect 27908 21180 27914 21192
rect 28037 21183 28095 21189
rect 28037 21180 28049 21183
rect 27908 21152 28049 21180
rect 27908 21140 27914 21152
rect 28037 21149 28049 21152
rect 28083 21149 28095 21183
rect 30150 21180 30156 21192
rect 30111 21152 30156 21180
rect 28037 21143 28095 21149
rect 30150 21140 30156 21152
rect 30208 21140 30214 21192
rect 22701 21115 22759 21121
rect 22701 21081 22713 21115
rect 22747 21112 22759 21115
rect 23342 21112 23348 21124
rect 22747 21084 23348 21112
rect 22747 21081 22759 21084
rect 22701 21075 22759 21081
rect 23342 21072 23348 21084
rect 23400 21072 23406 21124
rect 23802 21112 23808 21124
rect 23763 21084 23808 21112
rect 23802 21072 23808 21084
rect 23860 21072 23866 21124
rect 26565 21115 26623 21121
rect 26565 21112 26577 21115
rect 25016 21084 26577 21112
rect 25016 21044 25044 21084
rect 26565 21081 26577 21084
rect 26611 21112 26623 21115
rect 26838 21112 26844 21124
rect 26611 21084 26844 21112
rect 26611 21081 26623 21084
rect 26565 21075 26623 21081
rect 26838 21072 26844 21084
rect 26896 21072 26902 21124
rect 27298 21112 27304 21124
rect 27211 21084 27304 21112
rect 27298 21072 27304 21084
rect 27356 21112 27362 21124
rect 28681 21115 28739 21121
rect 28681 21112 28693 21115
rect 27356 21084 28693 21112
rect 27356 21072 27362 21084
rect 28681 21081 28693 21084
rect 28727 21081 28739 21115
rect 28681 21075 28739 21081
rect 29506 21072 29512 21124
rect 29564 21112 29570 21124
rect 29601 21115 29659 21121
rect 29601 21112 29613 21115
rect 29564 21084 29613 21112
rect 29564 21072 29570 21084
rect 29601 21081 29613 21084
rect 29647 21081 29659 21115
rect 30058 21112 30064 21124
rect 30019 21084 30064 21112
rect 29601 21075 29659 21081
rect 30058 21072 30064 21084
rect 30116 21072 30122 21124
rect 25182 21044 25188 21056
rect 22348 21016 25044 21044
rect 25143 21016 25188 21044
rect 25182 21004 25188 21016
rect 25240 21004 25246 21056
rect 25274 21004 25280 21056
rect 25332 21044 25338 21056
rect 25737 21047 25795 21053
rect 25737 21044 25749 21047
rect 25332 21016 25749 21044
rect 25332 21004 25338 21016
rect 25737 21013 25749 21016
rect 25783 21013 25795 21047
rect 25737 21007 25795 21013
rect 25642 20976 25648 20988
rect 21468 20948 21732 20976
rect 25603 20948 25648 20976
rect 21468 20936 21474 20948
rect 25642 20936 25648 20948
rect 25700 20936 25706 20988
rect 15338 20868 15344 20920
rect 15396 20908 15402 20920
rect 15433 20911 15491 20917
rect 15433 20908 15445 20911
rect 15396 20880 15445 20908
rect 15396 20868 15402 20880
rect 15433 20877 15445 20880
rect 15479 20877 15491 20911
rect 15433 20871 15491 20877
rect 15614 20868 15620 20920
rect 15672 20908 15678 20920
rect 17454 20908 17460 20920
rect 15672 20880 17460 20908
rect 15672 20868 15678 20880
rect 17454 20868 17460 20880
rect 17512 20908 17518 20920
rect 19849 20911 19907 20917
rect 19849 20908 19861 20911
rect 17512 20880 19861 20908
rect 17512 20868 17518 20880
rect 19849 20877 19861 20880
rect 19895 20877 19907 20911
rect 23986 20908 23992 20920
rect 23947 20880 23992 20908
rect 19849 20871 19907 20877
rect 23986 20868 23992 20880
rect 24044 20868 24050 20920
rect 26378 20868 26384 20920
rect 26436 20908 26442 20920
rect 28129 20911 28187 20917
rect 28129 20908 28141 20911
rect 26436 20880 28141 20908
rect 26436 20868 26442 20880
rect 28129 20877 28141 20880
rect 28175 20877 28187 20911
rect 28129 20871 28187 20877
rect 11000 20818 34368 20840
rect 11000 20766 14142 20818
rect 14194 20766 14206 20818
rect 14258 20766 14270 20818
rect 14322 20766 14334 20818
rect 14386 20766 24142 20818
rect 24194 20766 24206 20818
rect 24258 20766 24270 20818
rect 24322 20766 24334 20818
rect 24386 20766 34368 20818
rect 11000 20744 34368 20766
rect 22146 20664 22152 20716
rect 22204 20704 22210 20716
rect 22333 20707 22391 20713
rect 22333 20704 22345 20707
rect 22204 20676 22345 20704
rect 22204 20664 22210 20676
rect 22333 20673 22345 20676
rect 22379 20673 22391 20707
rect 22333 20667 22391 20673
rect 18006 20636 18012 20648
rect 17472 20608 18012 20636
rect 15522 20568 15528 20580
rect 15172 20540 15528 20568
rect 14970 20500 14976 20512
rect 14931 20472 14976 20500
rect 14970 20460 14976 20472
rect 15028 20460 15034 20512
rect 15172 20509 15200 20540
rect 15522 20528 15528 20540
rect 15580 20528 15586 20580
rect 15709 20571 15767 20577
rect 15709 20537 15721 20571
rect 15755 20568 15767 20571
rect 15982 20568 15988 20580
rect 15755 20540 15988 20568
rect 15755 20537 15767 20540
rect 15709 20531 15767 20537
rect 15982 20528 15988 20540
rect 16040 20568 16046 20580
rect 17472 20577 17500 20608
rect 18006 20596 18012 20608
rect 18064 20596 18070 20648
rect 24630 20596 24636 20648
rect 24688 20636 24694 20648
rect 27298 20636 27304 20648
rect 24688 20608 24860 20636
rect 27259 20608 27304 20636
rect 24688 20596 24694 20608
rect 17457 20571 17515 20577
rect 16040 20540 16856 20568
rect 16040 20528 16046 20540
rect 15157 20503 15215 20509
rect 15157 20469 15169 20503
rect 15203 20469 15215 20503
rect 15157 20463 15215 20469
rect 15246 20460 15252 20512
rect 15304 20500 15310 20512
rect 15341 20503 15399 20509
rect 15341 20500 15353 20503
rect 15304 20472 15353 20500
rect 15304 20460 15310 20472
rect 15341 20469 15353 20472
rect 15387 20469 15399 20503
rect 15341 20463 15399 20469
rect 14234 20392 14240 20444
rect 14292 20432 14298 20444
rect 14421 20435 14479 20441
rect 14421 20432 14433 20435
rect 14292 20404 14433 20432
rect 14292 20392 14298 20404
rect 14421 20401 14433 20404
rect 14467 20401 14479 20435
rect 15356 20432 15384 20463
rect 15614 20460 15620 20512
rect 15672 20500 15678 20512
rect 16828 20509 16856 20540
rect 17457 20537 17469 20571
rect 17503 20537 17515 20571
rect 17457 20531 17515 20537
rect 21410 20528 21416 20580
rect 21468 20528 21474 20580
rect 23710 20528 23716 20580
rect 23768 20568 23774 20580
rect 24722 20568 24728 20580
rect 23768 20540 24216 20568
rect 23768 20528 23774 20540
rect 15801 20503 15859 20509
rect 15801 20500 15813 20503
rect 15672 20472 15813 20500
rect 15672 20460 15678 20472
rect 15801 20469 15813 20472
rect 15847 20469 15859 20503
rect 15801 20463 15859 20469
rect 16813 20503 16871 20509
rect 16813 20469 16825 20503
rect 16859 20469 16871 20503
rect 18006 20500 18012 20512
rect 17967 20472 18012 20500
rect 16813 20463 16871 20469
rect 18006 20460 18012 20472
rect 18064 20460 18070 20512
rect 21134 20500 21140 20512
rect 21095 20472 21140 20500
rect 21134 20460 21140 20472
rect 21192 20500 21198 20512
rect 21428 20500 21456 20528
rect 21192 20472 21456 20500
rect 21192 20460 21198 20472
rect 21594 20460 21600 20512
rect 21652 20500 21658 20512
rect 21781 20503 21839 20509
rect 21781 20500 21793 20503
rect 21652 20472 21793 20500
rect 21652 20460 21658 20472
rect 21781 20469 21793 20472
rect 21827 20500 21839 20503
rect 22609 20503 22667 20509
rect 22609 20500 22621 20503
rect 21827 20472 22621 20500
rect 21827 20469 21839 20472
rect 21781 20463 21839 20469
rect 22609 20469 22621 20472
rect 22655 20469 22667 20503
rect 23986 20500 23992 20512
rect 23947 20472 23992 20500
rect 22609 20463 22667 20469
rect 23986 20460 23992 20472
rect 24044 20460 24050 20512
rect 24188 20509 24216 20540
rect 24464 20540 24728 20568
rect 24464 20509 24492 20540
rect 24722 20528 24728 20540
rect 24780 20528 24786 20580
rect 24832 20577 24860 20608
rect 27298 20596 27304 20608
rect 27356 20596 27362 20648
rect 29877 20639 29935 20645
rect 29877 20605 29889 20639
rect 29923 20636 29935 20639
rect 30242 20636 30248 20648
rect 29923 20608 30248 20636
rect 29923 20605 29935 20608
rect 29877 20599 29935 20605
rect 30242 20596 30248 20608
rect 30300 20596 30306 20648
rect 24817 20571 24875 20577
rect 24817 20537 24829 20571
rect 24863 20568 24875 20571
rect 24998 20568 25004 20580
rect 24863 20540 25004 20568
rect 24863 20537 24875 20540
rect 24817 20531 24875 20537
rect 24998 20528 25004 20540
rect 25056 20528 25062 20580
rect 26838 20568 26844 20580
rect 26799 20540 26844 20568
rect 26838 20528 26844 20540
rect 26896 20528 26902 20580
rect 27393 20571 27451 20577
rect 27393 20537 27405 20571
rect 27439 20568 27451 20571
rect 27942 20568 27948 20580
rect 27439 20540 27948 20568
rect 27439 20537 27451 20540
rect 27393 20531 27451 20537
rect 27942 20528 27948 20540
rect 28000 20528 28006 20580
rect 24173 20503 24231 20509
rect 24173 20469 24185 20503
rect 24219 20469 24231 20503
rect 24173 20463 24231 20469
rect 24449 20503 24507 20509
rect 24449 20469 24461 20503
rect 24495 20469 24507 20503
rect 24906 20500 24912 20512
rect 24867 20472 24912 20500
rect 24449 20463 24507 20469
rect 24906 20460 24912 20472
rect 24964 20460 24970 20512
rect 25461 20503 25519 20509
rect 25461 20469 25473 20503
rect 25507 20469 25519 20503
rect 26378 20500 26384 20512
rect 26339 20472 26384 20500
rect 25461 20463 25519 20469
rect 17270 20432 17276 20444
rect 15356 20404 17276 20432
rect 14421 20395 14479 20401
rect 17270 20392 17276 20404
rect 17328 20392 17334 20444
rect 18282 20432 18288 20444
rect 18243 20404 18288 20432
rect 18282 20392 18288 20404
rect 18340 20392 18346 20444
rect 19938 20432 19944 20444
rect 19510 20404 19944 20432
rect 19938 20392 19944 20404
rect 19996 20392 20002 20444
rect 20033 20435 20091 20441
rect 20033 20401 20045 20435
rect 20079 20401 20091 20435
rect 20033 20395 20091 20401
rect 19018 20324 19024 20376
rect 19076 20364 19082 20376
rect 20048 20364 20076 20395
rect 21410 20392 21416 20444
rect 21468 20432 21474 20444
rect 22517 20435 22575 20441
rect 22517 20432 22529 20435
rect 21468 20404 22529 20432
rect 21468 20392 21474 20404
rect 22517 20401 22529 20404
rect 22563 20401 22575 20435
rect 22517 20395 22575 20401
rect 23069 20435 23127 20441
rect 23069 20401 23081 20435
rect 23115 20401 23127 20435
rect 23069 20395 23127 20401
rect 23529 20435 23587 20441
rect 23529 20401 23541 20435
rect 23575 20432 23587 20435
rect 25182 20432 25188 20444
rect 23575 20404 25188 20432
rect 23575 20401 23587 20404
rect 23529 20395 23587 20401
rect 19076 20336 20076 20364
rect 23084 20364 23112 20395
rect 25182 20392 25188 20404
rect 25240 20432 25246 20444
rect 25476 20432 25504 20463
rect 26378 20460 26384 20472
rect 26436 20460 26442 20512
rect 25240 20404 25504 20432
rect 25240 20392 25246 20404
rect 25642 20392 25648 20444
rect 25700 20432 25706 20444
rect 26105 20435 26163 20441
rect 26105 20432 26117 20435
rect 25700 20404 26117 20432
rect 25700 20392 25706 20404
rect 26105 20401 26117 20404
rect 26151 20401 26163 20435
rect 26105 20395 26163 20401
rect 29598 20392 29604 20444
rect 29656 20432 29662 20444
rect 29693 20435 29751 20441
rect 29693 20432 29705 20435
rect 29656 20404 29705 20432
rect 29656 20392 29662 20404
rect 29693 20401 29705 20404
rect 29739 20401 29751 20435
rect 29693 20395 29751 20401
rect 23986 20364 23992 20376
rect 23084 20336 23992 20364
rect 19076 20324 19082 20336
rect 23986 20324 23992 20336
rect 24044 20324 24050 20376
rect 11000 20274 34368 20296
rect 11000 20222 19142 20274
rect 19194 20222 19206 20274
rect 19258 20222 19270 20274
rect 19322 20222 19334 20274
rect 19386 20222 29142 20274
rect 29194 20222 29206 20274
rect 29258 20222 29270 20274
rect 29322 20222 29334 20274
rect 29386 20222 34368 20274
rect 11000 20200 34368 20222
rect 14970 20120 14976 20172
rect 15028 20160 15034 20172
rect 16721 20163 16779 20169
rect 16721 20160 16733 20163
rect 15028 20132 16733 20160
rect 15028 20120 15034 20132
rect 16721 20129 16733 20132
rect 16767 20129 16779 20163
rect 16721 20123 16779 20129
rect 24449 20163 24507 20169
rect 24449 20129 24461 20163
rect 24495 20160 24507 20163
rect 25274 20160 25280 20172
rect 24495 20132 25280 20160
rect 24495 20129 24507 20132
rect 24449 20123 24507 20129
rect 25274 20120 25280 20132
rect 25332 20120 25338 20172
rect 28497 20163 28555 20169
rect 28497 20129 28509 20163
rect 28543 20160 28555 20163
rect 28543 20132 29644 20160
rect 28543 20129 28555 20132
rect 28497 20123 28555 20129
rect 14234 20092 14240 20104
rect 14195 20064 14240 20092
rect 14234 20052 14240 20064
rect 14292 20052 14298 20104
rect 14510 20052 14516 20104
rect 14568 20092 14574 20104
rect 15982 20092 15988 20104
rect 14568 20064 14726 20092
rect 15943 20064 15988 20092
rect 14568 20052 14574 20064
rect 15982 20052 15988 20064
rect 16040 20052 16046 20104
rect 19018 20092 19024 20104
rect 16644 20064 19024 20092
rect 13774 19984 13780 20036
rect 13832 20024 13838 20036
rect 13961 20027 14019 20033
rect 13961 20024 13973 20027
rect 13832 19996 13973 20024
rect 13832 19984 13838 19996
rect 13961 19993 13973 19996
rect 14007 19993 14019 20027
rect 13961 19987 14019 19993
rect 16445 20027 16503 20033
rect 16445 19993 16457 20027
rect 16491 19993 16503 20027
rect 16445 19987 16503 19993
rect 15338 19848 15344 19900
rect 15396 19888 15402 19900
rect 16460 19888 16488 19987
rect 16534 19984 16540 20036
rect 16592 20024 16598 20036
rect 16644 20033 16672 20064
rect 19018 20052 19024 20064
rect 19076 20052 19082 20104
rect 26841 20095 26899 20101
rect 24648 20064 26424 20092
rect 16629 20027 16687 20033
rect 16629 20024 16641 20027
rect 16592 19996 16641 20024
rect 16592 19984 16598 19996
rect 16629 19993 16641 19996
rect 16675 19993 16687 20027
rect 16629 19987 16687 19993
rect 17270 19984 17276 20036
rect 17328 20024 17334 20036
rect 18009 20027 18067 20033
rect 18009 20024 18021 20027
rect 17328 19996 18021 20024
rect 17328 19984 17334 19996
rect 18009 19993 18021 19996
rect 18055 19993 18067 20027
rect 18558 20024 18564 20036
rect 18519 19996 18564 20024
rect 18009 19987 18067 19993
rect 18558 19984 18564 19996
rect 18616 19984 18622 20036
rect 21410 20024 21416 20036
rect 21371 19996 21416 20024
rect 21410 19984 21416 19996
rect 21468 19984 21474 20036
rect 22146 20024 22152 20036
rect 22107 19996 22152 20024
rect 22146 19984 22152 19996
rect 22204 19984 22210 20036
rect 23621 20027 23679 20033
rect 23621 19993 23633 20027
rect 23667 20024 23679 20027
rect 23894 20024 23900 20036
rect 23667 19996 23900 20024
rect 23667 19993 23679 19996
rect 23621 19987 23679 19993
rect 23894 19984 23900 19996
rect 23952 19984 23958 20036
rect 24648 20033 24676 20064
rect 26396 20036 26424 20064
rect 26841 20061 26853 20095
rect 26887 20092 26899 20095
rect 27758 20092 27764 20104
rect 26887 20064 27764 20092
rect 26887 20061 26899 20064
rect 26841 20055 26899 20061
rect 27758 20052 27764 20064
rect 27816 20052 27822 20104
rect 29616 20036 29644 20132
rect 24633 20027 24691 20033
rect 24633 19993 24645 20027
rect 24679 19993 24691 20027
rect 24633 19987 24691 19993
rect 25090 19984 25096 20036
rect 25148 20024 25154 20036
rect 25277 20027 25335 20033
rect 25277 20024 25289 20027
rect 25148 19996 25289 20024
rect 25148 19984 25154 19996
rect 25277 19993 25289 19996
rect 25323 19993 25335 20027
rect 26378 20024 26384 20036
rect 26339 19996 26384 20024
rect 25277 19987 25335 19993
rect 26378 19984 26384 19996
rect 26436 19984 26442 20036
rect 27298 20024 27304 20036
rect 27259 19996 27304 20024
rect 27298 19984 27304 19996
rect 27356 19984 27362 20036
rect 27485 20027 27543 20033
rect 27485 19993 27497 20027
rect 27531 19993 27543 20027
rect 29598 20024 29604 20036
rect 29559 19996 29604 20024
rect 27485 19987 27543 19993
rect 17825 19959 17883 19965
rect 17825 19925 17837 19959
rect 17871 19956 17883 19959
rect 17914 19956 17920 19968
rect 17871 19928 17920 19956
rect 17871 19925 17883 19928
rect 17825 19919 17883 19925
rect 17914 19916 17920 19928
rect 17972 19916 17978 19968
rect 21781 19959 21839 19965
rect 21781 19925 21793 19959
rect 21827 19956 21839 19959
rect 27500 19956 27528 19987
rect 29598 19984 29604 19996
rect 29656 19984 29662 20036
rect 28129 19959 28187 19965
rect 28129 19956 28141 19959
rect 21827 19928 28141 19956
rect 21827 19925 21839 19928
rect 21781 19919 21839 19925
rect 28129 19925 28141 19928
rect 28175 19925 28187 19959
rect 28129 19919 28187 19925
rect 15396 19860 16488 19888
rect 15396 19848 15402 19860
rect 18282 19848 18288 19900
rect 18340 19888 18346 19900
rect 18469 19891 18527 19897
rect 18469 19888 18481 19891
rect 18340 19860 18481 19888
rect 18340 19848 18346 19860
rect 18469 19857 18481 19860
rect 18515 19857 18527 19891
rect 18469 19851 18527 19857
rect 27669 19891 27727 19897
rect 27669 19857 27681 19891
rect 27715 19888 27727 19891
rect 27942 19888 27948 19900
rect 27715 19860 27948 19888
rect 27715 19857 27727 19860
rect 27669 19851 27727 19857
rect 27942 19848 27948 19860
rect 28000 19848 28006 19900
rect 28494 19888 28500 19900
rect 28455 19860 28500 19888
rect 28494 19848 28500 19860
rect 28552 19848 28558 19900
rect 23250 19820 23256 19832
rect 23211 19792 23256 19820
rect 23250 19780 23256 19792
rect 23308 19780 23314 19832
rect 29690 19820 29696 19832
rect 29651 19792 29696 19820
rect 29690 19780 29696 19792
rect 29748 19780 29754 19832
rect 11000 19730 34368 19752
rect 11000 19678 14142 19730
rect 14194 19678 14206 19730
rect 14258 19678 14270 19730
rect 14322 19678 14334 19730
rect 14386 19678 24142 19730
rect 24194 19678 24206 19730
rect 24258 19678 24270 19730
rect 24322 19678 24334 19730
rect 24386 19678 34368 19730
rect 11000 19656 34368 19678
rect 14510 19616 14516 19628
rect 14471 19588 14516 19616
rect 14510 19576 14516 19588
rect 14568 19576 14574 19628
rect 17914 19616 17920 19628
rect 17875 19588 17920 19616
rect 17914 19576 17920 19588
rect 17972 19576 17978 19628
rect 18558 19576 18564 19628
rect 18616 19616 18622 19628
rect 19113 19619 19171 19625
rect 19113 19616 19125 19619
rect 18616 19588 19125 19616
rect 18616 19576 18622 19588
rect 19113 19585 19125 19588
rect 19159 19585 19171 19619
rect 19113 19579 19171 19585
rect 19938 19576 19944 19628
rect 19996 19616 20002 19628
rect 20033 19619 20091 19625
rect 20033 19616 20045 19619
rect 19996 19588 20045 19616
rect 19996 19576 20002 19588
rect 20033 19585 20045 19588
rect 20079 19585 20091 19619
rect 20033 19579 20091 19585
rect 29233 19551 29291 19557
rect 29233 19517 29245 19551
rect 29279 19548 29291 19551
rect 29598 19548 29604 19560
rect 29279 19520 29604 19548
rect 29279 19517 29291 19520
rect 29233 19511 29291 19517
rect 29598 19508 29604 19520
rect 29656 19508 29662 19560
rect 15522 19480 15528 19492
rect 15483 19452 15528 19480
rect 15522 19440 15528 19452
rect 15580 19440 15586 19492
rect 25001 19483 25059 19489
rect 25001 19449 25013 19483
rect 25047 19480 25059 19483
rect 26105 19483 26163 19489
rect 26105 19480 26117 19483
rect 25047 19452 26117 19480
rect 25047 19449 25059 19452
rect 25001 19443 25059 19449
rect 26105 19449 26117 19452
rect 26151 19449 26163 19483
rect 26105 19443 26163 19449
rect 14329 19415 14387 19421
rect 14329 19381 14341 19415
rect 14375 19412 14387 19415
rect 14602 19412 14608 19424
rect 14375 19384 14608 19412
rect 14375 19381 14387 19384
rect 14329 19375 14387 19381
rect 14602 19372 14608 19384
rect 14660 19372 14666 19424
rect 15338 19412 15344 19424
rect 15299 19384 15344 19412
rect 15338 19372 15344 19384
rect 15396 19372 15402 19424
rect 15893 19415 15951 19421
rect 15893 19381 15905 19415
rect 15939 19412 15951 19415
rect 16534 19412 16540 19424
rect 15939 19384 16540 19412
rect 15939 19381 15951 19384
rect 15893 19375 15951 19381
rect 16534 19372 16540 19384
rect 16592 19372 16598 19424
rect 18285 19415 18343 19421
rect 18285 19381 18297 19415
rect 18331 19412 18343 19415
rect 19018 19412 19024 19424
rect 18331 19384 19024 19412
rect 18331 19381 18343 19384
rect 18285 19375 18343 19381
rect 19018 19372 19024 19384
rect 19076 19372 19082 19424
rect 19570 19372 19576 19424
rect 19628 19412 19634 19424
rect 19849 19415 19907 19421
rect 19849 19412 19861 19415
rect 19628 19384 19861 19412
rect 19628 19372 19634 19384
rect 19849 19381 19861 19384
rect 19895 19381 19907 19415
rect 19849 19375 19907 19381
rect 22238 19372 22244 19424
rect 22296 19412 22302 19424
rect 22333 19415 22391 19421
rect 22333 19412 22345 19415
rect 22296 19384 22345 19412
rect 22296 19372 22302 19384
rect 22333 19381 22345 19384
rect 22379 19381 22391 19415
rect 22514 19412 22520 19424
rect 22475 19384 22520 19412
rect 22333 19375 22391 19381
rect 22514 19372 22520 19384
rect 22572 19412 22578 19424
rect 23069 19415 23127 19421
rect 23069 19412 23081 19415
rect 22572 19384 23081 19412
rect 22572 19372 22578 19384
rect 23069 19381 23081 19384
rect 23115 19381 23127 19415
rect 23250 19412 23256 19424
rect 23211 19384 23256 19412
rect 23069 19375 23127 19381
rect 23250 19372 23256 19384
rect 23308 19372 23314 19424
rect 25090 19372 25096 19424
rect 25148 19412 25154 19424
rect 25553 19415 25611 19421
rect 25553 19412 25565 19415
rect 25148 19384 25565 19412
rect 25148 19372 25154 19384
rect 25553 19381 25565 19384
rect 25599 19381 25611 19415
rect 27942 19412 27948 19424
rect 27903 19384 27948 19412
rect 25553 19375 25611 19381
rect 27942 19372 27948 19384
rect 28000 19372 28006 19424
rect 28865 19415 28923 19421
rect 28865 19381 28877 19415
rect 28911 19381 28923 19415
rect 28865 19375 28923 19381
rect 18837 19347 18895 19353
rect 18837 19313 18849 19347
rect 18883 19344 18895 19347
rect 19754 19344 19760 19356
rect 18883 19316 19760 19344
rect 18883 19313 18895 19316
rect 18837 19307 18895 19313
rect 19754 19304 19760 19316
rect 19812 19304 19818 19356
rect 24909 19347 24967 19353
rect 24909 19313 24921 19347
rect 24955 19344 24967 19347
rect 25642 19344 25648 19356
rect 24955 19316 25648 19344
rect 24955 19313 24967 19316
rect 24909 19307 24967 19313
rect 25642 19304 25648 19316
rect 25700 19304 25706 19356
rect 26013 19347 26071 19353
rect 26013 19313 26025 19347
rect 26059 19344 26071 19347
rect 27758 19344 27764 19356
rect 26059 19316 27764 19344
rect 26059 19313 26071 19316
rect 26013 19307 26071 19313
rect 27758 19304 27764 19316
rect 27816 19344 27822 19356
rect 28880 19344 28908 19375
rect 29690 19372 29696 19424
rect 29748 19412 29754 19424
rect 30061 19415 30119 19421
rect 30061 19412 30073 19415
rect 29748 19384 30073 19412
rect 29748 19372 29754 19384
rect 30061 19381 30073 19384
rect 30107 19381 30119 19415
rect 30061 19375 30119 19381
rect 27816 19316 28908 19344
rect 29969 19347 30027 19353
rect 27816 19304 27822 19316
rect 29969 19313 29981 19347
rect 30015 19313 30027 19347
rect 29969 19307 30027 19313
rect 23342 19236 23348 19288
rect 23400 19276 23406 19288
rect 23529 19279 23587 19285
rect 23529 19276 23541 19279
rect 23400 19248 23541 19276
rect 23400 19236 23406 19248
rect 23529 19245 23541 19248
rect 23575 19245 23587 19279
rect 23529 19239 23587 19245
rect 23618 19236 23624 19288
rect 23676 19276 23682 19288
rect 29984 19276 30012 19307
rect 23676 19248 30012 19276
rect 23676 19236 23682 19248
rect 11000 19186 34368 19208
rect 11000 19134 19142 19186
rect 19194 19134 19206 19186
rect 19258 19134 19270 19186
rect 19322 19134 19334 19186
rect 19386 19134 29142 19186
rect 29194 19134 29206 19186
rect 29258 19134 29270 19186
rect 29322 19134 29334 19186
rect 29386 19134 34368 19186
rect 11000 19112 34368 19134
rect 23618 19072 23624 19084
rect 19956 19044 23624 19072
rect 18006 18964 18012 19016
rect 18064 19004 18070 19016
rect 19021 19007 19079 19013
rect 18064 18976 18696 19004
rect 18064 18964 18070 18976
rect 18285 18939 18343 18945
rect 18285 18905 18297 18939
rect 18331 18936 18343 18939
rect 18374 18936 18380 18948
rect 18331 18908 18380 18936
rect 18331 18905 18343 18908
rect 18285 18899 18343 18905
rect 18374 18896 18380 18908
rect 18432 18896 18438 18948
rect 18561 18939 18619 18945
rect 18561 18905 18573 18939
rect 18607 18905 18619 18939
rect 18668 18936 18696 18976
rect 19021 18973 19033 19007
rect 19067 19004 19079 19007
rect 19754 19004 19760 19016
rect 19067 18976 19760 19004
rect 19067 18973 19079 18976
rect 19021 18967 19079 18973
rect 19754 18964 19760 18976
rect 19812 18964 19818 19016
rect 19956 18945 19984 19044
rect 23618 19032 23624 19044
rect 23676 19032 23682 19084
rect 27206 19072 27212 19084
rect 26672 19044 27212 19072
rect 21778 19004 21784 19016
rect 21442 18976 21784 19004
rect 21778 18964 21784 18976
rect 21836 18964 21842 19016
rect 22514 18964 22520 19016
rect 22572 19004 22578 19016
rect 26672 19013 26700 19044
rect 27206 19032 27212 19044
rect 27264 19072 27270 19084
rect 27264 19044 27528 19072
rect 27264 19032 27270 19044
rect 26657 19007 26715 19013
rect 22572 18976 23204 19004
rect 22572 18964 22578 18976
rect 19941 18939 19999 18945
rect 19941 18936 19953 18939
rect 18668 18908 19953 18936
rect 18561 18899 18619 18905
rect 19941 18905 19953 18908
rect 19987 18905 19999 18939
rect 22425 18939 22483 18945
rect 22425 18936 22437 18939
rect 19941 18899 19999 18905
rect 22348 18908 22437 18936
rect 18576 18868 18604 18899
rect 18300 18840 18604 18868
rect 20217 18871 20275 18877
rect 18300 18812 18328 18840
rect 20217 18837 20229 18871
rect 20263 18868 20275 18871
rect 20950 18868 20956 18880
rect 20263 18840 20956 18868
rect 20263 18837 20275 18840
rect 20217 18831 20275 18837
rect 20950 18828 20956 18840
rect 21008 18828 21014 18880
rect 21502 18828 21508 18880
rect 21560 18868 21566 18880
rect 21965 18871 22023 18877
rect 21965 18868 21977 18871
rect 21560 18840 21977 18868
rect 21560 18828 21566 18840
rect 21965 18837 21977 18840
rect 22011 18868 22023 18871
rect 22238 18868 22244 18880
rect 22011 18840 22244 18868
rect 22011 18837 22023 18840
rect 21965 18831 22023 18837
rect 22238 18828 22244 18840
rect 22296 18868 22302 18880
rect 22348 18868 22376 18908
rect 22425 18905 22437 18908
rect 22471 18905 22483 18939
rect 23066 18936 23072 18948
rect 23027 18908 23072 18936
rect 22425 18899 22483 18905
rect 23066 18896 23072 18908
rect 23124 18896 23130 18948
rect 23176 18945 23204 18976
rect 26657 18973 26669 19007
rect 26703 18973 26715 19007
rect 26657 18967 26715 18973
rect 27298 18964 27304 19016
rect 27356 19004 27362 19016
rect 27393 19007 27451 19013
rect 27393 19004 27405 19007
rect 27356 18976 27405 19004
rect 27356 18964 27362 18976
rect 27393 18973 27405 18976
rect 27439 18973 27451 19007
rect 27500 19004 27528 19044
rect 28494 19032 28500 19084
rect 28552 19072 28558 19084
rect 28773 19075 28831 19081
rect 28773 19072 28785 19075
rect 28552 19044 28785 19072
rect 28552 19032 28558 19044
rect 28773 19041 28785 19044
rect 28819 19041 28831 19075
rect 28773 19035 28831 19041
rect 29417 19007 29475 19013
rect 29417 19004 29429 19007
rect 27500 18976 29429 19004
rect 27393 18967 27451 18973
rect 29417 18973 29429 18976
rect 29463 18973 29475 19007
rect 29417 18967 29475 18973
rect 23161 18939 23219 18945
rect 23161 18905 23173 18939
rect 23207 18905 23219 18939
rect 23894 18936 23900 18948
rect 23855 18908 23900 18936
rect 23161 18899 23219 18905
rect 23894 18896 23900 18908
rect 23952 18896 23958 18948
rect 23986 18896 23992 18948
rect 24044 18936 24050 18948
rect 24357 18939 24415 18945
rect 24357 18936 24369 18939
rect 24044 18908 24369 18936
rect 24044 18896 24050 18908
rect 24357 18905 24369 18908
rect 24403 18905 24415 18939
rect 24357 18899 24415 18905
rect 26286 18896 26292 18948
rect 26344 18936 26350 18948
rect 26749 18939 26807 18945
rect 26344 18908 26700 18936
rect 26344 18896 26350 18908
rect 22296 18840 22376 18868
rect 26197 18871 26255 18877
rect 22296 18828 22302 18840
rect 26197 18837 26209 18871
rect 26243 18868 26255 18871
rect 26470 18868 26476 18880
rect 26243 18840 26476 18868
rect 26243 18837 26255 18840
rect 26197 18831 26255 18837
rect 26470 18828 26476 18840
rect 26528 18828 26534 18880
rect 26672 18868 26700 18908
rect 26749 18905 26761 18939
rect 26795 18936 26807 18939
rect 28034 18936 28040 18948
rect 26795 18908 28040 18936
rect 26795 18905 26807 18908
rect 26749 18899 26807 18905
rect 28034 18896 28040 18908
rect 28092 18896 28098 18948
rect 28129 18939 28187 18945
rect 28129 18905 28141 18939
rect 28175 18936 28187 18939
rect 28770 18936 28776 18948
rect 28175 18908 28776 18936
rect 28175 18905 28187 18908
rect 28129 18899 28187 18905
rect 28770 18896 28776 18908
rect 28828 18896 28834 18948
rect 27301 18871 27359 18877
rect 27301 18868 27313 18871
rect 26672 18840 27313 18868
rect 27301 18837 27313 18840
rect 27347 18837 27359 18871
rect 27301 18831 27359 18837
rect 28221 18871 28279 18877
rect 28221 18837 28233 18871
rect 28267 18868 28279 18871
rect 30702 18868 30708 18880
rect 28267 18840 30708 18868
rect 28267 18837 28279 18840
rect 28221 18831 28279 18837
rect 30702 18828 30708 18840
rect 30760 18828 30766 18880
rect 18282 18760 18288 18812
rect 18340 18760 18346 18812
rect 18377 18803 18435 18809
rect 18377 18769 18389 18803
rect 18423 18769 18435 18803
rect 18377 18763 18435 18769
rect 18392 18732 18420 18763
rect 22517 18735 22575 18741
rect 22517 18732 22529 18735
rect 18392 18704 22529 18732
rect 22517 18701 22529 18704
rect 22563 18701 22575 18735
rect 22517 18695 22575 18701
rect 24446 18692 24452 18744
rect 24504 18732 24510 18744
rect 24541 18735 24599 18741
rect 24541 18732 24553 18735
rect 24504 18704 24553 18732
rect 24504 18692 24510 18704
rect 24541 18701 24553 18704
rect 24587 18701 24599 18735
rect 29506 18732 29512 18744
rect 29467 18704 29512 18732
rect 24541 18695 24599 18701
rect 29506 18692 29512 18704
rect 29564 18692 29570 18744
rect 11000 18642 34368 18664
rect 11000 18590 14142 18642
rect 14194 18590 14206 18642
rect 14258 18590 14270 18642
rect 14322 18590 14334 18642
rect 14386 18590 24142 18642
rect 24194 18590 24206 18642
rect 24258 18590 24270 18642
rect 24322 18590 24334 18642
rect 24386 18590 34368 18642
rect 11000 18568 34368 18590
rect 13774 18488 13780 18540
rect 13832 18528 13838 18540
rect 18006 18528 18012 18540
rect 13832 18500 18012 18528
rect 13832 18488 13838 18500
rect 17656 18392 17684 18500
rect 18006 18488 18012 18500
rect 18064 18488 18070 18540
rect 20861 18531 20919 18537
rect 20861 18497 20873 18531
rect 20907 18528 20919 18531
rect 20950 18528 20956 18540
rect 20907 18500 20956 18528
rect 20907 18497 20919 18500
rect 20861 18491 20919 18497
rect 20950 18488 20956 18500
rect 21008 18488 21014 18540
rect 21612 18500 21916 18528
rect 21612 18460 21640 18500
rect 21888 18472 21916 18500
rect 21778 18460 21784 18472
rect 20600 18432 21640 18460
rect 21739 18432 21784 18460
rect 17733 18395 17791 18401
rect 17733 18392 17745 18395
rect 17656 18364 17745 18392
rect 17733 18361 17745 18364
rect 17779 18361 17791 18395
rect 17733 18355 17791 18361
rect 18374 18352 18380 18404
rect 18432 18392 18438 18404
rect 19757 18395 19815 18401
rect 19757 18392 19769 18395
rect 18432 18364 19769 18392
rect 18432 18352 18438 18364
rect 19757 18361 19769 18364
rect 19803 18361 19815 18395
rect 19757 18355 19815 18361
rect 14421 18327 14479 18333
rect 14421 18293 14433 18327
rect 14467 18324 14479 18327
rect 14602 18324 14608 18336
rect 14467 18296 14608 18324
rect 14467 18293 14479 18296
rect 14421 18287 14479 18293
rect 14602 18284 14608 18296
rect 14660 18284 14666 18336
rect 15801 18327 15859 18333
rect 15801 18293 15813 18327
rect 15847 18324 15859 18327
rect 15982 18324 15988 18336
rect 15847 18296 15988 18324
rect 15847 18293 15859 18296
rect 15801 18287 15859 18293
rect 15982 18284 15988 18296
rect 16040 18284 16046 18336
rect 14620 18256 14648 18284
rect 16902 18256 16908 18268
rect 14620 18228 16908 18256
rect 16902 18216 16908 18228
rect 16960 18216 16966 18268
rect 18006 18256 18012 18268
rect 17967 18228 18012 18256
rect 18006 18216 18012 18228
rect 18064 18216 18070 18268
rect 19662 18256 19668 18268
rect 19234 18228 19668 18256
rect 19662 18216 19668 18228
rect 19720 18216 19726 18268
rect 19846 18216 19852 18268
rect 19904 18256 19910 18268
rect 20600 18265 20628 18432
rect 21778 18420 21784 18432
rect 21836 18420 21842 18472
rect 21870 18420 21876 18472
rect 21928 18420 21934 18472
rect 28405 18463 28463 18469
rect 28405 18429 28417 18463
rect 28451 18460 28463 18463
rect 29598 18460 29604 18472
rect 28451 18432 29604 18460
rect 28451 18429 28463 18432
rect 28405 18423 28463 18429
rect 29598 18420 29604 18432
rect 29656 18420 29662 18472
rect 20858 18352 20864 18404
rect 20916 18392 20922 18404
rect 23342 18392 23348 18404
rect 20916 18364 21640 18392
rect 23303 18364 23348 18392
rect 20916 18352 20922 18364
rect 20769 18327 20827 18333
rect 20769 18293 20781 18327
rect 20815 18324 20827 18327
rect 21502 18324 21508 18336
rect 20815 18296 21508 18324
rect 20815 18293 20827 18296
rect 20769 18287 20827 18293
rect 21502 18284 21508 18296
rect 21560 18284 21566 18336
rect 21612 18333 21640 18364
rect 23342 18352 23348 18364
rect 23400 18352 23406 18404
rect 23894 18352 23900 18404
rect 23952 18392 23958 18404
rect 25093 18395 25151 18401
rect 25093 18392 25105 18395
rect 23952 18364 25105 18392
rect 23952 18352 23958 18364
rect 25093 18361 25105 18364
rect 25139 18361 25151 18395
rect 25093 18355 25151 18361
rect 27298 18352 27304 18404
rect 27356 18392 27362 18404
rect 27945 18395 28003 18401
rect 27945 18392 27957 18395
rect 27356 18364 27957 18392
rect 27356 18352 27362 18364
rect 27945 18361 27957 18364
rect 27991 18361 28003 18395
rect 27945 18355 28003 18361
rect 28497 18395 28555 18401
rect 28497 18361 28509 18395
rect 28543 18392 28555 18395
rect 29506 18392 29512 18404
rect 28543 18364 29512 18392
rect 28543 18361 28555 18364
rect 28497 18355 28555 18361
rect 29506 18352 29512 18364
rect 29564 18352 29570 18404
rect 21597 18327 21655 18333
rect 21597 18293 21609 18327
rect 21643 18293 21655 18327
rect 21597 18287 21655 18293
rect 21870 18284 21876 18336
rect 21928 18324 21934 18336
rect 22514 18324 22520 18336
rect 21928 18296 22520 18324
rect 21928 18284 21934 18296
rect 22514 18284 22520 18296
rect 22572 18284 22578 18336
rect 23069 18327 23127 18333
rect 23069 18293 23081 18327
rect 23115 18293 23127 18327
rect 23069 18287 23127 18293
rect 20585 18259 20643 18265
rect 20585 18256 20597 18259
rect 19904 18228 20597 18256
rect 19904 18216 19910 18228
rect 20585 18225 20597 18228
rect 20631 18225 20643 18259
rect 23084 18256 23112 18287
rect 24446 18284 24452 18336
rect 24504 18284 24510 18336
rect 26470 18324 26476 18336
rect 26431 18296 26476 18324
rect 26470 18284 26476 18296
rect 26528 18284 26534 18336
rect 27206 18324 27212 18336
rect 27167 18296 27212 18324
rect 27206 18284 27212 18296
rect 27264 18284 27270 18336
rect 27393 18327 27451 18333
rect 27393 18293 27405 18327
rect 27439 18324 27451 18327
rect 27758 18324 27764 18336
rect 27439 18296 27764 18324
rect 27439 18293 27451 18296
rect 27393 18287 27451 18293
rect 27758 18284 27764 18296
rect 27816 18284 27822 18336
rect 23618 18256 23624 18268
rect 23084 18228 23624 18256
rect 20585 18219 20643 18225
rect 23618 18216 23624 18228
rect 23676 18216 23682 18268
rect 14605 18191 14663 18197
rect 14605 18157 14617 18191
rect 14651 18188 14663 18191
rect 14694 18188 14700 18200
rect 14651 18160 14700 18188
rect 14651 18157 14663 18160
rect 14605 18151 14663 18157
rect 14694 18148 14700 18160
rect 14752 18148 14758 18200
rect 15614 18188 15620 18200
rect 15575 18160 15620 18188
rect 15614 18148 15620 18160
rect 15672 18148 15678 18200
rect 16920 18188 16948 18216
rect 19570 18188 19576 18200
rect 16920 18160 19576 18188
rect 19570 18148 19576 18160
rect 19628 18148 19634 18200
rect 20858 18148 20864 18200
rect 20916 18188 20922 18200
rect 23986 18188 23992 18200
rect 20916 18160 23992 18188
rect 20916 18148 20922 18160
rect 23986 18148 23992 18160
rect 24044 18148 24050 18200
rect 11000 18098 34368 18120
rect 11000 18046 19142 18098
rect 19194 18046 19206 18098
rect 19258 18046 19270 18098
rect 19322 18046 19334 18098
rect 19386 18046 29142 18098
rect 29194 18046 29206 18098
rect 29258 18046 29270 18098
rect 29322 18046 29334 18098
rect 29386 18046 34368 18098
rect 11000 18024 34368 18046
rect 19662 17944 19668 17996
rect 19720 17984 19726 17996
rect 21137 17987 21195 17993
rect 21137 17984 21149 17987
rect 19720 17956 21149 17984
rect 19720 17944 19726 17956
rect 21137 17953 21149 17956
rect 21183 17953 21195 17987
rect 21137 17947 21195 17953
rect 28034 17944 28040 17996
rect 28092 17984 28098 17996
rect 28129 17987 28187 17993
rect 28129 17984 28141 17987
rect 28092 17956 28141 17984
rect 28092 17944 28098 17956
rect 28129 17953 28141 17956
rect 28175 17953 28187 17987
rect 28129 17947 28187 17953
rect 14694 17876 14700 17928
rect 14752 17876 14758 17928
rect 15982 17916 15988 17928
rect 15943 17888 15988 17916
rect 15982 17876 15988 17888
rect 16040 17916 16046 17928
rect 16040 17888 16488 17916
rect 16040 17876 16046 17888
rect 13774 17808 13780 17860
rect 13832 17848 13838 17860
rect 16460 17857 16488 17888
rect 16644 17888 18788 17916
rect 16644 17857 16672 17888
rect 17196 17857 17224 17888
rect 13961 17851 14019 17857
rect 13961 17848 13973 17851
rect 13832 17820 13973 17848
rect 13832 17808 13838 17820
rect 13961 17817 13973 17820
rect 14007 17817 14019 17851
rect 13961 17811 14019 17817
rect 16445 17851 16503 17857
rect 16445 17817 16457 17851
rect 16491 17817 16503 17851
rect 16445 17811 16503 17817
rect 16629 17851 16687 17857
rect 16629 17817 16641 17851
rect 16675 17817 16687 17851
rect 16629 17811 16687 17817
rect 17181 17851 17239 17857
rect 17181 17817 17193 17851
rect 17227 17848 17239 17851
rect 17365 17851 17423 17857
rect 17227 17820 17261 17848
rect 17227 17817 17239 17820
rect 17181 17811 17239 17817
rect 17365 17817 17377 17851
rect 17411 17848 17423 17851
rect 18374 17848 18380 17860
rect 17411 17820 17960 17848
rect 18335 17820 18380 17848
rect 17411 17817 17423 17820
rect 17365 17811 17423 17817
rect 17932 17792 17960 17820
rect 18374 17808 18380 17820
rect 18432 17808 18438 17860
rect 18760 17792 18788 17888
rect 19570 17876 19576 17928
rect 19628 17916 19634 17928
rect 20858 17916 20864 17928
rect 19628 17888 20864 17916
rect 19628 17876 19634 17888
rect 20858 17876 20864 17888
rect 20916 17916 20922 17928
rect 20916 17888 20996 17916
rect 20916 17876 20922 17888
rect 19846 17848 19852 17860
rect 19807 17820 19852 17848
rect 19846 17808 19852 17820
rect 19904 17808 19910 17860
rect 20968 17857 20996 17888
rect 26470 17876 26476 17928
rect 26528 17916 26534 17928
rect 26749 17919 26807 17925
rect 26749 17916 26761 17919
rect 26528 17888 26761 17916
rect 26528 17876 26534 17888
rect 26749 17885 26761 17888
rect 26795 17885 26807 17919
rect 28402 17916 28408 17928
rect 26749 17879 26807 17885
rect 27408 17888 28408 17916
rect 20953 17851 21011 17857
rect 20953 17817 20965 17851
rect 20999 17817 21011 17851
rect 20953 17811 21011 17817
rect 22422 17808 22428 17860
rect 22480 17848 22486 17860
rect 22517 17851 22575 17857
rect 22517 17848 22529 17851
rect 22480 17820 22529 17848
rect 22480 17808 22486 17820
rect 22517 17817 22529 17820
rect 22563 17848 22575 17851
rect 23069 17851 23127 17857
rect 23069 17848 23081 17851
rect 22563 17820 23081 17848
rect 22563 17817 22575 17820
rect 22517 17811 22575 17817
rect 23069 17817 23081 17820
rect 23115 17817 23127 17851
rect 23250 17848 23256 17860
rect 23211 17820 23256 17848
rect 23069 17811 23127 17817
rect 23250 17808 23256 17820
rect 23308 17808 23314 17860
rect 23986 17808 23992 17860
rect 24044 17848 24050 17860
rect 24449 17851 24507 17857
rect 24449 17848 24461 17851
rect 24044 17820 24461 17848
rect 24044 17808 24050 17820
rect 24449 17817 24461 17820
rect 24495 17817 24507 17851
rect 24449 17811 24507 17817
rect 26657 17851 26715 17857
rect 26657 17817 26669 17851
rect 26703 17848 26715 17851
rect 27408 17848 27436 17888
rect 28402 17876 28408 17888
rect 28460 17876 28466 17928
rect 26703 17820 27436 17848
rect 27485 17851 27543 17857
rect 26703 17817 26715 17820
rect 26657 17811 26715 17817
rect 27485 17817 27497 17851
rect 27531 17817 27543 17851
rect 27485 17811 27543 17817
rect 14237 17783 14295 17789
rect 14237 17749 14249 17783
rect 14283 17780 14295 17783
rect 14283 17752 15936 17780
rect 14283 17749 14295 17752
rect 14237 17743 14295 17749
rect 15908 17712 15936 17752
rect 17914 17740 17920 17792
rect 17972 17780 17978 17792
rect 18285 17783 18343 17789
rect 18285 17780 18297 17783
rect 17972 17752 18297 17780
rect 17972 17740 17978 17752
rect 18285 17749 18297 17752
rect 18331 17749 18343 17783
rect 18285 17743 18343 17749
rect 18742 17740 18748 17792
rect 18800 17780 18806 17792
rect 19757 17783 19815 17789
rect 19757 17780 19769 17783
rect 18800 17752 19769 17780
rect 18800 17740 18806 17752
rect 19757 17749 19769 17752
rect 19803 17749 19815 17783
rect 19757 17743 19815 17749
rect 22330 17740 22336 17792
rect 22388 17780 22394 17792
rect 22388 17752 22433 17780
rect 22388 17740 22394 17752
rect 24998 17740 25004 17792
rect 25056 17780 25062 17792
rect 27500 17780 27528 17811
rect 27758 17808 27764 17860
rect 27816 17848 27822 17860
rect 28313 17851 28371 17857
rect 28313 17848 28325 17851
rect 27816 17820 28325 17848
rect 27816 17808 27822 17820
rect 28313 17817 28325 17820
rect 28359 17817 28371 17851
rect 28313 17811 28371 17817
rect 25056 17752 27528 17780
rect 27577 17783 27635 17789
rect 25056 17740 25062 17752
rect 27577 17749 27589 17783
rect 27623 17780 27635 17783
rect 28954 17780 28960 17792
rect 27623 17752 28960 17780
rect 27623 17749 27635 17752
rect 27577 17743 27635 17749
rect 28954 17740 28960 17752
rect 29012 17740 29018 17792
rect 17549 17715 17607 17721
rect 17549 17712 17561 17715
rect 15908 17684 17561 17712
rect 17549 17681 17561 17684
rect 17595 17681 17607 17715
rect 17549 17675 17607 17681
rect 23529 17647 23587 17653
rect 23529 17613 23541 17647
rect 23575 17644 23587 17647
rect 23802 17644 23808 17656
rect 23575 17616 23808 17644
rect 23575 17613 23587 17616
rect 23529 17607 23587 17613
rect 23802 17604 23808 17616
rect 23860 17604 23866 17656
rect 24538 17604 24544 17656
rect 24596 17644 24602 17656
rect 24633 17647 24691 17653
rect 24633 17644 24645 17647
rect 24596 17616 24645 17644
rect 24596 17604 24602 17616
rect 24633 17613 24645 17616
rect 24679 17613 24691 17647
rect 24633 17607 24691 17613
rect 11000 17554 34368 17576
rect 11000 17502 14142 17554
rect 14194 17502 14206 17554
rect 14258 17502 14270 17554
rect 14322 17502 14334 17554
rect 14386 17502 24142 17554
rect 24194 17502 24206 17554
rect 24258 17502 24270 17554
rect 24322 17502 24334 17554
rect 24386 17502 34368 17554
rect 11000 17480 34368 17502
rect 15338 17400 15344 17452
rect 15396 17440 15402 17452
rect 17362 17440 17368 17452
rect 15396 17412 17368 17440
rect 15396 17400 15402 17412
rect 17362 17400 17368 17412
rect 17420 17400 17426 17452
rect 18006 17400 18012 17452
rect 18064 17440 18070 17452
rect 19941 17443 19999 17449
rect 19941 17440 19953 17443
rect 18064 17412 19953 17440
rect 18064 17400 18070 17412
rect 19941 17409 19953 17412
rect 19987 17409 19999 17443
rect 19941 17403 19999 17409
rect 22330 17400 22336 17452
rect 22388 17440 22394 17452
rect 23066 17440 23072 17452
rect 22388 17412 23072 17440
rect 22388 17400 22394 17412
rect 23066 17400 23072 17412
rect 23124 17440 23130 17452
rect 23124 17412 25596 17440
rect 23124 17400 23130 17412
rect 12394 17332 12400 17384
rect 12452 17372 12458 17384
rect 15893 17375 15951 17381
rect 15893 17372 15905 17375
rect 12452 17344 15905 17372
rect 12452 17332 12458 17344
rect 15893 17341 15905 17344
rect 15939 17341 15951 17375
rect 15893 17335 15951 17341
rect 18561 17375 18619 17381
rect 18561 17341 18573 17375
rect 18607 17372 18619 17375
rect 20766 17372 20772 17384
rect 18607 17344 20772 17372
rect 18607 17341 18619 17344
rect 18561 17335 18619 17341
rect 20766 17332 20772 17344
rect 20824 17332 20830 17384
rect 11937 17307 11995 17313
rect 11937 17273 11949 17307
rect 11983 17304 11995 17307
rect 12670 17304 12676 17316
rect 11983 17276 12676 17304
rect 11983 17273 11995 17276
rect 11937 17267 11995 17273
rect 12670 17264 12676 17276
rect 12728 17264 12734 17316
rect 16997 17307 17055 17313
rect 14988 17276 15200 17304
rect 12029 17239 12087 17245
rect 12029 17205 12041 17239
rect 12075 17236 12087 17239
rect 12394 17236 12400 17248
rect 12075 17208 12400 17236
rect 12075 17205 12087 17208
rect 12029 17199 12087 17205
rect 12394 17196 12400 17208
rect 12452 17196 12458 17248
rect 14988 17245 15016 17276
rect 14973 17239 15031 17245
rect 14973 17205 14985 17239
rect 15019 17205 15031 17239
rect 14973 17199 15031 17205
rect 15065 17239 15123 17245
rect 15065 17205 15077 17239
rect 15111 17205 15123 17239
rect 15172 17236 15200 17276
rect 16997 17273 17009 17307
rect 17043 17304 17055 17307
rect 21226 17304 21232 17316
rect 17043 17276 21232 17304
rect 17043 17273 17055 17276
rect 16997 17267 17055 17273
rect 21226 17264 21232 17276
rect 21284 17264 21290 17316
rect 23250 17264 23256 17316
rect 23308 17304 23314 17316
rect 23526 17304 23532 17316
rect 23308 17276 23532 17304
rect 23308 17264 23314 17276
rect 23526 17264 23532 17276
rect 23584 17264 23590 17316
rect 23802 17304 23808 17316
rect 23763 17276 23808 17304
rect 23802 17264 23808 17276
rect 23860 17264 23866 17316
rect 25568 17313 25596 17412
rect 25553 17307 25611 17313
rect 25553 17273 25565 17307
rect 25599 17273 25611 17307
rect 25553 17267 25611 17273
rect 15338 17236 15344 17248
rect 15172 17208 15344 17236
rect 15065 17199 15123 17205
rect 12486 17168 12492 17180
rect 12447 17140 12492 17168
rect 12486 17128 12492 17140
rect 12544 17128 12550 17180
rect 15080 17168 15108 17199
rect 15338 17196 15344 17208
rect 15396 17236 15402 17248
rect 15525 17239 15583 17245
rect 15525 17236 15537 17239
rect 15396 17208 15537 17236
rect 15396 17196 15402 17208
rect 15525 17205 15537 17208
rect 15571 17205 15583 17239
rect 15525 17199 15583 17205
rect 15709 17239 15767 17245
rect 15709 17205 15721 17239
rect 15755 17236 15767 17239
rect 16718 17236 16724 17248
rect 15755 17208 16724 17236
rect 15755 17205 15767 17208
rect 15709 17199 15767 17205
rect 15724 17168 15752 17199
rect 16718 17196 16724 17208
rect 16776 17236 16782 17248
rect 17181 17239 17239 17245
rect 17181 17236 17193 17239
rect 16776 17208 17193 17236
rect 16776 17196 16782 17208
rect 17181 17205 17193 17208
rect 17227 17205 17239 17239
rect 17362 17236 17368 17248
rect 17323 17208 17368 17236
rect 17181 17199 17239 17205
rect 17362 17196 17368 17208
rect 17420 17196 17426 17248
rect 17733 17239 17791 17245
rect 17733 17205 17745 17239
rect 17779 17205 17791 17239
rect 17914 17236 17920 17248
rect 17875 17208 17920 17236
rect 17733 17199 17791 17205
rect 17748 17168 17776 17199
rect 17914 17196 17920 17208
rect 17972 17196 17978 17248
rect 18561 17239 18619 17245
rect 18561 17205 18573 17239
rect 18607 17236 18619 17239
rect 18653 17239 18711 17245
rect 18653 17236 18665 17239
rect 18607 17208 18665 17236
rect 18607 17205 18619 17208
rect 18561 17199 18619 17205
rect 18653 17205 18665 17208
rect 18699 17205 18711 17239
rect 18653 17199 18711 17205
rect 18745 17239 18803 17245
rect 18745 17205 18757 17239
rect 18791 17205 18803 17239
rect 18745 17199 18803 17205
rect 15080 17140 15752 17168
rect 16736 17140 17776 17168
rect 15614 17060 15620 17112
rect 15672 17100 15678 17112
rect 16736 17100 16764 17140
rect 18190 17128 18196 17180
rect 18248 17168 18254 17180
rect 18760 17168 18788 17199
rect 19478 17196 19484 17248
rect 19536 17236 19542 17248
rect 19849 17239 19907 17245
rect 19849 17236 19861 17239
rect 19536 17208 19861 17236
rect 19536 17196 19542 17208
rect 19849 17205 19861 17208
rect 19895 17205 19907 17239
rect 19849 17199 19907 17205
rect 18248 17140 18788 17168
rect 18248 17128 18254 17140
rect 19018 17128 19024 17180
rect 19076 17168 19082 17180
rect 19205 17171 19263 17177
rect 19205 17168 19217 17171
rect 19076 17140 19217 17168
rect 19076 17128 19082 17140
rect 19205 17137 19217 17140
rect 19251 17137 19263 17171
rect 19662 17168 19668 17180
rect 19623 17140 19668 17168
rect 19205 17131 19263 17137
rect 19662 17128 19668 17140
rect 19720 17128 19726 17180
rect 24538 17128 24544 17180
rect 24596 17128 24602 17180
rect 15672 17072 16764 17100
rect 15672 17060 15678 17072
rect 28954 17060 28960 17112
rect 29012 17100 29018 17112
rect 30610 17100 30616 17112
rect 29012 17072 30616 17100
rect 29012 17060 29018 17072
rect 30610 17060 30616 17072
rect 30668 17060 30674 17112
rect 11000 17010 34368 17032
rect 11000 16958 19142 17010
rect 19194 16958 19206 17010
rect 19258 16958 19270 17010
rect 19322 16958 19334 17010
rect 19386 16958 29142 17010
rect 29194 16958 29206 17010
rect 29258 16958 29270 17010
rect 29322 16958 29334 17010
rect 29386 16958 34368 17010
rect 11000 16936 34368 16958
rect 19849 16899 19907 16905
rect 19849 16896 19861 16899
rect 18300 16868 19861 16896
rect 12670 16828 12676 16840
rect 12136 16800 12676 16828
rect 12136 16769 12164 16800
rect 12670 16788 12676 16800
rect 12728 16788 12734 16840
rect 16718 16828 16724 16840
rect 15448 16800 16396 16828
rect 16679 16800 16724 16828
rect 12121 16763 12179 16769
rect 12121 16729 12133 16763
rect 12167 16729 12179 16763
rect 12394 16760 12400 16772
rect 12355 16732 12400 16760
rect 12121 16723 12179 16729
rect 12394 16720 12400 16732
rect 12452 16720 12458 16772
rect 15448 16769 15476 16800
rect 15433 16763 15491 16769
rect 15433 16729 15445 16763
rect 15479 16729 15491 16763
rect 15614 16760 15620 16772
rect 15575 16732 15620 16760
rect 15433 16723 15491 16729
rect 15614 16720 15620 16732
rect 15672 16760 15678 16772
rect 16368 16769 16396 16800
rect 16718 16788 16724 16800
rect 16776 16788 16782 16840
rect 18300 16837 18328 16868
rect 19849 16865 19861 16868
rect 19895 16865 19907 16899
rect 19849 16859 19907 16865
rect 18285 16831 18343 16837
rect 18285 16797 18297 16831
rect 18331 16797 18343 16831
rect 18742 16828 18748 16840
rect 18285 16791 18343 16797
rect 18392 16800 18748 16828
rect 16169 16763 16227 16769
rect 16169 16760 16181 16763
rect 15672 16732 16181 16760
rect 15672 16720 15678 16732
rect 16169 16729 16181 16732
rect 16215 16729 16227 16763
rect 16169 16723 16227 16729
rect 16353 16763 16411 16769
rect 16353 16729 16365 16763
rect 16399 16760 16411 16763
rect 17914 16760 17920 16772
rect 16399 16732 17920 16760
rect 16399 16729 16411 16732
rect 16353 16723 16411 16729
rect 17914 16720 17920 16732
rect 17972 16720 17978 16772
rect 18190 16760 18196 16772
rect 18151 16732 18196 16760
rect 18190 16720 18196 16732
rect 18248 16720 18254 16772
rect 18392 16769 18420 16800
rect 18742 16788 18748 16800
rect 18800 16788 18806 16840
rect 18837 16831 18895 16837
rect 18837 16797 18849 16831
rect 18883 16828 18895 16831
rect 19662 16828 19668 16840
rect 18883 16800 19668 16828
rect 18883 16797 18895 16800
rect 18837 16791 18895 16797
rect 19662 16788 19668 16800
rect 19720 16788 19726 16840
rect 21060 16800 23020 16828
rect 18377 16763 18435 16769
rect 18377 16729 18389 16763
rect 18423 16729 18435 16763
rect 18377 16723 18435 16729
rect 18466 16720 18472 16772
rect 18524 16760 18530 16772
rect 19573 16763 19631 16769
rect 19573 16760 19585 16763
rect 18524 16732 19585 16760
rect 18524 16720 18530 16732
rect 19573 16729 19585 16732
rect 19619 16729 19631 16763
rect 19573 16723 19631 16729
rect 19757 16763 19815 16769
rect 19757 16729 19769 16763
rect 19803 16729 19815 16763
rect 19757 16723 19815 16729
rect 12581 16695 12639 16701
rect 12581 16661 12593 16695
rect 12627 16692 12639 16695
rect 12762 16692 12768 16704
rect 12627 16664 12768 16692
rect 12627 16661 12639 16664
rect 12581 16655 12639 16661
rect 12762 16652 12768 16664
rect 12820 16652 12826 16704
rect 19772 16692 19800 16723
rect 20766 16720 20772 16772
rect 20824 16760 20830 16772
rect 21060 16769 21088 16800
rect 21045 16763 21103 16769
rect 21045 16760 21057 16763
rect 20824 16732 21057 16760
rect 20824 16720 20830 16732
rect 21045 16729 21057 16732
rect 21091 16729 21103 16763
rect 21045 16723 21103 16729
rect 21137 16763 21195 16769
rect 21137 16729 21149 16763
rect 21183 16729 21195 16763
rect 21137 16723 21195 16729
rect 22241 16763 22299 16769
rect 22241 16729 22253 16763
rect 22287 16760 22299 16763
rect 22422 16760 22428 16772
rect 22287 16732 22428 16760
rect 22287 16729 22299 16732
rect 22241 16723 22299 16729
rect 18392 16664 19800 16692
rect 18392 16636 18420 16664
rect 18374 16584 18380 16636
rect 18432 16584 18438 16636
rect 21152 16624 21180 16723
rect 22422 16720 22428 16732
rect 22480 16760 22486 16772
rect 22992 16769 23020 16800
rect 22793 16763 22851 16769
rect 22793 16760 22805 16763
rect 22480 16732 22805 16760
rect 22480 16720 22486 16732
rect 22793 16729 22805 16732
rect 22839 16729 22851 16763
rect 22793 16723 22851 16729
rect 22977 16763 23035 16769
rect 22977 16729 22989 16763
rect 23023 16729 23035 16763
rect 22977 16723 23035 16729
rect 23986 16720 23992 16772
rect 24044 16760 24050 16772
rect 24265 16763 24323 16769
rect 24265 16760 24277 16763
rect 24044 16732 24277 16760
rect 24044 16720 24050 16732
rect 24265 16729 24277 16732
rect 24311 16729 24323 16763
rect 24265 16723 24323 16729
rect 22146 16692 22152 16704
rect 22107 16664 22152 16692
rect 22146 16652 22152 16664
rect 22204 16652 22210 16704
rect 22330 16624 22336 16636
rect 21152 16596 22336 16624
rect 22330 16584 22336 16596
rect 22388 16584 22394 16636
rect 13958 16516 13964 16568
rect 14016 16556 14022 16568
rect 21042 16556 21048 16568
rect 14016 16528 21048 16556
rect 14016 16516 14022 16528
rect 21042 16516 21048 16528
rect 21100 16516 21106 16568
rect 21318 16556 21324 16568
rect 21279 16528 21324 16556
rect 21318 16516 21324 16528
rect 21376 16516 21382 16568
rect 23253 16559 23311 16565
rect 23253 16525 23265 16559
rect 23299 16556 23311 16559
rect 23526 16556 23532 16568
rect 23299 16528 23532 16556
rect 23299 16525 23311 16528
rect 23253 16519 23311 16525
rect 23526 16516 23532 16528
rect 23584 16516 23590 16568
rect 24449 16559 24507 16565
rect 24449 16525 24461 16559
rect 24495 16556 24507 16559
rect 24538 16556 24544 16568
rect 24495 16528 24544 16556
rect 24495 16525 24507 16528
rect 24449 16519 24507 16525
rect 24538 16516 24544 16528
rect 24596 16516 24602 16568
rect 11000 16466 34368 16488
rect 11000 16414 14142 16466
rect 14194 16414 14206 16466
rect 14258 16414 14270 16466
rect 14322 16414 14334 16466
rect 14386 16414 24142 16466
rect 24194 16414 24206 16466
rect 24258 16414 24270 16466
rect 24322 16414 24334 16466
rect 24386 16414 34368 16466
rect 11000 16392 34368 16414
rect 22146 16312 22152 16364
rect 22204 16352 22210 16364
rect 22204 16324 25320 16352
rect 22204 16312 22210 16324
rect 18190 16284 18196 16296
rect 17748 16256 18196 16284
rect 12486 16176 12492 16228
rect 12544 16216 12550 16228
rect 12857 16219 12915 16225
rect 12857 16216 12869 16219
rect 12544 16188 12869 16216
rect 12544 16176 12550 16188
rect 12857 16185 12869 16188
rect 12903 16185 12915 16219
rect 15338 16216 15344 16228
rect 15299 16188 15344 16216
rect 12857 16179 12915 16185
rect 15338 16176 15344 16188
rect 15396 16176 15402 16228
rect 17748 16225 17776 16256
rect 18190 16244 18196 16256
rect 18248 16244 18254 16296
rect 20766 16244 20772 16296
rect 20824 16284 20830 16296
rect 20824 16256 21548 16284
rect 20824 16244 20830 16256
rect 17733 16219 17791 16225
rect 17733 16185 17745 16219
rect 17779 16185 17791 16219
rect 18926 16216 18932 16228
rect 18887 16188 18932 16216
rect 17733 16179 17791 16185
rect 18926 16176 18932 16188
rect 18984 16176 18990 16228
rect 21318 16216 21324 16228
rect 21279 16188 21324 16216
rect 21318 16176 21324 16188
rect 21376 16176 21382 16228
rect 21520 16225 21548 16256
rect 21505 16219 21563 16225
rect 21505 16185 21517 16219
rect 21551 16185 21563 16219
rect 23250 16216 23256 16228
rect 23211 16188 23256 16216
rect 21505 16179 21563 16185
rect 23250 16176 23256 16188
rect 23308 16176 23314 16228
rect 23526 16216 23532 16228
rect 23487 16188 23532 16216
rect 23526 16176 23532 16188
rect 23584 16176 23590 16228
rect 25292 16225 25320 16324
rect 25277 16219 25335 16225
rect 25277 16185 25289 16219
rect 25323 16185 25335 16219
rect 25277 16179 25335 16185
rect 12394 16148 12400 16160
rect 12355 16120 12400 16148
rect 12394 16108 12400 16120
rect 12452 16108 12458 16160
rect 12670 16108 12676 16160
rect 12728 16148 12734 16160
rect 15614 16148 15620 16160
rect 12728 16120 12773 16148
rect 15575 16120 15620 16148
rect 12728 16108 12734 16120
rect 15614 16108 15620 16120
rect 15672 16108 15678 16160
rect 15801 16151 15859 16157
rect 15801 16117 15813 16151
rect 15847 16148 15859 16151
rect 17365 16151 17423 16157
rect 15847 16120 16672 16148
rect 15847 16117 15859 16120
rect 15801 16111 15859 16117
rect 11845 16083 11903 16089
rect 11845 16049 11857 16083
rect 11891 16049 11903 16083
rect 14786 16080 14792 16092
rect 14747 16052 14792 16080
rect 11845 16043 11903 16049
rect 11860 16012 11888 16043
rect 14786 16040 14792 16052
rect 14844 16040 14850 16092
rect 14510 16012 14516 16024
rect 11860 15984 14516 16012
rect 14510 15972 14516 15984
rect 14568 15972 14574 16024
rect 16644 16012 16672 16120
rect 17365 16117 17377 16151
rect 17411 16148 17423 16151
rect 17914 16148 17920 16160
rect 17411 16120 17920 16148
rect 17411 16117 17423 16120
rect 17365 16111 17423 16117
rect 17914 16108 17920 16120
rect 17972 16108 17978 16160
rect 18190 16148 18196 16160
rect 18151 16120 18196 16148
rect 18190 16108 18196 16120
rect 18248 16108 18254 16160
rect 19018 16148 19024 16160
rect 18979 16120 19024 16148
rect 19018 16108 19024 16120
rect 19076 16108 19082 16160
rect 19570 16108 19576 16160
rect 19628 16148 19634 16160
rect 19941 16151 19999 16157
rect 19941 16148 19953 16151
rect 19628 16120 19953 16148
rect 19628 16108 19634 16120
rect 19941 16117 19953 16120
rect 19987 16117 19999 16151
rect 21226 16148 21232 16160
rect 21187 16120 21232 16148
rect 19941 16111 19999 16117
rect 21226 16108 21232 16120
rect 21284 16108 21290 16160
rect 21597 16151 21655 16157
rect 21597 16117 21609 16151
rect 21643 16117 21655 16151
rect 21597 16111 21655 16117
rect 17181 16083 17239 16089
rect 17181 16049 17193 16083
rect 17227 16080 17239 16083
rect 17454 16080 17460 16092
rect 17227 16052 17460 16080
rect 17227 16049 17239 16052
rect 17181 16043 17239 16049
rect 17454 16040 17460 16052
rect 17512 16040 17518 16092
rect 18208 16080 18236 16108
rect 19846 16080 19852 16092
rect 18208 16052 19852 16080
rect 19846 16040 19852 16052
rect 19904 16040 19910 16092
rect 18466 16012 18472 16024
rect 16644 15984 18472 16012
rect 18466 15972 18472 15984
rect 18524 15972 18530 16024
rect 18834 15972 18840 16024
rect 18892 16012 18898 16024
rect 19113 16015 19171 16021
rect 19113 16012 19125 16015
rect 18892 15984 19125 16012
rect 18892 15972 18898 15984
rect 19113 15981 19125 15984
rect 19159 15981 19171 16015
rect 20122 16012 20128 16024
rect 20083 15984 20128 16012
rect 19113 15975 19171 15981
rect 20122 15972 20128 15984
rect 20180 15972 20186 16024
rect 20674 16012 20680 16024
rect 20635 15984 20680 16012
rect 20674 15972 20680 15984
rect 20732 15972 20738 16024
rect 21244 16012 21272 16108
rect 21612 16080 21640 16111
rect 22330 16080 22336 16092
rect 21612 16052 22336 16080
rect 22330 16040 22336 16052
rect 22388 16040 22394 16092
rect 24538 16040 24544 16092
rect 24596 16040 24602 16092
rect 22238 16012 22244 16024
rect 21244 15984 22244 16012
rect 22238 15972 22244 15984
rect 22296 15972 22302 16024
rect 11000 15922 34368 15944
rect 11000 15870 19142 15922
rect 19194 15870 19206 15922
rect 19258 15870 19270 15922
rect 19322 15870 19334 15922
rect 19386 15870 29142 15922
rect 29194 15870 29206 15922
rect 29258 15870 29270 15922
rect 29322 15870 29334 15922
rect 29386 15870 34368 15922
rect 11000 15848 34368 15870
rect 18742 15768 18748 15820
rect 18800 15808 18806 15820
rect 22422 15808 22428 15820
rect 18800 15780 22428 15808
rect 18800 15768 18806 15780
rect 22422 15768 22428 15780
rect 22480 15768 22486 15820
rect 17564 15712 18512 15740
rect 12213 15675 12271 15681
rect 12213 15641 12225 15675
rect 12259 15672 12271 15675
rect 12486 15672 12492 15684
rect 12259 15644 12492 15672
rect 12259 15641 12271 15644
rect 12213 15635 12271 15641
rect 12486 15632 12492 15644
rect 12544 15632 12550 15684
rect 12762 15672 12768 15684
rect 12723 15644 12768 15672
rect 12762 15632 12768 15644
rect 12820 15632 12826 15684
rect 12946 15672 12952 15684
rect 12907 15644 12952 15672
rect 12946 15632 12952 15644
rect 13004 15632 13010 15684
rect 13774 15632 13780 15684
rect 13832 15672 13838 15684
rect 14329 15675 14387 15681
rect 14329 15672 14341 15675
rect 13832 15644 14341 15672
rect 13832 15632 13838 15644
rect 14329 15641 14341 15644
rect 14375 15641 14387 15675
rect 14329 15635 14387 15641
rect 12762 15536 12768 15548
rect 12723 15508 12768 15536
rect 12762 15496 12768 15508
rect 12820 15496 12826 15548
rect 14344 15468 14372 15635
rect 15706 15632 15712 15684
rect 15764 15632 15770 15684
rect 16813 15675 16871 15681
rect 16813 15641 16825 15675
rect 16859 15641 16871 15675
rect 16813 15635 16871 15641
rect 17181 15675 17239 15681
rect 17181 15641 17193 15675
rect 17227 15672 17239 15675
rect 17362 15672 17368 15684
rect 17227 15644 17368 15672
rect 17227 15641 17239 15644
rect 17181 15635 17239 15641
rect 14605 15607 14663 15613
rect 14605 15573 14617 15607
rect 14651 15604 14663 15607
rect 15982 15604 15988 15616
rect 14651 15576 15988 15604
rect 14651 15573 14663 15576
rect 14605 15567 14663 15573
rect 15982 15564 15988 15576
rect 16040 15564 16046 15616
rect 16353 15607 16411 15613
rect 16353 15573 16365 15607
rect 16399 15604 16411 15607
rect 16828 15604 16856 15635
rect 17362 15632 17368 15644
rect 17420 15632 17426 15684
rect 17564 15681 17592 15712
rect 18484 15684 18512 15712
rect 18926 15700 18932 15752
rect 18984 15740 18990 15752
rect 19021 15743 19079 15749
rect 19021 15740 19033 15743
rect 18984 15712 19033 15740
rect 18984 15700 18990 15712
rect 19021 15709 19033 15712
rect 19067 15709 19079 15743
rect 19021 15703 19079 15709
rect 20122 15700 20128 15752
rect 20180 15740 20186 15752
rect 20180 15712 20338 15740
rect 20180 15700 20186 15712
rect 22238 15700 22244 15752
rect 22296 15700 22302 15752
rect 17549 15675 17607 15681
rect 17549 15641 17561 15675
rect 17595 15641 17607 15675
rect 18466 15672 18472 15684
rect 18427 15644 18472 15672
rect 17549 15635 17607 15641
rect 18466 15632 18472 15644
rect 18524 15632 18530 15684
rect 18558 15632 18564 15684
rect 18616 15672 18622 15684
rect 18616 15644 18661 15672
rect 18616 15632 18622 15644
rect 21410 15632 21416 15684
rect 21468 15672 21474 15684
rect 22149 15675 22207 15681
rect 22149 15672 22161 15675
rect 21468 15644 22161 15672
rect 21468 15632 21474 15644
rect 22149 15641 22161 15644
rect 22195 15641 22207 15675
rect 22256 15672 22284 15700
rect 22517 15675 22575 15681
rect 22517 15672 22529 15675
rect 22256 15644 22529 15672
rect 22149 15635 22207 15641
rect 22517 15641 22529 15644
rect 22563 15641 22575 15675
rect 22517 15635 22575 15641
rect 16399 15576 16856 15604
rect 18285 15607 18343 15613
rect 16399 15573 16411 15576
rect 16353 15567 16411 15573
rect 18285 15573 18297 15607
rect 18331 15604 18343 15607
rect 18374 15604 18380 15616
rect 18331 15576 18380 15604
rect 18331 15573 18343 15576
rect 18285 15567 18343 15573
rect 15614 15496 15620 15548
rect 15672 15536 15678 15548
rect 16368 15536 16396 15567
rect 18374 15564 18380 15576
rect 18432 15564 18438 15616
rect 19570 15564 19576 15616
rect 19628 15604 19634 15616
rect 21594 15604 21600 15616
rect 19628 15576 19673 15604
rect 21555 15576 21600 15604
rect 19628 15564 19634 15576
rect 21594 15564 21600 15576
rect 21652 15564 21658 15616
rect 15672 15508 16396 15536
rect 15672 15496 15678 15508
rect 16718 15468 16724 15480
rect 14344 15440 16724 15468
rect 16718 15428 16724 15440
rect 16776 15428 16782 15480
rect 19662 15428 19668 15480
rect 19720 15468 19726 15480
rect 19830 15471 19888 15477
rect 19830 15468 19842 15471
rect 19720 15440 19842 15468
rect 19720 15428 19726 15440
rect 19830 15437 19842 15440
rect 19876 15437 19888 15471
rect 23986 15468 23992 15480
rect 23947 15440 23992 15468
rect 19830 15431 19888 15437
rect 23986 15428 23992 15440
rect 24044 15428 24050 15480
rect 11000 15378 34368 15400
rect 11000 15326 14142 15378
rect 14194 15326 14206 15378
rect 14258 15326 14270 15378
rect 14322 15326 14334 15378
rect 14386 15326 24142 15378
rect 24194 15326 24206 15378
rect 24258 15326 24270 15378
rect 24322 15326 24334 15378
rect 24386 15326 34368 15378
rect 11000 15304 34368 15326
rect 15982 15264 15988 15276
rect 13884 15236 15752 15264
rect 15943 15236 15988 15264
rect 13884 15205 13912 15236
rect 13869 15199 13927 15205
rect 13869 15165 13881 15199
rect 13915 15165 13927 15199
rect 15614 15196 15620 15208
rect 13869 15159 13927 15165
rect 14896 15168 15620 15196
rect 12029 15131 12087 15137
rect 12029 15097 12041 15131
rect 12075 15128 12087 15131
rect 12394 15128 12400 15140
rect 12075 15100 12400 15128
rect 12075 15097 12087 15100
rect 12029 15091 12087 15097
rect 12394 15088 12400 15100
rect 12452 15088 12458 15140
rect 14896 15137 14924 15168
rect 15614 15156 15620 15168
rect 15672 15156 15678 15208
rect 15724 15196 15752 15236
rect 15982 15224 15988 15236
rect 16040 15224 16046 15276
rect 20677 15267 20735 15273
rect 20677 15233 20689 15267
rect 20723 15264 20735 15267
rect 20766 15264 20772 15276
rect 20723 15236 20772 15264
rect 20723 15233 20735 15236
rect 20677 15227 20735 15233
rect 20766 15224 20772 15236
rect 20824 15224 20830 15276
rect 18282 15196 18288 15208
rect 15724 15168 18288 15196
rect 18282 15156 18288 15168
rect 18340 15156 18346 15208
rect 18558 15156 18564 15208
rect 18616 15196 18622 15208
rect 21594 15196 21600 15208
rect 18616 15168 21600 15196
rect 18616 15156 18622 15168
rect 14881 15131 14939 15137
rect 14881 15097 14893 15131
rect 14927 15097 14939 15131
rect 18466 15128 18472 15140
rect 14881 15091 14939 15097
rect 17380 15100 18472 15128
rect 11937 15063 11995 15069
rect 11937 15029 11949 15063
rect 11983 15060 11995 15063
rect 12765 15063 12823 15069
rect 12765 15060 12777 15063
rect 11983 15032 12777 15060
rect 11983 15029 11995 15032
rect 11937 15023 11995 15029
rect 12765 15029 12777 15032
rect 12811 15060 12823 15063
rect 13038 15060 13044 15072
rect 12811 15032 12900 15060
rect 12999 15032 13044 15060
rect 12811 15029 12823 15032
rect 12765 15023 12823 15029
rect 12872 14924 12900 15032
rect 13038 15020 13044 15032
rect 13096 15020 13102 15072
rect 13406 15060 13412 15072
rect 13367 15032 13412 15060
rect 13406 15020 13412 15032
rect 13464 15020 13470 15072
rect 13498 15020 13504 15072
rect 13556 15060 13562 15072
rect 13685 15063 13743 15069
rect 13685 15060 13697 15063
rect 13556 15032 13697 15060
rect 13556 15020 13562 15032
rect 13685 15029 13697 15032
rect 13731 15029 13743 15063
rect 13685 15023 13743 15029
rect 14973 15063 15031 15069
rect 14973 15029 14985 15063
rect 15019 15060 15031 15063
rect 15062 15060 15068 15072
rect 15019 15032 15068 15060
rect 15019 15029 15031 15032
rect 14973 15023 15031 15029
rect 15062 15020 15068 15032
rect 15120 15060 15126 15072
rect 17380 15069 17408 15100
rect 18466 15088 18472 15100
rect 18524 15088 18530 15140
rect 19389 15131 19447 15137
rect 19389 15097 19401 15131
rect 19435 15128 19447 15131
rect 19662 15128 19668 15140
rect 19435 15100 19668 15128
rect 19435 15097 19447 15100
rect 19389 15091 19447 15097
rect 19662 15088 19668 15100
rect 19720 15088 19726 15140
rect 15525 15063 15583 15069
rect 15525 15060 15537 15063
rect 15120 15032 15537 15060
rect 15120 15020 15126 15032
rect 15525 15029 15537 15032
rect 15571 15029 15583 15063
rect 15525 15023 15583 15029
rect 15709 15063 15767 15069
rect 15709 15029 15721 15063
rect 15755 15029 15767 15063
rect 15709 15023 15767 15029
rect 17365 15063 17423 15069
rect 17365 15029 17377 15063
rect 17411 15029 17423 15063
rect 17365 15023 17423 15029
rect 17917 15063 17975 15069
rect 17917 15029 17929 15063
rect 17963 15029 17975 15063
rect 18834 15060 18840 15072
rect 18795 15032 18840 15060
rect 17917 15023 17975 15029
rect 15724 14992 15752 15023
rect 17454 14992 17460 15004
rect 15724 14964 17460 14992
rect 17454 14952 17460 14964
rect 17512 14952 17518 15004
rect 15890 14924 15896 14936
rect 12872 14896 15896 14924
rect 15890 14884 15896 14896
rect 15948 14884 15954 14936
rect 16902 14884 16908 14936
rect 16960 14924 16966 14936
rect 17932 14924 17960 15023
rect 18834 15020 18840 15032
rect 18892 15020 18898 15072
rect 19021 15063 19079 15069
rect 19021 15029 19033 15063
rect 19067 15060 19079 15063
rect 19478 15060 19484 15072
rect 19067 15032 19484 15060
rect 19067 15029 19079 15032
rect 19021 15023 19079 15029
rect 19478 15020 19484 15032
rect 19536 15020 19542 15072
rect 20232 15060 20260 15168
rect 21594 15156 21600 15168
rect 21652 15156 21658 15208
rect 22330 15088 22336 15140
rect 22388 15128 22394 15140
rect 22388 15100 22433 15128
rect 22388 15088 22394 15100
rect 20309 15063 20367 15069
rect 20309 15060 20321 15063
rect 20232 15032 20321 15060
rect 20309 15029 20321 15032
rect 20355 15029 20367 15063
rect 20309 15023 20367 15029
rect 22146 15020 22152 15072
rect 22204 15060 22210 15072
rect 22425 15063 22483 15069
rect 22425 15060 22437 15063
rect 22204 15032 22437 15060
rect 22204 15020 22210 15032
rect 22425 15029 22437 15032
rect 22471 15029 22483 15063
rect 22425 15023 22483 15029
rect 24081 15063 24139 15069
rect 24081 15029 24093 15063
rect 24127 15029 24139 15063
rect 24081 15023 24139 15029
rect 24357 15063 24415 15069
rect 24357 15029 24369 15063
rect 24403 15060 24415 15063
rect 24538 15060 24544 15072
rect 24403 15032 24544 15060
rect 24403 15029 24415 15032
rect 24357 15023 24415 15029
rect 24096 14992 24124 15023
rect 24538 15020 24544 15032
rect 24596 15020 24602 15072
rect 24446 14992 24452 15004
rect 24096 14964 24452 14992
rect 24446 14952 24452 14964
rect 24504 14952 24510 15004
rect 18098 14924 18104 14936
rect 16960 14896 17960 14924
rect 18059 14896 18104 14924
rect 16960 14884 16966 14896
rect 18098 14884 18104 14896
rect 18156 14884 18162 14936
rect 23894 14924 23900 14936
rect 23855 14896 23900 14924
rect 23894 14884 23900 14896
rect 23952 14884 23958 14936
rect 11000 14834 34368 14856
rect 11000 14782 19142 14834
rect 19194 14782 19206 14834
rect 19258 14782 19270 14834
rect 19322 14782 19334 14834
rect 19386 14782 29142 14834
rect 29194 14782 29206 14834
rect 29258 14782 29270 14834
rect 29322 14782 29334 14834
rect 29386 14782 34368 14834
rect 11000 14760 34368 14782
rect 12854 14720 12860 14732
rect 12504 14692 12860 14720
rect 12504 14593 12532 14692
rect 12854 14680 12860 14692
rect 12912 14720 12918 14732
rect 14786 14720 14792 14732
rect 12912 14692 14792 14720
rect 12912 14680 12918 14692
rect 14786 14680 14792 14692
rect 14844 14680 14850 14732
rect 15706 14720 15712 14732
rect 15667 14692 15712 14720
rect 15706 14680 15712 14692
rect 15764 14680 15770 14732
rect 15890 14680 15896 14732
rect 15948 14720 15954 14732
rect 21410 14720 21416 14732
rect 15948 14692 18328 14720
rect 21371 14692 21416 14720
rect 15948 14680 15954 14692
rect 13038 14652 13044 14664
rect 12999 14624 13044 14652
rect 13038 14612 13044 14624
rect 13096 14612 13102 14664
rect 16902 14652 16908 14664
rect 15540 14624 16908 14652
rect 12489 14587 12547 14593
rect 12489 14553 12501 14587
rect 12535 14553 12547 14587
rect 12762 14584 12768 14596
rect 12723 14556 12768 14584
rect 12489 14547 12547 14553
rect 12762 14544 12768 14556
rect 12820 14544 12826 14596
rect 13406 14544 13412 14596
rect 13464 14584 13470 14596
rect 13961 14587 14019 14593
rect 13961 14584 13973 14587
rect 13464 14556 13973 14584
rect 13464 14544 13470 14556
rect 13961 14553 13973 14556
rect 14007 14553 14019 14587
rect 13961 14547 14019 14553
rect 14510 14544 14516 14596
rect 14568 14584 14574 14596
rect 15540 14593 15568 14624
rect 16902 14612 16908 14624
rect 16960 14612 16966 14664
rect 18300 14652 18328 14692
rect 21410 14680 21416 14692
rect 21468 14680 21474 14732
rect 23161 14655 23219 14661
rect 23161 14652 23173 14655
rect 18300 14624 23173 14652
rect 23161 14621 23173 14624
rect 23207 14621 23219 14655
rect 23161 14615 23219 14621
rect 23986 14612 23992 14664
rect 24044 14652 24050 14664
rect 25185 14655 25243 14661
rect 25185 14652 25197 14655
rect 24044 14624 25197 14652
rect 24044 14612 24050 14624
rect 14789 14587 14847 14593
rect 14789 14584 14801 14587
rect 14568 14556 14801 14584
rect 14568 14544 14574 14556
rect 14789 14553 14801 14556
rect 14835 14553 14847 14587
rect 14789 14547 14847 14553
rect 15525 14587 15583 14593
rect 15525 14553 15537 14587
rect 15571 14553 15583 14587
rect 16718 14584 16724 14596
rect 16679 14556 16724 14584
rect 15525 14547 15583 14553
rect 16718 14544 16724 14556
rect 16776 14544 16782 14596
rect 18098 14544 18104 14596
rect 18156 14544 18162 14596
rect 18466 14544 18472 14596
rect 18524 14584 18530 14596
rect 18745 14587 18803 14593
rect 18745 14584 18757 14587
rect 18524 14556 18757 14584
rect 18524 14544 18530 14556
rect 18745 14553 18757 14556
rect 18791 14553 18803 14587
rect 21318 14584 21324 14596
rect 21279 14556 21324 14584
rect 18745 14547 18803 14553
rect 21318 14544 21324 14556
rect 21376 14544 21382 14596
rect 21594 14544 21600 14596
rect 21652 14584 21658 14596
rect 21873 14587 21931 14593
rect 21873 14584 21885 14587
rect 21652 14556 21885 14584
rect 21652 14544 21658 14556
rect 21873 14553 21885 14556
rect 21919 14553 21931 14587
rect 22146 14584 22152 14596
rect 22107 14556 22152 14584
rect 21873 14547 21931 14553
rect 22146 14544 22152 14556
rect 22204 14544 22210 14596
rect 23802 14584 23808 14596
rect 23763 14556 23808 14584
rect 23802 14544 23808 14556
rect 23860 14544 23866 14596
rect 23894 14544 23900 14596
rect 23952 14584 23958 14596
rect 24280 14593 24308 14624
rect 25185 14621 25197 14624
rect 25231 14621 25243 14655
rect 25185 14615 25243 14621
rect 24173 14587 24231 14593
rect 23952 14556 23997 14584
rect 23952 14544 23958 14556
rect 24173 14553 24185 14587
rect 24219 14553 24231 14587
rect 24173 14547 24231 14553
rect 24265 14587 24323 14593
rect 24265 14553 24277 14587
rect 24311 14553 24323 14587
rect 25366 14584 25372 14596
rect 25327 14556 25372 14584
rect 24265 14547 24323 14553
rect 12026 14516 12032 14528
rect 11987 14488 12032 14516
rect 12026 14476 12032 14488
rect 12084 14476 12090 14528
rect 14881 14519 14939 14525
rect 14881 14485 14893 14519
rect 14927 14516 14939 14519
rect 16994 14516 17000 14528
rect 14927 14488 16672 14516
rect 16955 14488 17000 14516
rect 14927 14485 14939 14488
rect 14881 14479 14939 14485
rect 14786 14448 14792 14460
rect 14747 14420 14792 14448
rect 14786 14408 14792 14420
rect 14844 14408 14850 14460
rect 16644 14380 16672 14488
rect 16994 14476 17000 14488
rect 17052 14476 17058 14528
rect 24188 14516 24216 14547
rect 25366 14544 25372 14556
rect 25424 14544 25430 14596
rect 25384 14516 25412 14544
rect 24188 14488 25412 14516
rect 23250 14380 23256 14392
rect 16644 14352 23256 14380
rect 23250 14340 23256 14352
rect 23308 14340 23314 14392
rect 23894 14340 23900 14392
rect 23952 14380 23958 14392
rect 25461 14383 25519 14389
rect 25461 14380 25473 14383
rect 23952 14352 25473 14380
rect 23952 14340 23958 14352
rect 25461 14349 25473 14352
rect 25507 14349 25519 14383
rect 25461 14343 25519 14349
rect 11000 14290 34368 14312
rect 11000 14238 14142 14290
rect 14194 14238 14206 14290
rect 14258 14238 14270 14290
rect 14322 14238 14334 14290
rect 14386 14238 24142 14290
rect 24194 14238 24206 14290
rect 24258 14238 24270 14290
rect 24322 14238 24334 14290
rect 24386 14238 34368 14290
rect 11000 14216 34368 14238
rect 12026 14176 12032 14188
rect 11987 14148 12032 14176
rect 12026 14136 12032 14148
rect 12084 14136 12090 14188
rect 12946 14136 12952 14188
rect 13004 14176 13010 14188
rect 13041 14179 13099 14185
rect 13041 14176 13053 14179
rect 13004 14148 13053 14176
rect 13004 14136 13010 14148
rect 13041 14145 13053 14148
rect 13087 14145 13099 14179
rect 13041 14139 13099 14145
rect 16994 14136 17000 14188
rect 17052 14176 17058 14188
rect 17181 14179 17239 14185
rect 17181 14176 17193 14179
rect 17052 14148 17193 14176
rect 17052 14136 17058 14148
rect 17181 14145 17193 14148
rect 17227 14145 17239 14179
rect 17181 14139 17239 14145
rect 12044 14040 12072 14136
rect 14694 14068 14700 14120
rect 14752 14108 14758 14120
rect 14752 14080 20076 14108
rect 14752 14068 14758 14080
rect 12765 14043 12823 14049
rect 12765 14040 12777 14043
rect 12044 14012 12777 14040
rect 12765 14009 12777 14012
rect 12811 14009 12823 14043
rect 12765 14003 12823 14009
rect 14513 14043 14571 14049
rect 14513 14009 14525 14043
rect 14559 14040 14571 14043
rect 16166 14040 16172 14052
rect 14559 14012 16172 14040
rect 14559 14009 14571 14012
rect 14513 14003 14571 14009
rect 16166 14000 16172 14012
rect 16224 14000 16230 14052
rect 17454 14000 17460 14052
rect 17512 14040 17518 14052
rect 17641 14043 17699 14049
rect 17641 14040 17653 14043
rect 17512 14012 17653 14040
rect 17512 14000 17518 14012
rect 17641 14009 17653 14012
rect 17687 14009 17699 14043
rect 18190 14040 18196 14052
rect 17641 14003 17699 14009
rect 17748 14012 18196 14040
rect 10462 13932 10468 13984
rect 10520 13972 10526 13984
rect 11661 13975 11719 13981
rect 11661 13972 11673 13975
rect 10520 13944 11673 13972
rect 10520 13932 10526 13944
rect 11661 13941 11673 13944
rect 11707 13941 11719 13975
rect 12854 13972 12860 13984
rect 12815 13944 12860 13972
rect 11661 13935 11719 13941
rect 12854 13932 12860 13944
rect 12912 13932 12918 13984
rect 14145 13975 14203 13981
rect 14145 13941 14157 13975
rect 14191 13972 14203 13975
rect 14786 13972 14792 13984
rect 14191 13944 14792 13972
rect 14191 13941 14203 13944
rect 14145 13935 14203 13941
rect 14786 13932 14792 13944
rect 14844 13932 14850 13984
rect 17748 13981 17776 14012
rect 18190 14000 18196 14012
rect 18248 14040 18254 14052
rect 19478 14040 19484 14052
rect 18248 14012 19340 14040
rect 19439 14012 19484 14040
rect 18248 14000 18254 14012
rect 17733 13975 17791 13981
rect 17733 13941 17745 13975
rect 17779 13941 17791 13975
rect 17733 13935 17791 13941
rect 17822 13932 17828 13984
rect 17880 13972 17886 13984
rect 18101 13975 18159 13981
rect 18101 13972 18113 13975
rect 17880 13944 18113 13972
rect 17880 13932 17886 13944
rect 18101 13941 18113 13944
rect 18147 13941 18159 13975
rect 18282 13972 18288 13984
rect 18243 13944 18288 13972
rect 18101 13935 18159 13941
rect 13498 13864 13504 13916
rect 13556 13904 13562 13916
rect 13961 13907 14019 13913
rect 13961 13904 13973 13907
rect 13556 13876 13973 13904
rect 13556 13864 13562 13876
rect 13961 13873 13973 13876
rect 14007 13873 14019 13907
rect 13961 13867 14019 13873
rect 18116 13836 18144 13935
rect 18282 13932 18288 13944
rect 18340 13932 18346 13984
rect 18926 13972 18932 13984
rect 18887 13944 18932 13972
rect 18926 13932 18932 13944
rect 18984 13932 18990 13984
rect 19312 13972 19340 14012
rect 19478 14000 19484 14012
rect 19536 14000 19542 14052
rect 20048 14049 20076 14080
rect 20508 14080 22836 14108
rect 20033 14043 20091 14049
rect 20033 14009 20045 14043
rect 20079 14009 20091 14043
rect 20033 14003 20091 14009
rect 20508 13972 20536 14080
rect 20769 14043 20827 14049
rect 20769 14009 20781 14043
rect 20815 14040 20827 14043
rect 21226 14040 21232 14052
rect 20815 14012 21232 14040
rect 20815 14009 20827 14012
rect 20769 14003 20827 14009
rect 21226 14000 21232 14012
rect 21284 14000 21290 14052
rect 20674 13972 20680 13984
rect 19312 13944 20536 13972
rect 20635 13944 20680 13972
rect 20674 13932 20680 13944
rect 20732 13932 20738 13984
rect 21045 13975 21103 13981
rect 21045 13941 21057 13975
rect 21091 13941 21103 13975
rect 21045 13935 21103 13941
rect 18650 13864 18656 13916
rect 18708 13904 18714 13916
rect 18745 13907 18803 13913
rect 18745 13904 18757 13907
rect 18708 13876 18757 13904
rect 18708 13864 18714 13876
rect 18745 13873 18757 13876
rect 18791 13873 18803 13907
rect 18745 13867 18803 13873
rect 18834 13864 18840 13916
rect 18892 13904 18898 13916
rect 19113 13907 19171 13913
rect 19113 13904 19125 13907
rect 18892 13876 19125 13904
rect 18892 13864 18898 13876
rect 19113 13873 19125 13876
rect 19159 13873 19171 13907
rect 21060 13904 21088 13935
rect 21134 13932 21140 13984
rect 21192 13972 21198 13984
rect 21192 13944 21237 13972
rect 21192 13932 21198 13944
rect 21318 13904 21324 13916
rect 21060 13876 21324 13904
rect 19113 13867 19171 13873
rect 21318 13864 21324 13876
rect 21376 13864 21382 13916
rect 22808 13904 22836 14080
rect 23713 14043 23771 14049
rect 23713 14009 23725 14043
rect 23759 14040 23771 14043
rect 23802 14040 23808 14052
rect 23759 14012 23808 14040
rect 23759 14009 23771 14012
rect 23713 14003 23771 14009
rect 23802 14000 23808 14012
rect 23860 14000 23866 14052
rect 23621 13975 23679 13981
rect 23621 13941 23633 13975
rect 23667 13972 23679 13975
rect 23894 13972 23900 13984
rect 23667 13944 23900 13972
rect 23667 13941 23679 13944
rect 23621 13935 23679 13941
rect 23894 13932 23900 13944
rect 23952 13932 23958 13984
rect 24446 13972 24452 13984
rect 24407 13944 24452 13972
rect 24446 13932 24452 13944
rect 24504 13932 24510 13984
rect 24538 13932 24544 13984
rect 24596 13972 24602 13984
rect 25550 13972 25556 13984
rect 24596 13944 24641 13972
rect 25511 13944 25556 13972
rect 24596 13932 24602 13944
rect 25550 13932 25556 13944
rect 25608 13932 25614 13984
rect 26013 13975 26071 13981
rect 26013 13941 26025 13975
rect 26059 13972 26071 13975
rect 27206 13972 27212 13984
rect 26059 13944 27212 13972
rect 26059 13941 26071 13944
rect 26013 13935 26071 13941
rect 27206 13932 27212 13944
rect 27264 13932 27270 13984
rect 22808 13876 26134 13904
rect 19021 13839 19079 13845
rect 19021 13836 19033 13839
rect 18116 13808 19033 13836
rect 19021 13805 19033 13808
rect 19067 13805 19079 13839
rect 19021 13799 19079 13805
rect 11000 13746 34368 13768
rect 11000 13694 19142 13746
rect 19194 13694 19206 13746
rect 19258 13694 19270 13746
rect 19322 13694 19334 13746
rect 19386 13694 29142 13746
rect 29194 13694 29206 13746
rect 29258 13694 29270 13746
rect 29322 13694 29334 13746
rect 29386 13694 34368 13746
rect 11000 13672 34368 13694
rect 12854 13592 12860 13644
rect 12912 13632 12918 13644
rect 14142 13632 14148 13644
rect 12912 13604 14148 13632
rect 12912 13592 12918 13604
rect 14142 13592 14148 13604
rect 14200 13632 14206 13644
rect 14694 13632 14700 13644
rect 14200 13604 14700 13632
rect 14200 13592 14206 13604
rect 14694 13592 14700 13604
rect 14752 13592 14758 13644
rect 21318 13632 21324 13644
rect 19772 13604 21324 13632
rect 13406 13564 13412 13576
rect 13367 13536 13412 13564
rect 13406 13524 13412 13536
rect 13464 13524 13470 13576
rect 15249 13567 15307 13573
rect 15249 13564 15261 13567
rect 13700 13536 15261 13564
rect 12949 13499 13007 13505
rect 12949 13465 12961 13499
rect 12995 13496 13007 13499
rect 13130 13496 13136 13508
rect 12995 13468 13136 13496
rect 12995 13465 13007 13468
rect 12949 13459 13007 13465
rect 13130 13456 13136 13468
rect 13188 13496 13194 13508
rect 13700 13496 13728 13536
rect 15249 13533 15261 13536
rect 15295 13533 15307 13567
rect 18282 13564 18288 13576
rect 15249 13527 15307 13533
rect 17840 13536 18288 13564
rect 14142 13505 14148 13508
rect 13188 13468 13728 13496
rect 14130 13499 14148 13505
rect 13188 13456 13194 13468
rect 14130 13465 14142 13499
rect 14130 13459 14148 13465
rect 14142 13456 14148 13459
rect 14200 13456 14206 13508
rect 14602 13496 14608 13508
rect 14563 13468 14608 13496
rect 14602 13456 14608 13468
rect 14660 13456 14666 13508
rect 14694 13456 14700 13508
rect 14752 13496 14758 13508
rect 14752 13468 14797 13496
rect 14752 13456 14758 13468
rect 15062 13456 15068 13508
rect 15120 13496 15126 13508
rect 17546 13496 17552 13508
rect 15120 13468 17552 13496
rect 15120 13456 15126 13468
rect 17546 13456 17552 13468
rect 17604 13456 17610 13508
rect 17840 13505 17868 13536
rect 18282 13524 18288 13536
rect 18340 13564 18346 13576
rect 18340 13536 19064 13564
rect 18340 13524 18346 13536
rect 17825 13499 17883 13505
rect 17825 13465 17837 13499
rect 17871 13465 17883 13499
rect 18558 13496 18564 13508
rect 18471 13468 18564 13496
rect 17825 13459 17883 13465
rect 18558 13456 18564 13468
rect 18616 13496 18622 13508
rect 18926 13496 18932 13508
rect 18616 13468 18932 13496
rect 18616 13456 18622 13468
rect 18926 13456 18932 13468
rect 18984 13456 18990 13508
rect 19036 13440 19064 13536
rect 19772 13505 19800 13604
rect 21318 13592 21324 13604
rect 21376 13592 21382 13644
rect 23250 13564 23256 13576
rect 20968 13536 21640 13564
rect 23211 13536 23256 13564
rect 19757 13499 19815 13505
rect 19757 13465 19769 13499
rect 19803 13465 19815 13499
rect 19757 13459 19815 13465
rect 20674 13456 20680 13508
rect 20732 13496 20738 13508
rect 20968 13505 20996 13536
rect 21612 13508 21640 13536
rect 23250 13524 23256 13536
rect 23308 13524 23314 13576
rect 25182 13524 25188 13576
rect 25240 13564 25246 13576
rect 27206 13564 27212 13576
rect 25240 13536 25950 13564
rect 27167 13536 27212 13564
rect 25240 13524 25246 13536
rect 27206 13524 27212 13536
rect 27264 13524 27270 13576
rect 20861 13499 20919 13505
rect 20861 13496 20873 13499
rect 20732 13468 20873 13496
rect 20732 13456 20738 13468
rect 20861 13465 20873 13468
rect 20907 13465 20919 13499
rect 20861 13459 20919 13465
rect 20953 13499 21011 13505
rect 20953 13465 20965 13499
rect 20999 13465 21011 13499
rect 21413 13499 21471 13505
rect 21413 13496 21425 13499
rect 20953 13459 21011 13465
rect 21060 13468 21425 13496
rect 12670 13388 12676 13440
rect 12728 13428 12734 13440
rect 12857 13431 12915 13437
rect 12857 13428 12869 13431
rect 12728 13400 12869 13428
rect 12728 13388 12734 13400
rect 12857 13397 12869 13400
rect 12903 13397 12915 13431
rect 12857 13391 12915 13397
rect 13038 13388 13044 13440
rect 13096 13428 13102 13440
rect 13961 13431 14019 13437
rect 13961 13428 13973 13431
rect 13096 13400 13973 13428
rect 13096 13388 13102 13400
rect 13961 13397 13973 13400
rect 14007 13397 14019 13431
rect 13961 13391 14019 13397
rect 13976 13292 14004 13391
rect 16902 13388 16908 13440
rect 16960 13428 16966 13440
rect 16997 13431 17055 13437
rect 16997 13428 17009 13431
rect 16960 13400 17009 13428
rect 16960 13388 16966 13400
rect 16997 13397 17009 13400
rect 17043 13397 17055 13431
rect 18009 13431 18067 13437
rect 18009 13428 18021 13431
rect 16997 13391 17055 13397
rect 17840 13400 18021 13428
rect 17840 13372 17868 13400
rect 18009 13397 18021 13400
rect 18055 13397 18067 13431
rect 18009 13391 18067 13397
rect 18469 13431 18527 13437
rect 18469 13397 18481 13431
rect 18515 13428 18527 13431
rect 18650 13428 18656 13440
rect 18515 13400 18656 13428
rect 18515 13397 18527 13400
rect 18469 13391 18527 13397
rect 18650 13388 18656 13400
rect 18708 13388 18714 13440
rect 19018 13428 19024 13440
rect 18979 13400 19024 13428
rect 19018 13388 19024 13400
rect 19076 13388 19082 13440
rect 19665 13431 19723 13437
rect 19665 13397 19677 13431
rect 19711 13397 19723 13431
rect 19665 13391 19723 13397
rect 20217 13431 20275 13437
rect 20217 13397 20229 13431
rect 20263 13397 20275 13431
rect 20876 13428 20904 13459
rect 21060 13428 21088 13468
rect 21413 13465 21425 13468
rect 21459 13465 21471 13499
rect 21594 13496 21600 13508
rect 21555 13468 21600 13496
rect 21413 13459 21471 13465
rect 21594 13456 21600 13468
rect 21652 13456 21658 13508
rect 23802 13496 23808 13508
rect 23763 13468 23808 13496
rect 23802 13456 23808 13468
rect 23860 13456 23866 13508
rect 24081 13499 24139 13505
rect 24081 13465 24093 13499
rect 24127 13496 24139 13499
rect 24538 13496 24544 13508
rect 24127 13468 24544 13496
rect 24127 13465 24139 13468
rect 24081 13459 24139 13465
rect 20876 13400 21088 13428
rect 21965 13431 22023 13437
rect 20217 13391 20275 13397
rect 21965 13397 21977 13431
rect 22011 13428 22023 13431
rect 24096 13428 24124 13459
rect 24538 13456 24544 13468
rect 24596 13456 24602 13508
rect 24814 13456 24820 13508
rect 24872 13496 24878 13508
rect 24872 13468 25228 13496
rect 24872 13456 24878 13468
rect 22011 13400 24124 13428
rect 24265 13431 24323 13437
rect 22011 13397 22023 13400
rect 21965 13391 22023 13397
rect 24265 13397 24277 13431
rect 24311 13428 24323 13431
rect 24446 13428 24452 13440
rect 24311 13400 24452 13428
rect 24311 13397 24323 13400
rect 24265 13391 24323 13397
rect 17822 13320 17828 13372
rect 17880 13320 17886 13372
rect 14602 13292 14608 13304
rect 13976 13264 14608 13292
rect 14602 13252 14608 13264
rect 14660 13252 14666 13304
rect 19680 13292 19708 13391
rect 20232 13360 20260 13391
rect 24446 13388 24452 13400
rect 24504 13428 24510 13440
rect 25200 13437 25228 13468
rect 25185 13431 25243 13437
rect 24504 13400 25136 13428
rect 24504 13388 24510 13400
rect 21226 13360 21232 13372
rect 20232 13332 21232 13360
rect 21226 13320 21232 13332
rect 21284 13320 21290 13372
rect 21134 13292 21140 13304
rect 19680 13264 21140 13292
rect 21134 13252 21140 13264
rect 21192 13252 21198 13304
rect 25108 13292 25136 13400
rect 25185 13397 25197 13431
rect 25231 13397 25243 13431
rect 25185 13391 25243 13397
rect 25461 13431 25519 13437
rect 25461 13397 25473 13431
rect 25507 13428 25519 13431
rect 25550 13428 25556 13440
rect 25507 13400 25556 13428
rect 25507 13397 25519 13400
rect 25461 13391 25519 13397
rect 25550 13388 25556 13400
rect 25608 13428 25614 13440
rect 26838 13428 26844 13440
rect 25608 13400 26844 13428
rect 25608 13388 25614 13400
rect 26838 13388 26844 13400
rect 26896 13388 26902 13440
rect 30610 13292 30616 13304
rect 25108 13264 30616 13292
rect 30610 13252 30616 13264
rect 30668 13252 30674 13304
rect 11000 13202 34368 13224
rect 11000 13150 14142 13202
rect 14194 13150 14206 13202
rect 14258 13150 14270 13202
rect 14322 13150 14334 13202
rect 14386 13150 24142 13202
rect 24194 13150 24206 13202
rect 24258 13150 24270 13202
rect 24322 13150 24334 13202
rect 24386 13150 34368 13202
rect 11000 13128 34368 13150
rect 14602 13048 14608 13100
rect 14660 13088 14666 13100
rect 15341 13091 15399 13097
rect 15341 13088 15353 13091
rect 14660 13060 15353 13088
rect 14660 13048 14666 13060
rect 15341 13057 15353 13060
rect 15387 13057 15399 13091
rect 25182 13088 25188 13100
rect 25143 13060 25188 13088
rect 15341 13051 15399 13057
rect 25182 13048 25188 13060
rect 25240 13048 25246 13100
rect 13498 13020 13504 13032
rect 13459 12992 13504 13020
rect 13498 12980 13504 12992
rect 13556 12980 13562 13032
rect 18837 13023 18895 13029
rect 14252 12992 15292 13020
rect 14252 12964 14280 12992
rect 12670 12912 12676 12964
rect 12728 12952 12734 12964
rect 14234 12952 14240 12964
rect 12728 12924 12773 12952
rect 14147 12924 14240 12952
rect 12728 12912 12734 12924
rect 14234 12912 14240 12924
rect 14292 12912 14298 12964
rect 13130 12884 13136 12896
rect 13091 12856 13136 12884
rect 13130 12844 13136 12856
rect 13188 12844 13194 12896
rect 13406 12884 13412 12896
rect 13367 12856 13412 12884
rect 13406 12844 13412 12856
rect 13464 12844 13470 12896
rect 14326 12884 14332 12896
rect 14239 12856 14332 12884
rect 14326 12844 14332 12856
rect 14384 12884 14390 12896
rect 14881 12887 14939 12893
rect 14881 12884 14893 12887
rect 14384 12856 14893 12884
rect 14384 12844 14390 12856
rect 14881 12853 14893 12856
rect 14927 12884 14939 12887
rect 14970 12884 14976 12896
rect 14927 12856 14976 12884
rect 14927 12853 14939 12856
rect 14881 12847 14939 12853
rect 14970 12844 14976 12856
rect 15028 12844 15034 12896
rect 15065 12887 15123 12893
rect 15065 12853 15077 12887
rect 15111 12884 15123 12887
rect 15264 12884 15292 12992
rect 18837 12989 18849 13023
rect 18883 13020 18895 13023
rect 19570 13020 19576 13032
rect 18883 12992 19576 13020
rect 18883 12989 18895 12992
rect 18837 12983 18895 12989
rect 19570 12980 19576 12992
rect 19628 12980 19634 13032
rect 21594 12980 21600 13032
rect 21652 13020 21658 13032
rect 22609 13023 22667 13029
rect 22609 13020 22621 13023
rect 21652 12992 22621 13020
rect 21652 12980 21658 12992
rect 22609 12989 22621 12992
rect 22655 12989 22667 13023
rect 22609 12983 22667 12989
rect 18101 12955 18159 12961
rect 18101 12921 18113 12955
rect 18147 12952 18159 12955
rect 18650 12952 18656 12964
rect 18147 12924 18656 12952
rect 18147 12921 18159 12924
rect 18101 12915 18159 12921
rect 18650 12912 18656 12924
rect 18708 12912 18714 12964
rect 20600 12924 20812 12952
rect 15430 12884 15436 12896
rect 15111 12856 15436 12884
rect 15111 12853 15123 12856
rect 15065 12847 15123 12853
rect 15430 12844 15436 12856
rect 15488 12844 15494 12896
rect 18469 12887 18527 12893
rect 18469 12853 18481 12887
rect 18515 12884 18527 12887
rect 18558 12884 18564 12896
rect 18515 12856 18564 12884
rect 18515 12853 18527 12856
rect 18469 12847 18527 12853
rect 18558 12844 18564 12856
rect 18616 12844 18622 12896
rect 18745 12887 18803 12893
rect 18745 12853 18757 12887
rect 18791 12884 18803 12887
rect 18834 12884 18840 12896
rect 18791 12856 18840 12884
rect 18791 12853 18803 12856
rect 18745 12847 18803 12853
rect 17546 12776 17552 12828
rect 17604 12816 17610 12828
rect 18760 12816 18788 12847
rect 18834 12844 18840 12856
rect 18892 12884 18898 12896
rect 20600 12893 20628 12924
rect 20585 12887 20643 12893
rect 20585 12884 20597 12887
rect 18892 12856 20597 12884
rect 18892 12844 18898 12856
rect 20585 12853 20597 12856
rect 20631 12853 20643 12887
rect 20585 12847 20643 12853
rect 20677 12887 20735 12893
rect 20677 12853 20689 12887
rect 20723 12853 20735 12887
rect 20677 12847 20735 12853
rect 17604 12788 18788 12816
rect 17604 12776 17610 12788
rect 15522 12708 15528 12760
rect 15580 12748 15586 12760
rect 20582 12748 20588 12760
rect 15580 12720 20588 12748
rect 15580 12708 15586 12720
rect 20582 12708 20588 12720
rect 20640 12708 20646 12760
rect 20692 12748 20720 12847
rect 20784 12816 20812 12924
rect 21778 12912 21784 12964
rect 21836 12952 21842 12964
rect 21836 12924 23204 12952
rect 21836 12912 21842 12924
rect 21042 12884 21048 12896
rect 21003 12856 21048 12884
rect 21042 12844 21048 12856
rect 21100 12844 21106 12896
rect 21137 12887 21195 12893
rect 21137 12853 21149 12887
rect 21183 12853 21195 12887
rect 21137 12847 21195 12853
rect 21152 12816 21180 12847
rect 21226 12844 21232 12896
rect 21284 12884 21290 12896
rect 23176 12893 23204 12924
rect 22793 12887 22851 12893
rect 22793 12884 22805 12887
rect 21284 12856 22805 12884
rect 21284 12844 21290 12856
rect 22793 12853 22805 12856
rect 22839 12853 22851 12887
rect 22793 12847 22851 12853
rect 23161 12887 23219 12893
rect 23161 12853 23173 12887
rect 23207 12853 23219 12887
rect 23161 12847 23219 12853
rect 23250 12844 23256 12896
rect 23308 12884 23314 12896
rect 24998 12884 25004 12896
rect 23308 12856 23353 12884
rect 24959 12856 25004 12884
rect 23308 12844 23314 12856
rect 24998 12844 25004 12856
rect 25056 12844 25062 12896
rect 25826 12884 25832 12896
rect 25787 12856 25832 12884
rect 25826 12844 25832 12856
rect 25884 12844 25890 12896
rect 21686 12816 21692 12828
rect 20784 12788 21180 12816
rect 21647 12788 21692 12816
rect 21686 12776 21692 12788
rect 21744 12776 21750 12828
rect 22698 12776 22704 12828
rect 22756 12816 22762 12828
rect 29966 12816 29972 12828
rect 22756 12788 29972 12816
rect 22756 12776 22762 12788
rect 29966 12776 29972 12788
rect 30024 12776 30030 12828
rect 20950 12748 20956 12760
rect 20692 12720 20956 12748
rect 20950 12708 20956 12720
rect 21008 12748 21014 12760
rect 23250 12748 23256 12760
rect 21008 12720 23256 12748
rect 21008 12708 21014 12720
rect 23250 12708 23256 12720
rect 23308 12708 23314 12760
rect 25826 12748 25832 12760
rect 25787 12720 25832 12748
rect 25826 12708 25832 12720
rect 25884 12708 25890 12760
rect 11000 12658 34368 12680
rect 11000 12606 19142 12658
rect 19194 12606 19206 12658
rect 19258 12606 19270 12658
rect 19322 12606 19334 12658
rect 19386 12606 29142 12658
rect 29194 12606 29206 12658
rect 29258 12606 29270 12658
rect 29322 12606 29334 12658
rect 29386 12606 34368 12658
rect 11000 12584 34368 12606
rect 12489 12547 12547 12553
rect 12489 12513 12501 12547
rect 12535 12544 12547 12547
rect 13406 12544 13412 12556
rect 12535 12516 13412 12544
rect 12535 12513 12547 12516
rect 12489 12507 12547 12513
rect 13406 12504 13412 12516
rect 13464 12504 13470 12556
rect 14878 12504 14884 12556
rect 14936 12544 14942 12556
rect 22698 12544 22704 12556
rect 14936 12516 22704 12544
rect 14936 12504 14942 12516
rect 22698 12504 22704 12516
rect 22756 12504 22762 12556
rect 23710 12544 23716 12556
rect 22900 12516 23716 12544
rect 15062 12476 15068 12488
rect 14712 12448 15068 12476
rect 12854 12408 12860 12420
rect 12815 12380 12860 12408
rect 12854 12368 12860 12380
rect 12912 12368 12918 12420
rect 13225 12411 13283 12417
rect 13225 12377 13237 12411
rect 13271 12408 13283 12411
rect 14326 12408 14332 12420
rect 13271 12380 14332 12408
rect 13271 12377 13283 12380
rect 13225 12371 13283 12377
rect 14326 12368 14332 12380
rect 14384 12368 14390 12420
rect 14418 12368 14424 12420
rect 14476 12408 14482 12420
rect 14712 12417 14740 12448
rect 15062 12436 15068 12448
rect 15120 12476 15126 12488
rect 16629 12479 16687 12485
rect 15120 12448 15292 12476
rect 15120 12436 15126 12448
rect 15264 12417 15292 12448
rect 16629 12445 16641 12479
rect 16675 12476 16687 12479
rect 16902 12476 16908 12488
rect 16675 12448 16908 12476
rect 16675 12445 16687 12448
rect 16629 12439 16687 12445
rect 16902 12436 16908 12448
rect 16960 12436 16966 12488
rect 17362 12436 17368 12488
rect 17420 12436 17426 12488
rect 18374 12436 18380 12488
rect 18432 12476 18438 12488
rect 19662 12476 19668 12488
rect 18432 12448 19668 12476
rect 18432 12436 18438 12448
rect 19662 12436 19668 12448
rect 19720 12476 19726 12488
rect 21686 12476 21692 12488
rect 19720 12448 21456 12476
rect 21647 12448 21692 12476
rect 19720 12436 19726 12448
rect 21428 12420 21456 12448
rect 21686 12436 21692 12448
rect 21744 12436 21750 12488
rect 22900 12462 22928 12516
rect 23710 12504 23716 12516
rect 23768 12544 23774 12556
rect 24998 12544 25004 12556
rect 23768 12516 25004 12544
rect 23768 12504 23774 12516
rect 24998 12504 25004 12516
rect 25056 12504 25062 12556
rect 23250 12436 23256 12488
rect 23308 12476 23314 12488
rect 23437 12479 23495 12485
rect 23437 12476 23449 12479
rect 23308 12448 23449 12476
rect 23308 12436 23314 12448
rect 23437 12445 23449 12448
rect 23483 12445 23495 12479
rect 23437 12439 23495 12445
rect 14513 12411 14571 12417
rect 14513 12408 14525 12411
rect 14476 12380 14525 12408
rect 14476 12368 14482 12380
rect 14513 12377 14525 12380
rect 14559 12377 14571 12411
rect 14513 12371 14571 12377
rect 14697 12411 14755 12417
rect 14697 12377 14709 12411
rect 14743 12377 14755 12411
rect 14697 12371 14755 12377
rect 15249 12411 15307 12417
rect 15249 12377 15261 12411
rect 15295 12377 15307 12411
rect 15430 12408 15436 12420
rect 15343 12380 15436 12408
rect 15249 12371 15307 12377
rect 15430 12368 15436 12380
rect 15488 12408 15494 12420
rect 16258 12408 16264 12420
rect 15488 12380 16264 12408
rect 15488 12368 15494 12380
rect 16258 12368 16264 12380
rect 16316 12368 16322 12420
rect 19570 12408 19576 12420
rect 19531 12380 19576 12408
rect 19570 12368 19576 12380
rect 19628 12368 19634 12420
rect 20122 12408 20128 12420
rect 20083 12380 20128 12408
rect 20122 12368 20128 12380
rect 20180 12368 20186 12420
rect 21410 12408 21416 12420
rect 21323 12380 21416 12408
rect 21410 12368 21416 12380
rect 21468 12368 21474 12420
rect 25826 12408 25832 12420
rect 25787 12380 25832 12408
rect 25826 12368 25832 12380
rect 25884 12368 25890 12420
rect 12949 12343 13007 12349
rect 12949 12309 12961 12343
rect 12995 12340 13007 12343
rect 13038 12340 13044 12352
rect 12995 12312 13044 12340
rect 12995 12309 13007 12312
rect 12949 12303 13007 12309
rect 13038 12300 13044 12312
rect 13096 12300 13102 12352
rect 13133 12343 13191 12349
rect 13133 12309 13145 12343
rect 13179 12340 13191 12343
rect 14234 12340 14240 12352
rect 13179 12312 14240 12340
rect 13179 12309 13191 12312
rect 13133 12303 13191 12309
rect 14234 12300 14240 12312
rect 14292 12300 14298 12352
rect 16353 12343 16411 12349
rect 16353 12309 16365 12343
rect 16399 12340 16411 12343
rect 16718 12340 16724 12352
rect 16399 12312 16724 12340
rect 16399 12309 16411 12312
rect 16353 12303 16411 12309
rect 16718 12300 16724 12312
rect 16776 12300 16782 12352
rect 17822 12300 17828 12352
rect 17880 12340 17886 12352
rect 18377 12343 18435 12349
rect 18377 12340 18389 12343
rect 17880 12312 18389 12340
rect 17880 12300 17886 12312
rect 18377 12309 18389 12312
rect 18423 12309 18435 12343
rect 18377 12303 18435 12309
rect 19018 12300 19024 12352
rect 19076 12340 19082 12352
rect 20401 12343 20459 12349
rect 20401 12340 20413 12343
rect 19076 12312 20413 12340
rect 19076 12300 19082 12312
rect 20401 12309 20413 12312
rect 20447 12309 20459 12343
rect 20401 12303 20459 12309
rect 21686 12300 21692 12352
rect 21744 12340 21750 12352
rect 24906 12340 24912 12352
rect 21744 12312 24912 12340
rect 21744 12300 21750 12312
rect 24906 12300 24912 12312
rect 24964 12300 24970 12352
rect 18650 12232 18656 12284
rect 18708 12272 18714 12284
rect 19665 12275 19723 12281
rect 19665 12272 19677 12275
rect 18708 12244 19677 12272
rect 18708 12232 18714 12244
rect 19665 12241 19677 12244
rect 19711 12241 19723 12275
rect 19665 12235 19723 12241
rect 12670 12164 12676 12216
rect 12728 12204 12734 12216
rect 15522 12204 15528 12216
rect 12728 12176 15528 12204
rect 12728 12164 12734 12176
rect 15522 12164 15528 12176
rect 15580 12164 15586 12216
rect 15706 12204 15712 12216
rect 15667 12176 15712 12204
rect 15706 12164 15712 12176
rect 15764 12164 15770 12216
rect 17270 12164 17276 12216
rect 17328 12204 17334 12216
rect 21502 12204 21508 12216
rect 17328 12176 21508 12204
rect 17328 12164 17334 12176
rect 21502 12164 21508 12176
rect 21560 12164 21566 12216
rect 23986 12164 23992 12216
rect 24044 12204 24050 12216
rect 25277 12207 25335 12213
rect 25277 12204 25289 12207
rect 24044 12176 25289 12204
rect 24044 12164 24050 12176
rect 25277 12173 25289 12176
rect 25323 12173 25335 12207
rect 25277 12167 25335 12173
rect 11000 12114 34368 12136
rect 11000 12062 14142 12114
rect 14194 12062 14206 12114
rect 14258 12062 14270 12114
rect 14322 12062 14334 12114
rect 14386 12062 24142 12114
rect 24194 12062 24206 12114
rect 24258 12062 24270 12114
rect 24322 12062 24334 12114
rect 24386 12062 34368 12114
rect 11000 12040 34368 12062
rect 14510 11960 14516 12012
rect 14568 12000 14574 12012
rect 14568 11972 16212 12000
rect 14568 11960 14574 11972
rect 14421 11867 14479 11873
rect 14421 11833 14433 11867
rect 14467 11864 14479 11867
rect 15706 11864 15712 11876
rect 14467 11836 15712 11864
rect 14467 11833 14479 11836
rect 14421 11827 14479 11833
rect 15706 11824 15712 11836
rect 15764 11824 15770 11876
rect 16184 11873 16212 11972
rect 16258 11960 16264 12012
rect 16316 12000 16322 12012
rect 17641 12003 17699 12009
rect 17641 12000 17653 12003
rect 16316 11972 17653 12000
rect 16316 11960 16322 11972
rect 17641 11969 17653 11972
rect 17687 12000 17699 12003
rect 20122 12000 20128 12012
rect 17687 11972 20128 12000
rect 17687 11969 17699 11972
rect 17641 11963 17699 11969
rect 20122 11960 20128 11972
rect 20180 11960 20186 12012
rect 21042 11960 21048 12012
rect 21100 12000 21106 12012
rect 21137 12003 21195 12009
rect 21137 12000 21149 12003
rect 21100 11972 21149 12000
rect 21100 11960 21106 11972
rect 21137 11969 21149 11972
rect 21183 11969 21195 12003
rect 21137 11963 21195 11969
rect 16169 11867 16227 11873
rect 16169 11833 16181 11867
rect 16215 11833 16227 11867
rect 16169 11827 16227 11833
rect 16718 11824 16724 11876
rect 16776 11864 16782 11876
rect 18374 11864 18380 11876
rect 16776 11836 18380 11864
rect 16776 11824 16782 11836
rect 18374 11824 18380 11836
rect 18432 11824 18438 11876
rect 18650 11864 18656 11876
rect 18611 11836 18656 11864
rect 18650 11824 18656 11836
rect 18708 11824 18714 11876
rect 18742 11824 18748 11876
rect 18800 11864 18806 11876
rect 18800 11836 20444 11864
rect 18800 11824 18806 11836
rect 14145 11799 14203 11805
rect 14145 11765 14157 11799
rect 14191 11765 14203 11799
rect 17822 11796 17828 11808
rect 17783 11768 17828 11796
rect 14145 11759 14203 11765
rect 14160 11660 14188 11759
rect 17822 11756 17828 11768
rect 17880 11756 17886 11808
rect 19754 11756 19760 11808
rect 19812 11756 19818 11808
rect 20416 11805 20444 11836
rect 21410 11824 21416 11876
rect 21468 11864 21474 11876
rect 26838 11864 26844 11876
rect 21468 11836 22192 11864
rect 21468 11824 21474 11836
rect 20401 11799 20459 11805
rect 20401 11765 20413 11799
rect 20447 11796 20459 11799
rect 21505 11799 21563 11805
rect 21505 11796 21517 11799
rect 20447 11768 21517 11796
rect 20447 11765 20459 11768
rect 20401 11759 20459 11765
rect 21505 11765 21517 11768
rect 21551 11796 21563 11799
rect 21778 11796 21784 11808
rect 21551 11768 21784 11796
rect 21551 11765 21563 11768
rect 21505 11759 21563 11765
rect 21778 11756 21784 11768
rect 21836 11756 21842 11808
rect 22164 11796 22192 11836
rect 22348 11836 23848 11864
rect 26799 11836 26844 11864
rect 22348 11805 22376 11836
rect 22333 11799 22391 11805
rect 22333 11796 22345 11799
rect 22164 11768 22345 11796
rect 22333 11765 22345 11768
rect 22379 11765 22391 11799
rect 23820 11796 23848 11836
rect 26838 11824 26844 11836
rect 26896 11824 26902 11876
rect 24814 11796 24820 11808
rect 23820 11768 24820 11796
rect 22333 11759 22391 11765
rect 24814 11756 24820 11768
rect 24872 11756 24878 11808
rect 16074 11728 16080 11740
rect 15646 11700 16080 11728
rect 16074 11688 16080 11700
rect 16132 11688 16138 11740
rect 22609 11731 22667 11737
rect 22609 11728 22621 11731
rect 20508 11700 22621 11728
rect 16718 11660 16724 11672
rect 14160 11632 16724 11660
rect 16718 11620 16724 11632
rect 16776 11620 16782 11672
rect 19478 11620 19484 11672
rect 19536 11660 19542 11672
rect 20508 11660 20536 11700
rect 22609 11697 22621 11700
rect 22655 11697 22667 11731
rect 22609 11691 22667 11697
rect 23158 11688 23164 11740
rect 23216 11688 23222 11740
rect 24357 11731 24415 11737
rect 24357 11697 24369 11731
rect 24403 11728 24415 11731
rect 25093 11731 25151 11737
rect 25093 11728 25105 11731
rect 24403 11700 25105 11728
rect 24403 11697 24415 11700
rect 24357 11691 24415 11697
rect 25093 11697 25105 11700
rect 25139 11697 25151 11731
rect 25093 11691 25151 11697
rect 25550 11688 25556 11740
rect 25608 11688 25614 11740
rect 19536 11632 20536 11660
rect 19536 11620 19542 11632
rect 11000 11570 34368 11592
rect 11000 11518 19142 11570
rect 19194 11518 19206 11570
rect 19258 11518 19270 11570
rect 19322 11518 19334 11570
rect 19386 11518 29142 11570
rect 29194 11518 29206 11570
rect 29258 11518 29270 11570
rect 29322 11518 29334 11570
rect 29386 11518 34368 11570
rect 11000 11496 34368 11518
rect 14970 11456 14976 11468
rect 14931 11428 14976 11456
rect 14970 11416 14976 11428
rect 15028 11416 15034 11468
rect 16074 11456 16080 11468
rect 16035 11428 16080 11456
rect 16074 11416 16080 11428
rect 16132 11416 16138 11468
rect 17362 11416 17368 11468
rect 17420 11456 17426 11468
rect 17457 11459 17515 11465
rect 17457 11456 17469 11459
rect 17420 11428 17469 11456
rect 17420 11416 17426 11428
rect 17457 11425 17469 11428
rect 17503 11425 17515 11459
rect 17457 11419 17515 11425
rect 19754 11416 19760 11468
rect 19812 11456 19818 11468
rect 19849 11459 19907 11465
rect 19849 11456 19861 11459
rect 19812 11428 19861 11456
rect 19812 11416 19818 11428
rect 19849 11425 19861 11428
rect 19895 11425 19907 11459
rect 21318 11456 21324 11468
rect 21279 11428 21324 11456
rect 19849 11419 19907 11425
rect 21318 11416 21324 11428
rect 21376 11416 21382 11468
rect 23158 11456 23164 11468
rect 23119 11428 23164 11456
rect 23158 11416 23164 11428
rect 23216 11416 23222 11468
rect 24725 11459 24783 11465
rect 24725 11425 24737 11459
rect 24771 11456 24783 11459
rect 25550 11456 25556 11468
rect 24771 11428 25556 11456
rect 24771 11425 24783 11428
rect 24725 11419 24783 11425
rect 25550 11416 25556 11428
rect 25608 11416 25614 11468
rect 25366 11388 25372 11400
rect 19680 11360 23020 11388
rect 25327 11360 25372 11388
rect 14510 11280 14516 11332
rect 14568 11320 14574 11332
rect 14789 11323 14847 11329
rect 14789 11320 14801 11323
rect 14568 11292 14801 11320
rect 14568 11280 14574 11292
rect 14789 11289 14801 11292
rect 14835 11289 14847 11323
rect 14789 11283 14847 11289
rect 15893 11323 15951 11329
rect 15893 11289 15905 11323
rect 15939 11320 15951 11323
rect 17086 11320 17092 11332
rect 15939 11292 17092 11320
rect 15939 11289 15951 11292
rect 15893 11283 15951 11289
rect 17086 11280 17092 11292
rect 17144 11320 17150 11332
rect 19680 11329 19708 11360
rect 17273 11323 17331 11329
rect 17273 11320 17285 11323
rect 17144 11292 17285 11320
rect 17144 11280 17150 11292
rect 17273 11289 17285 11292
rect 17319 11320 17331 11323
rect 19665 11323 19723 11329
rect 19665 11320 19677 11323
rect 17319 11292 19677 11320
rect 17319 11289 17331 11292
rect 17273 11283 17331 11289
rect 19665 11289 19677 11292
rect 19711 11289 19723 11323
rect 20950 11320 20956 11332
rect 20911 11292 20956 11320
rect 19665 11283 19723 11289
rect 20950 11280 20956 11292
rect 21008 11280 21014 11332
rect 22992 11329 23020 11360
rect 25366 11348 25372 11360
rect 25424 11348 25430 11400
rect 22977 11323 23035 11329
rect 22977 11289 22989 11323
rect 23023 11320 23035 11323
rect 23710 11320 23716 11332
rect 23023 11292 23716 11320
rect 23023 11289 23035 11292
rect 22977 11283 23035 11289
rect 23710 11280 23716 11292
rect 23768 11320 23774 11332
rect 24541 11323 24599 11329
rect 24541 11320 24553 11323
rect 23768 11292 24553 11320
rect 23768 11280 23774 11292
rect 24541 11289 24553 11292
rect 24587 11289 24599 11323
rect 24541 11283 24599 11289
rect 26013 11323 26071 11329
rect 26013 11289 26025 11323
rect 26059 11320 26071 11323
rect 30886 11320 30892 11332
rect 26059 11292 30892 11320
rect 26059 11289 26071 11292
rect 26013 11283 26071 11289
rect 30886 11280 30892 11292
rect 30944 11280 30950 11332
rect 11000 11026 34368 11048
rect 11000 10974 14142 11026
rect 14194 10974 14206 11026
rect 14258 10974 14270 11026
rect 14322 10974 14334 11026
rect 14386 10974 24142 11026
rect 24194 10974 24206 11026
rect 24258 10974 24270 11026
rect 24322 10974 24334 11026
rect 24386 10974 34368 11026
rect 11000 10952 34368 10974
<< via1 >>
rect 19142 34366 19194 34418
rect 19206 34366 19258 34418
rect 19270 34366 19322 34418
rect 19334 34366 19386 34418
rect 29142 34366 29194 34418
rect 29206 34366 29258 34418
rect 29270 34366 29322 34418
rect 29334 34366 29386 34418
rect 23624 34171 23676 34180
rect 23624 34137 23633 34171
rect 23633 34137 23667 34171
rect 23667 34137 23676 34171
rect 23624 34128 23676 34137
rect 26384 34128 26436 34180
rect 23440 33967 23492 33976
rect 23440 33933 23449 33967
rect 23449 33933 23483 33967
rect 23483 33933 23492 33967
rect 23440 33924 23492 33933
rect 25556 33967 25608 33976
rect 25556 33933 25565 33967
rect 25565 33933 25599 33967
rect 25599 33933 25608 33967
rect 25556 33924 25608 33933
rect 14142 33822 14194 33874
rect 14206 33822 14258 33874
rect 14270 33822 14322 33874
rect 14334 33822 14386 33874
rect 24142 33822 24194 33874
rect 24206 33822 24258 33874
rect 24270 33822 24322 33874
rect 24334 33822 24386 33874
rect 20128 33584 20180 33636
rect 20036 33516 20088 33568
rect 11020 33380 11072 33432
rect 20496 33448 20548 33500
rect 15436 33380 15488 33432
rect 16540 33380 16592 33432
rect 21508 33448 21560 33500
rect 21416 33423 21468 33432
rect 21416 33389 21425 33423
rect 21425 33389 21459 33423
rect 21459 33389 21468 33423
rect 25096 33584 25148 33636
rect 22428 33559 22480 33568
rect 22428 33525 22437 33559
rect 22437 33525 22471 33559
rect 22471 33525 22480 33559
rect 22428 33516 22480 33525
rect 23532 33516 23584 33568
rect 24176 33559 24228 33568
rect 24176 33525 24185 33559
rect 24185 33525 24219 33559
rect 24219 33525 24228 33559
rect 24176 33516 24228 33525
rect 22520 33491 22572 33500
rect 22520 33457 22529 33491
rect 22529 33457 22563 33491
rect 22563 33457 22572 33491
rect 22520 33448 22572 33457
rect 25004 33559 25056 33568
rect 25004 33525 25013 33559
rect 25013 33525 25047 33559
rect 25047 33525 25056 33559
rect 25004 33516 25056 33525
rect 33652 33584 33704 33636
rect 28040 33559 28092 33568
rect 28040 33525 28049 33559
rect 28049 33525 28083 33559
rect 28083 33525 28092 33559
rect 28040 33516 28092 33525
rect 28776 33516 28828 33568
rect 26200 33448 26252 33500
rect 26476 33448 26528 33500
rect 28132 33491 28184 33500
rect 28132 33457 28141 33491
rect 28141 33457 28175 33491
rect 28175 33457 28184 33491
rect 28132 33448 28184 33457
rect 21416 33380 21468 33389
rect 27120 33423 27172 33432
rect 27120 33389 27129 33423
rect 27129 33389 27163 33423
rect 27163 33389 27172 33423
rect 27120 33380 27172 33389
rect 27396 33380 27448 33432
rect 29512 33380 29564 33432
rect 19142 33278 19194 33330
rect 19206 33278 19258 33330
rect 19270 33278 19322 33330
rect 19334 33278 19386 33330
rect 29142 33278 29194 33330
rect 29206 33278 29258 33330
rect 29270 33278 29322 33330
rect 29334 33278 29386 33330
rect 24452 33176 24504 33228
rect 31444 33176 31496 33228
rect 20036 32972 20088 33024
rect 13964 32904 14016 32956
rect 20588 33040 20640 33092
rect 21508 33040 21560 33092
rect 22520 33108 22572 33160
rect 23624 33040 23676 33092
rect 27120 33108 27172 33160
rect 24176 33040 24228 33092
rect 24912 33040 24964 33092
rect 26292 33040 26344 33092
rect 28868 33040 28920 33092
rect 29052 33083 29104 33092
rect 29052 33049 29061 33083
rect 29061 33049 29095 33083
rect 29095 33049 29104 33083
rect 29052 33040 29104 33049
rect 30616 33040 30668 33092
rect 23716 32972 23768 33024
rect 25188 33015 25240 33024
rect 25188 32981 25197 33015
rect 25197 32981 25231 33015
rect 25231 32981 25240 33015
rect 25188 32972 25240 32981
rect 23072 32947 23124 32956
rect 23072 32913 23081 32947
rect 23081 32913 23115 32947
rect 23115 32913 23124 32947
rect 23072 32904 23124 32913
rect 25464 32904 25516 32956
rect 27120 32904 27172 32956
rect 21140 32879 21192 32888
rect 21140 32845 21149 32879
rect 21149 32845 21183 32879
rect 21183 32845 21192 32879
rect 21140 32836 21192 32845
rect 28408 32879 28460 32888
rect 28408 32845 28417 32879
rect 28417 32845 28451 32879
rect 28451 32845 28460 32879
rect 28408 32836 28460 32845
rect 29144 32879 29196 32888
rect 29144 32845 29153 32879
rect 29153 32845 29187 32879
rect 29187 32845 29196 32879
rect 29144 32836 29196 32845
rect 14142 32734 14194 32786
rect 14206 32734 14258 32786
rect 14270 32734 14322 32786
rect 14334 32734 14386 32786
rect 24142 32734 24194 32786
rect 24206 32734 24258 32786
rect 24270 32734 24322 32786
rect 24334 32734 24386 32786
rect 13228 32632 13280 32684
rect 21692 32632 21744 32684
rect 21324 32607 21376 32616
rect 21324 32573 21333 32607
rect 21333 32573 21367 32607
rect 21367 32573 21376 32607
rect 21324 32564 21376 32573
rect 22244 32564 22296 32616
rect 23532 32564 23584 32616
rect 21416 32496 21468 32548
rect 19760 32428 19812 32480
rect 21508 32471 21560 32480
rect 21508 32437 21517 32471
rect 21517 32437 21551 32471
rect 21551 32437 21560 32471
rect 21508 32428 21560 32437
rect 22888 32471 22940 32480
rect 22888 32437 22897 32471
rect 22897 32437 22931 32471
rect 22931 32437 22940 32471
rect 22888 32428 22940 32437
rect 25004 32564 25056 32616
rect 25464 32564 25516 32616
rect 24636 32496 24688 32548
rect 25924 32496 25976 32548
rect 27120 32539 27172 32548
rect 27120 32505 27129 32539
rect 27129 32505 27163 32539
rect 27163 32505 27172 32539
rect 27120 32496 27172 32505
rect 29144 32496 29196 32548
rect 25188 32428 25240 32480
rect 26292 32428 26344 32480
rect 28132 32428 28184 32480
rect 26476 32360 26528 32412
rect 27856 32360 27908 32412
rect 29052 32428 29104 32480
rect 28868 32403 28920 32412
rect 28868 32369 28877 32403
rect 28877 32369 28911 32403
rect 28911 32369 28920 32403
rect 28868 32360 28920 32369
rect 19142 32190 19194 32242
rect 19206 32190 19258 32242
rect 19270 32190 19322 32242
rect 19334 32190 19386 32242
rect 29142 32190 29194 32242
rect 29206 32190 29258 32242
rect 29270 32190 29322 32242
rect 29334 32190 29386 32242
rect 18196 32088 18248 32140
rect 19760 32063 19812 32072
rect 19760 32029 19769 32063
rect 19769 32029 19803 32063
rect 19803 32029 19812 32063
rect 19760 32020 19812 32029
rect 21508 32088 21560 32140
rect 23072 32020 23124 32072
rect 25464 32020 25516 32072
rect 25556 32020 25608 32072
rect 25924 32020 25976 32072
rect 26476 32063 26528 32072
rect 26476 32029 26485 32063
rect 26485 32029 26519 32063
rect 26519 32029 26528 32063
rect 26476 32020 26528 32029
rect 27856 32063 27908 32072
rect 27856 32029 27865 32063
rect 27865 32029 27899 32063
rect 27899 32029 27908 32063
rect 27856 32020 27908 32029
rect 28408 32020 28460 32072
rect 28868 32020 28920 32072
rect 20588 31995 20640 32004
rect 20588 31961 20597 31995
rect 20597 31961 20631 31995
rect 20631 31961 20640 31995
rect 20588 31952 20640 31961
rect 22244 31952 22296 32004
rect 23532 31995 23584 32004
rect 23532 31961 23541 31995
rect 23541 31961 23575 31995
rect 23575 31961 23584 31995
rect 23532 31952 23584 31961
rect 23624 31952 23676 32004
rect 25096 31952 25148 32004
rect 26200 31952 26252 32004
rect 28132 31952 28184 32004
rect 28592 31995 28644 32004
rect 28592 31961 28601 31995
rect 28601 31961 28635 31995
rect 28635 31961 28644 31995
rect 28592 31952 28644 31961
rect 23808 31884 23860 31936
rect 24728 31816 24780 31868
rect 14142 31646 14194 31698
rect 14206 31646 14258 31698
rect 14270 31646 14322 31698
rect 14334 31646 14386 31698
rect 24142 31646 24194 31698
rect 24206 31646 24258 31698
rect 24270 31646 24322 31698
rect 24334 31646 24386 31698
rect 23716 31544 23768 31596
rect 20496 31519 20548 31528
rect 20496 31485 20505 31519
rect 20505 31485 20539 31519
rect 20539 31485 20548 31519
rect 20496 31476 20548 31485
rect 21324 31476 21376 31528
rect 20036 31451 20088 31460
rect 20036 31417 20045 31451
rect 20045 31417 20079 31451
rect 20079 31417 20088 31451
rect 20036 31408 20088 31417
rect 21140 31408 21192 31460
rect 23348 31408 23400 31460
rect 23440 31408 23492 31460
rect 23808 31340 23860 31392
rect 25464 31340 25516 31392
rect 28960 31340 29012 31392
rect 20956 31272 21008 31324
rect 23532 31272 23584 31324
rect 24084 31272 24136 31324
rect 24544 31315 24596 31324
rect 24544 31281 24553 31315
rect 24553 31281 24587 31315
rect 24587 31281 24596 31315
rect 24544 31272 24596 31281
rect 29788 31272 29840 31324
rect 31260 31272 31312 31324
rect 21140 31204 21192 31256
rect 29604 31204 29656 31256
rect 29696 31204 29748 31256
rect 19142 31102 19194 31154
rect 19206 31102 19258 31154
rect 19270 31102 19322 31154
rect 19334 31102 19386 31154
rect 29142 31102 29194 31154
rect 29206 31102 29258 31154
rect 29270 31102 29322 31154
rect 29334 31102 29386 31154
rect 22428 31000 22480 31052
rect 21140 30932 21192 30984
rect 20128 30907 20180 30916
rect 20128 30873 20137 30907
rect 20137 30873 20171 30907
rect 20171 30873 20180 30907
rect 20128 30864 20180 30873
rect 22244 30864 22296 30916
rect 22520 30864 22572 30916
rect 22888 30932 22940 30984
rect 23256 30864 23308 30916
rect 26752 30864 26804 30916
rect 28500 30864 28552 30916
rect 29696 30907 29748 30916
rect 29696 30873 29705 30907
rect 29705 30873 29739 30907
rect 29739 30873 29748 30907
rect 29696 30864 29748 30873
rect 29972 30864 30024 30916
rect 31260 30907 31312 30916
rect 31260 30873 31269 30907
rect 31269 30873 31303 30907
rect 31303 30873 31312 30907
rect 31260 30864 31312 30873
rect 21140 30796 21192 30848
rect 21600 30796 21652 30848
rect 21692 30796 21744 30848
rect 22428 30796 22480 30848
rect 23348 30796 23400 30848
rect 25372 30796 25424 30848
rect 26200 30839 26252 30848
rect 26200 30805 26209 30839
rect 26209 30805 26243 30839
rect 26243 30805 26252 30839
rect 26200 30796 26252 30805
rect 26844 30796 26896 30848
rect 30800 30839 30852 30848
rect 30800 30805 30809 30839
rect 30809 30805 30843 30839
rect 30843 30805 30852 30839
rect 30800 30796 30852 30805
rect 32640 30796 32692 30848
rect 24084 30728 24136 30780
rect 26384 30728 26436 30780
rect 28592 30728 28644 30780
rect 29052 30728 29104 30780
rect 21232 30660 21284 30712
rect 23992 30660 24044 30712
rect 14142 30558 14194 30610
rect 14206 30558 14258 30610
rect 14270 30558 14322 30610
rect 14334 30558 14386 30610
rect 24142 30558 24194 30610
rect 24206 30558 24258 30610
rect 24270 30558 24322 30610
rect 24334 30558 24386 30610
rect 32640 30499 32692 30508
rect 32640 30465 32649 30499
rect 32649 30465 32683 30499
rect 32683 30465 32692 30499
rect 32640 30456 32692 30465
rect 16816 30388 16868 30440
rect 30616 30388 30668 30440
rect 31260 30388 31312 30440
rect 20128 30320 20180 30372
rect 26292 30320 26344 30372
rect 28500 30363 28552 30372
rect 28500 30329 28509 30363
rect 28509 30329 28543 30363
rect 28543 30329 28552 30363
rect 28500 30320 28552 30329
rect 28960 30320 29012 30372
rect 16172 30252 16224 30304
rect 17828 30116 17880 30168
rect 18472 30116 18524 30168
rect 20220 30252 20272 30304
rect 19944 30184 19996 30236
rect 20588 30184 20640 30236
rect 21600 30252 21652 30304
rect 25096 30295 25148 30304
rect 22336 30227 22388 30236
rect 22336 30193 22345 30227
rect 22345 30193 22379 30227
rect 22379 30193 22388 30227
rect 22336 30184 22388 30193
rect 23072 30227 23124 30236
rect 20404 30159 20456 30168
rect 20404 30125 20413 30159
rect 20413 30125 20447 30159
rect 20447 30125 20456 30159
rect 20404 30116 20456 30125
rect 22244 30116 22296 30168
rect 22612 30159 22664 30168
rect 22612 30125 22621 30159
rect 22621 30125 22655 30159
rect 22655 30125 22664 30159
rect 23072 30193 23081 30227
rect 23081 30193 23115 30227
rect 23115 30193 23124 30227
rect 23072 30184 23124 30193
rect 25096 30261 25105 30295
rect 25105 30261 25139 30295
rect 25139 30261 25148 30295
rect 25096 30252 25148 30261
rect 25832 30252 25884 30304
rect 26752 30295 26804 30304
rect 26752 30261 26761 30295
rect 26761 30261 26795 30295
rect 26795 30261 26804 30295
rect 26752 30252 26804 30261
rect 27120 30252 27172 30304
rect 30800 30252 30852 30304
rect 31444 30252 31496 30304
rect 29052 30184 29104 30236
rect 22612 30116 22664 30125
rect 22980 30116 23032 30168
rect 24728 30159 24780 30168
rect 24728 30125 24737 30159
rect 24737 30125 24771 30159
rect 24771 30125 24780 30159
rect 24728 30116 24780 30125
rect 31904 30159 31956 30168
rect 31904 30125 31913 30159
rect 31913 30125 31947 30159
rect 31947 30125 31956 30159
rect 31904 30116 31956 30125
rect 32824 30116 32876 30168
rect 19142 30014 19194 30066
rect 19206 30014 19258 30066
rect 19270 30014 19322 30066
rect 19334 30014 19386 30066
rect 29142 30014 29194 30066
rect 29206 30014 29258 30066
rect 29270 30014 29322 30066
rect 29334 30014 29386 30066
rect 17828 29844 17880 29896
rect 20220 29844 20272 29896
rect 20956 29887 21008 29896
rect 14516 29776 14568 29828
rect 16172 29819 16224 29828
rect 16172 29785 16181 29819
rect 16181 29785 16215 29819
rect 16215 29785 16224 29819
rect 16172 29776 16224 29785
rect 16816 29819 16868 29828
rect 16816 29785 16825 29819
rect 16825 29785 16859 29819
rect 16859 29785 16868 29819
rect 16816 29776 16868 29785
rect 17092 29751 17144 29760
rect 17092 29717 17101 29751
rect 17101 29717 17135 29751
rect 17135 29717 17144 29751
rect 17092 29708 17144 29717
rect 18472 29708 18524 29760
rect 19944 29708 19996 29760
rect 20680 29776 20732 29828
rect 20956 29853 20965 29887
rect 20965 29853 20999 29887
rect 20999 29853 21008 29887
rect 20956 29844 21008 29853
rect 23072 29912 23124 29964
rect 24452 29912 24504 29964
rect 25096 29912 25148 29964
rect 26936 29912 26988 29964
rect 20864 29776 20916 29828
rect 22520 29844 22572 29896
rect 22704 29887 22756 29896
rect 22704 29853 22713 29887
rect 22713 29853 22747 29887
rect 22747 29853 22756 29887
rect 22704 29844 22756 29853
rect 22244 29776 22296 29828
rect 23256 29844 23308 29896
rect 25280 29844 25332 29896
rect 23348 29776 23400 29828
rect 23992 29776 24044 29828
rect 25188 29819 25240 29828
rect 25188 29785 25197 29819
rect 25197 29785 25231 29819
rect 25231 29785 25240 29819
rect 25188 29776 25240 29785
rect 16356 29615 16408 29624
rect 16356 29581 16365 29615
rect 16365 29581 16399 29615
rect 16399 29581 16408 29615
rect 16356 29572 16408 29581
rect 22336 29708 22388 29760
rect 22888 29708 22940 29760
rect 24636 29708 24688 29760
rect 24544 29640 24596 29692
rect 25464 29776 25516 29828
rect 25832 29776 25884 29828
rect 26384 29819 26436 29828
rect 26384 29785 26393 29819
rect 26393 29785 26427 29819
rect 26427 29785 26436 29819
rect 26384 29776 26436 29785
rect 27396 29819 27448 29828
rect 27396 29785 27405 29819
rect 27405 29785 27439 29819
rect 27439 29785 27448 29819
rect 27396 29776 27448 29785
rect 27856 29819 27908 29828
rect 27856 29785 27865 29819
rect 27865 29785 27899 29819
rect 27899 29785 27908 29819
rect 27856 29776 27908 29785
rect 31812 29912 31864 29964
rect 28500 29887 28552 29896
rect 28500 29853 28509 29887
rect 28509 29853 28543 29887
rect 28543 29853 28552 29887
rect 28500 29844 28552 29853
rect 29604 29844 29656 29896
rect 31168 29844 31220 29896
rect 28960 29776 29012 29828
rect 29972 29819 30024 29828
rect 29972 29785 29981 29819
rect 29981 29785 30015 29819
rect 30015 29785 30024 29819
rect 29972 29776 30024 29785
rect 31904 29844 31956 29896
rect 26752 29708 26804 29760
rect 28868 29640 28920 29692
rect 30892 29751 30944 29760
rect 30892 29717 30901 29751
rect 30901 29717 30935 29751
rect 30935 29717 30944 29751
rect 30892 29708 30944 29717
rect 31168 29708 31220 29760
rect 32824 29683 32876 29692
rect 32824 29649 32833 29683
rect 32833 29649 32867 29683
rect 32867 29649 32876 29683
rect 32824 29640 32876 29649
rect 26108 29572 26160 29624
rect 14142 29470 14194 29522
rect 14206 29470 14258 29522
rect 14270 29470 14322 29522
rect 14334 29470 14386 29522
rect 24142 29470 24194 29522
rect 24206 29470 24258 29522
rect 24270 29470 24322 29522
rect 24334 29470 24386 29522
rect 23992 29368 24044 29420
rect 28040 29368 28092 29420
rect 13964 29300 14016 29352
rect 27948 29300 28000 29352
rect 29604 29300 29656 29352
rect 21232 29232 21284 29284
rect 21876 29232 21928 29284
rect 25832 29275 25884 29284
rect 25832 29241 25841 29275
rect 25841 29241 25875 29275
rect 25875 29241 25884 29275
rect 25832 29232 25884 29241
rect 17000 29207 17052 29216
rect 17000 29173 17009 29207
rect 17009 29173 17043 29207
rect 17043 29173 17052 29207
rect 17000 29164 17052 29173
rect 17184 29164 17236 29216
rect 17276 29207 17328 29216
rect 17276 29173 17285 29207
rect 17285 29173 17319 29207
rect 17319 29173 17328 29207
rect 17276 29164 17328 29173
rect 17736 29164 17788 29216
rect 21416 29164 21468 29216
rect 22704 29164 22756 29216
rect 24452 29207 24504 29216
rect 24452 29173 24461 29207
rect 24461 29173 24495 29207
rect 24495 29173 24504 29207
rect 24452 29164 24504 29173
rect 25096 29164 25148 29216
rect 25464 29207 25516 29216
rect 25464 29173 25474 29207
rect 25474 29173 25508 29207
rect 25508 29173 25516 29207
rect 25464 29164 25516 29173
rect 19944 29096 19996 29148
rect 20956 29139 21008 29148
rect 20956 29105 20965 29139
rect 20965 29105 20999 29139
rect 20999 29105 21008 29139
rect 20956 29096 21008 29105
rect 22888 29096 22940 29148
rect 23348 29139 23400 29148
rect 23348 29105 23357 29139
rect 23357 29105 23391 29139
rect 23391 29105 23400 29139
rect 23348 29096 23400 29105
rect 23716 29139 23768 29148
rect 23716 29105 23725 29139
rect 23725 29105 23759 29139
rect 23759 29105 23768 29139
rect 23716 29096 23768 29105
rect 23900 29096 23952 29148
rect 25556 29096 25608 29148
rect 26568 29164 26620 29216
rect 28960 29207 29012 29216
rect 28960 29173 28969 29207
rect 28969 29173 29003 29207
rect 29003 29173 29012 29207
rect 28960 29164 29012 29173
rect 31168 29164 31220 29216
rect 32824 29164 32876 29216
rect 26292 29139 26344 29148
rect 26292 29105 26301 29139
rect 26301 29105 26335 29139
rect 26335 29105 26344 29139
rect 26292 29096 26344 29105
rect 26660 29096 26712 29148
rect 29512 29139 29564 29148
rect 29512 29105 29521 29139
rect 29521 29105 29555 29139
rect 29555 29105 29564 29139
rect 31444 29139 31496 29148
rect 29512 29096 29564 29105
rect 31444 29105 31453 29139
rect 31453 29105 31487 29139
rect 31487 29105 31496 29139
rect 31444 29096 31496 29105
rect 20496 29028 20548 29080
rect 22704 29028 22756 29080
rect 23164 29071 23216 29080
rect 23164 29037 23173 29071
rect 23173 29037 23207 29071
rect 23207 29037 23216 29071
rect 23164 29028 23216 29037
rect 25096 29028 25148 29080
rect 26384 29028 26436 29080
rect 19142 28926 19194 28978
rect 19206 28926 19258 28978
rect 19270 28926 19322 28978
rect 19334 28926 19386 28978
rect 29142 28926 29194 28978
rect 29206 28926 29258 28978
rect 29270 28926 29322 28978
rect 29334 28926 29386 28978
rect 16908 28824 16960 28876
rect 23164 28824 23216 28876
rect 24452 28824 24504 28876
rect 25464 28867 25516 28876
rect 25464 28833 25473 28867
rect 25473 28833 25507 28867
rect 25507 28833 25516 28867
rect 25464 28824 25516 28833
rect 29512 28824 29564 28876
rect 31444 28824 31496 28876
rect 16356 28756 16408 28808
rect 17276 28756 17328 28808
rect 14516 28688 14568 28740
rect 14792 28688 14844 28740
rect 15344 28731 15396 28740
rect 15344 28697 15353 28731
rect 15353 28697 15387 28731
rect 15387 28697 15396 28731
rect 15344 28688 15396 28697
rect 17000 28688 17052 28740
rect 20956 28756 21008 28808
rect 21416 28799 21468 28808
rect 21416 28765 21425 28799
rect 21425 28765 21459 28799
rect 21459 28765 21468 28799
rect 21416 28756 21468 28765
rect 21692 28756 21744 28808
rect 22888 28799 22940 28808
rect 22888 28765 22897 28799
rect 22897 28765 22931 28799
rect 22931 28765 22940 28799
rect 22888 28756 22940 28765
rect 22980 28756 23032 28808
rect 23716 28756 23768 28808
rect 16816 28620 16868 28672
rect 17736 28620 17788 28672
rect 18288 28663 18340 28672
rect 18288 28629 18297 28663
rect 18297 28629 18331 28663
rect 18331 28629 18340 28663
rect 18288 28620 18340 28629
rect 20496 28552 20548 28604
rect 21508 28688 21560 28740
rect 22612 28688 22664 28740
rect 22704 28688 22756 28740
rect 21784 28663 21836 28672
rect 21784 28629 21793 28663
rect 21793 28629 21827 28663
rect 21827 28629 21836 28663
rect 21784 28620 21836 28629
rect 21876 28620 21928 28672
rect 25096 28688 25148 28740
rect 28960 28756 29012 28808
rect 24452 28620 24504 28672
rect 27028 28663 27080 28672
rect 27028 28629 27037 28663
rect 27037 28629 27071 28663
rect 27071 28629 27080 28663
rect 27028 28620 27080 28629
rect 27948 28731 28000 28740
rect 27948 28697 27957 28731
rect 27957 28697 27991 28731
rect 27991 28697 28000 28731
rect 27948 28688 28000 28697
rect 29972 28688 30024 28740
rect 31352 28688 31404 28740
rect 28960 28620 29012 28672
rect 23072 28552 23124 28604
rect 14516 28484 14568 28536
rect 26752 28484 26804 28536
rect 14142 28382 14194 28434
rect 14206 28382 14258 28434
rect 14270 28382 14322 28434
rect 14334 28382 14386 28434
rect 24142 28382 24194 28434
rect 24206 28382 24258 28434
rect 24270 28382 24322 28434
rect 24334 28382 24386 28434
rect 22428 28280 22480 28332
rect 25832 28280 25884 28332
rect 14148 28144 14200 28196
rect 16816 28144 16868 28196
rect 23348 28212 23400 28264
rect 17184 28119 17236 28128
rect 17184 28085 17193 28119
rect 17193 28085 17227 28119
rect 17227 28085 17236 28119
rect 17184 28076 17236 28085
rect 17644 28119 17696 28128
rect 14516 28008 14568 28060
rect 15436 28008 15488 28060
rect 17644 28085 17653 28119
rect 17653 28085 17687 28119
rect 17687 28085 17696 28119
rect 17644 28076 17696 28085
rect 17736 28076 17788 28128
rect 18196 28119 18248 28128
rect 18196 28085 18205 28119
rect 18205 28085 18239 28119
rect 18239 28085 18248 28119
rect 18196 28076 18248 28085
rect 13780 27940 13832 27992
rect 15344 27940 15396 27992
rect 18288 28008 18340 28060
rect 20036 28119 20088 28128
rect 20036 28085 20045 28119
rect 20045 28085 20079 28119
rect 20079 28085 20088 28119
rect 20036 28076 20088 28085
rect 22336 28119 22388 28128
rect 20496 28008 20548 28060
rect 22336 28085 22345 28119
rect 22345 28085 22379 28119
rect 22379 28085 22388 28119
rect 22336 28076 22388 28085
rect 22612 28144 22664 28196
rect 20404 27940 20456 27992
rect 22612 28008 22664 28060
rect 27120 28212 27172 28264
rect 25096 28144 25148 28196
rect 22888 28051 22940 28060
rect 22888 28017 22897 28051
rect 22897 28017 22931 28051
rect 22931 28017 22940 28051
rect 22888 28008 22940 28017
rect 23348 28051 23400 28060
rect 23348 28017 23357 28051
rect 23357 28017 23391 28051
rect 23391 28017 23400 28051
rect 23348 28008 23400 28017
rect 25464 28076 25516 28128
rect 26844 28144 26896 28196
rect 31076 28144 31128 28196
rect 28592 28119 28644 28128
rect 28592 28085 28601 28119
rect 28601 28085 28635 28119
rect 28635 28085 28644 28119
rect 28592 28076 28644 28085
rect 28960 28076 29012 28128
rect 23624 27983 23676 27992
rect 23624 27949 23633 27983
rect 23633 27949 23667 27983
rect 23667 27949 23676 27983
rect 23624 27940 23676 27949
rect 25924 28008 25976 28060
rect 26292 28051 26344 28060
rect 26292 28017 26301 28051
rect 26301 28017 26335 28051
rect 26335 28017 26344 28051
rect 26292 28008 26344 28017
rect 25004 27940 25056 27992
rect 25648 27940 25700 27992
rect 29512 27940 29564 27992
rect 19142 27838 19194 27890
rect 19206 27838 19258 27890
rect 19270 27838 19322 27890
rect 19334 27838 19386 27890
rect 29142 27838 29194 27890
rect 29206 27838 29258 27890
rect 29270 27838 29322 27890
rect 29334 27838 29386 27890
rect 20220 27779 20272 27788
rect 20220 27745 20229 27779
rect 20229 27745 20263 27779
rect 20263 27745 20272 27779
rect 20220 27736 20272 27745
rect 20588 27736 20640 27788
rect 14148 27668 14200 27720
rect 17092 27668 17144 27720
rect 20404 27711 20456 27720
rect 20404 27677 20413 27711
rect 20413 27677 20447 27711
rect 20447 27677 20456 27711
rect 20404 27668 20456 27677
rect 20496 27668 20548 27720
rect 21416 27668 21468 27720
rect 24820 27736 24872 27788
rect 14700 27643 14752 27652
rect 14700 27609 14709 27643
rect 14709 27609 14743 27643
rect 14743 27609 14752 27643
rect 14700 27600 14752 27609
rect 15068 27600 15120 27652
rect 14608 27532 14660 27584
rect 15344 27575 15396 27584
rect 15344 27541 15353 27575
rect 15353 27541 15387 27575
rect 15387 27541 15396 27575
rect 15344 27532 15396 27541
rect 15528 27532 15580 27584
rect 16908 27600 16960 27652
rect 17552 27643 17604 27652
rect 17552 27609 17561 27643
rect 17561 27609 17595 27643
rect 17595 27609 17604 27643
rect 17552 27600 17604 27609
rect 17644 27643 17696 27652
rect 17644 27609 17653 27643
rect 17653 27609 17687 27643
rect 17687 27609 17696 27643
rect 18104 27643 18156 27652
rect 17644 27600 17696 27609
rect 18104 27609 18113 27643
rect 18113 27609 18147 27643
rect 18147 27609 18156 27643
rect 18104 27600 18156 27609
rect 18472 27600 18524 27652
rect 20312 27643 20364 27652
rect 20312 27609 20321 27643
rect 20321 27609 20355 27643
rect 20355 27609 20364 27643
rect 20312 27600 20364 27609
rect 20588 27600 20640 27652
rect 21692 27643 21744 27652
rect 21692 27609 21701 27643
rect 21701 27609 21735 27643
rect 21735 27609 21744 27643
rect 21692 27600 21744 27609
rect 22612 27668 22664 27720
rect 22796 27668 22848 27720
rect 23072 27711 23124 27720
rect 23072 27677 23081 27711
rect 23081 27677 23115 27711
rect 23115 27677 23124 27711
rect 23072 27668 23124 27677
rect 24544 27668 24596 27720
rect 26568 27668 26620 27720
rect 24452 27600 24504 27652
rect 25372 27643 25424 27652
rect 25372 27609 25381 27643
rect 25381 27609 25415 27643
rect 25415 27609 25424 27643
rect 25372 27600 25424 27609
rect 25556 27643 25608 27652
rect 25556 27609 25565 27643
rect 25565 27609 25599 27643
rect 25599 27609 25608 27643
rect 25556 27600 25608 27609
rect 18196 27575 18248 27584
rect 18196 27541 18205 27575
rect 18205 27541 18239 27575
rect 18239 27541 18248 27575
rect 18196 27532 18248 27541
rect 19944 27532 19996 27584
rect 20956 27532 21008 27584
rect 21508 27575 21560 27584
rect 21508 27541 21517 27575
rect 21517 27541 21551 27575
rect 21551 27541 21560 27575
rect 21508 27532 21560 27541
rect 23532 27532 23584 27584
rect 25648 27532 25700 27584
rect 26292 27532 26344 27584
rect 26476 27532 26528 27584
rect 30892 27736 30944 27788
rect 27856 27600 27908 27652
rect 28500 27600 28552 27652
rect 27856 27464 27908 27516
rect 28592 27464 28644 27516
rect 21692 27396 21744 27448
rect 22796 27396 22848 27448
rect 25372 27396 25424 27448
rect 27304 27396 27356 27448
rect 28500 27396 28552 27448
rect 30340 27532 30392 27584
rect 14142 27294 14194 27346
rect 14206 27294 14258 27346
rect 14270 27294 14322 27346
rect 14334 27294 14386 27346
rect 24142 27294 24194 27346
rect 24206 27294 24258 27346
rect 24270 27294 24322 27346
rect 24334 27294 24386 27346
rect 22428 27192 22480 27244
rect 23440 27192 23492 27244
rect 25464 27192 25516 27244
rect 26660 27192 26712 27244
rect 14700 27056 14752 27108
rect 17000 27056 17052 27108
rect 17552 27124 17604 27176
rect 18012 27056 18064 27108
rect 21232 27056 21284 27108
rect 14516 27031 14568 27040
rect 14516 26997 14525 27031
rect 14525 26997 14559 27031
rect 14559 26997 14568 27031
rect 14516 26988 14568 26997
rect 14976 27031 15028 27040
rect 14976 26997 14985 27031
rect 14985 26997 15019 27031
rect 15019 26997 15028 27031
rect 14976 26988 15028 26997
rect 17276 26988 17328 27040
rect 17644 27031 17696 27040
rect 17644 26997 17653 27031
rect 17653 26997 17687 27031
rect 17687 26997 17696 27031
rect 17644 26988 17696 26997
rect 17920 26988 17972 27040
rect 20956 27031 21008 27040
rect 16632 26920 16684 26972
rect 20956 26997 20965 27031
rect 20965 26997 20999 27031
rect 20999 26997 21008 27031
rect 20956 26988 21008 26997
rect 21324 27031 21376 27040
rect 21324 26997 21333 27031
rect 21333 26997 21367 27031
rect 21367 26997 21376 27031
rect 21324 26988 21376 26997
rect 22612 26988 22664 27040
rect 23808 27056 23860 27108
rect 26108 27099 26160 27108
rect 26108 27065 26117 27099
rect 26117 27065 26151 27099
rect 26151 27065 26160 27099
rect 26108 27056 26160 27065
rect 23256 26988 23308 27040
rect 21784 26920 21836 26972
rect 22428 26963 22480 26972
rect 22428 26929 22437 26963
rect 22437 26929 22471 26963
rect 22471 26929 22480 26963
rect 22428 26920 22480 26929
rect 22980 26920 23032 26972
rect 23440 26920 23492 26972
rect 17092 26852 17144 26904
rect 20220 26852 20272 26904
rect 21968 26852 22020 26904
rect 25648 26920 25700 26972
rect 29604 26988 29656 27040
rect 29788 27056 29840 27108
rect 30340 27099 30392 27108
rect 30340 27065 30349 27099
rect 30349 27065 30383 27099
rect 30383 27065 30392 27099
rect 30340 27056 30392 27065
rect 31260 27099 31312 27108
rect 31260 27065 31269 27099
rect 31269 27065 31303 27099
rect 31303 27065 31312 27099
rect 31260 27056 31312 27065
rect 29512 26920 29564 26972
rect 29788 26963 29840 26972
rect 29788 26929 29797 26963
rect 29797 26929 29831 26963
rect 29831 26929 29840 26963
rect 29788 26920 29840 26929
rect 29880 26920 29932 26972
rect 25924 26852 25976 26904
rect 28960 26852 29012 26904
rect 19142 26750 19194 26802
rect 19206 26750 19258 26802
rect 19270 26750 19322 26802
rect 19334 26750 19386 26802
rect 29142 26750 29194 26802
rect 29206 26750 29258 26802
rect 29270 26750 29322 26802
rect 29334 26750 29386 26802
rect 17552 26648 17604 26700
rect 17920 26648 17972 26700
rect 20404 26648 20456 26700
rect 22612 26691 22664 26700
rect 22612 26657 22621 26691
rect 22621 26657 22655 26691
rect 22655 26657 22664 26691
rect 22612 26648 22664 26657
rect 25004 26648 25056 26700
rect 27580 26648 27632 26700
rect 27856 26648 27908 26700
rect 14516 26580 14568 26632
rect 17644 26580 17696 26632
rect 17828 26512 17880 26564
rect 19944 26580 19996 26632
rect 22428 26580 22480 26632
rect 23072 26580 23124 26632
rect 23624 26580 23676 26632
rect 26292 26580 26344 26632
rect 27028 26580 27080 26632
rect 19576 26555 19628 26564
rect 19576 26521 19585 26555
rect 19585 26521 19619 26555
rect 19619 26521 19628 26555
rect 19576 26512 19628 26521
rect 20220 26555 20272 26564
rect 20220 26521 20229 26555
rect 20229 26521 20263 26555
rect 20263 26521 20272 26555
rect 20220 26512 20272 26521
rect 20404 26555 20456 26564
rect 20404 26521 20413 26555
rect 20413 26521 20447 26555
rect 20447 26521 20456 26555
rect 20404 26512 20456 26521
rect 20496 26512 20548 26564
rect 21692 26512 21744 26564
rect 22244 26512 22296 26564
rect 23348 26512 23400 26564
rect 29788 26580 29840 26632
rect 27304 26555 27356 26564
rect 27304 26521 27313 26555
rect 27313 26521 27347 26555
rect 27347 26521 27356 26555
rect 27304 26512 27356 26521
rect 15436 26444 15488 26496
rect 18012 26487 18064 26496
rect 18012 26453 18021 26487
rect 18021 26453 18055 26487
rect 18055 26453 18064 26487
rect 18012 26444 18064 26453
rect 19668 26444 19720 26496
rect 26476 26487 26528 26496
rect 18104 26376 18156 26428
rect 18472 26376 18524 26428
rect 22612 26376 22664 26428
rect 26476 26453 26485 26487
rect 26485 26453 26519 26487
rect 26519 26453 26528 26487
rect 26476 26444 26528 26453
rect 23992 26376 24044 26428
rect 27580 26419 27632 26428
rect 27580 26385 27589 26419
rect 27589 26385 27623 26419
rect 27623 26385 27632 26419
rect 27580 26376 27632 26385
rect 19852 26308 19904 26360
rect 23256 26308 23308 26360
rect 25648 26308 25700 26360
rect 26752 26308 26804 26360
rect 29512 26555 29564 26564
rect 29512 26521 29521 26555
rect 29521 26521 29555 26555
rect 29555 26521 29564 26555
rect 29512 26512 29564 26521
rect 29604 26512 29656 26564
rect 31444 26555 31496 26564
rect 31444 26521 31453 26555
rect 31453 26521 31487 26555
rect 31487 26521 31496 26555
rect 31444 26512 31496 26521
rect 28408 26308 28460 26360
rect 30248 26308 30300 26360
rect 14142 26206 14194 26258
rect 14206 26206 14258 26258
rect 14270 26206 14322 26258
rect 14334 26206 14386 26258
rect 24142 26206 24194 26258
rect 24206 26206 24258 26258
rect 24270 26206 24322 26258
rect 24334 26206 24386 26258
rect 14608 26104 14660 26156
rect 22612 26147 22664 26156
rect 22612 26113 22621 26147
rect 22621 26113 22655 26147
rect 22655 26113 22664 26147
rect 22612 26104 22664 26113
rect 23992 26104 24044 26156
rect 21324 26036 21376 26088
rect 25464 26104 25516 26156
rect 25556 26036 25608 26088
rect 26476 26104 26528 26156
rect 14792 25968 14844 26020
rect 16908 25968 16960 26020
rect 17828 26011 17880 26020
rect 17828 25977 17837 26011
rect 17837 25977 17871 26011
rect 17871 25977 17880 26011
rect 17828 25968 17880 25977
rect 14516 25900 14568 25952
rect 14976 25900 15028 25952
rect 16632 25900 16684 25952
rect 17276 25900 17328 25952
rect 17552 25943 17604 25952
rect 17552 25909 17561 25943
rect 17561 25909 17595 25943
rect 17595 25909 17604 25943
rect 17552 25900 17604 25909
rect 19484 25968 19536 26020
rect 20312 25968 20364 26020
rect 22704 26011 22756 26020
rect 22704 25977 22713 26011
rect 22713 25977 22747 26011
rect 22747 25977 22756 26011
rect 22704 25968 22756 25977
rect 25188 25968 25240 26020
rect 26108 25968 26160 26020
rect 13964 25807 14016 25816
rect 13964 25773 13973 25807
rect 13973 25773 14007 25807
rect 14007 25773 14016 25807
rect 13964 25764 14016 25773
rect 20404 25900 20456 25952
rect 20956 25943 21008 25952
rect 20956 25909 20965 25943
rect 20965 25909 20999 25943
rect 20999 25909 21008 25943
rect 20956 25900 21008 25909
rect 21600 25900 21652 25952
rect 24544 25900 24596 25952
rect 25832 25900 25884 25952
rect 20312 25832 20364 25884
rect 22336 25875 22388 25884
rect 22336 25841 22345 25875
rect 22345 25841 22379 25875
rect 22379 25841 22388 25875
rect 22336 25832 22388 25841
rect 23808 25764 23860 25816
rect 24084 25832 24136 25884
rect 26384 25832 26436 25884
rect 26936 25943 26988 25952
rect 26936 25909 26945 25943
rect 26945 25909 26979 25943
rect 26979 25909 26988 25943
rect 26936 25900 26988 25909
rect 28316 25943 28368 25952
rect 28316 25909 28325 25943
rect 28325 25909 28359 25943
rect 28359 25909 28368 25943
rect 28316 25900 28368 25909
rect 25280 25764 25332 25816
rect 28224 25764 28276 25816
rect 29604 25832 29656 25884
rect 31444 26036 31496 26088
rect 30248 26011 30300 26020
rect 30248 25977 30257 26011
rect 30257 25977 30291 26011
rect 30291 25977 30300 26011
rect 30248 25968 30300 25977
rect 30524 25900 30576 25952
rect 31536 25900 31588 25952
rect 32180 25832 32232 25884
rect 31904 25807 31956 25816
rect 31904 25773 31913 25807
rect 31913 25773 31947 25807
rect 31947 25773 31956 25807
rect 31904 25764 31956 25773
rect 19142 25662 19194 25714
rect 19206 25662 19258 25714
rect 19270 25662 19322 25714
rect 19334 25662 19386 25714
rect 29142 25662 29194 25714
rect 29206 25662 29258 25714
rect 29270 25662 29322 25714
rect 29334 25662 29386 25714
rect 13964 25492 14016 25544
rect 17092 25535 17144 25544
rect 17092 25501 17101 25535
rect 17101 25501 17135 25535
rect 17135 25501 17144 25535
rect 17092 25492 17144 25501
rect 19484 25492 19536 25544
rect 13780 25424 13832 25476
rect 16724 25424 16776 25476
rect 17644 25424 17696 25476
rect 17828 25424 17880 25476
rect 19024 25424 19076 25476
rect 19576 25424 19628 25476
rect 19852 25467 19904 25476
rect 19852 25433 19861 25467
rect 19861 25433 19895 25467
rect 19895 25433 19904 25467
rect 19852 25424 19904 25433
rect 15988 25399 16040 25408
rect 15988 25365 15997 25399
rect 15997 25365 16031 25399
rect 16031 25365 16040 25399
rect 15988 25356 16040 25365
rect 20404 25467 20456 25476
rect 20404 25433 20413 25467
rect 20413 25433 20447 25467
rect 20447 25433 20456 25467
rect 20404 25424 20456 25433
rect 21416 25467 21468 25476
rect 21416 25433 21425 25467
rect 21425 25433 21459 25467
rect 21459 25433 21468 25467
rect 21416 25424 21468 25433
rect 21600 25467 21652 25476
rect 21600 25433 21609 25467
rect 21609 25433 21643 25467
rect 21643 25433 21652 25467
rect 21600 25424 21652 25433
rect 22704 25492 22756 25544
rect 22888 25492 22940 25544
rect 23532 25467 23584 25476
rect 23532 25433 23541 25467
rect 23541 25433 23575 25467
rect 23575 25433 23584 25467
rect 23532 25424 23584 25433
rect 25280 25492 25332 25544
rect 29512 25560 29564 25612
rect 32180 25603 32232 25612
rect 32180 25569 32189 25603
rect 32189 25569 32223 25603
rect 32223 25569 32232 25603
rect 32180 25560 32232 25569
rect 28316 25535 28368 25544
rect 28316 25501 28325 25535
rect 28325 25501 28359 25535
rect 28359 25501 28368 25535
rect 28316 25492 28368 25501
rect 29788 25535 29840 25544
rect 29788 25501 29797 25535
rect 29797 25501 29831 25535
rect 29831 25501 29840 25535
rect 29788 25492 29840 25501
rect 30524 25492 30576 25544
rect 31536 25535 31588 25544
rect 25832 25424 25884 25476
rect 22704 25399 22756 25408
rect 22704 25365 22713 25399
rect 22713 25365 22747 25399
rect 22747 25365 22756 25399
rect 22704 25356 22756 25365
rect 24636 25356 24688 25408
rect 26108 25424 26160 25476
rect 26384 25424 26436 25476
rect 17736 25288 17788 25340
rect 18656 25288 18708 25340
rect 28960 25424 29012 25476
rect 30616 25424 30668 25476
rect 31536 25501 31545 25535
rect 31545 25501 31579 25535
rect 31579 25501 31588 25535
rect 31536 25492 31588 25501
rect 32364 25467 32416 25476
rect 32364 25433 32373 25467
rect 32373 25433 32407 25467
rect 32407 25433 32416 25467
rect 32364 25424 32416 25433
rect 28592 25356 28644 25408
rect 13964 25220 14016 25272
rect 22612 25263 22664 25272
rect 22612 25229 22621 25263
rect 22621 25229 22655 25263
rect 22655 25229 22664 25263
rect 22612 25220 22664 25229
rect 25924 25220 25976 25272
rect 14142 25118 14194 25170
rect 14206 25118 14258 25170
rect 14270 25118 14322 25170
rect 14334 25118 14386 25170
rect 24142 25118 24194 25170
rect 24206 25118 24258 25170
rect 24270 25118 24322 25170
rect 24334 25118 24386 25170
rect 13964 24880 14016 24932
rect 15988 24880 16040 24932
rect 19484 24880 19536 24932
rect 14700 24855 14752 24864
rect 14700 24821 14709 24855
rect 14709 24821 14743 24855
rect 14743 24821 14752 24855
rect 14700 24812 14752 24821
rect 15068 24855 15120 24864
rect 13412 24744 13464 24796
rect 15068 24821 15077 24855
rect 15077 24821 15111 24855
rect 15111 24821 15120 24855
rect 15068 24812 15120 24821
rect 15528 24855 15580 24864
rect 15528 24821 15537 24855
rect 15537 24821 15571 24855
rect 15571 24821 15580 24855
rect 15528 24812 15580 24821
rect 16908 24855 16960 24864
rect 16908 24821 16917 24855
rect 16917 24821 16951 24855
rect 16951 24821 16960 24855
rect 16908 24812 16960 24821
rect 19576 24855 19628 24864
rect 17460 24787 17512 24796
rect 17460 24753 17469 24787
rect 17469 24753 17503 24787
rect 17503 24753 17512 24787
rect 17460 24744 17512 24753
rect 19576 24821 19585 24855
rect 19585 24821 19619 24855
rect 19619 24821 19628 24855
rect 19576 24812 19628 24821
rect 21048 25016 21100 25068
rect 23072 25016 23124 25068
rect 23900 25016 23952 25068
rect 25556 25016 25608 25068
rect 21600 24880 21652 24932
rect 21232 24855 21284 24864
rect 21232 24821 21241 24855
rect 21241 24821 21275 24855
rect 21275 24821 21284 24855
rect 21232 24812 21284 24821
rect 21324 24812 21376 24864
rect 22336 24855 22388 24864
rect 22336 24821 22345 24855
rect 22345 24821 22379 24855
rect 22379 24821 22388 24855
rect 22336 24812 22388 24821
rect 22704 24948 22756 25000
rect 23440 24948 23492 25000
rect 23072 24880 23124 24932
rect 25648 24923 25700 24932
rect 23440 24855 23492 24864
rect 23440 24821 23449 24855
rect 23449 24821 23483 24855
rect 23483 24821 23492 24855
rect 23440 24812 23492 24821
rect 25648 24889 25657 24923
rect 25657 24889 25691 24923
rect 25691 24889 25700 24923
rect 25648 24880 25700 24889
rect 26752 24880 26804 24932
rect 26384 24855 26436 24864
rect 26384 24821 26393 24855
rect 26393 24821 26427 24855
rect 26427 24821 26436 24855
rect 26384 24812 26436 24821
rect 28224 25059 28276 25068
rect 28224 25025 28233 25059
rect 28233 25025 28267 25059
rect 28267 25025 28276 25059
rect 28224 25016 28276 25025
rect 30708 24991 30760 25000
rect 30708 24957 30717 24991
rect 30717 24957 30751 24991
rect 30751 24957 30760 24991
rect 30708 24948 30760 24957
rect 31352 24948 31404 25000
rect 29880 24812 29932 24864
rect 30340 24855 30392 24864
rect 30340 24821 30349 24855
rect 30349 24821 30383 24855
rect 30383 24821 30392 24855
rect 30340 24812 30392 24821
rect 31168 24812 31220 24864
rect 32364 24855 32416 24864
rect 32364 24821 32373 24855
rect 32373 24821 32407 24855
rect 32407 24821 32416 24855
rect 32364 24812 32416 24821
rect 18656 24676 18708 24728
rect 19668 24744 19720 24796
rect 21508 24676 21560 24728
rect 23256 24744 23308 24796
rect 23348 24744 23400 24796
rect 25280 24744 25332 24796
rect 27028 24744 27080 24796
rect 27948 24787 28000 24796
rect 27948 24753 27957 24787
rect 27957 24753 27991 24787
rect 27991 24753 28000 24787
rect 27948 24744 28000 24753
rect 30248 24744 30300 24796
rect 22520 24676 22572 24728
rect 22980 24676 23032 24728
rect 24360 24676 24412 24728
rect 19142 24574 19194 24626
rect 19206 24574 19258 24626
rect 19270 24574 19322 24626
rect 19334 24574 19386 24626
rect 29142 24574 29194 24626
rect 29206 24574 29258 24626
rect 29270 24574 29322 24626
rect 29334 24574 29386 24626
rect 22612 24472 22664 24524
rect 25096 24472 25148 24524
rect 13412 24447 13464 24456
rect 13412 24413 13421 24447
rect 13421 24413 13455 24447
rect 13455 24413 13464 24447
rect 13412 24404 13464 24413
rect 16632 24404 16684 24456
rect 14608 24336 14660 24388
rect 14700 24336 14752 24388
rect 16908 24336 16960 24388
rect 17460 24379 17512 24388
rect 16632 24268 16684 24320
rect 17460 24345 17469 24379
rect 17469 24345 17503 24379
rect 17503 24345 17512 24379
rect 17460 24336 17512 24345
rect 17828 24379 17880 24388
rect 17828 24345 17837 24379
rect 17837 24345 17871 24379
rect 17871 24345 17880 24379
rect 17828 24336 17880 24345
rect 19576 24404 19628 24456
rect 18472 24379 18524 24388
rect 18472 24345 18481 24379
rect 18481 24345 18515 24379
rect 18515 24345 18524 24379
rect 18472 24336 18524 24345
rect 18656 24379 18708 24388
rect 18656 24345 18665 24379
rect 18665 24345 18699 24379
rect 18699 24345 18708 24379
rect 18656 24336 18708 24345
rect 19208 24336 19260 24388
rect 19484 24336 19536 24388
rect 19668 24379 19720 24388
rect 19668 24345 19677 24379
rect 19677 24345 19711 24379
rect 19711 24345 19720 24379
rect 19668 24336 19720 24345
rect 20036 24336 20088 24388
rect 22520 24379 22572 24388
rect 22520 24345 22529 24379
rect 22529 24345 22563 24379
rect 22563 24345 22572 24379
rect 22520 24336 22572 24345
rect 18932 24268 18984 24320
rect 19852 24268 19904 24320
rect 22428 24311 22480 24320
rect 22428 24277 22437 24311
rect 22437 24277 22471 24311
rect 22471 24277 22480 24311
rect 22888 24379 22940 24388
rect 22888 24345 22897 24379
rect 22897 24345 22931 24379
rect 22931 24345 22940 24379
rect 22888 24336 22940 24345
rect 23808 24336 23860 24388
rect 23992 24336 24044 24388
rect 24360 24379 24412 24388
rect 24360 24345 24369 24379
rect 24369 24345 24403 24379
rect 24403 24345 24412 24379
rect 24360 24336 24412 24345
rect 24820 24336 24872 24388
rect 25924 24447 25976 24456
rect 25924 24413 25933 24447
rect 25933 24413 25967 24447
rect 25967 24413 25976 24447
rect 25924 24404 25976 24413
rect 28868 24404 28920 24456
rect 25464 24379 25516 24388
rect 22428 24268 22480 24277
rect 23440 24268 23492 24320
rect 25464 24345 25473 24379
rect 25473 24345 25507 24379
rect 25507 24345 25516 24379
rect 25464 24336 25516 24345
rect 27028 24379 27080 24388
rect 27028 24345 27037 24379
rect 27037 24345 27071 24379
rect 27071 24345 27080 24379
rect 27028 24336 27080 24345
rect 27856 24379 27908 24388
rect 27856 24345 27865 24379
rect 27865 24345 27899 24379
rect 27899 24345 27908 24379
rect 28592 24379 28644 24388
rect 27856 24336 27908 24345
rect 26384 24268 26436 24320
rect 27948 24311 28000 24320
rect 27948 24277 27957 24311
rect 27957 24277 27991 24311
rect 27991 24277 28000 24311
rect 27948 24268 28000 24277
rect 28592 24345 28601 24379
rect 28601 24345 28635 24379
rect 28635 24345 28644 24379
rect 28592 24336 28644 24345
rect 30524 24404 30576 24456
rect 31352 24404 31404 24456
rect 31904 24404 31956 24456
rect 32364 24404 32416 24456
rect 28960 24268 29012 24320
rect 29788 24336 29840 24388
rect 30340 24336 30392 24388
rect 30708 24336 30760 24388
rect 29972 24268 30024 24320
rect 31168 24268 31220 24320
rect 25464 24200 25516 24252
rect 20404 24132 20456 24184
rect 23072 24132 23124 24184
rect 31812 24132 31864 24184
rect 14142 24030 14194 24082
rect 14206 24030 14258 24082
rect 14270 24030 14322 24082
rect 14334 24030 14386 24082
rect 24142 24030 24194 24082
rect 24206 24030 24258 24082
rect 24270 24030 24322 24082
rect 24334 24030 24386 24082
rect 13136 23928 13188 23980
rect 27948 23928 28000 23980
rect 16540 23860 16592 23912
rect 27304 23860 27356 23912
rect 30708 23903 30760 23912
rect 30708 23869 30717 23903
rect 30717 23869 30751 23903
rect 30751 23869 30760 23903
rect 30708 23860 30760 23869
rect 14608 23792 14660 23844
rect 14792 23724 14844 23776
rect 16724 23792 16776 23844
rect 18932 23792 18984 23844
rect 16080 23724 16132 23776
rect 18380 23724 18432 23776
rect 19024 23767 19076 23776
rect 19024 23733 19033 23767
rect 19033 23733 19067 23767
rect 19067 23733 19076 23767
rect 19024 23724 19076 23733
rect 19208 23792 19260 23844
rect 19576 23724 19628 23776
rect 19852 23724 19904 23776
rect 18012 23699 18064 23708
rect 18012 23665 18021 23699
rect 18021 23665 18055 23699
rect 18055 23665 18064 23699
rect 18012 23656 18064 23665
rect 19668 23656 19720 23708
rect 20128 23724 20180 23776
rect 21416 23724 21468 23776
rect 22980 23792 23032 23844
rect 23808 23792 23860 23844
rect 31812 23835 31864 23844
rect 31812 23801 31821 23835
rect 31821 23801 31855 23835
rect 31855 23801 31864 23835
rect 31812 23792 31864 23801
rect 22888 23767 22940 23776
rect 22888 23733 22897 23767
rect 22897 23733 22931 23767
rect 22931 23733 22940 23767
rect 22888 23724 22940 23733
rect 23992 23724 24044 23776
rect 24636 23767 24688 23776
rect 24636 23733 24645 23767
rect 24645 23733 24679 23767
rect 24679 23733 24688 23767
rect 24636 23724 24688 23733
rect 25004 23767 25056 23776
rect 25004 23733 25013 23767
rect 25013 23733 25047 23767
rect 25047 23733 25056 23767
rect 25004 23724 25056 23733
rect 26752 23724 26804 23776
rect 28868 23767 28920 23776
rect 28868 23733 28877 23767
rect 28877 23733 28911 23767
rect 28911 23733 28920 23767
rect 28868 23724 28920 23733
rect 23164 23656 23216 23708
rect 26292 23699 26344 23708
rect 26292 23665 26301 23699
rect 26301 23665 26335 23699
rect 26335 23665 26344 23699
rect 26292 23656 26344 23665
rect 28132 23656 28184 23708
rect 29788 23699 29840 23708
rect 23716 23631 23768 23640
rect 23716 23597 23725 23631
rect 23725 23597 23759 23631
rect 23759 23597 23768 23631
rect 23716 23588 23768 23597
rect 29788 23665 29797 23699
rect 29797 23665 29831 23699
rect 29831 23665 29840 23699
rect 29788 23656 29840 23665
rect 30248 23767 30300 23776
rect 30248 23733 30257 23767
rect 30257 23733 30291 23767
rect 30291 23733 30300 23767
rect 30248 23724 30300 23733
rect 19142 23486 19194 23538
rect 19206 23486 19258 23538
rect 19270 23486 19322 23538
rect 19334 23486 19386 23538
rect 29142 23486 29194 23538
rect 29206 23486 29258 23538
rect 29270 23486 29322 23538
rect 29334 23486 29386 23538
rect 16908 23427 16960 23436
rect 16908 23393 16917 23427
rect 16917 23393 16951 23427
rect 16951 23393 16960 23427
rect 16908 23384 16960 23393
rect 21048 23427 21100 23436
rect 21048 23393 21057 23427
rect 21057 23393 21091 23427
rect 21091 23393 21100 23427
rect 21048 23384 21100 23393
rect 21416 23384 21468 23436
rect 14700 23291 14752 23300
rect 14700 23257 14709 23291
rect 14709 23257 14743 23291
rect 14743 23257 14752 23291
rect 14700 23248 14752 23257
rect 14792 23291 14844 23300
rect 14792 23257 14801 23291
rect 14801 23257 14835 23291
rect 14835 23257 14844 23291
rect 15068 23291 15120 23300
rect 14792 23248 14844 23257
rect 15068 23257 15077 23291
rect 15077 23257 15111 23291
rect 15111 23257 15120 23291
rect 15068 23248 15120 23257
rect 15252 23248 15304 23300
rect 15436 23316 15488 23368
rect 18012 23316 18064 23368
rect 16724 23248 16776 23300
rect 17828 23291 17880 23300
rect 17828 23257 17837 23291
rect 17837 23257 17871 23291
rect 17871 23257 17880 23291
rect 17828 23248 17880 23257
rect 18380 23248 18432 23300
rect 13412 23180 13464 23232
rect 15528 23223 15580 23232
rect 15528 23189 15537 23223
rect 15537 23189 15571 23223
rect 15571 23189 15580 23223
rect 15528 23180 15580 23189
rect 15988 23180 16040 23232
rect 19208 23248 19260 23300
rect 19484 23316 19536 23368
rect 19760 23316 19812 23368
rect 20588 23316 20640 23368
rect 21968 23316 22020 23368
rect 22980 23384 23032 23436
rect 25464 23384 25516 23436
rect 28500 23384 28552 23436
rect 29788 23384 29840 23436
rect 22520 23316 22572 23368
rect 23072 23359 23124 23368
rect 23072 23325 23081 23359
rect 23081 23325 23115 23359
rect 23115 23325 23124 23359
rect 23072 23316 23124 23325
rect 25280 23316 25332 23368
rect 19576 23248 19628 23300
rect 20772 23291 20824 23300
rect 20772 23257 20781 23291
rect 20781 23257 20815 23291
rect 20815 23257 20824 23291
rect 20772 23248 20824 23257
rect 19484 23180 19536 23232
rect 23164 23248 23216 23300
rect 23900 23248 23952 23300
rect 27304 23291 27356 23300
rect 27304 23257 27313 23291
rect 27313 23257 27347 23291
rect 27347 23257 27356 23291
rect 27304 23248 27356 23257
rect 28040 23291 28092 23300
rect 28040 23257 28049 23291
rect 28049 23257 28083 23291
rect 28083 23257 28092 23291
rect 28040 23248 28092 23257
rect 28132 23248 28184 23300
rect 30892 23291 30944 23300
rect 30892 23257 30901 23291
rect 30901 23257 30935 23291
rect 30935 23257 30944 23291
rect 30892 23248 30944 23257
rect 21416 23180 21468 23232
rect 21508 23180 21560 23232
rect 22612 23180 22664 23232
rect 26108 23180 26160 23232
rect 27212 23180 27264 23232
rect 27396 23223 27448 23232
rect 27396 23189 27405 23223
rect 27405 23189 27439 23223
rect 27439 23189 27448 23223
rect 27396 23180 27448 23189
rect 27856 23180 27908 23232
rect 11940 23112 11992 23164
rect 19576 23112 19628 23164
rect 23992 23112 24044 23164
rect 18932 23044 18984 23096
rect 19484 23044 19536 23096
rect 23624 23044 23676 23096
rect 24912 23044 24964 23096
rect 25464 23087 25516 23096
rect 25464 23053 25473 23087
rect 25473 23053 25507 23087
rect 25507 23053 25516 23087
rect 25464 23044 25516 23053
rect 29604 23087 29656 23096
rect 29604 23053 29613 23087
rect 29613 23053 29647 23087
rect 29647 23053 29656 23087
rect 29604 23044 29656 23053
rect 14142 22942 14194 22994
rect 14206 22942 14258 22994
rect 14270 22942 14322 22994
rect 14334 22942 14386 22994
rect 24142 22942 24194 22994
rect 24206 22942 24258 22994
rect 24270 22942 24322 22994
rect 24334 22942 24386 22994
rect 13780 22840 13832 22892
rect 14700 22840 14752 22892
rect 19852 22883 19904 22892
rect 19852 22849 19861 22883
rect 19861 22849 19895 22883
rect 19895 22849 19904 22883
rect 19852 22840 19904 22849
rect 22336 22840 22388 22892
rect 22704 22840 22756 22892
rect 18472 22815 18524 22824
rect 18472 22781 18481 22815
rect 18481 22781 18515 22815
rect 18515 22781 18524 22815
rect 18472 22772 18524 22781
rect 13412 22747 13464 22756
rect 13412 22713 13421 22747
rect 13421 22713 13455 22747
rect 13455 22713 13464 22747
rect 13412 22704 13464 22713
rect 15436 22704 15488 22756
rect 16080 22704 16132 22756
rect 15620 22679 15672 22688
rect 15620 22645 15629 22679
rect 15629 22645 15663 22679
rect 15663 22645 15672 22679
rect 15620 22636 15672 22645
rect 15896 22636 15948 22688
rect 16632 22636 16684 22688
rect 18012 22636 18064 22688
rect 18380 22679 18432 22688
rect 18380 22645 18389 22679
rect 18389 22645 18423 22679
rect 18423 22645 18432 22679
rect 18380 22636 18432 22645
rect 20772 22704 20824 22756
rect 21508 22704 21560 22756
rect 23164 22704 23216 22756
rect 23992 22747 24044 22756
rect 23992 22713 24001 22747
rect 24001 22713 24035 22747
rect 24035 22713 24044 22747
rect 23992 22704 24044 22713
rect 25464 22704 25516 22756
rect 25924 22747 25976 22756
rect 25924 22713 25933 22747
rect 25933 22713 25967 22747
rect 25967 22713 25976 22747
rect 25924 22704 25976 22713
rect 14700 22568 14752 22620
rect 18840 22543 18892 22552
rect 18840 22509 18849 22543
rect 18849 22509 18883 22543
rect 18883 22509 18892 22543
rect 18840 22500 18892 22509
rect 19760 22679 19812 22688
rect 19760 22645 19769 22679
rect 19769 22645 19803 22679
rect 19803 22645 19812 22679
rect 19760 22636 19812 22645
rect 19944 22636 19996 22688
rect 21968 22636 22020 22688
rect 19484 22568 19536 22620
rect 21140 22568 21192 22620
rect 21416 22611 21468 22620
rect 21416 22577 21425 22611
rect 21425 22577 21459 22611
rect 21459 22577 21468 22611
rect 21416 22568 21468 22577
rect 22888 22636 22940 22688
rect 23348 22636 23400 22688
rect 23624 22679 23676 22688
rect 23624 22645 23633 22679
rect 23633 22645 23667 22679
rect 23667 22645 23676 22679
rect 23624 22636 23676 22645
rect 20128 22500 20180 22552
rect 20956 22500 21008 22552
rect 21508 22500 21560 22552
rect 22704 22611 22756 22620
rect 22704 22577 22713 22611
rect 22713 22577 22747 22611
rect 22747 22577 22756 22611
rect 22704 22568 22756 22577
rect 25096 22679 25148 22688
rect 25096 22645 25105 22679
rect 25105 22645 25139 22679
rect 25139 22645 25148 22679
rect 25096 22636 25148 22645
rect 24452 22568 24504 22620
rect 25004 22568 25056 22620
rect 27396 22704 27448 22756
rect 28776 22704 28828 22756
rect 26384 22636 26436 22688
rect 27212 22636 27264 22688
rect 30248 22679 30300 22688
rect 30248 22645 30257 22679
rect 30257 22645 30291 22679
rect 30291 22645 30300 22679
rect 30248 22636 30300 22645
rect 30892 22704 30944 22756
rect 31260 22704 31312 22756
rect 30800 22636 30852 22688
rect 26476 22611 26528 22620
rect 26476 22577 26485 22611
rect 26485 22577 26519 22611
rect 26519 22577 26528 22611
rect 26476 22568 26528 22577
rect 23808 22500 23860 22552
rect 19142 22398 19194 22450
rect 19206 22398 19258 22450
rect 19270 22398 19322 22450
rect 19334 22398 19386 22450
rect 29142 22398 29194 22450
rect 29206 22398 29258 22450
rect 29270 22398 29322 22450
rect 29334 22398 29386 22450
rect 17828 22296 17880 22348
rect 18380 22296 18432 22348
rect 20588 22296 20640 22348
rect 21416 22296 21468 22348
rect 21508 22339 21560 22348
rect 21508 22305 21517 22339
rect 21517 22305 21551 22339
rect 21551 22305 21560 22339
rect 21508 22296 21560 22305
rect 22704 22296 22756 22348
rect 25280 22296 25332 22348
rect 15620 22228 15672 22280
rect 19944 22271 19996 22280
rect 19944 22237 19953 22271
rect 19953 22237 19987 22271
rect 19987 22237 19996 22271
rect 19944 22228 19996 22237
rect 20128 22271 20180 22280
rect 20128 22237 20137 22271
rect 20137 22237 20171 22271
rect 20171 22237 20180 22271
rect 20128 22228 20180 22237
rect 21140 22228 21192 22280
rect 14792 22092 14844 22144
rect 15436 22092 15488 22144
rect 16172 22203 16224 22212
rect 16172 22169 16181 22203
rect 16181 22169 16215 22203
rect 16215 22169 16224 22203
rect 16172 22160 16224 22169
rect 16724 22160 16776 22212
rect 17920 22160 17972 22212
rect 15896 22092 15948 22144
rect 16080 22135 16132 22144
rect 16080 22101 16089 22135
rect 16089 22101 16123 22135
rect 16123 22101 16132 22135
rect 16080 22092 16132 22101
rect 18288 22092 18340 22144
rect 19024 22092 19076 22144
rect 22980 22228 23032 22280
rect 24636 22228 24688 22280
rect 20496 22135 20548 22144
rect 20496 22101 20505 22135
rect 20505 22101 20539 22135
rect 20539 22101 20548 22135
rect 20496 22092 20548 22101
rect 22244 22160 22296 22212
rect 22336 22160 22388 22212
rect 22888 22160 22940 22212
rect 23164 22092 23216 22144
rect 25464 22160 25516 22212
rect 26200 22160 26252 22212
rect 27764 22203 27816 22212
rect 27764 22169 27773 22203
rect 27773 22169 27807 22203
rect 27807 22169 27816 22203
rect 29512 22296 29564 22348
rect 27764 22160 27816 22169
rect 23992 22092 24044 22144
rect 27856 22135 27908 22144
rect 27856 22101 27865 22135
rect 27865 22101 27899 22135
rect 27899 22101 27908 22135
rect 27856 22092 27908 22101
rect 29512 22160 29564 22212
rect 30248 22203 30300 22212
rect 30248 22169 30257 22203
rect 30257 22169 30291 22203
rect 30291 22169 30300 22203
rect 30248 22160 30300 22169
rect 30800 22203 30852 22212
rect 30800 22169 30809 22203
rect 30809 22169 30843 22203
rect 30843 22169 30852 22203
rect 30800 22160 30852 22169
rect 31260 22203 31312 22212
rect 31260 22169 31269 22203
rect 31269 22169 31303 22203
rect 31303 22169 31312 22203
rect 31260 22160 31312 22169
rect 30064 22092 30116 22144
rect 22336 22024 22388 22076
rect 22428 22024 22480 22076
rect 29880 22024 29932 22076
rect 18012 21999 18064 22008
rect 18012 21965 18036 21999
rect 18036 21965 18064 21999
rect 18012 21956 18064 21965
rect 21968 21956 22020 22008
rect 29328 21956 29380 22008
rect 30248 21956 30300 22008
rect 14142 21854 14194 21906
rect 14206 21854 14258 21906
rect 14270 21854 14322 21906
rect 14334 21854 14386 21906
rect 24142 21854 24194 21906
rect 24206 21854 24258 21906
rect 24270 21854 24322 21906
rect 24334 21854 24386 21906
rect 14700 21752 14752 21804
rect 15896 21727 15948 21736
rect 15896 21693 15905 21727
rect 15905 21693 15939 21727
rect 15939 21693 15948 21727
rect 15896 21684 15948 21693
rect 14608 21548 14660 21600
rect 14884 21548 14936 21600
rect 16172 21616 16224 21668
rect 19760 21616 19812 21668
rect 22704 21752 22756 21804
rect 21416 21684 21468 21736
rect 22244 21684 22296 21736
rect 22980 21727 23032 21736
rect 22980 21693 22989 21727
rect 22989 21693 23023 21727
rect 23023 21693 23032 21727
rect 22980 21684 23032 21693
rect 15528 21548 15580 21600
rect 17460 21591 17512 21600
rect 17460 21557 17469 21591
rect 17469 21557 17503 21591
rect 17503 21557 17512 21591
rect 17460 21548 17512 21557
rect 17828 21548 17880 21600
rect 18104 21548 18156 21600
rect 18288 21591 18340 21600
rect 18288 21557 18297 21591
rect 18297 21557 18331 21591
rect 18331 21557 18340 21591
rect 18288 21548 18340 21557
rect 18840 21591 18892 21600
rect 16080 21480 16132 21532
rect 18840 21557 18849 21591
rect 18849 21557 18883 21591
rect 18883 21557 18892 21591
rect 18840 21548 18892 21557
rect 22336 21616 22388 21668
rect 28040 21752 28092 21804
rect 28868 21752 28920 21804
rect 27856 21684 27908 21736
rect 24452 21616 24504 21668
rect 28316 21616 28368 21668
rect 20496 21548 20548 21600
rect 21416 21591 21468 21600
rect 21416 21557 21425 21591
rect 21425 21557 21459 21591
rect 21459 21557 21468 21591
rect 21416 21548 21468 21557
rect 22152 21548 22204 21600
rect 22888 21591 22940 21600
rect 22888 21557 22897 21591
rect 22897 21557 22931 21591
rect 22931 21557 22940 21591
rect 22888 21548 22940 21557
rect 23164 21591 23216 21600
rect 23164 21557 23173 21591
rect 23173 21557 23207 21591
rect 23207 21557 23216 21591
rect 23164 21548 23216 21557
rect 23900 21548 23952 21600
rect 24636 21548 24688 21600
rect 25004 21591 25056 21600
rect 25004 21557 25013 21591
rect 25013 21557 25047 21591
rect 25047 21557 25056 21591
rect 25004 21548 25056 21557
rect 26200 21548 26252 21600
rect 27764 21548 27816 21600
rect 29328 21548 29380 21600
rect 29604 21548 29656 21600
rect 29880 21591 29932 21600
rect 26108 21480 26160 21532
rect 28500 21480 28552 21532
rect 29512 21480 29564 21532
rect 29880 21557 29889 21591
rect 29889 21557 29923 21591
rect 29923 21557 29932 21591
rect 29880 21548 29932 21557
rect 31996 21684 32048 21736
rect 32180 21616 32232 21668
rect 31168 21591 31220 21600
rect 31168 21557 31177 21591
rect 31177 21557 31211 21591
rect 31211 21557 31220 21591
rect 31168 21548 31220 21557
rect 31996 21591 32048 21600
rect 31996 21557 32005 21591
rect 32005 21557 32039 21591
rect 32039 21557 32048 21591
rect 31996 21548 32048 21557
rect 32088 21591 32140 21600
rect 32088 21557 32097 21591
rect 32097 21557 32131 21591
rect 32131 21557 32140 21591
rect 32088 21548 32140 21557
rect 17276 21455 17328 21464
rect 17276 21421 17285 21455
rect 17285 21421 17319 21455
rect 17319 21421 17328 21455
rect 17276 21412 17328 21421
rect 19576 21412 19628 21464
rect 21416 21412 21468 21464
rect 24636 21412 24688 21464
rect 27948 21455 28000 21464
rect 27948 21421 27957 21455
rect 27957 21421 27991 21455
rect 27991 21421 28000 21455
rect 27948 21412 28000 21421
rect 30156 21412 30208 21464
rect 19142 21310 19194 21362
rect 19206 21310 19258 21362
rect 19270 21310 19322 21362
rect 19334 21310 19386 21362
rect 29142 21310 29194 21362
rect 29206 21310 29258 21362
rect 29270 21310 29322 21362
rect 29334 21310 29386 21362
rect 20496 21208 20548 21260
rect 17828 21140 17880 21192
rect 18012 21183 18064 21192
rect 18012 21149 18021 21183
rect 18021 21149 18055 21183
rect 18055 21149 18064 21183
rect 18012 21140 18064 21149
rect 18104 21140 18156 21192
rect 19576 21183 19628 21192
rect 19576 21149 19585 21183
rect 19585 21149 19619 21183
rect 19619 21149 19628 21183
rect 19576 21140 19628 21149
rect 22612 21208 22664 21260
rect 28500 21208 28552 21260
rect 16172 21115 16224 21124
rect 16172 21081 16181 21115
rect 16181 21081 16215 21115
rect 16215 21081 16224 21115
rect 16172 21072 16224 21081
rect 15988 21004 16040 21056
rect 16080 21004 16132 21056
rect 16448 21072 16500 21124
rect 17920 21072 17972 21124
rect 19760 21115 19812 21124
rect 19760 21081 19769 21115
rect 19769 21081 19803 21115
rect 19803 21081 19812 21115
rect 19760 21072 19812 21081
rect 21048 21072 21100 21124
rect 18012 21004 18064 21056
rect 18380 21004 18432 21056
rect 21600 21047 21652 21056
rect 21600 21013 21609 21047
rect 21609 21013 21643 21047
rect 21643 21013 21652 21047
rect 21600 21004 21652 21013
rect 21416 20936 21468 20988
rect 22152 21072 22204 21124
rect 22428 21140 22480 21192
rect 27764 21140 27816 21192
rect 27856 21140 27908 21192
rect 30156 21183 30208 21192
rect 30156 21149 30165 21183
rect 30165 21149 30199 21183
rect 30199 21149 30208 21183
rect 30156 21140 30208 21149
rect 23348 21072 23400 21124
rect 23808 21115 23860 21124
rect 23808 21081 23817 21115
rect 23817 21081 23851 21115
rect 23851 21081 23860 21115
rect 23808 21072 23860 21081
rect 26844 21072 26896 21124
rect 27304 21115 27356 21124
rect 27304 21081 27313 21115
rect 27313 21081 27347 21115
rect 27347 21081 27356 21115
rect 27304 21072 27356 21081
rect 29512 21072 29564 21124
rect 30064 21115 30116 21124
rect 30064 21081 30073 21115
rect 30073 21081 30107 21115
rect 30107 21081 30116 21115
rect 30064 21072 30116 21081
rect 25188 21047 25240 21056
rect 25188 21013 25197 21047
rect 25197 21013 25231 21047
rect 25231 21013 25240 21047
rect 25188 21004 25240 21013
rect 25280 21004 25332 21056
rect 25648 20979 25700 20988
rect 25648 20945 25657 20979
rect 25657 20945 25691 20979
rect 25691 20945 25700 20979
rect 25648 20936 25700 20945
rect 15344 20868 15396 20920
rect 15620 20868 15672 20920
rect 17460 20868 17512 20920
rect 23992 20911 24044 20920
rect 23992 20877 24001 20911
rect 24001 20877 24035 20911
rect 24035 20877 24044 20911
rect 23992 20868 24044 20877
rect 26384 20868 26436 20920
rect 14142 20766 14194 20818
rect 14206 20766 14258 20818
rect 14270 20766 14322 20818
rect 14334 20766 14386 20818
rect 24142 20766 24194 20818
rect 24206 20766 24258 20818
rect 24270 20766 24322 20818
rect 24334 20766 24386 20818
rect 22152 20664 22204 20716
rect 14976 20503 15028 20512
rect 14976 20469 14985 20503
rect 14985 20469 15019 20503
rect 15019 20469 15028 20503
rect 14976 20460 15028 20469
rect 15528 20528 15580 20580
rect 15988 20528 16040 20580
rect 18012 20596 18064 20648
rect 24636 20596 24688 20648
rect 27304 20639 27356 20648
rect 15252 20460 15304 20512
rect 14240 20392 14292 20444
rect 15620 20460 15672 20512
rect 21416 20528 21468 20580
rect 23716 20528 23768 20580
rect 18012 20503 18064 20512
rect 18012 20469 18021 20503
rect 18021 20469 18055 20503
rect 18055 20469 18064 20503
rect 18012 20460 18064 20469
rect 21140 20503 21192 20512
rect 21140 20469 21149 20503
rect 21149 20469 21183 20503
rect 21183 20469 21192 20503
rect 21140 20460 21192 20469
rect 21600 20460 21652 20512
rect 23992 20503 24044 20512
rect 23992 20469 24001 20503
rect 24001 20469 24035 20503
rect 24035 20469 24044 20503
rect 23992 20460 24044 20469
rect 24728 20528 24780 20580
rect 27304 20605 27313 20639
rect 27313 20605 27347 20639
rect 27347 20605 27356 20639
rect 27304 20596 27356 20605
rect 30248 20596 30300 20648
rect 25004 20528 25056 20580
rect 26844 20571 26896 20580
rect 26844 20537 26853 20571
rect 26853 20537 26887 20571
rect 26887 20537 26896 20571
rect 26844 20528 26896 20537
rect 27948 20528 28000 20580
rect 24912 20503 24964 20512
rect 24912 20469 24921 20503
rect 24921 20469 24955 20503
rect 24955 20469 24964 20503
rect 24912 20460 24964 20469
rect 26384 20503 26436 20512
rect 17276 20392 17328 20444
rect 18288 20435 18340 20444
rect 18288 20401 18297 20435
rect 18297 20401 18331 20435
rect 18331 20401 18340 20435
rect 18288 20392 18340 20401
rect 19944 20392 19996 20444
rect 19024 20324 19076 20376
rect 21416 20392 21468 20444
rect 25188 20392 25240 20444
rect 26384 20469 26393 20503
rect 26393 20469 26427 20503
rect 26427 20469 26436 20503
rect 26384 20460 26436 20469
rect 25648 20392 25700 20444
rect 29604 20392 29656 20444
rect 23992 20324 24044 20376
rect 19142 20222 19194 20274
rect 19206 20222 19258 20274
rect 19270 20222 19322 20274
rect 19334 20222 19386 20274
rect 29142 20222 29194 20274
rect 29206 20222 29258 20274
rect 29270 20222 29322 20274
rect 29334 20222 29386 20274
rect 14976 20120 15028 20172
rect 25280 20120 25332 20172
rect 14240 20095 14292 20104
rect 14240 20061 14249 20095
rect 14249 20061 14283 20095
rect 14283 20061 14292 20095
rect 14240 20052 14292 20061
rect 14516 20052 14568 20104
rect 15988 20095 16040 20104
rect 15988 20061 15997 20095
rect 15997 20061 16031 20095
rect 16031 20061 16040 20095
rect 15988 20052 16040 20061
rect 13780 19984 13832 20036
rect 15344 19848 15396 19900
rect 16540 19984 16592 20036
rect 19024 20052 19076 20104
rect 17276 19984 17328 20036
rect 18564 20027 18616 20036
rect 18564 19993 18573 20027
rect 18573 19993 18607 20027
rect 18607 19993 18616 20027
rect 18564 19984 18616 19993
rect 21416 20027 21468 20036
rect 21416 19993 21425 20027
rect 21425 19993 21459 20027
rect 21459 19993 21468 20027
rect 21416 19984 21468 19993
rect 22152 20027 22204 20036
rect 22152 19993 22161 20027
rect 22161 19993 22195 20027
rect 22195 19993 22204 20027
rect 22152 19984 22204 19993
rect 23900 19984 23952 20036
rect 27764 20052 27816 20104
rect 25096 19984 25148 20036
rect 26384 20027 26436 20036
rect 26384 19993 26393 20027
rect 26393 19993 26427 20027
rect 26427 19993 26436 20027
rect 26384 19984 26436 19993
rect 27304 20027 27356 20036
rect 27304 19993 27313 20027
rect 27313 19993 27347 20027
rect 27347 19993 27356 20027
rect 27304 19984 27356 19993
rect 29604 20027 29656 20036
rect 17920 19916 17972 19968
rect 29604 19993 29613 20027
rect 29613 19993 29647 20027
rect 29647 19993 29656 20027
rect 29604 19984 29656 19993
rect 18288 19848 18340 19900
rect 27948 19848 28000 19900
rect 28500 19891 28552 19900
rect 28500 19857 28509 19891
rect 28509 19857 28543 19891
rect 28543 19857 28552 19891
rect 28500 19848 28552 19857
rect 23256 19823 23308 19832
rect 23256 19789 23265 19823
rect 23265 19789 23299 19823
rect 23299 19789 23308 19823
rect 23256 19780 23308 19789
rect 29696 19823 29748 19832
rect 29696 19789 29705 19823
rect 29705 19789 29739 19823
rect 29739 19789 29748 19823
rect 29696 19780 29748 19789
rect 14142 19678 14194 19730
rect 14206 19678 14258 19730
rect 14270 19678 14322 19730
rect 14334 19678 14386 19730
rect 24142 19678 24194 19730
rect 24206 19678 24258 19730
rect 24270 19678 24322 19730
rect 24334 19678 24386 19730
rect 14516 19619 14568 19628
rect 14516 19585 14525 19619
rect 14525 19585 14559 19619
rect 14559 19585 14568 19619
rect 14516 19576 14568 19585
rect 17920 19619 17972 19628
rect 17920 19585 17929 19619
rect 17929 19585 17963 19619
rect 17963 19585 17972 19619
rect 17920 19576 17972 19585
rect 18564 19576 18616 19628
rect 19944 19576 19996 19628
rect 29604 19508 29656 19560
rect 15528 19483 15580 19492
rect 15528 19449 15537 19483
rect 15537 19449 15571 19483
rect 15571 19449 15580 19483
rect 15528 19440 15580 19449
rect 14608 19372 14660 19424
rect 15344 19415 15396 19424
rect 15344 19381 15353 19415
rect 15353 19381 15387 19415
rect 15387 19381 15396 19415
rect 15344 19372 15396 19381
rect 16540 19372 16592 19424
rect 19024 19415 19076 19424
rect 19024 19381 19033 19415
rect 19033 19381 19067 19415
rect 19067 19381 19076 19415
rect 19024 19372 19076 19381
rect 19576 19372 19628 19424
rect 22244 19372 22296 19424
rect 22520 19415 22572 19424
rect 22520 19381 22529 19415
rect 22529 19381 22563 19415
rect 22563 19381 22572 19415
rect 22520 19372 22572 19381
rect 23256 19415 23308 19424
rect 23256 19381 23265 19415
rect 23265 19381 23299 19415
rect 23299 19381 23308 19415
rect 23256 19372 23308 19381
rect 25096 19372 25148 19424
rect 27948 19415 28000 19424
rect 27948 19381 27957 19415
rect 27957 19381 27991 19415
rect 27991 19381 28000 19415
rect 27948 19372 28000 19381
rect 19760 19304 19812 19356
rect 25648 19304 25700 19356
rect 27764 19304 27816 19356
rect 29696 19372 29748 19424
rect 23348 19236 23400 19288
rect 23624 19236 23676 19288
rect 19142 19134 19194 19186
rect 19206 19134 19258 19186
rect 19270 19134 19322 19186
rect 19334 19134 19386 19186
rect 29142 19134 29194 19186
rect 29206 19134 29258 19186
rect 29270 19134 29322 19186
rect 29334 19134 29386 19186
rect 18012 18964 18064 19016
rect 18380 18896 18432 18948
rect 19760 18964 19812 19016
rect 23624 19032 23676 19084
rect 21784 18964 21836 19016
rect 22520 18964 22572 19016
rect 27212 19032 27264 19084
rect 20956 18828 21008 18880
rect 21508 18828 21560 18880
rect 22244 18828 22296 18880
rect 23072 18939 23124 18948
rect 23072 18905 23081 18939
rect 23081 18905 23115 18939
rect 23115 18905 23124 18939
rect 23072 18896 23124 18905
rect 27304 18964 27356 19016
rect 28500 19032 28552 19084
rect 23900 18939 23952 18948
rect 23900 18905 23909 18939
rect 23909 18905 23943 18939
rect 23943 18905 23952 18939
rect 23900 18896 23952 18905
rect 23992 18896 24044 18948
rect 26292 18896 26344 18948
rect 26476 18828 26528 18880
rect 28040 18896 28092 18948
rect 28776 18896 28828 18948
rect 30708 18828 30760 18880
rect 18288 18760 18340 18812
rect 24452 18692 24504 18744
rect 29512 18735 29564 18744
rect 29512 18701 29521 18735
rect 29521 18701 29555 18735
rect 29555 18701 29564 18735
rect 29512 18692 29564 18701
rect 14142 18590 14194 18642
rect 14206 18590 14258 18642
rect 14270 18590 14322 18642
rect 14334 18590 14386 18642
rect 24142 18590 24194 18642
rect 24206 18590 24258 18642
rect 24270 18590 24322 18642
rect 24334 18590 24386 18642
rect 13780 18488 13832 18540
rect 18012 18488 18064 18540
rect 20956 18488 21008 18540
rect 21784 18463 21836 18472
rect 18380 18352 18432 18404
rect 14608 18284 14660 18336
rect 15988 18284 16040 18336
rect 16908 18216 16960 18268
rect 18012 18259 18064 18268
rect 18012 18225 18021 18259
rect 18021 18225 18055 18259
rect 18055 18225 18064 18259
rect 18012 18216 18064 18225
rect 19668 18216 19720 18268
rect 19852 18216 19904 18268
rect 21784 18429 21793 18463
rect 21793 18429 21827 18463
rect 21827 18429 21836 18463
rect 21784 18420 21836 18429
rect 21876 18420 21928 18472
rect 29604 18420 29656 18472
rect 20864 18352 20916 18404
rect 23348 18395 23400 18404
rect 21508 18284 21560 18336
rect 23348 18361 23357 18395
rect 23357 18361 23391 18395
rect 23391 18361 23400 18395
rect 23348 18352 23400 18361
rect 23900 18352 23952 18404
rect 27304 18352 27356 18404
rect 29512 18352 29564 18404
rect 21876 18284 21928 18336
rect 22520 18284 22572 18336
rect 24452 18284 24504 18336
rect 26476 18327 26528 18336
rect 26476 18293 26485 18327
rect 26485 18293 26519 18327
rect 26519 18293 26528 18327
rect 26476 18284 26528 18293
rect 27212 18327 27264 18336
rect 27212 18293 27221 18327
rect 27221 18293 27255 18327
rect 27255 18293 27264 18327
rect 27212 18284 27264 18293
rect 27764 18284 27816 18336
rect 23624 18216 23676 18268
rect 14700 18148 14752 18200
rect 15620 18191 15672 18200
rect 15620 18157 15629 18191
rect 15629 18157 15663 18191
rect 15663 18157 15672 18191
rect 15620 18148 15672 18157
rect 19576 18148 19628 18200
rect 20864 18148 20916 18200
rect 23992 18148 24044 18200
rect 19142 18046 19194 18098
rect 19206 18046 19258 18098
rect 19270 18046 19322 18098
rect 19334 18046 19386 18098
rect 29142 18046 29194 18098
rect 29206 18046 29258 18098
rect 29270 18046 29322 18098
rect 29334 18046 29386 18098
rect 19668 17944 19720 17996
rect 28040 17944 28092 17996
rect 14700 17876 14752 17928
rect 15988 17919 16040 17928
rect 15988 17885 15997 17919
rect 15997 17885 16031 17919
rect 16031 17885 16040 17919
rect 15988 17876 16040 17885
rect 13780 17808 13832 17860
rect 18380 17851 18432 17860
rect 18380 17817 18389 17851
rect 18389 17817 18423 17851
rect 18423 17817 18432 17851
rect 18380 17808 18432 17817
rect 19576 17876 19628 17928
rect 20864 17876 20916 17928
rect 19852 17851 19904 17860
rect 19852 17817 19861 17851
rect 19861 17817 19895 17851
rect 19895 17817 19904 17851
rect 19852 17808 19904 17817
rect 26476 17876 26528 17928
rect 22428 17808 22480 17860
rect 23256 17851 23308 17860
rect 23256 17817 23265 17851
rect 23265 17817 23299 17851
rect 23299 17817 23308 17851
rect 23256 17808 23308 17817
rect 23992 17808 24044 17860
rect 28408 17876 28460 17928
rect 17920 17740 17972 17792
rect 18748 17740 18800 17792
rect 22336 17783 22388 17792
rect 22336 17749 22345 17783
rect 22345 17749 22379 17783
rect 22379 17749 22388 17783
rect 22336 17740 22388 17749
rect 25004 17740 25056 17792
rect 27764 17808 27816 17860
rect 28960 17740 29012 17792
rect 23808 17604 23860 17656
rect 24544 17604 24596 17656
rect 14142 17502 14194 17554
rect 14206 17502 14258 17554
rect 14270 17502 14322 17554
rect 14334 17502 14386 17554
rect 24142 17502 24194 17554
rect 24206 17502 24258 17554
rect 24270 17502 24322 17554
rect 24334 17502 24386 17554
rect 15344 17400 15396 17452
rect 17368 17400 17420 17452
rect 18012 17400 18064 17452
rect 22336 17400 22388 17452
rect 23072 17400 23124 17452
rect 12400 17332 12452 17384
rect 20772 17332 20824 17384
rect 12676 17264 12728 17316
rect 12400 17196 12452 17248
rect 21232 17264 21284 17316
rect 23256 17264 23308 17316
rect 23532 17307 23584 17316
rect 23532 17273 23541 17307
rect 23541 17273 23575 17307
rect 23575 17273 23584 17307
rect 23532 17264 23584 17273
rect 23808 17307 23860 17316
rect 23808 17273 23817 17307
rect 23817 17273 23851 17307
rect 23851 17273 23860 17307
rect 23808 17264 23860 17273
rect 12492 17171 12544 17180
rect 12492 17137 12501 17171
rect 12501 17137 12535 17171
rect 12535 17137 12544 17171
rect 12492 17128 12544 17137
rect 15344 17196 15396 17248
rect 16724 17196 16776 17248
rect 17368 17239 17420 17248
rect 17368 17205 17377 17239
rect 17377 17205 17411 17239
rect 17411 17205 17420 17239
rect 17368 17196 17420 17205
rect 17920 17239 17972 17248
rect 17920 17205 17929 17239
rect 17929 17205 17963 17239
rect 17963 17205 17972 17239
rect 17920 17196 17972 17205
rect 15620 17060 15672 17112
rect 18196 17128 18248 17180
rect 19484 17196 19536 17248
rect 19024 17128 19076 17180
rect 19668 17171 19720 17180
rect 19668 17137 19677 17171
rect 19677 17137 19711 17171
rect 19711 17137 19720 17171
rect 19668 17128 19720 17137
rect 24544 17128 24596 17180
rect 28960 17060 29012 17112
rect 30616 17060 30668 17112
rect 19142 16958 19194 17010
rect 19206 16958 19258 17010
rect 19270 16958 19322 17010
rect 19334 16958 19386 17010
rect 29142 16958 29194 17010
rect 29206 16958 29258 17010
rect 29270 16958 29322 17010
rect 29334 16958 29386 17010
rect 12676 16788 12728 16840
rect 16724 16831 16776 16840
rect 12400 16763 12452 16772
rect 12400 16729 12409 16763
rect 12409 16729 12443 16763
rect 12443 16729 12452 16763
rect 12400 16720 12452 16729
rect 15620 16763 15672 16772
rect 15620 16729 15629 16763
rect 15629 16729 15663 16763
rect 15663 16729 15672 16763
rect 16724 16797 16733 16831
rect 16733 16797 16767 16831
rect 16767 16797 16776 16831
rect 16724 16788 16776 16797
rect 15620 16720 15672 16729
rect 17920 16720 17972 16772
rect 18196 16763 18248 16772
rect 18196 16729 18205 16763
rect 18205 16729 18239 16763
rect 18239 16729 18248 16763
rect 18196 16720 18248 16729
rect 18748 16788 18800 16840
rect 19668 16788 19720 16840
rect 18472 16720 18524 16772
rect 12768 16652 12820 16704
rect 20772 16720 20824 16772
rect 18380 16584 18432 16636
rect 22428 16720 22480 16772
rect 23992 16720 24044 16772
rect 22152 16695 22204 16704
rect 22152 16661 22161 16695
rect 22161 16661 22195 16695
rect 22195 16661 22204 16695
rect 22152 16652 22204 16661
rect 22336 16584 22388 16636
rect 13964 16516 14016 16568
rect 21048 16516 21100 16568
rect 21324 16559 21376 16568
rect 21324 16525 21333 16559
rect 21333 16525 21367 16559
rect 21367 16525 21376 16559
rect 21324 16516 21376 16525
rect 23532 16516 23584 16568
rect 24544 16516 24596 16568
rect 14142 16414 14194 16466
rect 14206 16414 14258 16466
rect 14270 16414 14322 16466
rect 14334 16414 14386 16466
rect 24142 16414 24194 16466
rect 24206 16414 24258 16466
rect 24270 16414 24322 16466
rect 24334 16414 24386 16466
rect 22152 16312 22204 16364
rect 12492 16176 12544 16228
rect 15344 16219 15396 16228
rect 15344 16185 15353 16219
rect 15353 16185 15387 16219
rect 15387 16185 15396 16219
rect 15344 16176 15396 16185
rect 18196 16244 18248 16296
rect 20772 16244 20824 16296
rect 18932 16219 18984 16228
rect 18932 16185 18941 16219
rect 18941 16185 18975 16219
rect 18975 16185 18984 16219
rect 18932 16176 18984 16185
rect 21324 16219 21376 16228
rect 21324 16185 21333 16219
rect 21333 16185 21367 16219
rect 21367 16185 21376 16219
rect 21324 16176 21376 16185
rect 23256 16219 23308 16228
rect 23256 16185 23265 16219
rect 23265 16185 23299 16219
rect 23299 16185 23308 16219
rect 23256 16176 23308 16185
rect 23532 16219 23584 16228
rect 23532 16185 23541 16219
rect 23541 16185 23575 16219
rect 23575 16185 23584 16219
rect 23532 16176 23584 16185
rect 12400 16151 12452 16160
rect 12400 16117 12409 16151
rect 12409 16117 12443 16151
rect 12443 16117 12452 16151
rect 12400 16108 12452 16117
rect 12676 16151 12728 16160
rect 12676 16117 12685 16151
rect 12685 16117 12719 16151
rect 12719 16117 12728 16151
rect 15620 16151 15672 16160
rect 12676 16108 12728 16117
rect 15620 16117 15629 16151
rect 15629 16117 15663 16151
rect 15663 16117 15672 16151
rect 15620 16108 15672 16117
rect 14792 16083 14844 16092
rect 14792 16049 14801 16083
rect 14801 16049 14835 16083
rect 14835 16049 14844 16083
rect 14792 16040 14844 16049
rect 14516 15972 14568 16024
rect 17920 16108 17972 16160
rect 18196 16151 18248 16160
rect 18196 16117 18205 16151
rect 18205 16117 18239 16151
rect 18239 16117 18248 16151
rect 18196 16108 18248 16117
rect 19024 16151 19076 16160
rect 19024 16117 19033 16151
rect 19033 16117 19067 16151
rect 19067 16117 19076 16151
rect 19024 16108 19076 16117
rect 19576 16108 19628 16160
rect 21232 16151 21284 16160
rect 21232 16117 21241 16151
rect 21241 16117 21275 16151
rect 21275 16117 21284 16151
rect 21232 16108 21284 16117
rect 17460 16040 17512 16092
rect 19852 16040 19904 16092
rect 18472 15972 18524 16024
rect 18840 15972 18892 16024
rect 20128 16015 20180 16024
rect 20128 15981 20137 16015
rect 20137 15981 20171 16015
rect 20171 15981 20180 16015
rect 20128 15972 20180 15981
rect 20680 16015 20732 16024
rect 20680 15981 20689 16015
rect 20689 15981 20723 16015
rect 20723 15981 20732 16015
rect 20680 15972 20732 15981
rect 22336 16040 22388 16092
rect 24544 16040 24596 16092
rect 22244 15972 22296 16024
rect 19142 15870 19194 15922
rect 19206 15870 19258 15922
rect 19270 15870 19322 15922
rect 19334 15870 19386 15922
rect 29142 15870 29194 15922
rect 29206 15870 29258 15922
rect 29270 15870 29322 15922
rect 29334 15870 29386 15922
rect 18748 15768 18800 15820
rect 22428 15768 22480 15820
rect 12492 15632 12544 15684
rect 12768 15675 12820 15684
rect 12768 15641 12777 15675
rect 12777 15641 12811 15675
rect 12811 15641 12820 15675
rect 12768 15632 12820 15641
rect 12952 15675 13004 15684
rect 12952 15641 12961 15675
rect 12961 15641 12995 15675
rect 12995 15641 13004 15675
rect 12952 15632 13004 15641
rect 13780 15632 13832 15684
rect 12768 15539 12820 15548
rect 12768 15505 12777 15539
rect 12777 15505 12811 15539
rect 12811 15505 12820 15539
rect 12768 15496 12820 15505
rect 15712 15632 15764 15684
rect 15988 15564 16040 15616
rect 17368 15632 17420 15684
rect 18932 15700 18984 15752
rect 20128 15700 20180 15752
rect 22244 15700 22296 15752
rect 18472 15675 18524 15684
rect 18472 15641 18481 15675
rect 18481 15641 18515 15675
rect 18515 15641 18524 15675
rect 18472 15632 18524 15641
rect 18564 15675 18616 15684
rect 18564 15641 18573 15675
rect 18573 15641 18607 15675
rect 18607 15641 18616 15675
rect 18564 15632 18616 15641
rect 21416 15632 21468 15684
rect 15620 15496 15672 15548
rect 18380 15564 18432 15616
rect 19576 15607 19628 15616
rect 19576 15573 19585 15607
rect 19585 15573 19619 15607
rect 19619 15573 19628 15607
rect 21600 15607 21652 15616
rect 19576 15564 19628 15573
rect 21600 15573 21609 15607
rect 21609 15573 21643 15607
rect 21643 15573 21652 15607
rect 21600 15564 21652 15573
rect 16724 15428 16776 15480
rect 19668 15428 19720 15480
rect 23992 15471 24044 15480
rect 23992 15437 24001 15471
rect 24001 15437 24035 15471
rect 24035 15437 24044 15471
rect 23992 15428 24044 15437
rect 14142 15326 14194 15378
rect 14206 15326 14258 15378
rect 14270 15326 14322 15378
rect 14334 15326 14386 15378
rect 24142 15326 24194 15378
rect 24206 15326 24258 15378
rect 24270 15326 24322 15378
rect 24334 15326 24386 15378
rect 15988 15267 16040 15276
rect 12400 15088 12452 15140
rect 15620 15156 15672 15208
rect 15988 15233 15997 15267
rect 15997 15233 16031 15267
rect 16031 15233 16040 15267
rect 15988 15224 16040 15233
rect 20772 15224 20824 15276
rect 18288 15156 18340 15208
rect 18564 15156 18616 15208
rect 13044 15063 13096 15072
rect 13044 15029 13053 15063
rect 13053 15029 13087 15063
rect 13087 15029 13096 15063
rect 13044 15020 13096 15029
rect 13412 15063 13464 15072
rect 13412 15029 13421 15063
rect 13421 15029 13455 15063
rect 13455 15029 13464 15063
rect 13412 15020 13464 15029
rect 13504 15020 13556 15072
rect 15068 15020 15120 15072
rect 18472 15088 18524 15140
rect 19668 15088 19720 15140
rect 18840 15063 18892 15072
rect 17460 14995 17512 15004
rect 17460 14961 17469 14995
rect 17469 14961 17503 14995
rect 17503 14961 17512 14995
rect 17460 14952 17512 14961
rect 15896 14884 15948 14936
rect 16908 14884 16960 14936
rect 18840 15029 18849 15063
rect 18849 15029 18883 15063
rect 18883 15029 18892 15063
rect 18840 15020 18892 15029
rect 19484 15020 19536 15072
rect 21600 15156 21652 15208
rect 22336 15131 22388 15140
rect 22336 15097 22345 15131
rect 22345 15097 22379 15131
rect 22379 15097 22388 15131
rect 22336 15088 22388 15097
rect 22152 15020 22204 15072
rect 24544 15020 24596 15072
rect 24452 14952 24504 15004
rect 18104 14927 18156 14936
rect 18104 14893 18113 14927
rect 18113 14893 18147 14927
rect 18147 14893 18156 14927
rect 18104 14884 18156 14893
rect 23900 14927 23952 14936
rect 23900 14893 23909 14927
rect 23909 14893 23943 14927
rect 23943 14893 23952 14927
rect 23900 14884 23952 14893
rect 19142 14782 19194 14834
rect 19206 14782 19258 14834
rect 19270 14782 19322 14834
rect 19334 14782 19386 14834
rect 29142 14782 29194 14834
rect 29206 14782 29258 14834
rect 29270 14782 29322 14834
rect 29334 14782 29386 14834
rect 12860 14680 12912 14732
rect 14792 14680 14844 14732
rect 15712 14723 15764 14732
rect 15712 14689 15721 14723
rect 15721 14689 15755 14723
rect 15755 14689 15764 14723
rect 15712 14680 15764 14689
rect 15896 14680 15948 14732
rect 21416 14723 21468 14732
rect 13044 14655 13096 14664
rect 13044 14621 13053 14655
rect 13053 14621 13087 14655
rect 13087 14621 13096 14655
rect 13044 14612 13096 14621
rect 12768 14587 12820 14596
rect 12768 14553 12777 14587
rect 12777 14553 12811 14587
rect 12811 14553 12820 14587
rect 12768 14544 12820 14553
rect 13412 14544 13464 14596
rect 14516 14544 14568 14596
rect 16908 14612 16960 14664
rect 21416 14689 21425 14723
rect 21425 14689 21459 14723
rect 21459 14689 21468 14723
rect 21416 14680 21468 14689
rect 23992 14612 24044 14664
rect 16724 14587 16776 14596
rect 16724 14553 16733 14587
rect 16733 14553 16767 14587
rect 16767 14553 16776 14587
rect 16724 14544 16776 14553
rect 18104 14544 18156 14596
rect 18472 14544 18524 14596
rect 21324 14587 21376 14596
rect 21324 14553 21333 14587
rect 21333 14553 21367 14587
rect 21367 14553 21376 14587
rect 21324 14544 21376 14553
rect 21600 14544 21652 14596
rect 22152 14587 22204 14596
rect 22152 14553 22161 14587
rect 22161 14553 22195 14587
rect 22195 14553 22204 14587
rect 22152 14544 22204 14553
rect 23808 14587 23860 14596
rect 23808 14553 23817 14587
rect 23817 14553 23851 14587
rect 23851 14553 23860 14587
rect 23808 14544 23860 14553
rect 23900 14587 23952 14596
rect 23900 14553 23909 14587
rect 23909 14553 23943 14587
rect 23943 14553 23952 14587
rect 23900 14544 23952 14553
rect 25372 14587 25424 14596
rect 12032 14519 12084 14528
rect 12032 14485 12041 14519
rect 12041 14485 12075 14519
rect 12075 14485 12084 14519
rect 12032 14476 12084 14485
rect 17000 14519 17052 14528
rect 14792 14451 14844 14460
rect 14792 14417 14801 14451
rect 14801 14417 14835 14451
rect 14835 14417 14844 14451
rect 14792 14408 14844 14417
rect 17000 14485 17009 14519
rect 17009 14485 17043 14519
rect 17043 14485 17052 14519
rect 17000 14476 17052 14485
rect 25372 14553 25381 14587
rect 25381 14553 25415 14587
rect 25415 14553 25424 14587
rect 25372 14544 25424 14553
rect 23256 14340 23308 14392
rect 23900 14340 23952 14392
rect 14142 14238 14194 14290
rect 14206 14238 14258 14290
rect 14270 14238 14322 14290
rect 14334 14238 14386 14290
rect 24142 14238 24194 14290
rect 24206 14238 24258 14290
rect 24270 14238 24322 14290
rect 24334 14238 24386 14290
rect 12032 14179 12084 14188
rect 12032 14145 12041 14179
rect 12041 14145 12075 14179
rect 12075 14145 12084 14179
rect 12032 14136 12084 14145
rect 12952 14136 13004 14188
rect 17000 14136 17052 14188
rect 14700 14068 14752 14120
rect 16172 14000 16224 14052
rect 17460 14000 17512 14052
rect 10468 13932 10520 13984
rect 12860 13975 12912 13984
rect 12860 13941 12869 13975
rect 12869 13941 12903 13975
rect 12903 13941 12912 13975
rect 12860 13932 12912 13941
rect 14792 13932 14844 13984
rect 18196 14000 18248 14052
rect 19484 14043 19536 14052
rect 17828 13932 17880 13984
rect 18288 13975 18340 13984
rect 13504 13864 13556 13916
rect 18288 13941 18297 13975
rect 18297 13941 18331 13975
rect 18331 13941 18340 13975
rect 18288 13932 18340 13941
rect 18932 13975 18984 13984
rect 18932 13941 18941 13975
rect 18941 13941 18975 13975
rect 18975 13941 18984 13975
rect 18932 13932 18984 13941
rect 19484 14009 19493 14043
rect 19493 14009 19527 14043
rect 19527 14009 19536 14043
rect 19484 14000 19536 14009
rect 21232 14000 21284 14052
rect 20680 13975 20732 13984
rect 20680 13941 20689 13975
rect 20689 13941 20723 13975
rect 20723 13941 20732 13975
rect 20680 13932 20732 13941
rect 18656 13864 18708 13916
rect 18840 13864 18892 13916
rect 21140 13975 21192 13984
rect 21140 13941 21149 13975
rect 21149 13941 21183 13975
rect 21183 13941 21192 13975
rect 21140 13932 21192 13941
rect 21324 13864 21376 13916
rect 23808 14000 23860 14052
rect 23900 13932 23952 13984
rect 24452 13975 24504 13984
rect 24452 13941 24461 13975
rect 24461 13941 24495 13975
rect 24495 13941 24504 13975
rect 24452 13932 24504 13941
rect 24544 13975 24596 13984
rect 24544 13941 24553 13975
rect 24553 13941 24587 13975
rect 24587 13941 24596 13975
rect 25556 13975 25608 13984
rect 24544 13932 24596 13941
rect 25556 13941 25565 13975
rect 25565 13941 25599 13975
rect 25599 13941 25608 13975
rect 25556 13932 25608 13941
rect 27212 13932 27264 13984
rect 19142 13694 19194 13746
rect 19206 13694 19258 13746
rect 19270 13694 19322 13746
rect 19334 13694 19386 13746
rect 29142 13694 29194 13746
rect 29206 13694 29258 13746
rect 29270 13694 29322 13746
rect 29334 13694 29386 13746
rect 12860 13592 12912 13644
rect 14148 13592 14200 13644
rect 14700 13592 14752 13644
rect 13412 13567 13464 13576
rect 13412 13533 13421 13567
rect 13421 13533 13455 13567
rect 13455 13533 13464 13567
rect 13412 13524 13464 13533
rect 13136 13456 13188 13508
rect 14148 13499 14200 13508
rect 14148 13465 14176 13499
rect 14176 13465 14200 13499
rect 14148 13456 14200 13465
rect 14608 13499 14660 13508
rect 14608 13465 14617 13499
rect 14617 13465 14651 13499
rect 14651 13465 14660 13499
rect 14608 13456 14660 13465
rect 14700 13499 14752 13508
rect 14700 13465 14709 13499
rect 14709 13465 14743 13499
rect 14743 13465 14752 13499
rect 14700 13456 14752 13465
rect 15068 13456 15120 13508
rect 17552 13499 17604 13508
rect 17552 13465 17561 13499
rect 17561 13465 17595 13499
rect 17595 13465 17604 13499
rect 17552 13456 17604 13465
rect 18288 13524 18340 13576
rect 18564 13499 18616 13508
rect 18564 13465 18573 13499
rect 18573 13465 18607 13499
rect 18607 13465 18616 13499
rect 18564 13456 18616 13465
rect 18932 13456 18984 13508
rect 21324 13592 21376 13644
rect 23256 13567 23308 13576
rect 20680 13456 20732 13508
rect 23256 13533 23265 13567
rect 23265 13533 23299 13567
rect 23299 13533 23308 13567
rect 23256 13524 23308 13533
rect 25188 13524 25240 13576
rect 27212 13567 27264 13576
rect 27212 13533 27221 13567
rect 27221 13533 27255 13567
rect 27255 13533 27264 13567
rect 27212 13524 27264 13533
rect 12676 13388 12728 13440
rect 13044 13388 13096 13440
rect 16908 13388 16960 13440
rect 18656 13388 18708 13440
rect 19024 13431 19076 13440
rect 19024 13397 19033 13431
rect 19033 13397 19067 13431
rect 19067 13397 19076 13431
rect 19024 13388 19076 13397
rect 21600 13499 21652 13508
rect 21600 13465 21609 13499
rect 21609 13465 21643 13499
rect 21643 13465 21652 13499
rect 21600 13456 21652 13465
rect 23808 13499 23860 13508
rect 23808 13465 23817 13499
rect 23817 13465 23851 13499
rect 23851 13465 23860 13499
rect 23808 13456 23860 13465
rect 24544 13456 24596 13508
rect 24820 13456 24872 13508
rect 17828 13320 17880 13372
rect 14608 13252 14660 13304
rect 24452 13388 24504 13440
rect 21232 13320 21284 13372
rect 21140 13252 21192 13304
rect 25556 13388 25608 13440
rect 26844 13388 26896 13440
rect 30616 13252 30668 13304
rect 14142 13150 14194 13202
rect 14206 13150 14258 13202
rect 14270 13150 14322 13202
rect 14334 13150 14386 13202
rect 24142 13150 24194 13202
rect 24206 13150 24258 13202
rect 24270 13150 24322 13202
rect 24334 13150 24386 13202
rect 14608 13048 14660 13100
rect 25188 13091 25240 13100
rect 25188 13057 25197 13091
rect 25197 13057 25231 13091
rect 25231 13057 25240 13091
rect 25188 13048 25240 13057
rect 13504 13023 13556 13032
rect 13504 12989 13513 13023
rect 13513 12989 13547 13023
rect 13547 12989 13556 13023
rect 13504 12980 13556 12989
rect 12676 12955 12728 12964
rect 12676 12921 12685 12955
rect 12685 12921 12719 12955
rect 12719 12921 12728 12955
rect 14240 12955 14292 12964
rect 12676 12912 12728 12921
rect 14240 12921 14249 12955
rect 14249 12921 14283 12955
rect 14283 12921 14292 12955
rect 14240 12912 14292 12921
rect 13136 12887 13188 12896
rect 13136 12853 13145 12887
rect 13145 12853 13179 12887
rect 13179 12853 13188 12887
rect 13136 12844 13188 12853
rect 13412 12887 13464 12896
rect 13412 12853 13421 12887
rect 13421 12853 13455 12887
rect 13455 12853 13464 12887
rect 13412 12844 13464 12853
rect 14332 12887 14384 12896
rect 14332 12853 14341 12887
rect 14341 12853 14375 12887
rect 14375 12853 14384 12887
rect 14332 12844 14384 12853
rect 14976 12844 15028 12896
rect 19576 12980 19628 13032
rect 21600 12980 21652 13032
rect 18656 12912 18708 12964
rect 15436 12844 15488 12896
rect 18564 12844 18616 12896
rect 17552 12776 17604 12828
rect 18840 12844 18892 12896
rect 15528 12708 15580 12760
rect 20588 12708 20640 12760
rect 21784 12912 21836 12964
rect 21048 12887 21100 12896
rect 21048 12853 21057 12887
rect 21057 12853 21091 12887
rect 21091 12853 21100 12887
rect 21048 12844 21100 12853
rect 21232 12844 21284 12896
rect 23256 12887 23308 12896
rect 23256 12853 23265 12887
rect 23265 12853 23299 12887
rect 23299 12853 23308 12887
rect 25004 12887 25056 12896
rect 23256 12844 23308 12853
rect 25004 12853 25013 12887
rect 25013 12853 25047 12887
rect 25047 12853 25056 12887
rect 25004 12844 25056 12853
rect 25832 12887 25884 12896
rect 25832 12853 25841 12887
rect 25841 12853 25875 12887
rect 25875 12853 25884 12887
rect 25832 12844 25884 12853
rect 21692 12819 21744 12828
rect 21692 12785 21701 12819
rect 21701 12785 21735 12819
rect 21735 12785 21744 12819
rect 21692 12776 21744 12785
rect 22704 12776 22756 12828
rect 29972 12776 30024 12828
rect 20956 12708 21008 12760
rect 23256 12708 23308 12760
rect 25832 12751 25884 12760
rect 25832 12717 25841 12751
rect 25841 12717 25875 12751
rect 25875 12717 25884 12751
rect 25832 12708 25884 12717
rect 19142 12606 19194 12658
rect 19206 12606 19258 12658
rect 19270 12606 19322 12658
rect 19334 12606 19386 12658
rect 29142 12606 29194 12658
rect 29206 12606 29258 12658
rect 29270 12606 29322 12658
rect 29334 12606 29386 12658
rect 13412 12504 13464 12556
rect 14884 12504 14936 12556
rect 22704 12504 22756 12556
rect 12860 12411 12912 12420
rect 12860 12377 12869 12411
rect 12869 12377 12903 12411
rect 12903 12377 12912 12411
rect 12860 12368 12912 12377
rect 14332 12368 14384 12420
rect 14424 12368 14476 12420
rect 15068 12436 15120 12488
rect 16908 12436 16960 12488
rect 17368 12436 17420 12488
rect 18380 12436 18432 12488
rect 19668 12436 19720 12488
rect 21692 12479 21744 12488
rect 21692 12445 21701 12479
rect 21701 12445 21735 12479
rect 21735 12445 21744 12479
rect 21692 12436 21744 12445
rect 23716 12504 23768 12556
rect 25004 12504 25056 12556
rect 23256 12436 23308 12488
rect 15436 12411 15488 12420
rect 15436 12377 15445 12411
rect 15445 12377 15479 12411
rect 15479 12377 15488 12411
rect 15436 12368 15488 12377
rect 16264 12368 16316 12420
rect 19576 12411 19628 12420
rect 19576 12377 19585 12411
rect 19585 12377 19619 12411
rect 19619 12377 19628 12411
rect 19576 12368 19628 12377
rect 20128 12411 20180 12420
rect 20128 12377 20137 12411
rect 20137 12377 20171 12411
rect 20171 12377 20180 12411
rect 20128 12368 20180 12377
rect 21416 12411 21468 12420
rect 21416 12377 21425 12411
rect 21425 12377 21459 12411
rect 21459 12377 21468 12411
rect 21416 12368 21468 12377
rect 25832 12411 25884 12420
rect 25832 12377 25841 12411
rect 25841 12377 25875 12411
rect 25875 12377 25884 12411
rect 25832 12368 25884 12377
rect 13044 12300 13096 12352
rect 14240 12300 14292 12352
rect 16724 12300 16776 12352
rect 17828 12300 17880 12352
rect 19024 12300 19076 12352
rect 21692 12300 21744 12352
rect 24912 12300 24964 12352
rect 18656 12232 18708 12284
rect 12676 12164 12728 12216
rect 15528 12164 15580 12216
rect 15712 12207 15764 12216
rect 15712 12173 15721 12207
rect 15721 12173 15755 12207
rect 15755 12173 15764 12207
rect 15712 12164 15764 12173
rect 17276 12164 17328 12216
rect 21508 12164 21560 12216
rect 23992 12164 24044 12216
rect 14142 12062 14194 12114
rect 14206 12062 14258 12114
rect 14270 12062 14322 12114
rect 14334 12062 14386 12114
rect 24142 12062 24194 12114
rect 24206 12062 24258 12114
rect 24270 12062 24322 12114
rect 24334 12062 24386 12114
rect 14516 11960 14568 12012
rect 15712 11824 15764 11876
rect 16264 11960 16316 12012
rect 20128 11960 20180 12012
rect 21048 11960 21100 12012
rect 16724 11824 16776 11876
rect 18380 11867 18432 11876
rect 18380 11833 18389 11867
rect 18389 11833 18423 11867
rect 18423 11833 18432 11867
rect 18380 11824 18432 11833
rect 18656 11867 18708 11876
rect 18656 11833 18665 11867
rect 18665 11833 18699 11867
rect 18699 11833 18708 11867
rect 18656 11824 18708 11833
rect 18748 11824 18800 11876
rect 17828 11799 17880 11808
rect 17828 11765 17837 11799
rect 17837 11765 17871 11799
rect 17871 11765 17880 11799
rect 17828 11756 17880 11765
rect 19760 11756 19812 11808
rect 21416 11824 21468 11876
rect 26844 11867 26896 11876
rect 21784 11756 21836 11808
rect 26844 11833 26853 11867
rect 26853 11833 26887 11867
rect 26887 11833 26896 11867
rect 26844 11824 26896 11833
rect 24820 11799 24872 11808
rect 24820 11765 24829 11799
rect 24829 11765 24863 11799
rect 24863 11765 24872 11799
rect 24820 11756 24872 11765
rect 16080 11688 16132 11740
rect 16724 11620 16776 11672
rect 19484 11620 19536 11672
rect 23164 11688 23216 11740
rect 25556 11688 25608 11740
rect 19142 11518 19194 11570
rect 19206 11518 19258 11570
rect 19270 11518 19322 11570
rect 19334 11518 19386 11570
rect 29142 11518 29194 11570
rect 29206 11518 29258 11570
rect 29270 11518 29322 11570
rect 29334 11518 29386 11570
rect 14976 11459 15028 11468
rect 14976 11425 14985 11459
rect 14985 11425 15019 11459
rect 15019 11425 15028 11459
rect 14976 11416 15028 11425
rect 16080 11459 16132 11468
rect 16080 11425 16089 11459
rect 16089 11425 16123 11459
rect 16123 11425 16132 11459
rect 16080 11416 16132 11425
rect 17368 11416 17420 11468
rect 19760 11416 19812 11468
rect 21324 11459 21376 11468
rect 21324 11425 21333 11459
rect 21333 11425 21367 11459
rect 21367 11425 21376 11459
rect 21324 11416 21376 11425
rect 23164 11459 23216 11468
rect 23164 11425 23173 11459
rect 23173 11425 23207 11459
rect 23207 11425 23216 11459
rect 23164 11416 23216 11425
rect 25556 11416 25608 11468
rect 25372 11391 25424 11400
rect 14516 11280 14568 11332
rect 17092 11280 17144 11332
rect 20956 11323 21008 11332
rect 20956 11289 20965 11323
rect 20965 11289 20999 11323
rect 20999 11289 21008 11323
rect 20956 11280 21008 11289
rect 25372 11357 25381 11391
rect 25381 11357 25415 11391
rect 25415 11357 25424 11391
rect 25372 11348 25424 11357
rect 23716 11280 23768 11332
rect 30892 11280 30944 11332
rect 14142 10974 14194 11026
rect 14206 10974 14258 11026
rect 14270 10974 14322 11026
rect 14334 10974 14386 11026
rect 24142 10974 24194 11026
rect 24206 10974 24258 11026
rect 24270 10974 24322 11026
rect 24334 10974 24386 11026
<< metal2 >>
rect 11018 35809 11074 36609
rect 13226 35809 13282 36609
rect 15434 35809 15490 36609
rect 17826 35809 17882 36609
rect 20034 35809 20090 36609
rect 22242 35809 22298 36609
rect 24634 35809 24690 36609
rect 26842 35809 26898 36609
rect 29234 35809 29290 36609
rect 31442 35809 31498 36609
rect 33650 35809 33706 36609
rect 11032 33438 11060 35809
rect 11020 33432 11072 33438
rect 11020 33374 11072 33380
rect 13240 32690 13268 35809
rect 14116 33876 14412 33896
rect 14172 33874 14196 33876
rect 14252 33874 14276 33876
rect 14332 33874 14356 33876
rect 14194 33822 14196 33874
rect 14258 33822 14270 33874
rect 14332 33822 14334 33874
rect 14172 33820 14196 33822
rect 14252 33820 14276 33822
rect 14332 33820 14356 33822
rect 14116 33800 14412 33820
rect 15448 33438 15476 35809
rect 15436 33432 15488 33438
rect 15436 33374 15488 33380
rect 16540 33432 16592 33438
rect 16540 33374 16592 33380
rect 13962 33128 14018 33137
rect 13962 33063 14018 33072
rect 13976 32962 14004 33063
rect 13964 32956 14016 32962
rect 13964 32898 14016 32904
rect 14116 32788 14412 32808
rect 14172 32786 14196 32788
rect 14252 32786 14276 32788
rect 14332 32786 14356 32788
rect 14194 32734 14196 32786
rect 14258 32734 14270 32786
rect 14332 32734 14334 32786
rect 14172 32732 14196 32734
rect 14252 32732 14276 32734
rect 14332 32732 14356 32734
rect 14116 32712 14412 32732
rect 13228 32684 13280 32690
rect 13228 32626 13280 32632
rect 14116 31700 14412 31720
rect 14172 31698 14196 31700
rect 14252 31698 14276 31700
rect 14332 31698 14356 31700
rect 14194 31646 14196 31698
rect 14258 31646 14270 31698
rect 14332 31646 14334 31698
rect 14172 31644 14196 31646
rect 14252 31644 14276 31646
rect 14332 31644 14356 31646
rect 14116 31624 14412 31644
rect 14116 30612 14412 30632
rect 14172 30610 14196 30612
rect 14252 30610 14276 30612
rect 14332 30610 14356 30612
rect 14194 30558 14196 30610
rect 14258 30558 14270 30610
rect 14332 30558 14334 30610
rect 14172 30556 14196 30558
rect 14252 30556 14276 30558
rect 14332 30556 14356 30558
rect 14116 30536 14412 30556
rect 16172 30304 16224 30310
rect 16172 30246 16224 30252
rect 13962 29864 14018 29873
rect 16184 29834 16212 30246
rect 13962 29799 14018 29808
rect 14516 29828 14568 29834
rect 13976 29358 14004 29799
rect 14516 29770 14568 29776
rect 16172 29828 16224 29834
rect 16172 29770 16224 29776
rect 14116 29524 14412 29544
rect 14172 29522 14196 29524
rect 14252 29522 14276 29524
rect 14332 29522 14356 29524
rect 14194 29470 14196 29522
rect 14258 29470 14270 29522
rect 14332 29470 14334 29522
rect 14172 29468 14196 29470
rect 14252 29468 14276 29470
rect 14332 29468 14356 29470
rect 14116 29448 14412 29468
rect 13964 29352 14016 29358
rect 13964 29294 14016 29300
rect 14528 28746 14556 29770
rect 16356 29624 16408 29630
rect 16356 29566 16408 29572
rect 16368 28814 16396 29566
rect 16356 28808 16408 28814
rect 16356 28750 16408 28756
rect 14516 28740 14568 28746
rect 14516 28682 14568 28688
rect 14792 28740 14844 28746
rect 14792 28682 14844 28688
rect 15344 28740 15396 28746
rect 15344 28682 15396 28688
rect 14516 28536 14568 28542
rect 14516 28478 14568 28484
rect 14116 28436 14412 28456
rect 14172 28434 14196 28436
rect 14252 28434 14276 28436
rect 14332 28434 14356 28436
rect 14194 28382 14196 28434
rect 14258 28382 14270 28434
rect 14332 28382 14334 28434
rect 14172 28380 14196 28382
rect 14252 28380 14276 28382
rect 14332 28380 14356 28382
rect 14116 28360 14412 28380
rect 14148 28196 14200 28202
rect 14148 28138 14200 28144
rect 13780 27992 13832 27998
rect 13780 27934 13832 27940
rect 11938 26328 11994 26337
rect 11938 26263 11994 26272
rect 11952 23170 11980 26263
rect 13792 25482 13820 27934
rect 14160 27726 14188 28138
rect 14528 28066 14556 28478
rect 14516 28060 14568 28066
rect 14516 28002 14568 28008
rect 14148 27720 14200 27726
rect 14148 27662 14200 27668
rect 14700 27652 14752 27658
rect 14700 27594 14752 27600
rect 14608 27584 14660 27590
rect 14608 27526 14660 27532
rect 14116 27348 14412 27368
rect 14172 27346 14196 27348
rect 14252 27346 14276 27348
rect 14332 27346 14356 27348
rect 14194 27294 14196 27346
rect 14258 27294 14270 27346
rect 14332 27294 14334 27346
rect 14172 27292 14196 27294
rect 14252 27292 14276 27294
rect 14332 27292 14356 27294
rect 14116 27272 14412 27292
rect 14516 27040 14568 27046
rect 14516 26982 14568 26988
rect 14528 26638 14556 26982
rect 14516 26632 14568 26638
rect 14516 26574 14568 26580
rect 14116 26260 14412 26280
rect 14172 26258 14196 26260
rect 14252 26258 14276 26260
rect 14332 26258 14356 26260
rect 14194 26206 14196 26258
rect 14258 26206 14270 26258
rect 14332 26206 14334 26258
rect 14172 26204 14196 26206
rect 14252 26204 14276 26206
rect 14332 26204 14356 26206
rect 14116 26184 14412 26204
rect 14528 25958 14556 26574
rect 14620 26162 14648 27526
rect 14712 27114 14740 27594
rect 14700 27108 14752 27114
rect 14700 27050 14752 27056
rect 14608 26156 14660 26162
rect 14608 26098 14660 26104
rect 14804 26026 14832 28682
rect 15356 27998 15384 28682
rect 15436 28060 15488 28066
rect 15436 28002 15488 28008
rect 15344 27992 15396 27998
rect 15344 27934 15396 27940
rect 15068 27652 15120 27658
rect 15068 27594 15120 27600
rect 14976 27040 15028 27046
rect 14976 26982 15028 26988
rect 14792 26020 14844 26026
rect 14792 25962 14844 25968
rect 14516 25952 14568 25958
rect 14516 25894 14568 25900
rect 13964 25816 14016 25822
rect 13964 25758 14016 25764
rect 13976 25550 14004 25758
rect 13964 25544 14016 25550
rect 13964 25486 14016 25492
rect 13780 25476 13832 25482
rect 13780 25418 13832 25424
rect 13412 24796 13464 24802
rect 13412 24738 13464 24744
rect 13424 24462 13452 24738
rect 13412 24456 13464 24462
rect 13412 24398 13464 24404
rect 13136 23980 13188 23986
rect 13136 23922 13188 23928
rect 11940 23164 11992 23170
rect 11940 23106 11992 23112
rect 13148 23073 13176 23922
rect 13412 23232 13464 23238
rect 13412 23174 13464 23180
rect 13134 23064 13190 23073
rect 13134 22999 13190 23008
rect 13424 22762 13452 23174
rect 13792 22898 13820 25418
rect 13964 25272 14016 25278
rect 13964 25214 14016 25220
rect 13976 24938 14004 25214
rect 14116 25172 14412 25192
rect 14172 25170 14196 25172
rect 14252 25170 14276 25172
rect 14332 25170 14356 25172
rect 14194 25118 14196 25170
rect 14258 25118 14270 25170
rect 14332 25118 14334 25170
rect 14172 25116 14196 25118
rect 14252 25116 14276 25118
rect 14332 25116 14356 25118
rect 14116 25096 14412 25116
rect 13964 24932 14016 24938
rect 13964 24874 14016 24880
rect 14700 24864 14752 24870
rect 14700 24806 14752 24812
rect 14712 24394 14740 24806
rect 14608 24388 14660 24394
rect 14608 24330 14660 24336
rect 14700 24388 14752 24394
rect 14700 24330 14752 24336
rect 14116 24084 14412 24104
rect 14172 24082 14196 24084
rect 14252 24082 14276 24084
rect 14332 24082 14356 24084
rect 14194 24030 14196 24082
rect 14258 24030 14270 24082
rect 14332 24030 14334 24082
rect 14172 24028 14196 24030
rect 14252 24028 14276 24030
rect 14332 24028 14356 24030
rect 14116 24008 14412 24028
rect 14620 23850 14648 24330
rect 14804 23866 14832 25962
rect 14988 25958 15016 26982
rect 14976 25952 15028 25958
rect 14976 25894 15028 25900
rect 15080 24870 15108 27594
rect 15344 27584 15396 27590
rect 15448 27538 15476 28002
rect 15396 27532 15476 27538
rect 15344 27526 15476 27532
rect 15528 27584 15580 27590
rect 15528 27526 15580 27532
rect 15356 27510 15476 27526
rect 15448 26502 15476 27510
rect 15436 26496 15488 26502
rect 15436 26438 15488 26444
rect 15540 24870 15568 27526
rect 15988 25408 16040 25414
rect 15988 25350 16040 25356
rect 16000 24938 16028 25350
rect 15988 24932 16040 24938
rect 15988 24874 16040 24880
rect 15068 24864 15120 24870
rect 15068 24806 15120 24812
rect 15528 24864 15580 24870
rect 15528 24806 15580 24812
rect 14608 23844 14660 23850
rect 14804 23838 14924 23866
rect 14608 23786 14660 23792
rect 14792 23776 14844 23782
rect 14792 23718 14844 23724
rect 14804 23306 14832 23718
rect 14700 23300 14752 23306
rect 14700 23242 14752 23248
rect 14792 23300 14844 23306
rect 14792 23242 14844 23248
rect 14116 22996 14412 23016
rect 14172 22994 14196 22996
rect 14252 22994 14276 22996
rect 14332 22994 14356 22996
rect 14194 22942 14196 22994
rect 14258 22942 14270 22994
rect 14332 22942 14334 22994
rect 14172 22940 14196 22942
rect 14252 22940 14276 22942
rect 14332 22940 14356 22942
rect 14116 22920 14412 22940
rect 14712 22898 14740 23242
rect 13780 22892 13832 22898
rect 13780 22834 13832 22840
rect 14700 22892 14752 22898
rect 14700 22834 14752 22840
rect 13412 22756 13464 22762
rect 13412 22698 13464 22704
rect 13792 20042 13820 22834
rect 14700 22620 14752 22626
rect 14700 22562 14752 22568
rect 14116 21908 14412 21928
rect 14172 21906 14196 21908
rect 14252 21906 14276 21908
rect 14332 21906 14356 21908
rect 14194 21854 14196 21906
rect 14258 21854 14270 21906
rect 14332 21854 14334 21906
rect 14172 21852 14196 21854
rect 14252 21852 14276 21854
rect 14332 21852 14356 21854
rect 14116 21832 14412 21852
rect 14712 21810 14740 22562
rect 14804 22150 14832 23242
rect 14792 22144 14844 22150
rect 14792 22086 14844 22092
rect 14700 21804 14752 21810
rect 14700 21746 14752 21752
rect 14896 21606 14924 23838
rect 15080 23306 15108 24806
rect 15436 23368 15488 23374
rect 15436 23310 15488 23316
rect 15068 23300 15120 23306
rect 15068 23242 15120 23248
rect 15252 23300 15304 23306
rect 15252 23242 15304 23248
rect 14608 21600 14660 21606
rect 14608 21542 14660 21548
rect 14884 21600 14936 21606
rect 14884 21542 14936 21548
rect 14116 20820 14412 20840
rect 14172 20818 14196 20820
rect 14252 20818 14276 20820
rect 14332 20818 14356 20820
rect 14194 20766 14196 20818
rect 14258 20766 14270 20818
rect 14332 20766 14334 20818
rect 14172 20764 14196 20766
rect 14252 20764 14276 20766
rect 14332 20764 14356 20766
rect 14116 20744 14412 20764
rect 14240 20444 14292 20450
rect 14240 20386 14292 20392
rect 14252 20110 14280 20386
rect 14240 20104 14292 20110
rect 14240 20046 14292 20052
rect 14516 20104 14568 20110
rect 14516 20046 14568 20052
rect 13780 20036 13832 20042
rect 13780 19978 13832 19984
rect 12674 19800 12730 19809
rect 12674 19735 12730 19744
rect 12400 17384 12452 17390
rect 12400 17326 12452 17332
rect 12412 17254 12440 17326
rect 12688 17322 12716 19735
rect 13792 18546 13820 19978
rect 14116 19732 14412 19752
rect 14172 19730 14196 19732
rect 14252 19730 14276 19732
rect 14332 19730 14356 19732
rect 14194 19678 14196 19730
rect 14258 19678 14270 19730
rect 14332 19678 14334 19730
rect 14172 19676 14196 19678
rect 14252 19676 14276 19678
rect 14332 19676 14356 19678
rect 14116 19656 14412 19676
rect 14528 19634 14556 20046
rect 14516 19628 14568 19634
rect 14516 19570 14568 19576
rect 14620 19430 14648 21542
rect 15264 20518 15292 23242
rect 15448 22762 15476 23310
rect 15540 23238 15568 24806
rect 16000 23238 16028 24874
rect 16552 23918 16580 33374
rect 17840 32978 17868 35809
rect 19116 34420 19412 34440
rect 19172 34418 19196 34420
rect 19252 34418 19276 34420
rect 19332 34418 19356 34420
rect 19194 34366 19196 34418
rect 19258 34366 19270 34418
rect 19332 34366 19334 34418
rect 19172 34364 19196 34366
rect 19252 34364 19276 34366
rect 19332 34364 19356 34366
rect 19116 34344 19412 34364
rect 20048 33658 20076 35809
rect 22256 35698 22284 35809
rect 22072 35670 22284 35698
rect 20048 33642 20168 33658
rect 20048 33636 20180 33642
rect 20048 33630 20128 33636
rect 20128 33578 20180 33584
rect 20036 33568 20088 33574
rect 20036 33510 20088 33516
rect 19116 33332 19412 33352
rect 19172 33330 19196 33332
rect 19252 33330 19276 33332
rect 19332 33330 19356 33332
rect 19194 33278 19196 33330
rect 19258 33278 19270 33330
rect 19332 33278 19334 33330
rect 19172 33276 19196 33278
rect 19252 33276 19276 33278
rect 19332 33276 19356 33278
rect 19116 33256 19412 33276
rect 20048 33030 20076 33510
rect 20496 33500 20548 33506
rect 20496 33442 20548 33448
rect 21508 33500 21560 33506
rect 21508 33442 21560 33448
rect 20036 33024 20088 33030
rect 17840 32950 18236 32978
rect 20036 32966 20088 32972
rect 18208 32146 18236 32950
rect 19760 32480 19812 32486
rect 19760 32422 19812 32428
rect 19116 32244 19412 32264
rect 19172 32242 19196 32244
rect 19252 32242 19276 32244
rect 19332 32242 19356 32244
rect 19194 32190 19196 32242
rect 19258 32190 19270 32242
rect 19332 32190 19334 32242
rect 19172 32188 19196 32190
rect 19252 32188 19276 32190
rect 19332 32188 19356 32190
rect 19116 32168 19412 32188
rect 18196 32140 18248 32146
rect 18196 32082 18248 32088
rect 19772 32078 19800 32422
rect 19760 32072 19812 32078
rect 19760 32014 19812 32020
rect 20048 31466 20076 32966
rect 20508 31534 20536 33442
rect 21416 33432 21468 33438
rect 21416 33374 21468 33380
rect 20588 33092 20640 33098
rect 20588 33034 20640 33040
rect 20600 32010 20628 33034
rect 21140 32888 21192 32894
rect 21140 32830 21192 32836
rect 20588 32004 20640 32010
rect 20588 31946 20640 31952
rect 20496 31528 20548 31534
rect 20496 31470 20548 31476
rect 21152 31466 21180 32830
rect 21324 32616 21376 32622
rect 21324 32558 21376 32564
rect 21336 31534 21364 32558
rect 21428 32554 21456 33374
rect 21520 33098 21548 33442
rect 21508 33092 21560 33098
rect 21508 33034 21560 33040
rect 21416 32548 21468 32554
rect 21416 32490 21468 32496
rect 21520 32486 21548 33034
rect 21692 32684 21744 32690
rect 21692 32626 21744 32632
rect 21508 32480 21560 32486
rect 21508 32422 21560 32428
rect 21520 32146 21548 32422
rect 21508 32140 21560 32146
rect 21508 32082 21560 32088
rect 21324 31528 21376 31534
rect 21324 31470 21376 31476
rect 20036 31460 20088 31466
rect 20036 31402 20088 31408
rect 21140 31460 21192 31466
rect 21140 31402 21192 31408
rect 20956 31324 21008 31330
rect 20956 31266 21008 31272
rect 19116 31156 19412 31176
rect 19172 31154 19196 31156
rect 19252 31154 19276 31156
rect 19332 31154 19356 31156
rect 19194 31102 19196 31154
rect 19258 31102 19270 31154
rect 19332 31102 19334 31154
rect 19172 31100 19196 31102
rect 19252 31100 19276 31102
rect 19332 31100 19356 31102
rect 19116 31080 19412 31100
rect 20128 30916 20180 30922
rect 20128 30858 20180 30864
rect 16816 30440 16868 30446
rect 16816 30382 16868 30388
rect 16828 29834 16856 30382
rect 20140 30378 20168 30858
rect 20128 30372 20180 30378
rect 20128 30314 20180 30320
rect 20220 30304 20272 30310
rect 20220 30246 20272 30252
rect 19944 30236 19996 30242
rect 19944 30178 19996 30184
rect 17828 30168 17880 30174
rect 17828 30110 17880 30116
rect 18472 30168 18524 30174
rect 18472 30110 18524 30116
rect 17840 29902 17868 30110
rect 17828 29896 17880 29902
rect 17828 29838 17880 29844
rect 16816 29828 16868 29834
rect 16816 29770 16868 29776
rect 16828 28898 16856 29770
rect 18484 29766 18512 30110
rect 19116 30068 19412 30088
rect 19172 30066 19196 30068
rect 19252 30066 19276 30068
rect 19332 30066 19356 30068
rect 19194 30014 19196 30066
rect 19258 30014 19270 30066
rect 19332 30014 19334 30066
rect 19172 30012 19196 30014
rect 19252 30012 19276 30014
rect 19332 30012 19356 30014
rect 19116 29992 19412 30012
rect 19956 29766 19984 30178
rect 20232 29902 20260 30246
rect 20588 30236 20640 30242
rect 20508 30196 20588 30224
rect 20404 30168 20456 30174
rect 20324 30128 20404 30156
rect 20220 29896 20272 29902
rect 20220 29838 20272 29844
rect 17092 29760 17144 29766
rect 17092 29702 17144 29708
rect 18472 29760 18524 29766
rect 18472 29702 18524 29708
rect 19944 29760 19996 29766
rect 19944 29702 19996 29708
rect 17000 29216 17052 29222
rect 17000 29158 17052 29164
rect 16828 28882 16948 28898
rect 16828 28876 16960 28882
rect 16828 28870 16908 28876
rect 16908 28818 16960 28824
rect 17012 28746 17040 29158
rect 17000 28740 17052 28746
rect 17000 28682 17052 28688
rect 16816 28672 16868 28678
rect 16816 28614 16868 28620
rect 16828 28202 16856 28614
rect 16816 28196 16868 28202
rect 16816 28138 16868 28144
rect 16908 27652 16960 27658
rect 16908 27594 16960 27600
rect 16632 26972 16684 26978
rect 16632 26914 16684 26920
rect 16644 25958 16672 26914
rect 16920 26026 16948 27594
rect 17012 27114 17040 28682
rect 17104 27726 17132 29702
rect 17184 29216 17236 29222
rect 17184 29158 17236 29164
rect 17276 29216 17328 29222
rect 17276 29158 17328 29164
rect 17736 29216 17788 29222
rect 17736 29158 17788 29164
rect 17196 28134 17224 29158
rect 17288 28814 17316 29158
rect 17276 28808 17328 28814
rect 17276 28750 17328 28756
rect 17184 28128 17236 28134
rect 17184 28070 17236 28076
rect 17092 27720 17144 27726
rect 17092 27662 17144 27668
rect 17288 27538 17316 28750
rect 17748 28678 17776 29158
rect 17736 28672 17788 28678
rect 17736 28614 17788 28620
rect 18288 28672 18340 28678
rect 18288 28614 18340 28620
rect 17748 28134 17776 28614
rect 17644 28128 17696 28134
rect 17644 28070 17696 28076
rect 17736 28128 17788 28134
rect 17736 28070 17788 28076
rect 18196 28128 18248 28134
rect 18196 28070 18248 28076
rect 17656 27658 17684 28070
rect 17552 27652 17604 27658
rect 17552 27594 17604 27600
rect 17644 27652 17696 27658
rect 17644 27594 17696 27600
rect 17104 27510 17316 27538
rect 17000 27108 17052 27114
rect 17000 27050 17052 27056
rect 17104 26910 17132 27510
rect 17564 27182 17592 27594
rect 17552 27176 17604 27182
rect 17552 27118 17604 27124
rect 17276 27040 17328 27046
rect 17276 26982 17328 26988
rect 17644 27040 17696 27046
rect 17644 26982 17696 26988
rect 17092 26904 17144 26910
rect 17092 26846 17144 26852
rect 16908 26020 16960 26026
rect 16908 25962 16960 25968
rect 16632 25952 16684 25958
rect 16632 25894 16684 25900
rect 16644 24462 16672 25894
rect 17104 25550 17132 26846
rect 17288 25958 17316 26982
rect 17552 26700 17604 26706
rect 17552 26642 17604 26648
rect 17564 25958 17592 26642
rect 17656 26638 17684 26982
rect 17644 26632 17696 26638
rect 17644 26574 17696 26580
rect 17276 25952 17328 25958
rect 17276 25894 17328 25900
rect 17552 25952 17604 25958
rect 17552 25894 17604 25900
rect 17092 25544 17144 25550
rect 17092 25486 17144 25492
rect 17656 25482 17684 26574
rect 16724 25476 16776 25482
rect 16724 25418 16776 25424
rect 17644 25476 17696 25482
rect 17644 25418 17696 25424
rect 16632 24456 16684 24462
rect 16632 24398 16684 24404
rect 16632 24320 16684 24326
rect 16632 24262 16684 24268
rect 16540 23912 16592 23918
rect 16540 23854 16592 23860
rect 16080 23776 16132 23782
rect 16080 23718 16132 23724
rect 15528 23232 15580 23238
rect 15528 23174 15580 23180
rect 15988 23232 16040 23238
rect 15988 23174 16040 23180
rect 15436 22756 15488 22762
rect 15436 22698 15488 22704
rect 15448 22150 15476 22698
rect 15436 22144 15488 22150
rect 15436 22086 15488 22092
rect 15540 22098 15568 23174
rect 16092 22762 16120 23718
rect 16080 22756 16132 22762
rect 16080 22698 16132 22704
rect 15620 22688 15672 22694
rect 15620 22630 15672 22636
rect 15896 22688 15948 22694
rect 15896 22630 15948 22636
rect 15632 22286 15660 22630
rect 15620 22280 15672 22286
rect 15620 22222 15672 22228
rect 15908 22150 15936 22630
rect 16092 22150 16120 22698
rect 16644 22694 16672 24262
rect 16736 23850 16764 25418
rect 17748 25346 17776 28070
rect 18104 27652 18156 27658
rect 18104 27594 18156 27600
rect 18012 27108 18064 27114
rect 18012 27050 18064 27056
rect 17920 27040 17972 27046
rect 17920 26982 17972 26988
rect 17932 26706 17960 26982
rect 17920 26700 17972 26706
rect 17920 26642 17972 26648
rect 17828 26564 17880 26570
rect 17828 26506 17880 26512
rect 17840 26026 17868 26506
rect 18024 26502 18052 27050
rect 18012 26496 18064 26502
rect 18012 26438 18064 26444
rect 18116 26434 18144 27594
rect 18208 27590 18236 28070
rect 18300 28066 18328 28614
rect 18288 28060 18340 28066
rect 18288 28002 18340 28008
rect 18484 27658 18512 29702
rect 19956 29154 19984 29702
rect 19944 29148 19996 29154
rect 19944 29090 19996 29096
rect 19116 28980 19412 29000
rect 19172 28978 19196 28980
rect 19252 28978 19276 28980
rect 19332 28978 19356 28980
rect 19194 28926 19196 28978
rect 19258 28926 19270 28978
rect 19332 28926 19334 28978
rect 19172 28924 19196 28926
rect 19252 28924 19276 28926
rect 19332 28924 19356 28926
rect 19116 28904 19412 28924
rect 19116 27892 19412 27912
rect 19172 27890 19196 27892
rect 19252 27890 19276 27892
rect 19332 27890 19356 27892
rect 19194 27838 19196 27890
rect 19258 27838 19270 27890
rect 19332 27838 19334 27890
rect 19172 27836 19196 27838
rect 19252 27836 19276 27838
rect 19332 27836 19356 27838
rect 19116 27816 19412 27836
rect 18472 27652 18524 27658
rect 18472 27594 18524 27600
rect 19956 27590 19984 29090
rect 20036 28128 20088 28134
rect 20036 28070 20088 28076
rect 18196 27584 18248 27590
rect 18196 27526 18248 27532
rect 19944 27584 19996 27590
rect 19944 27526 19996 27532
rect 19116 26804 19412 26824
rect 19172 26802 19196 26804
rect 19252 26802 19276 26804
rect 19332 26802 19356 26804
rect 19194 26750 19196 26802
rect 19258 26750 19270 26802
rect 19332 26750 19334 26802
rect 19172 26748 19196 26750
rect 19252 26748 19276 26750
rect 19332 26748 19356 26750
rect 19116 26728 19412 26748
rect 19956 26638 19984 27526
rect 19944 26632 19996 26638
rect 19944 26574 19996 26580
rect 19576 26564 19628 26570
rect 19576 26506 19628 26512
rect 18104 26428 18156 26434
rect 18104 26370 18156 26376
rect 18472 26428 18524 26434
rect 18472 26370 18524 26376
rect 17828 26020 17880 26026
rect 17828 25962 17880 25968
rect 17840 25482 17868 25962
rect 17828 25476 17880 25482
rect 17828 25418 17880 25424
rect 17736 25340 17788 25346
rect 17736 25282 17788 25288
rect 16908 24864 16960 24870
rect 16908 24806 16960 24812
rect 16920 24394 16948 24806
rect 17460 24796 17512 24802
rect 17460 24738 17512 24744
rect 17472 24394 17500 24738
rect 17840 24394 17868 25418
rect 18484 24394 18512 26370
rect 19484 26020 19536 26026
rect 19484 25962 19536 25968
rect 19116 25716 19412 25736
rect 19172 25714 19196 25716
rect 19252 25714 19276 25716
rect 19332 25714 19356 25716
rect 19194 25662 19196 25714
rect 19258 25662 19270 25714
rect 19332 25662 19334 25714
rect 19172 25660 19196 25662
rect 19252 25660 19276 25662
rect 19332 25660 19356 25662
rect 19116 25640 19412 25660
rect 19496 25550 19524 25962
rect 19484 25544 19536 25550
rect 19484 25486 19536 25492
rect 19024 25476 19076 25482
rect 19024 25418 19076 25424
rect 18656 25340 18708 25346
rect 18656 25282 18708 25288
rect 18668 24734 18696 25282
rect 18656 24728 18708 24734
rect 18656 24670 18708 24676
rect 18668 24394 18696 24670
rect 16908 24388 16960 24394
rect 16908 24330 16960 24336
rect 17460 24388 17512 24394
rect 17460 24330 17512 24336
rect 17828 24388 17880 24394
rect 17828 24330 17880 24336
rect 18472 24388 18524 24394
rect 18472 24330 18524 24336
rect 18656 24388 18708 24394
rect 18656 24330 18708 24336
rect 16724 23844 16776 23850
rect 16724 23786 16776 23792
rect 16736 23306 16764 23786
rect 16920 23442 16948 24330
rect 16908 23436 16960 23442
rect 16908 23378 16960 23384
rect 17840 23306 17868 24330
rect 18932 24320 18984 24326
rect 18932 24262 18984 24268
rect 18944 23850 18972 24262
rect 18932 23844 18984 23850
rect 18932 23786 18984 23792
rect 18380 23776 18432 23782
rect 18380 23718 18432 23724
rect 18012 23708 18064 23714
rect 18012 23650 18064 23656
rect 18024 23374 18052 23650
rect 18012 23368 18064 23374
rect 18012 23310 18064 23316
rect 16724 23300 16776 23306
rect 16724 23242 16776 23248
rect 17828 23300 17880 23306
rect 17828 23242 17880 23248
rect 16632 22688 16684 22694
rect 16632 22630 16684 22636
rect 16736 22218 16764 23242
rect 17840 22354 17868 23242
rect 18024 22694 18052 23310
rect 18392 23306 18420 23718
rect 18380 23300 18432 23306
rect 18432 23260 18512 23288
rect 18380 23242 18432 23248
rect 18484 23209 18512 23260
rect 18470 23200 18526 23209
rect 18470 23135 18526 23144
rect 18484 22830 18512 23135
rect 18944 23102 18972 23786
rect 19036 23782 19064 25418
rect 19496 24938 19524 25486
rect 19588 25482 19616 26506
rect 19668 26496 19720 26502
rect 19668 26438 19720 26444
rect 19576 25476 19628 25482
rect 19576 25418 19628 25424
rect 19484 24932 19536 24938
rect 19484 24874 19536 24880
rect 19116 24628 19412 24648
rect 19172 24626 19196 24628
rect 19252 24626 19276 24628
rect 19332 24626 19356 24628
rect 19194 24574 19196 24626
rect 19258 24574 19270 24626
rect 19332 24574 19334 24626
rect 19172 24572 19196 24574
rect 19252 24572 19276 24574
rect 19332 24572 19356 24574
rect 19116 24552 19412 24572
rect 19496 24394 19524 24874
rect 19576 24864 19628 24870
rect 19576 24806 19628 24812
rect 19588 24462 19616 24806
rect 19680 24802 19708 26438
rect 19852 26360 19904 26366
rect 19852 26302 19904 26308
rect 19864 25482 19892 26302
rect 19852 25476 19904 25482
rect 19852 25418 19904 25424
rect 19668 24796 19720 24802
rect 19668 24738 19720 24744
rect 19576 24456 19628 24462
rect 19576 24398 19628 24404
rect 19208 24388 19260 24394
rect 19208 24330 19260 24336
rect 19484 24388 19536 24394
rect 19484 24330 19536 24336
rect 19220 23850 19248 24330
rect 19208 23844 19260 23850
rect 19208 23786 19260 23792
rect 19588 23782 19616 24398
rect 20048 24394 20076 28070
rect 20232 27794 20260 29838
rect 20220 27788 20272 27794
rect 20220 27730 20272 27736
rect 20232 26910 20260 27730
rect 20324 27658 20352 30128
rect 20404 30110 20456 30116
rect 20508 29850 20536 30196
rect 20588 30178 20640 30184
rect 20968 29902 20996 31266
rect 21140 31256 21192 31262
rect 21140 31198 21192 31204
rect 21152 30990 21180 31198
rect 21140 30984 21192 30990
rect 21140 30926 21192 30932
rect 21152 30854 21180 30926
rect 21704 30854 21732 32626
rect 21140 30848 21192 30854
rect 21140 30790 21192 30796
rect 21600 30848 21652 30854
rect 21600 30790 21652 30796
rect 21692 30848 21744 30854
rect 21692 30790 21744 30796
rect 21232 30712 21284 30718
rect 21232 30654 21284 30660
rect 20956 29896 21008 29902
rect 20508 29834 20720 29850
rect 20956 29838 21008 29844
rect 20508 29828 20732 29834
rect 20508 29822 20680 29828
rect 20508 29086 20536 29822
rect 20680 29770 20732 29776
rect 20864 29828 20916 29834
rect 20864 29770 20916 29776
rect 20876 29136 20904 29770
rect 21244 29290 21272 30654
rect 21612 30310 21640 30790
rect 21600 30304 21652 30310
rect 21600 30246 21652 30252
rect 21232 29284 21284 29290
rect 21232 29226 21284 29232
rect 21876 29284 21928 29290
rect 21876 29226 21928 29232
rect 21416 29216 21468 29222
rect 21416 29158 21468 29164
rect 20956 29148 21008 29154
rect 20876 29108 20956 29136
rect 20956 29090 21008 29096
rect 20496 29080 20548 29086
rect 20496 29022 20548 29028
rect 20508 28610 20536 29022
rect 20968 28814 20996 29090
rect 21428 28814 21456 29158
rect 20956 28808 21008 28814
rect 20956 28750 21008 28756
rect 21416 28808 21468 28814
rect 21416 28750 21468 28756
rect 21692 28808 21744 28814
rect 21692 28750 21744 28756
rect 21508 28740 21560 28746
rect 21508 28682 21560 28688
rect 20496 28604 20548 28610
rect 20496 28546 20548 28552
rect 20508 28066 20536 28546
rect 20496 28060 20548 28066
rect 20496 28002 20548 28008
rect 20404 27992 20456 27998
rect 20404 27934 20456 27940
rect 20416 27726 20444 27934
rect 20508 27726 20536 28002
rect 20588 27788 20640 27794
rect 20588 27730 20640 27736
rect 20404 27720 20456 27726
rect 20404 27662 20456 27668
rect 20496 27720 20548 27726
rect 20496 27662 20548 27668
rect 20312 27652 20364 27658
rect 20312 27594 20364 27600
rect 20220 26904 20272 26910
rect 20220 26846 20272 26852
rect 20232 26570 20260 26846
rect 20416 26706 20444 27662
rect 20600 27658 20628 27730
rect 21416 27720 21468 27726
rect 21416 27662 21468 27668
rect 20588 27652 20640 27658
rect 20588 27594 20640 27600
rect 20404 26700 20456 26706
rect 20404 26642 20456 26648
rect 20416 26570 20444 26642
rect 20220 26564 20272 26570
rect 20404 26564 20456 26570
rect 20220 26506 20272 26512
rect 20324 26524 20404 26552
rect 20324 26026 20352 26524
rect 20404 26506 20456 26512
rect 20496 26564 20548 26570
rect 20496 26506 20548 26512
rect 20508 26450 20536 26506
rect 20416 26422 20536 26450
rect 20312 26020 20364 26026
rect 20312 25962 20364 25968
rect 20324 25890 20352 25962
rect 20416 25958 20444 26422
rect 20404 25952 20456 25958
rect 20404 25894 20456 25900
rect 20312 25884 20364 25890
rect 20312 25826 20364 25832
rect 20416 25482 20444 25894
rect 20404 25476 20456 25482
rect 20404 25418 20456 25424
rect 19668 24388 19720 24394
rect 19668 24330 19720 24336
rect 20036 24388 20088 24394
rect 20036 24330 20088 24336
rect 19024 23776 19076 23782
rect 19024 23718 19076 23724
rect 19576 23776 19628 23782
rect 19576 23718 19628 23724
rect 18932 23096 18984 23102
rect 18932 23038 18984 23044
rect 18472 22824 18524 22830
rect 18472 22766 18524 22772
rect 18012 22688 18064 22694
rect 18012 22630 18064 22636
rect 18380 22688 18432 22694
rect 18380 22630 18432 22636
rect 18392 22354 18420 22630
rect 18840 22552 18892 22558
rect 18840 22494 18892 22500
rect 17828 22348 17880 22354
rect 17828 22290 17880 22296
rect 18380 22348 18432 22354
rect 18380 22290 18432 22296
rect 16172 22212 16224 22218
rect 16172 22154 16224 22160
rect 16724 22212 16776 22218
rect 16724 22154 16776 22160
rect 15896 22144 15948 22150
rect 15540 22070 15660 22098
rect 15896 22086 15948 22092
rect 16080 22144 16132 22150
rect 16080 22086 16132 22092
rect 15528 21600 15580 21606
rect 15528 21542 15580 21548
rect 15344 20920 15396 20926
rect 15344 20862 15396 20868
rect 14976 20512 15028 20518
rect 14976 20454 15028 20460
rect 15252 20512 15304 20518
rect 15252 20454 15304 20460
rect 14988 20178 15016 20454
rect 14976 20172 15028 20178
rect 14976 20114 15028 20120
rect 15356 19906 15384 20862
rect 15540 20586 15568 21542
rect 15632 20926 15660 22070
rect 15908 21742 15936 22086
rect 15896 21736 15948 21742
rect 15896 21678 15948 21684
rect 16184 21674 16212 22154
rect 16172 21668 16224 21674
rect 16172 21610 16224 21616
rect 16080 21532 16132 21538
rect 16080 21474 16132 21480
rect 16092 21062 16120 21474
rect 16184 21146 16212 21610
rect 17840 21606 17868 22290
rect 17920 22212 17972 22218
rect 17920 22154 17972 22160
rect 17460 21600 17512 21606
rect 17460 21542 17512 21548
rect 17828 21600 17880 21606
rect 17828 21542 17880 21548
rect 17276 21464 17328 21470
rect 17276 21406 17328 21412
rect 16184 21130 16488 21146
rect 16172 21124 16500 21130
rect 16224 21118 16448 21124
rect 16172 21066 16224 21072
rect 16448 21066 16500 21072
rect 15988 21056 16040 21062
rect 15988 20998 16040 21004
rect 16080 21056 16132 21062
rect 16080 20998 16132 21004
rect 15620 20920 15672 20926
rect 15620 20862 15672 20868
rect 15528 20580 15580 20586
rect 15528 20522 15580 20528
rect 15344 19900 15396 19906
rect 15344 19842 15396 19848
rect 15356 19430 15384 19842
rect 15540 19498 15568 20522
rect 15632 20518 15660 20862
rect 16000 20586 16028 20998
rect 15988 20580 16040 20586
rect 15988 20522 16040 20528
rect 15620 20512 15672 20518
rect 15620 20454 15672 20460
rect 16000 20110 16028 20522
rect 15988 20104 16040 20110
rect 15988 20046 16040 20052
rect 15528 19492 15580 19498
rect 15528 19434 15580 19440
rect 14608 19424 14660 19430
rect 14608 19366 14660 19372
rect 15344 19424 15396 19430
rect 15344 19366 15396 19372
rect 14116 18644 14412 18664
rect 14172 18642 14196 18644
rect 14252 18642 14276 18644
rect 14332 18642 14356 18644
rect 14194 18590 14196 18642
rect 14258 18590 14270 18642
rect 14332 18590 14334 18642
rect 14172 18588 14196 18590
rect 14252 18588 14276 18590
rect 14332 18588 14356 18590
rect 14116 18568 14412 18588
rect 13780 18540 13832 18546
rect 13780 18482 13832 18488
rect 13792 17866 13820 18482
rect 14620 18342 14648 19366
rect 14608 18336 14660 18342
rect 14608 18278 14660 18284
rect 15988 18336 16040 18342
rect 15988 18278 16040 18284
rect 14700 18200 14752 18206
rect 14700 18142 14752 18148
rect 15620 18200 15672 18206
rect 15620 18142 15672 18148
rect 14712 17934 14740 18142
rect 14700 17928 14752 17934
rect 14700 17870 14752 17876
rect 13780 17860 13832 17866
rect 13780 17802 13832 17808
rect 12676 17316 12728 17322
rect 12676 17258 12728 17264
rect 12400 17248 12452 17254
rect 12400 17190 12452 17196
rect 12412 16778 12440 17190
rect 12492 17180 12544 17186
rect 12492 17122 12544 17128
rect 12400 16772 12452 16778
rect 12400 16714 12452 16720
rect 12504 16234 12532 17122
rect 12688 16846 12716 17258
rect 12676 16840 12728 16846
rect 12676 16782 12728 16788
rect 12768 16704 12820 16710
rect 12768 16646 12820 16652
rect 12492 16228 12544 16234
rect 12492 16170 12544 16176
rect 12400 16160 12452 16166
rect 12400 16102 12452 16108
rect 12412 15146 12440 16102
rect 12504 15690 12532 16170
rect 12676 16160 12728 16166
rect 12676 16102 12728 16108
rect 12492 15684 12544 15690
rect 12492 15626 12544 15632
rect 12688 15536 12716 16102
rect 12780 15690 12808 16646
rect 13792 15690 13820 17802
rect 14116 17556 14412 17576
rect 14172 17554 14196 17556
rect 14252 17554 14276 17556
rect 14332 17554 14356 17556
rect 14194 17502 14196 17554
rect 14258 17502 14270 17554
rect 14332 17502 14334 17554
rect 14172 17500 14196 17502
rect 14252 17500 14276 17502
rect 14332 17500 14356 17502
rect 14116 17480 14412 17500
rect 15344 17452 15396 17458
rect 15344 17394 15396 17400
rect 15356 17254 15384 17394
rect 15344 17248 15396 17254
rect 15344 17190 15396 17196
rect 13964 16568 14016 16574
rect 13964 16510 14016 16516
rect 13976 16273 14004 16510
rect 14116 16468 14412 16488
rect 14172 16466 14196 16468
rect 14252 16466 14276 16468
rect 14332 16466 14356 16468
rect 14194 16414 14196 16466
rect 14258 16414 14270 16466
rect 14332 16414 14334 16466
rect 14172 16412 14196 16414
rect 14252 16412 14276 16414
rect 14332 16412 14356 16414
rect 14116 16392 14412 16412
rect 13962 16264 14018 16273
rect 15356 16234 15384 17190
rect 15632 17118 15660 18142
rect 16000 17934 16028 18278
rect 15988 17928 16040 17934
rect 15988 17870 16040 17876
rect 15620 17112 15672 17118
rect 15620 17054 15672 17060
rect 15632 16778 15660 17054
rect 15620 16772 15672 16778
rect 15620 16714 15672 16720
rect 13962 16199 14018 16208
rect 15344 16228 15396 16234
rect 15344 16170 15396 16176
rect 15620 16160 15672 16166
rect 15620 16102 15672 16108
rect 14792 16092 14844 16098
rect 14792 16034 14844 16040
rect 14516 16024 14568 16030
rect 14516 15966 14568 15972
rect 12768 15684 12820 15690
rect 12768 15626 12820 15632
rect 12952 15684 13004 15690
rect 12952 15626 13004 15632
rect 13780 15684 13832 15690
rect 13780 15626 13832 15632
rect 12768 15548 12820 15554
rect 12688 15508 12768 15536
rect 12768 15490 12820 15496
rect 12400 15140 12452 15146
rect 12400 15082 12452 15088
rect 12780 14602 12808 15490
rect 12860 14732 12912 14738
rect 12860 14674 12912 14680
rect 12768 14596 12820 14602
rect 12768 14538 12820 14544
rect 12032 14528 12084 14534
rect 12032 14470 12084 14476
rect 12044 14194 12072 14470
rect 12032 14188 12084 14194
rect 12032 14130 12084 14136
rect 12872 13990 12900 14674
rect 12964 14194 12992 15626
rect 14116 15380 14412 15400
rect 14172 15378 14196 15380
rect 14252 15378 14276 15380
rect 14332 15378 14356 15380
rect 14194 15326 14196 15378
rect 14258 15326 14270 15378
rect 14332 15326 14334 15378
rect 14172 15324 14196 15326
rect 14252 15324 14276 15326
rect 14332 15324 14356 15326
rect 14116 15304 14412 15324
rect 13044 15072 13096 15078
rect 13044 15014 13096 15020
rect 13412 15072 13464 15078
rect 13412 15014 13464 15020
rect 13504 15072 13556 15078
rect 13504 15014 13556 15020
rect 13056 14670 13084 15014
rect 13044 14664 13096 14670
rect 13044 14606 13096 14612
rect 13424 14602 13452 15014
rect 13412 14596 13464 14602
rect 13412 14538 13464 14544
rect 12952 14188 13004 14194
rect 12952 14130 13004 14136
rect 10468 13984 10520 13990
rect 10468 13926 10520 13932
rect 12860 13984 12912 13990
rect 12860 13926 12912 13932
rect 10480 9624 10508 13926
rect 12860 13644 12912 13650
rect 12860 13586 12912 13592
rect 12676 13440 12728 13446
rect 12676 13382 12728 13388
rect 12688 13009 12716 13382
rect 12674 13000 12730 13009
rect 12674 12935 12676 12944
rect 12728 12935 12730 12944
rect 12676 12906 12728 12912
rect 12872 12426 12900 13586
rect 13424 13582 13452 14538
rect 13516 13922 13544 15014
rect 14528 14602 14556 15966
rect 14804 14738 14832 16034
rect 15632 15554 15660 16102
rect 15712 15684 15764 15690
rect 15712 15626 15764 15632
rect 15620 15548 15672 15554
rect 15620 15490 15672 15496
rect 15632 15214 15660 15490
rect 15620 15208 15672 15214
rect 15620 15150 15672 15156
rect 15068 15072 15120 15078
rect 15068 15014 15120 15020
rect 14792 14732 14844 14738
rect 14792 14674 14844 14680
rect 14516 14596 14568 14602
rect 14516 14538 14568 14544
rect 14792 14460 14844 14466
rect 14792 14402 14844 14408
rect 14116 14292 14412 14312
rect 14172 14290 14196 14292
rect 14252 14290 14276 14292
rect 14332 14290 14356 14292
rect 14194 14238 14196 14290
rect 14258 14238 14270 14290
rect 14332 14238 14334 14290
rect 14172 14236 14196 14238
rect 14252 14236 14276 14238
rect 14332 14236 14356 14238
rect 14116 14216 14412 14236
rect 14700 14120 14752 14126
rect 14700 14062 14752 14068
rect 13504 13916 13556 13922
rect 13504 13858 13556 13864
rect 13412 13576 13464 13582
rect 13412 13518 13464 13524
rect 13136 13508 13188 13514
rect 13136 13450 13188 13456
rect 13044 13440 13096 13446
rect 13044 13382 13096 13388
rect 12860 12420 12912 12426
rect 12860 12362 12912 12368
rect 13056 12358 13084 13382
rect 13148 12902 13176 13450
rect 13516 13038 13544 13858
rect 14712 13650 14740 14062
rect 14804 13990 14832 14402
rect 14792 13984 14844 13990
rect 14792 13926 14844 13932
rect 14148 13644 14200 13650
rect 14148 13586 14200 13592
rect 14700 13644 14752 13650
rect 14700 13586 14752 13592
rect 14160 13514 14188 13586
rect 14712 13514 14740 13586
rect 15080 13514 15108 15014
rect 15724 14738 15752 15626
rect 15988 15616 16040 15622
rect 15988 15558 16040 15564
rect 16000 15282 16028 15558
rect 15988 15276 16040 15282
rect 15988 15218 16040 15224
rect 15896 14936 15948 14942
rect 15896 14878 15948 14884
rect 15908 14738 15936 14878
rect 15712 14732 15764 14738
rect 15712 14674 15764 14680
rect 15896 14732 15948 14738
rect 15896 14674 15948 14680
rect 16184 14058 16212 21066
rect 17288 20450 17316 21406
rect 17472 20926 17500 21542
rect 17840 21198 17868 21542
rect 17828 21192 17880 21198
rect 17828 21134 17880 21140
rect 17932 21130 17960 22154
rect 18288 22144 18340 22150
rect 18288 22086 18340 22092
rect 18012 22008 18064 22014
rect 18012 21950 18064 21956
rect 18024 21198 18052 21950
rect 18300 21606 18328 22086
rect 18852 21606 18880 22494
rect 19036 22150 19064 23718
rect 19116 23540 19412 23560
rect 19172 23538 19196 23540
rect 19252 23538 19276 23540
rect 19332 23538 19356 23540
rect 19194 23486 19196 23538
rect 19258 23486 19270 23538
rect 19332 23486 19334 23538
rect 19172 23484 19196 23486
rect 19252 23484 19276 23486
rect 19332 23484 19356 23486
rect 19116 23464 19412 23484
rect 19484 23368 19536 23374
rect 19220 23316 19484 23322
rect 19220 23310 19536 23316
rect 19220 23306 19524 23310
rect 19588 23306 19616 23718
rect 19680 23714 19708 24330
rect 19852 24320 19904 24326
rect 19852 24262 19904 24268
rect 19864 23782 19892 24262
rect 20416 24190 20444 25418
rect 20404 24184 20456 24190
rect 20404 24126 20456 24132
rect 19852 23776 19904 23782
rect 19852 23718 19904 23724
rect 20128 23776 20180 23782
rect 20128 23718 20180 23724
rect 19668 23708 19720 23714
rect 19668 23650 19720 23656
rect 19760 23368 19812 23374
rect 19760 23310 19812 23316
rect 19208 23300 19524 23306
rect 19260 23294 19524 23300
rect 19576 23300 19628 23306
rect 19208 23242 19260 23248
rect 19576 23242 19628 23248
rect 19484 23232 19536 23238
rect 19482 23200 19484 23209
rect 19536 23200 19538 23209
rect 19482 23135 19538 23144
rect 19576 23164 19628 23170
rect 19576 23106 19628 23112
rect 19484 23096 19536 23102
rect 19484 23038 19536 23044
rect 19496 22626 19524 23038
rect 19588 22801 19616 23106
rect 19574 22792 19630 22801
rect 19574 22727 19630 22736
rect 19772 22694 19800 23310
rect 19864 22898 19892 23718
rect 19852 22892 19904 22898
rect 19852 22834 19904 22840
rect 19760 22688 19812 22694
rect 19760 22630 19812 22636
rect 19944 22688 19996 22694
rect 19944 22630 19996 22636
rect 19484 22620 19536 22626
rect 19484 22562 19536 22568
rect 19116 22452 19412 22472
rect 19172 22450 19196 22452
rect 19252 22450 19276 22452
rect 19332 22450 19356 22452
rect 19194 22398 19196 22450
rect 19258 22398 19270 22450
rect 19332 22398 19334 22450
rect 19172 22396 19196 22398
rect 19252 22396 19276 22398
rect 19332 22396 19356 22398
rect 19116 22376 19412 22396
rect 19024 22144 19076 22150
rect 19024 22086 19076 22092
rect 19772 21674 19800 22630
rect 19956 22286 19984 22630
rect 20140 22558 20168 23718
rect 20600 23374 20628 27594
rect 20956 27584 21008 27590
rect 20956 27526 21008 27532
rect 20968 27046 20996 27526
rect 21232 27108 21284 27114
rect 21232 27050 21284 27056
rect 20956 27040 21008 27046
rect 20956 26982 21008 26988
rect 20956 25952 21008 25958
rect 20956 25894 21008 25900
rect 20588 23368 20640 23374
rect 20588 23310 20640 23316
rect 20128 22552 20180 22558
rect 20128 22494 20180 22500
rect 20140 22286 20168 22494
rect 20600 22354 20628 23310
rect 20772 23300 20824 23306
rect 20772 23242 20824 23248
rect 20784 22762 20812 23242
rect 20772 22756 20824 22762
rect 20772 22698 20824 22704
rect 20968 22558 20996 25894
rect 21048 25068 21100 25074
rect 21048 25010 21100 25016
rect 21060 23442 21088 25010
rect 21244 24870 21272 27050
rect 21324 27040 21376 27046
rect 21324 26982 21376 26988
rect 21336 26094 21364 26982
rect 21324 26088 21376 26094
rect 21324 26030 21376 26036
rect 21336 24870 21364 26030
rect 21428 25482 21456 27662
rect 21520 27590 21548 28682
rect 21704 27658 21732 28750
rect 21888 28678 21916 29226
rect 21784 28672 21836 28678
rect 21784 28614 21836 28620
rect 21876 28672 21928 28678
rect 21876 28614 21928 28620
rect 21692 27652 21744 27658
rect 21692 27594 21744 27600
rect 21508 27584 21560 27590
rect 21508 27526 21560 27532
rect 21416 25476 21468 25482
rect 21416 25418 21468 25424
rect 21232 24864 21284 24870
rect 21232 24806 21284 24812
rect 21324 24864 21376 24870
rect 21324 24806 21376 24812
rect 21428 23782 21456 25418
rect 21520 24734 21548 27526
rect 21704 27454 21732 27594
rect 21692 27448 21744 27454
rect 21692 27390 21744 27396
rect 21704 26570 21732 27390
rect 21796 26978 21824 28614
rect 21784 26972 21836 26978
rect 21784 26914 21836 26920
rect 21968 26904 22020 26910
rect 21968 26846 22020 26852
rect 21692 26564 21744 26570
rect 21692 26506 21744 26512
rect 21600 25952 21652 25958
rect 21600 25894 21652 25900
rect 21612 25482 21640 25894
rect 21600 25476 21652 25482
rect 21600 25418 21652 25424
rect 21612 24938 21640 25418
rect 21600 24932 21652 24938
rect 21600 24874 21652 24880
rect 21508 24728 21560 24734
rect 21508 24670 21560 24676
rect 21416 23776 21468 23782
rect 21416 23718 21468 23724
rect 21428 23442 21456 23718
rect 21048 23436 21100 23442
rect 21048 23378 21100 23384
rect 21416 23436 21468 23442
rect 21416 23378 21468 23384
rect 21520 23238 21548 24670
rect 21980 23374 22008 26846
rect 21968 23368 22020 23374
rect 21968 23310 22020 23316
rect 21416 23232 21468 23238
rect 21416 23174 21468 23180
rect 21508 23232 21560 23238
rect 21508 23174 21560 23180
rect 21428 22626 21456 23174
rect 21520 22762 21548 23174
rect 21508 22756 21560 22762
rect 21508 22698 21560 22704
rect 21980 22694 22008 23310
rect 21968 22688 22020 22694
rect 21968 22630 22020 22636
rect 21140 22620 21192 22626
rect 21140 22562 21192 22568
rect 21416 22620 21468 22626
rect 21416 22562 21468 22568
rect 20956 22552 21008 22558
rect 20956 22494 21008 22500
rect 20588 22348 20640 22354
rect 20588 22290 20640 22296
rect 21152 22286 21180 22562
rect 21428 22354 21456 22562
rect 21508 22552 21560 22558
rect 21508 22494 21560 22500
rect 21520 22354 21548 22494
rect 21416 22348 21468 22354
rect 21416 22290 21468 22296
rect 21508 22348 21560 22354
rect 21508 22290 21560 22296
rect 19944 22280 19996 22286
rect 19944 22222 19996 22228
rect 20128 22280 20180 22286
rect 20128 22222 20180 22228
rect 21140 22280 21192 22286
rect 21140 22222 21192 22228
rect 20496 22144 20548 22150
rect 20496 22086 20548 22092
rect 19760 21668 19812 21674
rect 19760 21610 19812 21616
rect 20508 21606 20536 22086
rect 21428 21742 21456 22290
rect 21980 22014 22008 22630
rect 21968 22008 22020 22014
rect 21968 21950 22020 21956
rect 21416 21736 21468 21742
rect 21416 21678 21468 21684
rect 18104 21600 18156 21606
rect 18104 21542 18156 21548
rect 18288 21600 18340 21606
rect 18288 21542 18340 21548
rect 18840 21600 18892 21606
rect 18840 21542 18892 21548
rect 20496 21600 20548 21606
rect 20496 21542 20548 21548
rect 21416 21600 21468 21606
rect 21416 21542 21468 21548
rect 18116 21198 18144 21542
rect 19576 21464 19628 21470
rect 19576 21406 19628 21412
rect 19116 21364 19412 21384
rect 19172 21362 19196 21364
rect 19252 21362 19276 21364
rect 19332 21362 19356 21364
rect 19194 21310 19196 21362
rect 19258 21310 19270 21362
rect 19332 21310 19334 21362
rect 19172 21308 19196 21310
rect 19252 21308 19276 21310
rect 19332 21308 19356 21310
rect 19116 21288 19412 21308
rect 19588 21198 19616 21406
rect 20508 21266 20536 21542
rect 21428 21470 21456 21542
rect 21416 21464 21468 21470
rect 21416 21406 21468 21412
rect 20496 21260 20548 21266
rect 20496 21202 20548 21208
rect 18012 21192 18064 21198
rect 18012 21134 18064 21140
rect 18104 21192 18156 21198
rect 18104 21134 18156 21140
rect 19576 21192 19628 21198
rect 19576 21134 19628 21140
rect 17920 21124 17972 21130
rect 17920 21066 17972 21072
rect 17460 20920 17512 20926
rect 17460 20862 17512 20868
rect 17276 20444 17328 20450
rect 17276 20386 17328 20392
rect 17288 20042 17316 20386
rect 16540 20036 16592 20042
rect 16540 19978 16592 19984
rect 17276 20036 17328 20042
rect 17276 19978 17328 19984
rect 16552 19430 16580 19978
rect 17932 19974 17960 21066
rect 18024 21062 18052 21134
rect 19760 21124 19812 21130
rect 19760 21066 19812 21072
rect 21048 21124 21100 21130
rect 21048 21066 21100 21072
rect 18012 21056 18064 21062
rect 18012 20998 18064 21004
rect 18380 21056 18432 21062
rect 18380 20998 18432 21004
rect 18024 20654 18052 20998
rect 18012 20648 18064 20654
rect 18012 20590 18064 20596
rect 18012 20512 18064 20518
rect 18012 20454 18064 20460
rect 17920 19968 17972 19974
rect 17920 19910 17972 19916
rect 17932 19634 17960 19910
rect 17920 19628 17972 19634
rect 17920 19570 17972 19576
rect 16540 19424 16592 19430
rect 16540 19366 16592 19372
rect 18024 19022 18052 20454
rect 18288 20444 18340 20450
rect 18288 20386 18340 20392
rect 18300 19906 18328 20386
rect 18288 19900 18340 19906
rect 18288 19842 18340 19848
rect 18012 19016 18064 19022
rect 18012 18958 18064 18964
rect 18024 18546 18052 18958
rect 18392 18954 18420 20998
rect 19024 20376 19076 20382
rect 19024 20318 19076 20324
rect 19036 20110 19064 20318
rect 19116 20276 19412 20296
rect 19172 20274 19196 20276
rect 19252 20274 19276 20276
rect 19332 20274 19356 20276
rect 19194 20222 19196 20274
rect 19258 20222 19270 20274
rect 19332 20222 19334 20274
rect 19172 20220 19196 20222
rect 19252 20220 19276 20222
rect 19332 20220 19356 20222
rect 19116 20200 19412 20220
rect 19024 20104 19076 20110
rect 19024 20046 19076 20052
rect 18564 20036 18616 20042
rect 18564 19978 18616 19984
rect 18576 19634 18604 19978
rect 18564 19628 18616 19634
rect 18564 19570 18616 19576
rect 19036 19430 19064 20046
rect 19024 19424 19076 19430
rect 19024 19366 19076 19372
rect 19576 19424 19628 19430
rect 19576 19366 19628 19372
rect 19116 19188 19412 19208
rect 19172 19186 19196 19188
rect 19252 19186 19276 19188
rect 19332 19186 19356 19188
rect 19194 19134 19196 19186
rect 19258 19134 19270 19186
rect 19332 19134 19334 19186
rect 19172 19132 19196 19134
rect 19252 19132 19276 19134
rect 19332 19132 19356 19134
rect 19116 19112 19412 19132
rect 18380 18948 18432 18954
rect 18380 18890 18432 18896
rect 18288 18812 18340 18818
rect 18288 18754 18340 18760
rect 18012 18540 18064 18546
rect 18012 18482 18064 18488
rect 16908 18268 16960 18274
rect 16908 18210 16960 18216
rect 18012 18268 18064 18274
rect 18012 18210 18064 18216
rect 16724 17248 16776 17254
rect 16724 17190 16776 17196
rect 16736 16846 16764 17190
rect 16724 16840 16776 16846
rect 16724 16782 16776 16788
rect 16724 15480 16776 15486
rect 16724 15422 16776 15428
rect 16736 14602 16764 15422
rect 16920 14942 16948 18210
rect 17920 17792 17972 17798
rect 17920 17734 17972 17740
rect 17368 17452 17420 17458
rect 17368 17394 17420 17400
rect 17380 17254 17408 17394
rect 17932 17254 17960 17734
rect 18024 17458 18052 18210
rect 18012 17452 18064 17458
rect 18012 17394 18064 17400
rect 17368 17248 17420 17254
rect 17368 17190 17420 17196
rect 17920 17248 17972 17254
rect 17920 17190 17972 17196
rect 17380 15690 17408 17190
rect 17932 16778 17960 17190
rect 18196 17180 18248 17186
rect 18196 17122 18248 17128
rect 18208 16778 18236 17122
rect 17920 16772 17972 16778
rect 17920 16714 17972 16720
rect 18196 16772 18248 16778
rect 18196 16714 18248 16720
rect 17932 16166 17960 16714
rect 18208 16302 18236 16714
rect 18196 16296 18248 16302
rect 18196 16238 18248 16244
rect 17920 16160 17972 16166
rect 17920 16102 17972 16108
rect 18196 16160 18248 16166
rect 18196 16102 18248 16108
rect 17460 16092 17512 16098
rect 17460 16034 17512 16040
rect 17368 15684 17420 15690
rect 17368 15626 17420 15632
rect 17472 15010 17500 16034
rect 17460 15004 17512 15010
rect 17460 14946 17512 14952
rect 16908 14936 16960 14942
rect 16908 14878 16960 14884
rect 16920 14670 16948 14878
rect 16908 14664 16960 14670
rect 16960 14612 17132 14618
rect 16908 14606 17132 14612
rect 16724 14596 16776 14602
rect 16920 14590 17132 14606
rect 16724 14538 16776 14544
rect 16172 14052 16224 14058
rect 16172 13994 16224 14000
rect 14148 13508 14200 13514
rect 14148 13450 14200 13456
rect 14608 13508 14660 13514
rect 14608 13450 14660 13456
rect 14700 13508 14752 13514
rect 14700 13450 14752 13456
rect 15068 13508 15120 13514
rect 15068 13450 15120 13456
rect 14620 13310 14648 13450
rect 14608 13304 14660 13310
rect 14608 13246 14660 13252
rect 14116 13204 14412 13224
rect 14172 13202 14196 13204
rect 14252 13202 14276 13204
rect 14332 13202 14356 13204
rect 14194 13150 14196 13202
rect 14258 13150 14270 13202
rect 14332 13150 14334 13202
rect 14172 13148 14196 13150
rect 14252 13148 14276 13150
rect 14332 13148 14356 13150
rect 14116 13128 14412 13148
rect 14620 13106 14648 13246
rect 14608 13100 14660 13106
rect 14608 13042 14660 13048
rect 13504 13032 13556 13038
rect 13504 12974 13556 12980
rect 14240 12964 14292 12970
rect 14240 12906 14292 12912
rect 13136 12896 13188 12902
rect 13136 12838 13188 12844
rect 13412 12896 13464 12902
rect 13412 12838 13464 12844
rect 13424 12562 13452 12838
rect 13412 12556 13464 12562
rect 13412 12498 13464 12504
rect 14252 12358 14280 12906
rect 14332 12896 14384 12902
rect 14332 12838 14384 12844
rect 14976 12896 15028 12902
rect 14976 12838 15028 12844
rect 14344 12426 14372 12838
rect 14884 12556 14936 12562
rect 14884 12498 14936 12504
rect 14332 12420 14384 12426
rect 14332 12362 14384 12368
rect 14424 12420 14476 12426
rect 14424 12362 14476 12368
rect 13044 12352 13096 12358
rect 13044 12294 13096 12300
rect 14240 12352 14292 12358
rect 14240 12294 14292 12300
rect 12676 12216 12728 12222
rect 14436 12204 14464 12362
rect 14436 12176 14556 12204
rect 12676 12158 12728 12164
rect 12688 9624 12716 12158
rect 14116 12116 14412 12136
rect 14172 12114 14196 12116
rect 14252 12114 14276 12116
rect 14332 12114 14356 12116
rect 14194 12062 14196 12114
rect 14258 12062 14270 12114
rect 14332 12062 14334 12114
rect 14172 12060 14196 12062
rect 14252 12060 14276 12062
rect 14332 12060 14356 12062
rect 14116 12040 14412 12060
rect 14528 12018 14556 12176
rect 14516 12012 14568 12018
rect 14516 11954 14568 11960
rect 14528 11338 14556 11954
rect 14516 11332 14568 11338
rect 14516 11274 14568 11280
rect 14116 11028 14412 11048
rect 14172 11026 14196 11028
rect 14252 11026 14276 11028
rect 14332 11026 14356 11028
rect 14194 10974 14196 11026
rect 14258 10974 14270 11026
rect 14332 10974 14334 11026
rect 14172 10972 14196 10974
rect 14252 10972 14276 10974
rect 14332 10972 14356 10974
rect 14116 10952 14412 10972
rect 14896 9624 14924 12498
rect 14988 11474 15016 12838
rect 15080 12494 15108 13450
rect 15436 12896 15488 12902
rect 15436 12838 15488 12844
rect 15068 12488 15120 12494
rect 15068 12430 15120 12436
rect 15448 12426 15476 12838
rect 15528 12760 15580 12766
rect 15528 12702 15580 12708
rect 15436 12420 15488 12426
rect 15436 12362 15488 12368
rect 15540 12222 15568 12702
rect 16264 12420 16316 12426
rect 16264 12362 16316 12368
rect 15528 12216 15580 12222
rect 15528 12158 15580 12164
rect 15712 12216 15764 12222
rect 15712 12158 15764 12164
rect 15724 11882 15752 12158
rect 16276 12018 16304 12362
rect 16736 12358 16764 14538
rect 17000 14528 17052 14534
rect 17000 14470 17052 14476
rect 17012 14194 17040 14470
rect 17000 14188 17052 14194
rect 17000 14130 17052 14136
rect 16908 13440 16960 13446
rect 16908 13382 16960 13388
rect 16920 12494 16948 13382
rect 16908 12488 16960 12494
rect 16908 12430 16960 12436
rect 16724 12352 16776 12358
rect 16724 12294 16776 12300
rect 16264 12012 16316 12018
rect 16264 11954 16316 11960
rect 16736 11882 16764 12294
rect 15712 11876 15764 11882
rect 15712 11818 15764 11824
rect 16724 11876 16776 11882
rect 16724 11818 16776 11824
rect 16080 11740 16132 11746
rect 16080 11682 16132 11688
rect 16092 11474 16120 11682
rect 16736 11678 16764 11818
rect 16724 11672 16776 11678
rect 16724 11614 16776 11620
rect 14976 11468 15028 11474
rect 14976 11410 15028 11416
rect 16080 11468 16132 11474
rect 16080 11410 16132 11416
rect 17104 11338 17132 14590
rect 17472 14058 17500 14946
rect 18104 14936 18156 14942
rect 18104 14878 18156 14884
rect 18116 14602 18144 14878
rect 18104 14596 18156 14602
rect 18104 14538 18156 14544
rect 18208 14058 18236 16102
rect 18300 15214 18328 18754
rect 18380 18404 18432 18410
rect 18380 18346 18432 18352
rect 18392 17866 18420 18346
rect 19588 18206 19616 19366
rect 19772 19362 19800 21066
rect 19944 20444 19996 20450
rect 19944 20386 19996 20392
rect 19956 19634 19984 20386
rect 19944 19628 19996 19634
rect 19944 19570 19996 19576
rect 19760 19356 19812 19362
rect 19760 19298 19812 19304
rect 19772 19022 19800 19298
rect 19760 19016 19812 19022
rect 19760 18958 19812 18964
rect 20956 18880 21008 18886
rect 20956 18822 21008 18828
rect 20968 18546 20996 18822
rect 20956 18540 21008 18546
rect 20956 18482 21008 18488
rect 20864 18404 20916 18410
rect 20864 18346 20916 18352
rect 19668 18268 19720 18274
rect 19668 18210 19720 18216
rect 19852 18268 19904 18274
rect 19852 18210 19904 18216
rect 19576 18200 19628 18206
rect 19576 18142 19628 18148
rect 19116 18100 19412 18120
rect 19172 18098 19196 18100
rect 19252 18098 19276 18100
rect 19332 18098 19356 18100
rect 19194 18046 19196 18098
rect 19258 18046 19270 18098
rect 19332 18046 19334 18098
rect 19172 18044 19196 18046
rect 19252 18044 19276 18046
rect 19332 18044 19356 18046
rect 19116 18024 19412 18044
rect 19588 17934 19616 18142
rect 19680 18002 19708 18210
rect 19668 17996 19720 18002
rect 19668 17938 19720 17944
rect 19576 17928 19628 17934
rect 19576 17870 19628 17876
rect 18380 17860 18432 17866
rect 18380 17802 18432 17808
rect 18392 16642 18420 17802
rect 18748 17792 18800 17798
rect 18748 17734 18800 17740
rect 18760 16846 18788 17734
rect 19484 17248 19536 17254
rect 19484 17190 19536 17196
rect 19024 17180 19076 17186
rect 19024 17122 19076 17128
rect 18748 16840 18800 16846
rect 18748 16782 18800 16788
rect 18472 16772 18524 16778
rect 18472 16714 18524 16720
rect 18380 16636 18432 16642
rect 18380 16578 18432 16584
rect 18392 15622 18420 16578
rect 18484 16030 18512 16714
rect 18472 16024 18524 16030
rect 18472 15966 18524 15972
rect 18484 15690 18512 15966
rect 18760 15826 18788 16782
rect 18932 16228 18984 16234
rect 18932 16170 18984 16176
rect 18840 16024 18892 16030
rect 18840 15966 18892 15972
rect 18748 15820 18800 15826
rect 18748 15762 18800 15768
rect 18472 15684 18524 15690
rect 18472 15626 18524 15632
rect 18564 15684 18616 15690
rect 18564 15626 18616 15632
rect 18380 15616 18432 15622
rect 18380 15558 18432 15564
rect 18288 15208 18340 15214
rect 18288 15150 18340 15156
rect 18484 15146 18512 15626
rect 18576 15214 18604 15626
rect 18564 15208 18616 15214
rect 18564 15150 18616 15156
rect 18472 15140 18524 15146
rect 18472 15082 18524 15088
rect 18484 14602 18512 15082
rect 18472 14596 18524 14602
rect 18472 14538 18524 14544
rect 17460 14052 17512 14058
rect 17460 13994 17512 14000
rect 18196 14052 18248 14058
rect 18196 13994 18248 14000
rect 17828 13984 17880 13990
rect 17828 13926 17880 13932
rect 18288 13984 18340 13990
rect 18288 13926 18340 13932
rect 17552 13508 17604 13514
rect 17552 13450 17604 13456
rect 17564 12834 17592 13450
rect 17840 13378 17868 13926
rect 18300 13582 18328 13926
rect 18656 13916 18708 13922
rect 18760 13904 18788 15762
rect 18852 15078 18880 15966
rect 18944 15758 18972 16170
rect 19036 16166 19064 17122
rect 19116 17012 19412 17032
rect 19172 17010 19196 17012
rect 19252 17010 19276 17012
rect 19332 17010 19356 17012
rect 19194 16958 19196 17010
rect 19258 16958 19270 17010
rect 19332 16958 19334 17010
rect 19172 16956 19196 16958
rect 19252 16956 19276 16958
rect 19332 16956 19356 16958
rect 19116 16936 19412 16956
rect 19024 16160 19076 16166
rect 19024 16102 19076 16108
rect 19116 15924 19412 15944
rect 19172 15922 19196 15924
rect 19252 15922 19276 15924
rect 19332 15922 19356 15924
rect 19194 15870 19196 15922
rect 19258 15870 19270 15922
rect 19332 15870 19334 15922
rect 19172 15868 19196 15870
rect 19252 15868 19276 15870
rect 19332 15868 19356 15870
rect 19116 15848 19412 15868
rect 18932 15752 18984 15758
rect 18932 15694 18984 15700
rect 18840 15072 18892 15078
rect 18840 15014 18892 15020
rect 18944 13990 18972 15694
rect 19496 15078 19524 17190
rect 19588 16166 19616 17870
rect 19864 17866 19892 18210
rect 20876 18206 20904 18346
rect 20864 18200 20916 18206
rect 20864 18142 20916 18148
rect 20876 17934 20904 18142
rect 20864 17928 20916 17934
rect 20864 17870 20916 17876
rect 19852 17860 19904 17866
rect 19852 17802 19904 17808
rect 19668 17180 19720 17186
rect 19668 17122 19720 17128
rect 19680 16846 19708 17122
rect 19668 16840 19720 16846
rect 19668 16782 19720 16788
rect 19576 16160 19628 16166
rect 19576 16102 19628 16108
rect 19864 16098 19892 17802
rect 20772 17384 20824 17390
rect 20772 17326 20824 17332
rect 20784 16778 20812 17326
rect 20772 16772 20824 16778
rect 20772 16714 20824 16720
rect 20784 16302 20812 16714
rect 21060 16574 21088 21066
rect 21428 20994 21456 21406
rect 21600 21056 21652 21062
rect 21600 20998 21652 21004
rect 21416 20988 21468 20994
rect 21416 20930 21468 20936
rect 21428 20586 21456 20930
rect 21416 20580 21468 20586
rect 21416 20522 21468 20528
rect 21612 20518 21640 20998
rect 22072 20738 22100 35670
rect 23624 34180 23676 34186
rect 23624 34122 23676 34128
rect 23440 33976 23492 33982
rect 23440 33918 23492 33924
rect 22428 33568 22480 33574
rect 22428 33510 22480 33516
rect 22244 32616 22296 32622
rect 22244 32558 22296 32564
rect 22256 32010 22284 32558
rect 22244 32004 22296 32010
rect 22244 31946 22296 31952
rect 22256 30922 22284 31946
rect 22440 31058 22468 33510
rect 22520 33500 22572 33506
rect 22520 33442 22572 33448
rect 22532 33166 22560 33442
rect 22520 33160 22572 33166
rect 22520 33102 22572 33108
rect 23072 32956 23124 32962
rect 23072 32898 23124 32904
rect 22888 32480 22940 32486
rect 22888 32422 22940 32428
rect 22428 31052 22480 31058
rect 22428 30994 22480 31000
rect 22900 30990 22928 32422
rect 23084 32078 23112 32898
rect 23072 32072 23124 32078
rect 23072 32014 23124 32020
rect 23452 31466 23480 33918
rect 23532 33568 23584 33574
rect 23532 33510 23584 33516
rect 23544 32622 23572 33510
rect 23636 33098 23664 34122
rect 24116 33876 24412 33896
rect 24172 33874 24196 33876
rect 24252 33874 24276 33876
rect 24332 33874 24356 33876
rect 24194 33822 24196 33874
rect 24258 33822 24270 33874
rect 24332 33822 24334 33874
rect 24172 33820 24196 33822
rect 24252 33820 24276 33822
rect 24332 33820 24356 33822
rect 24116 33800 24412 33820
rect 24176 33568 24228 33574
rect 24176 33510 24228 33516
rect 24188 33098 24216 33510
rect 24452 33228 24504 33234
rect 24452 33170 24504 33176
rect 23624 33092 23676 33098
rect 23624 33034 23676 33040
rect 24176 33092 24228 33098
rect 24176 33034 24228 33040
rect 23532 32616 23584 32622
rect 23532 32558 23584 32564
rect 23636 32010 23664 33034
rect 23716 33024 23768 33030
rect 23716 32966 23768 32972
rect 23532 32004 23584 32010
rect 23532 31946 23584 31952
rect 23624 32004 23676 32010
rect 23624 31946 23676 31952
rect 23348 31460 23400 31466
rect 23348 31402 23400 31408
rect 23440 31460 23492 31466
rect 23440 31402 23492 31408
rect 22888 30984 22940 30990
rect 22888 30926 22940 30932
rect 22244 30916 22296 30922
rect 22244 30858 22296 30864
rect 22520 30916 22572 30922
rect 22520 30858 22572 30864
rect 23256 30916 23308 30922
rect 23256 30858 23308 30864
rect 22428 30848 22480 30854
rect 22428 30790 22480 30796
rect 22336 30236 22388 30242
rect 22336 30178 22388 30184
rect 22244 30168 22296 30174
rect 22244 30110 22296 30116
rect 22256 29834 22284 30110
rect 22244 29828 22296 29834
rect 22244 29770 22296 29776
rect 22348 29766 22376 30178
rect 22336 29760 22388 29766
rect 22336 29702 22388 29708
rect 22440 28338 22468 30790
rect 22532 29902 22560 30858
rect 23072 30236 23124 30242
rect 23072 30178 23124 30184
rect 22612 30168 22664 30174
rect 22980 30168 23032 30174
rect 22664 30128 22744 30156
rect 22612 30110 22664 30116
rect 22716 29902 22744 30128
rect 22980 30110 23032 30116
rect 22520 29896 22572 29902
rect 22520 29838 22572 29844
rect 22704 29896 22756 29902
rect 22704 29838 22756 29844
rect 22716 29222 22744 29838
rect 22888 29760 22940 29766
rect 22888 29702 22940 29708
rect 22704 29216 22756 29222
rect 22704 29158 22756 29164
rect 22716 29086 22744 29158
rect 22900 29154 22928 29702
rect 22888 29148 22940 29154
rect 22888 29090 22940 29096
rect 22704 29080 22756 29086
rect 22704 29022 22756 29028
rect 22716 28746 22744 29022
rect 22900 28814 22928 29090
rect 22992 28814 23020 30110
rect 23084 29970 23112 30178
rect 23072 29964 23124 29970
rect 23072 29906 23124 29912
rect 23268 29902 23296 30858
rect 23360 30854 23388 31402
rect 23544 31330 23572 31946
rect 23728 31602 23756 32966
rect 24116 32788 24412 32808
rect 24172 32786 24196 32788
rect 24252 32786 24276 32788
rect 24332 32786 24356 32788
rect 24194 32734 24196 32786
rect 24258 32734 24270 32786
rect 24332 32734 24334 32786
rect 24172 32732 24196 32734
rect 24252 32732 24276 32734
rect 24332 32732 24356 32734
rect 24116 32712 24412 32732
rect 23808 31936 23860 31942
rect 23808 31878 23860 31884
rect 23716 31596 23768 31602
rect 23716 31538 23768 31544
rect 23820 31398 23848 31878
rect 24116 31700 24412 31720
rect 24172 31698 24196 31700
rect 24252 31698 24276 31700
rect 24332 31698 24356 31700
rect 24194 31646 24196 31698
rect 24258 31646 24270 31698
rect 24332 31646 24334 31698
rect 24172 31644 24196 31646
rect 24252 31644 24276 31646
rect 24332 31644 24356 31646
rect 24116 31624 24412 31644
rect 23808 31392 23860 31398
rect 23808 31334 23860 31340
rect 23532 31324 23584 31330
rect 23532 31266 23584 31272
rect 23348 30848 23400 30854
rect 23348 30790 23400 30796
rect 23256 29896 23308 29902
rect 23256 29838 23308 29844
rect 23348 29828 23400 29834
rect 23348 29770 23400 29776
rect 23360 29154 23388 29770
rect 23348 29148 23400 29154
rect 23348 29090 23400 29096
rect 23716 29148 23768 29154
rect 23716 29090 23768 29096
rect 23164 29080 23216 29086
rect 23164 29022 23216 29028
rect 23176 28882 23204 29022
rect 23164 28876 23216 28882
rect 23164 28818 23216 28824
rect 22888 28808 22940 28814
rect 22888 28750 22940 28756
rect 22980 28808 23032 28814
rect 22980 28750 23032 28756
rect 22612 28740 22664 28746
rect 22612 28682 22664 28688
rect 22704 28740 22756 28746
rect 22704 28682 22756 28688
rect 22428 28332 22480 28338
rect 22428 28274 22480 28280
rect 22440 28218 22468 28274
rect 22256 28190 22468 28218
rect 22624 28202 22652 28682
rect 22612 28196 22664 28202
rect 22256 27946 22284 28190
rect 22612 28138 22664 28144
rect 22336 28128 22388 28134
rect 22388 28088 22468 28116
rect 22336 28070 22388 28076
rect 22256 27918 22376 27946
rect 22244 26564 22296 26570
rect 22244 26506 22296 26512
rect 22256 22218 22284 26506
rect 22348 25890 22376 27918
rect 22440 27250 22468 28088
rect 22612 28060 22664 28066
rect 22612 28002 22664 28008
rect 22888 28060 22940 28066
rect 22888 28002 22940 28008
rect 22624 27726 22652 28002
rect 22612 27720 22664 27726
rect 22612 27662 22664 27668
rect 22796 27720 22848 27726
rect 22796 27662 22848 27668
rect 22808 27454 22836 27662
rect 22796 27448 22848 27454
rect 22796 27390 22848 27396
rect 22428 27244 22480 27250
rect 22428 27186 22480 27192
rect 22612 27040 22664 27046
rect 22612 26982 22664 26988
rect 22428 26972 22480 26978
rect 22428 26914 22480 26920
rect 22440 26638 22468 26914
rect 22624 26706 22652 26982
rect 22612 26700 22664 26706
rect 22612 26642 22664 26648
rect 22428 26632 22480 26638
rect 22428 26574 22480 26580
rect 22612 26428 22664 26434
rect 22612 26370 22664 26376
rect 22624 26162 22652 26370
rect 22612 26156 22664 26162
rect 22612 26098 22664 26104
rect 22704 26020 22756 26026
rect 22704 25962 22756 25968
rect 22336 25884 22388 25890
rect 22336 25826 22388 25832
rect 22716 25550 22744 25962
rect 22900 25550 22928 28002
rect 22992 26978 23020 28750
rect 23072 28604 23124 28610
rect 23072 28546 23124 28552
rect 23084 27726 23112 28546
rect 23360 28270 23388 29090
rect 23728 28814 23756 29090
rect 23716 28808 23768 28814
rect 23716 28750 23768 28756
rect 23348 28264 23400 28270
rect 23348 28206 23400 28212
rect 23348 28060 23400 28066
rect 23348 28002 23400 28008
rect 23072 27720 23124 27726
rect 23072 27662 23124 27668
rect 22980 26972 23032 26978
rect 22980 26914 23032 26920
rect 22704 25544 22756 25550
rect 22704 25486 22756 25492
rect 22888 25544 22940 25550
rect 22888 25486 22940 25492
rect 22704 25408 22756 25414
rect 22704 25350 22756 25356
rect 22612 25272 22664 25278
rect 22612 25214 22664 25220
rect 22336 24864 22388 24870
rect 22336 24806 22388 24812
rect 22518 24832 22574 24841
rect 22348 22898 22376 24806
rect 22518 24767 22574 24776
rect 22532 24734 22560 24767
rect 22520 24728 22572 24734
rect 22520 24670 22572 24676
rect 22624 24530 22652 25214
rect 22716 25006 22744 25350
rect 22704 25000 22756 25006
rect 22704 24942 22756 24948
rect 22992 24734 23020 26914
rect 23084 26638 23112 27662
rect 23256 27040 23308 27046
rect 23256 26982 23308 26988
rect 23072 26632 23124 26638
rect 23072 26574 23124 26580
rect 23084 25074 23112 26574
rect 23268 26366 23296 26982
rect 23360 26570 23388 28002
rect 23624 27992 23676 27998
rect 23624 27934 23676 27940
rect 23532 27584 23584 27590
rect 23532 27526 23584 27532
rect 23440 27244 23492 27250
rect 23440 27186 23492 27192
rect 23452 26978 23480 27186
rect 23440 26972 23492 26978
rect 23440 26914 23492 26920
rect 23348 26564 23400 26570
rect 23348 26506 23400 26512
rect 23256 26360 23308 26366
rect 23256 26302 23308 26308
rect 23072 25068 23124 25074
rect 23072 25010 23124 25016
rect 23084 24938 23112 25010
rect 23360 24954 23388 26506
rect 23452 25006 23480 26914
rect 23544 25482 23572 27526
rect 23636 26638 23664 27934
rect 23820 27266 23848 31334
rect 24084 31324 24136 31330
rect 24084 31266 24136 31272
rect 24096 30786 24124 31266
rect 24084 30780 24136 30786
rect 24084 30722 24136 30728
rect 23992 30712 24044 30718
rect 23992 30654 24044 30660
rect 24004 29834 24032 30654
rect 24116 30612 24412 30632
rect 24172 30610 24196 30612
rect 24252 30610 24276 30612
rect 24332 30610 24356 30612
rect 24194 30558 24196 30610
rect 24258 30558 24270 30610
rect 24332 30558 24334 30610
rect 24172 30556 24196 30558
rect 24252 30556 24276 30558
rect 24332 30556 24356 30558
rect 24116 30536 24412 30556
rect 24464 29970 24492 33170
rect 24648 32554 24676 35809
rect 26384 34180 26436 34186
rect 26384 34122 26436 34128
rect 25556 33976 25608 33982
rect 25556 33918 25608 33924
rect 25096 33636 25148 33642
rect 25096 33578 25148 33584
rect 25004 33568 25056 33574
rect 25004 33510 25056 33516
rect 24912 33092 24964 33098
rect 24912 33034 24964 33040
rect 24636 32548 24688 32554
rect 24636 32490 24688 32496
rect 24728 31868 24780 31874
rect 24728 31810 24780 31816
rect 24544 31324 24596 31330
rect 24544 31266 24596 31272
rect 24452 29964 24504 29970
rect 24452 29906 24504 29912
rect 23992 29828 24044 29834
rect 23992 29770 24044 29776
rect 24004 29426 24032 29770
rect 24556 29698 24584 31266
rect 24740 30174 24768 31810
rect 24728 30168 24780 30174
rect 24728 30110 24780 30116
rect 24636 29760 24688 29766
rect 24636 29702 24688 29708
rect 24544 29692 24596 29698
rect 24544 29634 24596 29640
rect 24116 29524 24412 29544
rect 24172 29522 24196 29524
rect 24252 29522 24276 29524
rect 24332 29522 24356 29524
rect 24194 29470 24196 29522
rect 24258 29470 24270 29522
rect 24332 29470 24334 29522
rect 24172 29468 24196 29470
rect 24252 29468 24276 29470
rect 24332 29468 24356 29470
rect 24116 29448 24412 29468
rect 23992 29420 24044 29426
rect 23992 29362 24044 29368
rect 24452 29216 24504 29222
rect 24452 29158 24504 29164
rect 23900 29148 23952 29154
rect 23900 29090 23952 29096
rect 23728 27238 23848 27266
rect 23624 26632 23676 26638
rect 23624 26574 23676 26580
rect 23532 25476 23584 25482
rect 23532 25418 23584 25424
rect 23072 24932 23124 24938
rect 23072 24874 23124 24880
rect 23268 24926 23388 24954
rect 23440 25000 23492 25006
rect 23440 24942 23492 24948
rect 23268 24802 23296 24926
rect 23452 24870 23480 24942
rect 23440 24864 23492 24870
rect 23440 24806 23492 24812
rect 23256 24796 23308 24802
rect 23256 24738 23308 24744
rect 23348 24796 23400 24802
rect 23348 24738 23400 24744
rect 22980 24728 23032 24734
rect 22980 24670 23032 24676
rect 22612 24524 22664 24530
rect 22612 24466 22664 24472
rect 22520 24388 22572 24394
rect 22520 24330 22572 24336
rect 22428 24320 22480 24326
rect 22428 24262 22480 24268
rect 22336 22892 22388 22898
rect 22336 22834 22388 22840
rect 22348 22218 22376 22834
rect 22440 22370 22468 24262
rect 22532 23374 22560 24330
rect 22520 23368 22572 23374
rect 22520 23310 22572 23316
rect 22624 23238 22652 24466
rect 22888 24388 22940 24394
rect 22888 24330 22940 24336
rect 22900 23782 22928 24330
rect 22992 23850 23020 24670
rect 23072 24184 23124 24190
rect 23072 24126 23124 24132
rect 22980 23844 23032 23850
rect 22980 23786 23032 23792
rect 22888 23776 22940 23782
rect 22888 23718 22940 23724
rect 22992 23442 23020 23786
rect 22980 23436 23032 23442
rect 22980 23378 23032 23384
rect 23084 23374 23112 24126
rect 23164 23708 23216 23714
rect 23164 23650 23216 23656
rect 23072 23368 23124 23374
rect 23072 23310 23124 23316
rect 23176 23306 23204 23650
rect 23164 23300 23216 23306
rect 23164 23242 23216 23248
rect 22612 23232 22664 23238
rect 22612 23174 22664 23180
rect 22704 22892 22756 22898
rect 22704 22834 22756 22840
rect 22716 22626 22744 22834
rect 23164 22756 23216 22762
rect 23164 22698 23216 22704
rect 22888 22688 22940 22694
rect 22888 22630 22940 22636
rect 22704 22620 22756 22626
rect 22704 22562 22756 22568
rect 22440 22342 22560 22370
rect 22716 22354 22744 22562
rect 22244 22212 22296 22218
rect 22244 22154 22296 22160
rect 22336 22212 22388 22218
rect 22336 22154 22388 22160
rect 22256 21742 22284 22154
rect 22336 22076 22388 22082
rect 22336 22018 22388 22024
rect 22428 22076 22480 22082
rect 22428 22018 22480 22024
rect 22244 21736 22296 21742
rect 22244 21678 22296 21684
rect 22348 21674 22376 22018
rect 22336 21668 22388 21674
rect 22336 21610 22388 21616
rect 22152 21600 22204 21606
rect 22152 21542 22204 21548
rect 22164 21130 22192 21542
rect 22440 21198 22468 22018
rect 22532 21962 22560 22342
rect 22704 22348 22756 22354
rect 22704 22290 22756 22296
rect 22532 21934 22652 21962
rect 22624 21266 22652 21934
rect 22716 21810 22744 22290
rect 22900 22218 22928 22630
rect 22980 22280 23032 22286
rect 22980 22222 23032 22228
rect 22888 22212 22940 22218
rect 22888 22154 22940 22160
rect 22704 21804 22756 21810
rect 22704 21746 22756 21752
rect 22900 21606 22928 22154
rect 22992 21742 23020 22222
rect 23176 22150 23204 22698
rect 23360 22694 23388 24738
rect 23452 24326 23480 24806
rect 23440 24320 23492 24326
rect 23440 24262 23492 24268
rect 23728 23730 23756 27238
rect 23808 27108 23860 27114
rect 23808 27050 23860 27056
rect 23820 25822 23848 27050
rect 23808 25816 23860 25822
rect 23808 25758 23860 25764
rect 23912 25074 23940 29090
rect 24464 28882 24492 29158
rect 24452 28876 24504 28882
rect 24452 28818 24504 28824
rect 24452 28672 24504 28678
rect 24452 28614 24504 28620
rect 24116 28436 24412 28456
rect 24172 28434 24196 28436
rect 24252 28434 24276 28436
rect 24332 28434 24356 28436
rect 24194 28382 24196 28434
rect 24258 28382 24270 28434
rect 24332 28382 24334 28434
rect 24172 28380 24196 28382
rect 24252 28380 24276 28382
rect 24332 28380 24356 28382
rect 24116 28360 24412 28380
rect 24464 27658 24492 28614
rect 24544 27720 24596 27726
rect 24544 27662 24596 27668
rect 24452 27652 24504 27658
rect 24452 27594 24504 27600
rect 24116 27348 24412 27368
rect 24172 27346 24196 27348
rect 24252 27346 24276 27348
rect 24332 27346 24356 27348
rect 24194 27294 24196 27346
rect 24258 27294 24270 27346
rect 24332 27294 24334 27346
rect 24172 27292 24196 27294
rect 24252 27292 24276 27294
rect 24332 27292 24356 27294
rect 24116 27272 24412 27292
rect 23992 26428 24044 26434
rect 23992 26370 24044 26376
rect 24004 26162 24032 26370
rect 24116 26260 24412 26280
rect 24172 26258 24196 26260
rect 24252 26258 24276 26260
rect 24332 26258 24356 26260
rect 24194 26206 24196 26258
rect 24258 26206 24270 26258
rect 24332 26206 24334 26258
rect 24172 26204 24196 26206
rect 24252 26204 24276 26206
rect 24332 26204 24356 26206
rect 24116 26184 24412 26204
rect 23992 26156 24044 26162
rect 23992 26098 24044 26104
rect 24556 25958 24584 27662
rect 24544 25952 24596 25958
rect 24544 25894 24596 25900
rect 24084 25884 24136 25890
rect 24004 25844 24084 25872
rect 23900 25068 23952 25074
rect 23900 25010 23952 25016
rect 23808 24388 23860 24394
rect 23808 24330 23860 24336
rect 23820 23850 23848 24330
rect 23808 23844 23860 23850
rect 23808 23786 23860 23792
rect 23728 23702 23848 23730
rect 23716 23640 23768 23646
rect 23716 23582 23768 23588
rect 23624 23096 23676 23102
rect 23624 23038 23676 23044
rect 23636 22694 23664 23038
rect 23348 22688 23400 22694
rect 23348 22630 23400 22636
rect 23624 22688 23676 22694
rect 23624 22630 23676 22636
rect 23164 22144 23216 22150
rect 23164 22086 23216 22092
rect 22980 21736 23032 21742
rect 22980 21678 23032 21684
rect 23176 21606 23204 22086
rect 22888 21600 22940 21606
rect 22888 21542 22940 21548
rect 23164 21600 23216 21606
rect 23164 21542 23216 21548
rect 22612 21260 22664 21266
rect 22612 21202 22664 21208
rect 22428 21192 22480 21198
rect 22428 21134 22480 21140
rect 23360 21130 23388 22630
rect 22152 21124 22204 21130
rect 22152 21066 22204 21072
rect 23348 21124 23400 21130
rect 23348 21066 23400 21072
rect 22072 20722 22192 20738
rect 22072 20716 22204 20722
rect 22072 20710 22152 20716
rect 22152 20658 22204 20664
rect 21140 20512 21192 20518
rect 21140 20454 21192 20460
rect 21600 20512 21652 20518
rect 21600 20454 21652 20460
rect 21048 16568 21100 16574
rect 21048 16510 21100 16516
rect 21152 16386 21180 20454
rect 21416 20444 21468 20450
rect 21416 20386 21468 20392
rect 21428 20042 21456 20386
rect 22164 20042 22192 20658
rect 23728 20586 23756 23582
rect 23820 22778 23848 23702
rect 23912 23306 23940 25010
rect 24004 24394 24032 25844
rect 24084 25826 24136 25832
rect 24648 25414 24676 29702
rect 24636 25408 24688 25414
rect 24636 25350 24688 25356
rect 24116 25172 24412 25192
rect 24172 25170 24196 25172
rect 24252 25170 24276 25172
rect 24332 25170 24356 25172
rect 24194 25118 24196 25170
rect 24258 25118 24270 25170
rect 24332 25118 24334 25170
rect 24172 25116 24196 25118
rect 24252 25116 24276 25118
rect 24332 25116 24356 25118
rect 24116 25096 24412 25116
rect 24360 24728 24412 24734
rect 24360 24670 24412 24676
rect 24372 24394 24400 24670
rect 23992 24388 24044 24394
rect 23992 24330 24044 24336
rect 24360 24388 24412 24394
rect 24360 24330 24412 24336
rect 24116 24084 24412 24104
rect 24172 24082 24196 24084
rect 24252 24082 24276 24084
rect 24332 24082 24356 24084
rect 24194 24030 24196 24082
rect 24258 24030 24270 24082
rect 24332 24030 24334 24082
rect 24172 24028 24196 24030
rect 24252 24028 24276 24030
rect 24332 24028 24356 24030
rect 24116 24008 24412 24028
rect 24648 23782 24676 25350
rect 23992 23776 24044 23782
rect 23992 23718 24044 23724
rect 24636 23776 24688 23782
rect 24636 23718 24688 23724
rect 23900 23300 23952 23306
rect 23900 23242 23952 23248
rect 24004 23170 24032 23718
rect 23992 23164 24044 23170
rect 23992 23106 24044 23112
rect 23820 22750 23940 22778
rect 24004 22762 24032 23106
rect 24116 22996 24412 23016
rect 24172 22994 24196 22996
rect 24252 22994 24276 22996
rect 24332 22994 24356 22996
rect 24194 22942 24196 22994
rect 24258 22942 24270 22994
rect 24332 22942 24334 22994
rect 24172 22940 24196 22942
rect 24252 22940 24276 22942
rect 24332 22940 24356 22942
rect 24116 22920 24412 22940
rect 23808 22552 23860 22558
rect 23808 22494 23860 22500
rect 23820 21130 23848 22494
rect 23912 21606 23940 22750
rect 23992 22756 24044 22762
rect 23992 22698 24044 22704
rect 24004 22150 24032 22698
rect 24452 22620 24504 22626
rect 24452 22562 24504 22568
rect 23992 22144 24044 22150
rect 23992 22086 24044 22092
rect 24116 21908 24412 21928
rect 24172 21906 24196 21908
rect 24252 21906 24276 21908
rect 24332 21906 24356 21908
rect 24194 21854 24196 21906
rect 24258 21854 24270 21906
rect 24332 21854 24334 21906
rect 24172 21852 24196 21854
rect 24252 21852 24276 21854
rect 24332 21852 24356 21854
rect 24116 21832 24412 21852
rect 24464 21674 24492 22562
rect 24648 22286 24676 23718
rect 24636 22280 24688 22286
rect 24636 22222 24688 22228
rect 24452 21668 24504 21674
rect 24452 21610 24504 21616
rect 23900 21600 23952 21606
rect 23900 21542 23952 21548
rect 24636 21600 24688 21606
rect 24636 21542 24688 21548
rect 24648 21470 24676 21542
rect 24636 21464 24688 21470
rect 24636 21406 24688 21412
rect 23808 21124 23860 21130
rect 23808 21066 23860 21072
rect 23992 20920 24044 20926
rect 23992 20862 24044 20868
rect 23716 20580 23768 20586
rect 23716 20522 23768 20528
rect 24004 20518 24032 20862
rect 24116 20820 24412 20840
rect 24172 20818 24196 20820
rect 24252 20818 24276 20820
rect 24332 20818 24356 20820
rect 24194 20766 24196 20818
rect 24258 20766 24270 20818
rect 24332 20766 24334 20818
rect 24172 20764 24196 20766
rect 24252 20764 24276 20766
rect 24332 20764 24356 20766
rect 24116 20744 24412 20764
rect 24648 20654 24676 21406
rect 24636 20648 24688 20654
rect 24636 20590 24688 20596
rect 24740 20586 24768 30110
rect 24820 27788 24872 27794
rect 24820 27730 24872 27736
rect 24832 24394 24860 27730
rect 24820 24388 24872 24394
rect 24820 24330 24872 24336
rect 24924 23102 24952 33034
rect 25016 32622 25044 33510
rect 25004 32616 25056 32622
rect 25004 32558 25056 32564
rect 25108 32010 25136 33578
rect 25188 33024 25240 33030
rect 25188 32966 25240 32972
rect 25200 32486 25228 32966
rect 25464 32956 25516 32962
rect 25464 32898 25516 32904
rect 25476 32622 25504 32898
rect 25464 32616 25516 32622
rect 25464 32558 25516 32564
rect 25188 32480 25240 32486
rect 25188 32422 25240 32428
rect 25476 32078 25504 32558
rect 25568 32078 25596 33918
rect 26396 33658 26424 34122
rect 26396 33630 26516 33658
rect 26488 33506 26516 33630
rect 26200 33500 26252 33506
rect 26200 33442 26252 33448
rect 26476 33500 26528 33506
rect 26476 33442 26528 33448
rect 25924 32548 25976 32554
rect 25924 32490 25976 32496
rect 25936 32078 25964 32490
rect 25464 32072 25516 32078
rect 25464 32014 25516 32020
rect 25556 32072 25608 32078
rect 25556 32014 25608 32020
rect 25924 32072 25976 32078
rect 25924 32014 25976 32020
rect 25096 32004 25148 32010
rect 25096 31946 25148 31952
rect 25464 31392 25516 31398
rect 25464 31334 25516 31340
rect 25372 30848 25424 30854
rect 25372 30790 25424 30796
rect 25096 30304 25148 30310
rect 25096 30246 25148 30252
rect 25108 29970 25136 30246
rect 25096 29964 25148 29970
rect 25096 29906 25148 29912
rect 25108 29222 25136 29906
rect 25280 29896 25332 29902
rect 25280 29838 25332 29844
rect 25188 29828 25240 29834
rect 25188 29770 25240 29776
rect 25096 29216 25148 29222
rect 25096 29158 25148 29164
rect 25096 29080 25148 29086
rect 25096 29022 25148 29028
rect 25108 28746 25136 29022
rect 25096 28740 25148 28746
rect 25096 28682 25148 28688
rect 25108 28202 25136 28682
rect 25096 28196 25148 28202
rect 25096 28138 25148 28144
rect 25004 27992 25056 27998
rect 25004 27934 25056 27940
rect 25016 26706 25044 27934
rect 25004 26700 25056 26706
rect 25004 26642 25056 26648
rect 25016 23782 25044 26642
rect 25108 24530 25136 28138
rect 25200 26026 25228 29770
rect 25188 26020 25240 26026
rect 25188 25962 25240 25968
rect 25292 25822 25320 29838
rect 25384 27658 25412 30790
rect 25476 29834 25504 31334
rect 25936 30904 25964 32014
rect 26212 32010 26240 33442
rect 26292 33092 26344 33098
rect 26292 33034 26344 33040
rect 26304 32486 26332 33034
rect 26292 32480 26344 32486
rect 26292 32422 26344 32428
rect 26200 32004 26252 32010
rect 26200 31946 26252 31952
rect 25752 30876 25964 30904
rect 25464 29828 25516 29834
rect 25464 29770 25516 29776
rect 25464 29216 25516 29222
rect 25464 29158 25516 29164
rect 25476 28882 25504 29158
rect 25556 29148 25608 29154
rect 25556 29090 25608 29096
rect 25464 28876 25516 28882
rect 25464 28818 25516 28824
rect 25476 28134 25504 28818
rect 25464 28128 25516 28134
rect 25464 28070 25516 28076
rect 25568 27658 25596 29090
rect 25648 27992 25700 27998
rect 25648 27934 25700 27940
rect 25372 27652 25424 27658
rect 25372 27594 25424 27600
rect 25556 27652 25608 27658
rect 25556 27594 25608 27600
rect 25384 27454 25412 27594
rect 25660 27590 25688 27934
rect 25648 27584 25700 27590
rect 25648 27526 25700 27532
rect 25372 27448 25424 27454
rect 25372 27390 25424 27396
rect 25464 27244 25516 27250
rect 25464 27186 25516 27192
rect 25476 26162 25504 27186
rect 25648 26972 25700 26978
rect 25648 26914 25700 26920
rect 25660 26366 25688 26914
rect 25648 26360 25700 26366
rect 25648 26302 25700 26308
rect 25464 26156 25516 26162
rect 25464 26098 25516 26104
rect 25556 26088 25608 26094
rect 25556 26030 25608 26036
rect 25280 25816 25332 25822
rect 25280 25758 25332 25764
rect 25292 25550 25320 25758
rect 25280 25544 25332 25550
rect 25280 25486 25332 25492
rect 25568 25074 25596 26030
rect 25556 25068 25608 25074
rect 25556 25010 25608 25016
rect 25660 24938 25688 26302
rect 25648 24932 25700 24938
rect 25648 24874 25700 24880
rect 25280 24796 25332 24802
rect 25280 24738 25332 24744
rect 25096 24524 25148 24530
rect 25096 24466 25148 24472
rect 25004 23776 25056 23782
rect 25004 23718 25056 23724
rect 25292 23374 25320 24738
rect 25464 24388 25516 24394
rect 25464 24330 25516 24336
rect 25476 24258 25504 24330
rect 25464 24252 25516 24258
rect 25464 24194 25516 24200
rect 25476 23442 25504 24194
rect 25464 23436 25516 23442
rect 25464 23378 25516 23384
rect 25280 23368 25332 23374
rect 25280 23310 25332 23316
rect 24912 23096 24964 23102
rect 24912 23038 24964 23044
rect 25464 23096 25516 23102
rect 25464 23038 25516 23044
rect 24924 22778 24952 23038
rect 24924 22750 25320 22778
rect 25476 22762 25504 23038
rect 25096 22688 25148 22694
rect 25096 22630 25148 22636
rect 25004 22620 25056 22626
rect 25004 22562 25056 22568
rect 25016 21606 25044 22562
rect 25004 21600 25056 21606
rect 25004 21542 25056 21548
rect 24728 20580 24780 20586
rect 24728 20522 24780 20528
rect 25004 20580 25056 20586
rect 25004 20522 25056 20528
rect 23992 20512 24044 20518
rect 23992 20454 24044 20460
rect 24912 20512 24964 20518
rect 24912 20454 24964 20460
rect 23992 20376 24044 20382
rect 23992 20318 24044 20324
rect 21416 20036 21468 20042
rect 21416 19978 21468 19984
rect 22152 20036 22204 20042
rect 22152 19978 22204 19984
rect 23900 20036 23952 20042
rect 23900 19978 23952 19984
rect 21428 17338 21456 19978
rect 23256 19832 23308 19838
rect 23256 19774 23308 19780
rect 23268 19430 23296 19774
rect 22244 19424 22296 19430
rect 22244 19366 22296 19372
rect 22520 19424 22572 19430
rect 22520 19366 22572 19372
rect 23256 19424 23308 19430
rect 23256 19366 23308 19372
rect 21784 19016 21836 19022
rect 21784 18958 21836 18964
rect 21508 18880 21560 18886
rect 21508 18822 21560 18828
rect 21520 18342 21548 18822
rect 21796 18478 21824 18958
rect 22256 18886 22284 19366
rect 22532 19022 22560 19366
rect 22520 19016 22572 19022
rect 22520 18958 22572 18964
rect 22244 18880 22296 18886
rect 22244 18822 22296 18828
rect 21784 18472 21836 18478
rect 21784 18414 21836 18420
rect 21876 18472 21928 18478
rect 21876 18414 21928 18420
rect 21888 18342 21916 18414
rect 22532 18342 22560 18958
rect 23072 18948 23124 18954
rect 23072 18890 23124 18896
rect 21508 18336 21560 18342
rect 21508 18278 21560 18284
rect 21876 18336 21928 18342
rect 21876 18278 21928 18284
rect 22520 18336 22572 18342
rect 22520 18278 22572 18284
rect 22428 17860 22480 17866
rect 22428 17802 22480 17808
rect 22336 17792 22388 17798
rect 22336 17734 22388 17740
rect 22348 17458 22376 17734
rect 22336 17452 22388 17458
rect 22336 17394 22388 17400
rect 21232 17316 21284 17322
rect 21428 17310 21548 17338
rect 21232 17258 21284 17264
rect 20968 16358 21180 16386
rect 20772 16296 20824 16302
rect 20772 16238 20824 16244
rect 19852 16092 19904 16098
rect 19852 16034 19904 16040
rect 20128 16024 20180 16030
rect 20128 15966 20180 15972
rect 20680 16024 20732 16030
rect 20680 15966 20732 15972
rect 20140 15758 20168 15966
rect 20128 15752 20180 15758
rect 20128 15694 20180 15700
rect 19576 15616 19628 15622
rect 19576 15558 19628 15564
rect 19484 15072 19536 15078
rect 19484 15014 19536 15020
rect 19116 14836 19412 14856
rect 19172 14834 19196 14836
rect 19252 14834 19276 14836
rect 19332 14834 19356 14836
rect 19194 14782 19196 14834
rect 19258 14782 19270 14834
rect 19332 14782 19334 14834
rect 19172 14780 19196 14782
rect 19252 14780 19276 14782
rect 19332 14780 19356 14782
rect 19116 14760 19412 14780
rect 19496 14058 19524 15014
rect 19484 14052 19536 14058
rect 19484 13994 19536 14000
rect 18932 13984 18984 13990
rect 18932 13926 18984 13932
rect 18840 13916 18892 13922
rect 18760 13876 18840 13904
rect 18656 13858 18708 13864
rect 18840 13858 18892 13864
rect 18288 13576 18340 13582
rect 18288 13518 18340 13524
rect 18564 13508 18616 13514
rect 18564 13450 18616 13456
rect 17828 13372 17880 13378
rect 17828 13314 17880 13320
rect 17552 12828 17604 12834
rect 17552 12770 17604 12776
rect 17368 12488 17420 12494
rect 17368 12430 17420 12436
rect 17276 12216 17328 12222
rect 17276 12158 17328 12164
rect 17092 11332 17144 11338
rect 17092 11274 17144 11280
rect 17288 9624 17316 12158
rect 17380 11474 17408 12430
rect 17840 12358 17868 13314
rect 18576 12902 18604 13450
rect 18668 13446 18696 13858
rect 18656 13440 18708 13446
rect 18656 13382 18708 13388
rect 18668 12970 18696 13382
rect 18656 12964 18708 12970
rect 18656 12906 18708 12912
rect 18564 12896 18616 12902
rect 18564 12838 18616 12844
rect 18668 12850 18696 12906
rect 18852 12902 18880 13858
rect 18944 13514 18972 13926
rect 19116 13748 19412 13768
rect 19172 13746 19196 13748
rect 19252 13746 19276 13748
rect 19332 13746 19356 13748
rect 19194 13694 19196 13746
rect 19258 13694 19270 13746
rect 19332 13694 19334 13746
rect 19172 13692 19196 13694
rect 19252 13692 19276 13694
rect 19332 13692 19356 13694
rect 19116 13672 19412 13692
rect 18932 13508 18984 13514
rect 18932 13450 18984 13456
rect 19024 13440 19076 13446
rect 19024 13382 19076 13388
rect 18840 12896 18892 12902
rect 18668 12822 18788 12850
rect 18840 12838 18892 12844
rect 18380 12488 18432 12494
rect 18380 12430 18432 12436
rect 17828 12352 17880 12358
rect 17828 12294 17880 12300
rect 17840 11814 17868 12294
rect 18392 11882 18420 12430
rect 18656 12284 18708 12290
rect 18656 12226 18708 12232
rect 18668 11882 18696 12226
rect 18760 11882 18788 12822
rect 19036 12358 19064 13382
rect 19588 13122 19616 15558
rect 19668 15480 19720 15486
rect 19668 15422 19720 15428
rect 19680 15146 19708 15422
rect 19668 15140 19720 15146
rect 19668 15082 19720 15088
rect 20692 13990 20720 15966
rect 20784 15282 20812 16238
rect 20772 15276 20824 15282
rect 20772 15218 20824 15224
rect 20680 13984 20732 13990
rect 20680 13926 20732 13932
rect 20692 13514 20720 13926
rect 20680 13508 20732 13514
rect 20680 13450 20732 13456
rect 19588 13094 19708 13122
rect 19576 13032 19628 13038
rect 19576 12974 19628 12980
rect 19116 12660 19412 12680
rect 19172 12658 19196 12660
rect 19252 12658 19276 12660
rect 19332 12658 19356 12660
rect 19194 12606 19196 12658
rect 19258 12606 19270 12658
rect 19332 12606 19334 12658
rect 19172 12604 19196 12606
rect 19252 12604 19276 12606
rect 19332 12604 19356 12606
rect 19116 12584 19412 12604
rect 19588 12426 19616 12974
rect 19680 12494 19708 13094
rect 20968 12850 20996 16358
rect 21244 16166 21272 17258
rect 21324 16568 21376 16574
rect 21324 16510 21376 16516
rect 21336 16234 21364 16510
rect 21324 16228 21376 16234
rect 21324 16170 21376 16176
rect 21232 16160 21284 16166
rect 21232 16102 21284 16108
rect 21336 14602 21364 16170
rect 21416 15684 21468 15690
rect 21416 15626 21468 15632
rect 21428 14738 21456 15626
rect 21416 14732 21468 14738
rect 21416 14674 21468 14680
rect 21324 14596 21376 14602
rect 21324 14538 21376 14544
rect 21232 14052 21284 14058
rect 21232 13994 21284 14000
rect 21140 13984 21192 13990
rect 21140 13926 21192 13932
rect 21152 13310 21180 13926
rect 21244 13378 21272 13994
rect 21324 13916 21376 13922
rect 21324 13858 21376 13864
rect 21336 13650 21364 13858
rect 21324 13644 21376 13650
rect 21324 13586 21376 13592
rect 21232 13372 21284 13378
rect 21232 13314 21284 13320
rect 21140 13304 21192 13310
rect 21140 13246 21192 13252
rect 21152 12986 21180 13246
rect 21060 12958 21180 12986
rect 21060 12902 21088 12958
rect 21244 12902 21272 13314
rect 20600 12822 20996 12850
rect 21048 12896 21100 12902
rect 21048 12838 21100 12844
rect 21232 12896 21284 12902
rect 21232 12838 21284 12844
rect 20600 12766 20628 12822
rect 20588 12760 20640 12766
rect 20588 12702 20640 12708
rect 20956 12760 21008 12766
rect 20956 12702 21008 12708
rect 19668 12488 19720 12494
rect 19668 12430 19720 12436
rect 19576 12420 19628 12426
rect 19576 12362 19628 12368
rect 20128 12420 20180 12426
rect 20128 12362 20180 12368
rect 19024 12352 19076 12358
rect 19024 12294 19076 12300
rect 20140 12018 20168 12362
rect 20128 12012 20180 12018
rect 20128 11954 20180 11960
rect 18380 11876 18432 11882
rect 18380 11818 18432 11824
rect 18656 11876 18708 11882
rect 18656 11818 18708 11824
rect 18748 11876 18800 11882
rect 18748 11818 18800 11824
rect 17828 11808 17880 11814
rect 17828 11750 17880 11756
rect 19760 11808 19812 11814
rect 19760 11750 19812 11756
rect 19484 11672 19536 11678
rect 19484 11614 19536 11620
rect 19116 11572 19412 11592
rect 19172 11570 19196 11572
rect 19252 11570 19276 11572
rect 19332 11570 19356 11572
rect 19194 11518 19196 11570
rect 19258 11518 19270 11570
rect 19332 11518 19334 11570
rect 19172 11516 19196 11518
rect 19252 11516 19276 11518
rect 19332 11516 19356 11518
rect 19116 11496 19412 11516
rect 17368 11468 17420 11474
rect 17368 11410 17420 11416
rect 19496 9624 19524 11614
rect 19772 11474 19800 11750
rect 19760 11468 19812 11474
rect 19760 11410 19812 11416
rect 20968 11338 20996 12702
rect 21060 12018 21088 12838
rect 21048 12012 21100 12018
rect 21048 11954 21100 11960
rect 21336 11474 21364 13586
rect 21416 12420 21468 12426
rect 21416 12362 21468 12368
rect 21428 11882 21456 12362
rect 21520 12222 21548 17310
rect 22440 16778 22468 17802
rect 23084 17458 23112 18890
rect 23268 17866 23296 19366
rect 23348 19288 23400 19294
rect 23348 19230 23400 19236
rect 23624 19288 23676 19294
rect 23624 19230 23676 19236
rect 23360 18410 23388 19230
rect 23636 19090 23664 19230
rect 23624 19084 23676 19090
rect 23624 19026 23676 19032
rect 23348 18404 23400 18410
rect 23348 18346 23400 18352
rect 23636 18274 23664 19026
rect 23912 18954 23940 19978
rect 24004 18954 24032 20318
rect 24116 19732 24412 19752
rect 24172 19730 24196 19732
rect 24252 19730 24276 19732
rect 24332 19730 24356 19732
rect 24194 19678 24196 19730
rect 24258 19678 24270 19730
rect 24332 19678 24334 19730
rect 24172 19676 24196 19678
rect 24252 19676 24276 19678
rect 24332 19676 24356 19678
rect 24116 19656 24412 19676
rect 23900 18948 23952 18954
rect 23900 18890 23952 18896
rect 23992 18948 24044 18954
rect 23992 18890 24044 18896
rect 23912 18410 23940 18890
rect 23900 18404 23952 18410
rect 23900 18346 23952 18352
rect 23624 18268 23676 18274
rect 23624 18210 23676 18216
rect 23256 17860 23308 17866
rect 23256 17802 23308 17808
rect 23072 17452 23124 17458
rect 23072 17394 23124 17400
rect 23256 17316 23308 17322
rect 23256 17258 23308 17264
rect 23532 17316 23584 17322
rect 23636 17304 23664 18210
rect 24004 18206 24032 18890
rect 24452 18744 24504 18750
rect 24452 18686 24504 18692
rect 24116 18644 24412 18664
rect 24172 18642 24196 18644
rect 24252 18642 24276 18644
rect 24332 18642 24356 18644
rect 24194 18590 24196 18642
rect 24258 18590 24270 18642
rect 24332 18590 24334 18642
rect 24172 18588 24196 18590
rect 24252 18588 24276 18590
rect 24332 18588 24356 18590
rect 24116 18568 24412 18588
rect 24464 18342 24492 18686
rect 24452 18336 24504 18342
rect 24452 18278 24504 18284
rect 23992 18200 24044 18206
rect 23992 18142 24044 18148
rect 24004 17866 24032 18142
rect 23992 17860 24044 17866
rect 23992 17802 24044 17808
rect 23808 17656 23860 17662
rect 23808 17598 23860 17604
rect 23820 17322 23848 17598
rect 23584 17276 23664 17304
rect 23808 17316 23860 17322
rect 23532 17258 23584 17264
rect 23808 17258 23860 17264
rect 22428 16772 22480 16778
rect 22428 16714 22480 16720
rect 22152 16704 22204 16710
rect 22152 16646 22204 16652
rect 22164 16370 22192 16646
rect 22336 16636 22388 16642
rect 22336 16578 22388 16584
rect 22152 16364 22204 16370
rect 22152 16306 22204 16312
rect 21600 15616 21652 15622
rect 21600 15558 21652 15564
rect 21612 15214 21640 15558
rect 21600 15208 21652 15214
rect 21600 15150 21652 15156
rect 21612 14602 21640 15150
rect 22164 15078 22192 16306
rect 22348 16098 22376 16578
rect 22336 16092 22388 16098
rect 22336 16034 22388 16040
rect 22244 16024 22296 16030
rect 22244 15966 22296 15972
rect 22256 15758 22284 15966
rect 22244 15752 22296 15758
rect 22244 15694 22296 15700
rect 22348 15146 22376 16034
rect 22440 15826 22468 16714
rect 23268 16234 23296 17258
rect 24004 16778 24032 17802
rect 24544 17656 24596 17662
rect 24544 17598 24596 17604
rect 24116 17556 24412 17576
rect 24172 17554 24196 17556
rect 24252 17554 24276 17556
rect 24332 17554 24356 17556
rect 24194 17502 24196 17554
rect 24258 17502 24270 17554
rect 24332 17502 24334 17554
rect 24172 17500 24196 17502
rect 24252 17500 24276 17502
rect 24332 17500 24356 17502
rect 24116 17480 24412 17500
rect 24556 17186 24584 17598
rect 24544 17180 24596 17186
rect 24544 17122 24596 17128
rect 23992 16772 24044 16778
rect 23992 16714 24044 16720
rect 23532 16568 23584 16574
rect 23532 16510 23584 16516
rect 24544 16568 24596 16574
rect 24544 16510 24596 16516
rect 23544 16234 23572 16510
rect 24116 16468 24412 16488
rect 24172 16466 24196 16468
rect 24252 16466 24276 16468
rect 24332 16466 24356 16468
rect 24194 16414 24196 16466
rect 24258 16414 24270 16466
rect 24332 16414 24334 16466
rect 24172 16412 24196 16414
rect 24252 16412 24276 16414
rect 24332 16412 24356 16414
rect 24116 16392 24412 16412
rect 23256 16228 23308 16234
rect 23256 16170 23308 16176
rect 23532 16228 23584 16234
rect 23532 16170 23584 16176
rect 24556 16098 24584 16510
rect 24544 16092 24596 16098
rect 24544 16034 24596 16040
rect 22428 15820 22480 15826
rect 22428 15762 22480 15768
rect 23992 15480 24044 15486
rect 23992 15422 24044 15428
rect 22336 15140 22388 15146
rect 22336 15082 22388 15088
rect 22152 15072 22204 15078
rect 22152 15014 22204 15020
rect 22164 14602 22192 15014
rect 23900 14936 23952 14942
rect 23900 14878 23952 14884
rect 23912 14602 23940 14878
rect 24004 14670 24032 15422
rect 24116 15380 24412 15400
rect 24172 15378 24196 15380
rect 24252 15378 24276 15380
rect 24332 15378 24356 15380
rect 24194 15326 24196 15378
rect 24258 15326 24270 15378
rect 24332 15326 24334 15378
rect 24172 15324 24196 15326
rect 24252 15324 24276 15326
rect 24332 15324 24356 15326
rect 24116 15304 24412 15324
rect 24544 15072 24596 15078
rect 24544 15014 24596 15020
rect 24452 15004 24504 15010
rect 24452 14946 24504 14952
rect 23992 14664 24044 14670
rect 23992 14606 24044 14612
rect 21600 14596 21652 14602
rect 21600 14538 21652 14544
rect 22152 14596 22204 14602
rect 22152 14538 22204 14544
rect 23808 14596 23860 14602
rect 23808 14538 23860 14544
rect 23900 14596 23952 14602
rect 23900 14538 23952 14544
rect 23256 14392 23308 14398
rect 23256 14334 23308 14340
rect 23268 13582 23296 14334
rect 23820 14058 23848 14538
rect 23900 14392 23952 14398
rect 23900 14334 23952 14340
rect 23808 14052 23860 14058
rect 23808 13994 23860 14000
rect 23256 13576 23308 13582
rect 23256 13518 23308 13524
rect 23820 13514 23848 13994
rect 23912 13990 23940 14334
rect 24116 14292 24412 14312
rect 24172 14290 24196 14292
rect 24252 14290 24276 14292
rect 24332 14290 24356 14292
rect 24194 14238 24196 14290
rect 24258 14238 24270 14290
rect 24332 14238 24334 14290
rect 24172 14236 24196 14238
rect 24252 14236 24276 14238
rect 24332 14236 24356 14238
rect 24116 14216 24412 14236
rect 24464 13990 24492 14946
rect 24556 13990 24584 15014
rect 23900 13984 23952 13990
rect 23900 13926 23952 13932
rect 24452 13984 24504 13990
rect 24452 13926 24504 13932
rect 24544 13984 24596 13990
rect 24544 13926 24596 13932
rect 21600 13508 21652 13514
rect 21600 13450 21652 13456
rect 23808 13508 23860 13514
rect 23808 13450 23860 13456
rect 21612 13038 21640 13450
rect 24464 13446 24492 13926
rect 24556 13514 24584 13926
rect 24544 13508 24596 13514
rect 24544 13450 24596 13456
rect 24820 13508 24872 13514
rect 24820 13450 24872 13456
rect 24452 13440 24504 13446
rect 24452 13382 24504 13388
rect 24116 13204 24412 13224
rect 24172 13202 24196 13204
rect 24252 13202 24276 13204
rect 24332 13202 24356 13204
rect 24194 13150 24196 13202
rect 24258 13150 24270 13202
rect 24332 13150 24334 13202
rect 24172 13148 24196 13150
rect 24252 13148 24276 13150
rect 24332 13148 24356 13150
rect 24116 13128 24412 13148
rect 21600 13032 21652 13038
rect 21600 12974 21652 12980
rect 21784 12964 21836 12970
rect 21784 12906 21836 12912
rect 21692 12828 21744 12834
rect 21692 12770 21744 12776
rect 21704 12494 21732 12770
rect 21692 12488 21744 12494
rect 21692 12430 21744 12436
rect 21692 12352 21744 12358
rect 21692 12294 21744 12300
rect 21508 12216 21560 12222
rect 21508 12158 21560 12164
rect 21416 11876 21468 11882
rect 21416 11818 21468 11824
rect 21324 11468 21376 11474
rect 21324 11410 21376 11416
rect 20956 11332 21008 11338
rect 20956 11274 21008 11280
rect 21704 9624 21732 12294
rect 21796 11814 21824 12906
rect 23256 12896 23308 12902
rect 23256 12838 23308 12844
rect 22704 12828 22756 12834
rect 22704 12770 22756 12776
rect 22716 12562 22744 12770
rect 23268 12766 23296 12838
rect 23256 12760 23308 12766
rect 23256 12702 23308 12708
rect 22704 12556 22756 12562
rect 22704 12498 22756 12504
rect 23268 12494 23296 12702
rect 23716 12556 23768 12562
rect 23716 12498 23768 12504
rect 23256 12488 23308 12494
rect 23256 12430 23308 12436
rect 21784 11808 21836 11814
rect 21784 11750 21836 11756
rect 23164 11740 23216 11746
rect 23164 11682 23216 11688
rect 23176 11474 23204 11682
rect 23164 11468 23216 11474
rect 23164 11410 23216 11416
rect 23728 11338 23756 12498
rect 23992 12216 24044 12222
rect 23992 12158 24044 12164
rect 23716 11332 23768 11338
rect 23716 11274 23768 11280
rect 24004 10538 24032 12158
rect 24116 12116 24412 12136
rect 24172 12114 24196 12116
rect 24252 12114 24276 12116
rect 24332 12114 24356 12116
rect 24194 12062 24196 12114
rect 24258 12062 24270 12114
rect 24332 12062 24334 12114
rect 24172 12060 24196 12062
rect 24252 12060 24276 12062
rect 24332 12060 24356 12062
rect 24116 12040 24412 12060
rect 24832 11814 24860 13450
rect 24924 12358 24952 20454
rect 25016 17798 25044 20522
rect 25108 20042 25136 22630
rect 25292 22354 25320 22750
rect 25464 22756 25516 22762
rect 25464 22698 25516 22704
rect 25280 22348 25332 22354
rect 25280 22290 25332 22296
rect 25476 22218 25504 22698
rect 25464 22212 25516 22218
rect 25464 22154 25516 22160
rect 25188 21056 25240 21062
rect 25188 20998 25240 21004
rect 25280 21056 25332 21062
rect 25280 20998 25332 21004
rect 25200 20450 25228 20998
rect 25188 20444 25240 20450
rect 25188 20386 25240 20392
rect 25292 20178 25320 20998
rect 25648 20988 25700 20994
rect 25648 20930 25700 20936
rect 25660 20450 25688 20930
rect 25648 20444 25700 20450
rect 25648 20386 25700 20392
rect 25280 20172 25332 20178
rect 25280 20114 25332 20120
rect 25096 20036 25148 20042
rect 25096 19978 25148 19984
rect 25108 19430 25136 19978
rect 25096 19424 25148 19430
rect 25096 19366 25148 19372
rect 25660 19362 25688 20386
rect 25648 19356 25700 19362
rect 25648 19298 25700 19304
rect 25752 18460 25780 30876
rect 26200 30848 26252 30854
rect 26200 30790 26252 30796
rect 25832 30304 25884 30310
rect 25832 30246 25884 30252
rect 25844 29834 25872 30246
rect 25832 29828 25884 29834
rect 25832 29770 25884 29776
rect 25844 29290 25872 29770
rect 26108 29624 26160 29630
rect 26108 29566 26160 29572
rect 25832 29284 25884 29290
rect 25832 29226 25884 29232
rect 25832 28332 25884 28338
rect 25832 28274 25884 28280
rect 25844 25958 25872 28274
rect 25924 28060 25976 28066
rect 25924 28002 25976 28008
rect 25936 26910 25964 28002
rect 26120 27114 26148 29566
rect 26108 27108 26160 27114
rect 26108 27050 26160 27056
rect 25924 26904 25976 26910
rect 25924 26846 25976 26852
rect 26120 26026 26148 27050
rect 26108 26020 26160 26026
rect 26108 25962 26160 25968
rect 25832 25952 25884 25958
rect 25832 25894 25884 25900
rect 25844 25482 25872 25894
rect 26120 25482 26148 25962
rect 25832 25476 25884 25482
rect 25832 25418 25884 25424
rect 26108 25476 26160 25482
rect 26108 25418 26160 25424
rect 25924 25272 25976 25278
rect 25924 25214 25976 25220
rect 25936 24462 25964 25214
rect 25924 24456 25976 24462
rect 25924 24398 25976 24404
rect 26120 23238 26148 25418
rect 26108 23232 26160 23238
rect 26108 23174 26160 23180
rect 25922 22792 25978 22801
rect 25922 22727 25924 22736
rect 25976 22727 25978 22736
rect 25924 22698 25976 22704
rect 26120 21538 26148 23174
rect 26212 22218 26240 30790
rect 26304 30378 26332 32422
rect 26488 32418 26516 33442
rect 26476 32412 26528 32418
rect 26476 32354 26528 32360
rect 26488 32078 26516 32354
rect 26476 32072 26528 32078
rect 26476 32014 26528 32020
rect 26752 30916 26804 30922
rect 26752 30858 26804 30864
rect 26384 30780 26436 30786
rect 26384 30722 26436 30728
rect 26292 30372 26344 30378
rect 26292 30314 26344 30320
rect 26396 29834 26424 30722
rect 26764 30310 26792 30858
rect 26856 30854 26884 35809
rect 29248 34610 29276 35809
rect 29248 34582 29552 34610
rect 29116 34420 29412 34440
rect 29172 34418 29196 34420
rect 29252 34418 29276 34420
rect 29332 34418 29356 34420
rect 29194 34366 29196 34418
rect 29258 34366 29270 34418
rect 29332 34366 29334 34418
rect 29172 34364 29196 34366
rect 29252 34364 29276 34366
rect 29332 34364 29356 34366
rect 29116 34344 29412 34364
rect 28040 33568 28092 33574
rect 28040 33510 28092 33516
rect 28776 33568 28828 33574
rect 28776 33510 28828 33516
rect 27120 33432 27172 33438
rect 27120 33374 27172 33380
rect 27396 33432 27448 33438
rect 27396 33374 27448 33380
rect 27132 33166 27160 33374
rect 27120 33160 27172 33166
rect 27120 33102 27172 33108
rect 27120 32956 27172 32962
rect 27120 32898 27172 32904
rect 27132 32554 27160 32898
rect 27120 32548 27172 32554
rect 27120 32490 27172 32496
rect 26844 30848 26896 30854
rect 26844 30790 26896 30796
rect 26752 30304 26804 30310
rect 26752 30246 26804 30252
rect 27120 30304 27172 30310
rect 27120 30246 27172 30252
rect 26384 29828 26436 29834
rect 26384 29770 26436 29776
rect 26292 29148 26344 29154
rect 26292 29090 26344 29096
rect 26304 28066 26332 29090
rect 26396 29086 26424 29770
rect 26764 29766 26792 30246
rect 26936 29964 26988 29970
rect 26936 29906 26988 29912
rect 26752 29760 26804 29766
rect 26752 29702 26804 29708
rect 26568 29216 26620 29222
rect 26568 29158 26620 29164
rect 26384 29080 26436 29086
rect 26384 29022 26436 29028
rect 26292 28060 26344 28066
rect 26292 28002 26344 28008
rect 26580 27726 26608 29158
rect 26660 29148 26712 29154
rect 26660 29090 26712 29096
rect 26568 27720 26620 27726
rect 26568 27662 26620 27668
rect 26292 27584 26344 27590
rect 26292 27526 26344 27532
rect 26476 27584 26528 27590
rect 26476 27526 26528 27532
rect 26304 26638 26332 27526
rect 26292 26632 26344 26638
rect 26292 26574 26344 26580
rect 26304 23714 26332 26574
rect 26488 26502 26516 27526
rect 26672 27250 26700 29090
rect 26752 28536 26804 28542
rect 26752 28478 26804 28484
rect 26660 27244 26712 27250
rect 26660 27186 26712 27192
rect 26476 26496 26528 26502
rect 26476 26438 26528 26444
rect 26488 26162 26516 26438
rect 26764 26366 26792 28478
rect 26844 28196 26896 28202
rect 26844 28138 26896 28144
rect 26752 26360 26804 26366
rect 26752 26302 26804 26308
rect 26476 26156 26528 26162
rect 26476 26098 26528 26104
rect 26384 25884 26436 25890
rect 26384 25826 26436 25832
rect 26396 25482 26424 25826
rect 26384 25476 26436 25482
rect 26384 25418 26436 25424
rect 26396 24870 26424 25418
rect 26764 24938 26792 26302
rect 26752 24932 26804 24938
rect 26752 24874 26804 24880
rect 26384 24864 26436 24870
rect 26384 24806 26436 24812
rect 26474 24832 26530 24841
rect 26474 24767 26530 24776
rect 26384 24320 26436 24326
rect 26384 24262 26436 24268
rect 26292 23708 26344 23714
rect 26292 23650 26344 23656
rect 26200 22212 26252 22218
rect 26200 22154 26252 22160
rect 26212 21606 26240 22154
rect 26200 21600 26252 21606
rect 26200 21542 26252 21548
rect 26108 21532 26160 21538
rect 26108 21474 26160 21480
rect 26304 18954 26332 23650
rect 26396 22694 26424 24262
rect 26384 22688 26436 22694
rect 26384 22630 26436 22636
rect 26488 22626 26516 24767
rect 26764 23782 26792 24874
rect 26752 23776 26804 23782
rect 26752 23718 26804 23724
rect 26856 23322 26884 28138
rect 26948 25958 26976 29906
rect 27028 28672 27080 28678
rect 27028 28614 27080 28620
rect 27040 26638 27068 28614
rect 27132 28270 27160 30246
rect 27408 29834 27436 33374
rect 27856 32412 27908 32418
rect 27856 32354 27908 32360
rect 27868 32078 27896 32354
rect 27856 32072 27908 32078
rect 27856 32014 27908 32020
rect 27396 29828 27448 29834
rect 27396 29770 27448 29776
rect 27856 29828 27908 29834
rect 27856 29770 27908 29776
rect 27120 28264 27172 28270
rect 27120 28206 27172 28212
rect 27868 27658 27896 29770
rect 28052 29426 28080 33510
rect 28132 33500 28184 33506
rect 28132 33442 28184 33448
rect 28144 32486 28172 33442
rect 28408 32888 28460 32894
rect 28408 32830 28460 32836
rect 28132 32480 28184 32486
rect 28132 32422 28184 32428
rect 28144 32010 28172 32422
rect 28420 32078 28448 32830
rect 28408 32072 28460 32078
rect 28408 32014 28460 32020
rect 28132 32004 28184 32010
rect 28132 31946 28184 31952
rect 28592 32004 28644 32010
rect 28592 31946 28644 31952
rect 28500 30916 28552 30922
rect 28500 30858 28552 30864
rect 28512 30378 28540 30858
rect 28604 30786 28632 31946
rect 28592 30780 28644 30786
rect 28592 30722 28644 30728
rect 28500 30372 28552 30378
rect 28500 30314 28552 30320
rect 28512 29902 28540 30314
rect 28500 29896 28552 29902
rect 28500 29838 28552 29844
rect 28788 29680 28816 33510
rect 29524 33438 29552 34582
rect 31074 33944 31130 33953
rect 31074 33879 31130 33888
rect 29512 33432 29564 33438
rect 29512 33374 29564 33380
rect 29116 33332 29412 33352
rect 29172 33330 29196 33332
rect 29252 33330 29276 33332
rect 29332 33330 29356 33332
rect 29194 33278 29196 33330
rect 29258 33278 29270 33330
rect 29332 33278 29334 33330
rect 29172 33276 29196 33278
rect 29252 33276 29276 33278
rect 29332 33276 29356 33278
rect 29116 33256 29412 33276
rect 28868 33092 28920 33098
rect 28868 33034 28920 33040
rect 29052 33092 29104 33098
rect 29052 33034 29104 33040
rect 30616 33092 30668 33098
rect 30616 33034 30668 33040
rect 28880 32418 28908 33034
rect 29064 32486 29092 33034
rect 29144 32888 29196 32894
rect 29144 32830 29196 32836
rect 29156 32554 29184 32830
rect 29144 32548 29196 32554
rect 29144 32490 29196 32496
rect 29052 32480 29104 32486
rect 29052 32422 29104 32428
rect 28868 32412 28920 32418
rect 28868 32354 28920 32360
rect 28880 32078 28908 32354
rect 29116 32244 29412 32264
rect 29172 32242 29196 32244
rect 29252 32242 29276 32244
rect 29332 32242 29356 32244
rect 29194 32190 29196 32242
rect 29258 32190 29270 32242
rect 29332 32190 29334 32242
rect 29172 32188 29196 32190
rect 29252 32188 29276 32190
rect 29332 32188 29356 32190
rect 29116 32168 29412 32188
rect 28868 32072 28920 32078
rect 28868 32014 28920 32020
rect 28960 31392 29012 31398
rect 28960 31334 29012 31340
rect 28972 30378 29000 31334
rect 29788 31324 29840 31330
rect 29788 31266 29840 31272
rect 29604 31256 29656 31262
rect 29604 31198 29656 31204
rect 29696 31256 29748 31262
rect 29696 31198 29748 31204
rect 29116 31156 29412 31176
rect 29172 31154 29196 31156
rect 29252 31154 29276 31156
rect 29332 31154 29356 31156
rect 29194 31102 29196 31154
rect 29258 31102 29270 31154
rect 29332 31102 29334 31154
rect 29172 31100 29196 31102
rect 29252 31100 29276 31102
rect 29332 31100 29356 31102
rect 29116 31080 29412 31100
rect 29052 30780 29104 30786
rect 29052 30722 29104 30728
rect 28960 30372 29012 30378
rect 28960 30314 29012 30320
rect 29064 30242 29092 30722
rect 29052 30236 29104 30242
rect 29052 30178 29104 30184
rect 29116 30068 29412 30088
rect 29172 30066 29196 30068
rect 29252 30066 29276 30068
rect 29332 30066 29356 30068
rect 29194 30014 29196 30066
rect 29258 30014 29270 30066
rect 29332 30014 29334 30066
rect 29172 30012 29196 30014
rect 29252 30012 29276 30014
rect 29332 30012 29356 30014
rect 29116 29992 29412 30012
rect 29616 29902 29644 31198
rect 29708 30922 29736 31198
rect 29696 30916 29748 30922
rect 29696 30858 29748 30864
rect 29604 29896 29656 29902
rect 29604 29838 29656 29844
rect 28960 29828 29012 29834
rect 28960 29770 29012 29776
rect 28868 29692 28920 29698
rect 28788 29652 28868 29680
rect 28868 29634 28920 29640
rect 28040 29420 28092 29426
rect 28040 29362 28092 29368
rect 27948 29352 28000 29358
rect 27948 29294 28000 29300
rect 27960 28746 27988 29294
rect 27948 28740 28000 28746
rect 27948 28682 28000 28688
rect 28880 28660 28908 29634
rect 28972 29222 29000 29770
rect 29616 29358 29644 29838
rect 29604 29352 29656 29358
rect 29604 29294 29656 29300
rect 28960 29216 29012 29222
rect 28960 29158 29012 29164
rect 28972 28814 29000 29158
rect 29512 29148 29564 29154
rect 29512 29090 29564 29096
rect 29116 28980 29412 29000
rect 29172 28978 29196 28980
rect 29252 28978 29276 28980
rect 29332 28978 29356 28980
rect 29194 28926 29196 28978
rect 29258 28926 29270 28978
rect 29332 28926 29334 28978
rect 29172 28924 29196 28926
rect 29252 28924 29276 28926
rect 29332 28924 29356 28926
rect 29116 28904 29412 28924
rect 29524 28882 29552 29090
rect 29512 28876 29564 28882
rect 29512 28818 29564 28824
rect 28960 28808 29012 28814
rect 28960 28750 29012 28756
rect 28960 28672 29012 28678
rect 28880 28632 28960 28660
rect 28960 28614 29012 28620
rect 28972 28134 29000 28614
rect 28592 28128 28644 28134
rect 28592 28070 28644 28076
rect 28960 28128 29012 28134
rect 28960 28070 29012 28076
rect 27856 27652 27908 27658
rect 27856 27594 27908 27600
rect 28500 27652 28552 27658
rect 28500 27594 28552 27600
rect 27856 27516 27908 27522
rect 27856 27458 27908 27464
rect 27304 27448 27356 27454
rect 27304 27390 27356 27396
rect 27028 26632 27080 26638
rect 27028 26574 27080 26580
rect 27316 26570 27344 27390
rect 27868 26706 27896 27458
rect 28512 27454 28540 27594
rect 28604 27522 28632 28070
rect 28592 27516 28644 27522
rect 28592 27458 28644 27464
rect 28500 27448 28552 27454
rect 28500 27390 28552 27396
rect 27580 26700 27632 26706
rect 27580 26642 27632 26648
rect 27856 26700 27908 26706
rect 27856 26642 27908 26648
rect 27304 26564 27356 26570
rect 27304 26506 27356 26512
rect 27592 26434 27620 26642
rect 27580 26428 27632 26434
rect 27580 26370 27632 26376
rect 28408 26360 28460 26366
rect 28408 26302 28460 26308
rect 26936 25952 26988 25958
rect 26936 25894 26988 25900
rect 28316 25952 28368 25958
rect 28316 25894 28368 25900
rect 28224 25816 28276 25822
rect 28224 25758 28276 25764
rect 28236 25074 28264 25758
rect 28328 25550 28356 25894
rect 28316 25544 28368 25550
rect 28316 25486 28368 25492
rect 28224 25068 28276 25074
rect 28224 25010 28276 25016
rect 27946 24832 28002 24841
rect 27028 24796 27080 24802
rect 27946 24767 27948 24776
rect 27028 24738 27080 24744
rect 28000 24767 28002 24776
rect 27948 24738 28000 24744
rect 27040 24394 27068 24738
rect 27028 24388 27080 24394
rect 27028 24330 27080 24336
rect 27856 24388 27908 24394
rect 27856 24330 27908 24336
rect 27304 23912 27356 23918
rect 27304 23854 27356 23860
rect 26580 23294 26884 23322
rect 27316 23306 27344 23854
rect 27304 23300 27356 23306
rect 26476 22620 26528 22626
rect 26476 22562 26528 22568
rect 26384 20920 26436 20926
rect 26384 20862 26436 20868
rect 26396 20518 26424 20862
rect 26384 20512 26436 20518
rect 26384 20454 26436 20460
rect 26396 20042 26424 20454
rect 26384 20036 26436 20042
rect 26384 19978 26436 19984
rect 26292 18948 26344 18954
rect 26292 18890 26344 18896
rect 26476 18880 26528 18886
rect 26476 18822 26528 18828
rect 25752 18432 25872 18460
rect 25004 17792 25056 17798
rect 25004 17734 25056 17740
rect 25372 14596 25424 14602
rect 25372 14538 25424 14544
rect 25188 13576 25240 13582
rect 25188 13518 25240 13524
rect 25200 13106 25228 13518
rect 25188 13100 25240 13106
rect 25188 13042 25240 13048
rect 25004 12896 25056 12902
rect 25004 12838 25056 12844
rect 25016 12562 25044 12838
rect 25004 12556 25056 12562
rect 25004 12498 25056 12504
rect 24912 12352 24964 12358
rect 24912 12294 24964 12300
rect 24820 11808 24872 11814
rect 24820 11750 24872 11756
rect 25384 11406 25412 14538
rect 25556 13984 25608 13990
rect 25556 13926 25608 13932
rect 25568 13446 25596 13926
rect 25556 13440 25608 13446
rect 25556 13382 25608 13388
rect 25844 12902 25872 18432
rect 26488 18342 26516 18822
rect 26476 18336 26528 18342
rect 26476 18278 26528 18284
rect 26488 17934 26516 18278
rect 26476 17928 26528 17934
rect 26476 17870 26528 17876
rect 26580 13666 26608 23294
rect 27304 23242 27356 23248
rect 27868 23238 27896 24330
rect 27948 24320 28000 24326
rect 27948 24262 28000 24268
rect 27960 23986 27988 24262
rect 27948 23980 28000 23986
rect 27948 23922 28000 23928
rect 28132 23708 28184 23714
rect 28132 23650 28184 23656
rect 28144 23306 28172 23650
rect 28040 23300 28092 23306
rect 28040 23242 28092 23248
rect 28132 23300 28184 23306
rect 28132 23242 28184 23248
rect 27212 23232 27264 23238
rect 27212 23174 27264 23180
rect 27396 23232 27448 23238
rect 27396 23174 27448 23180
rect 27856 23232 27908 23238
rect 27856 23174 27908 23180
rect 27224 22694 27252 23174
rect 27408 22762 27436 23174
rect 27396 22756 27448 22762
rect 27396 22698 27448 22704
rect 27212 22688 27264 22694
rect 27212 22630 27264 22636
rect 27764 22212 27816 22218
rect 27764 22154 27816 22160
rect 27776 21606 27804 22154
rect 27856 22144 27908 22150
rect 27856 22086 27908 22092
rect 27868 21742 27896 22086
rect 28052 21810 28080 23242
rect 28040 21804 28092 21810
rect 28040 21746 28092 21752
rect 27856 21736 27908 21742
rect 27856 21678 27908 21684
rect 27764 21600 27816 21606
rect 27764 21542 27816 21548
rect 27776 21198 27804 21542
rect 27868 21198 27896 21678
rect 28316 21668 28368 21674
rect 28316 21610 28368 21616
rect 27948 21464 28000 21470
rect 27948 21406 28000 21412
rect 27764 21192 27816 21198
rect 27764 21134 27816 21140
rect 27856 21192 27908 21198
rect 27856 21134 27908 21140
rect 26844 21124 26896 21130
rect 26844 21066 26896 21072
rect 27304 21124 27356 21130
rect 27304 21066 27356 21072
rect 26856 20586 26884 21066
rect 27316 20654 27344 21066
rect 27304 20648 27356 20654
rect 27304 20590 27356 20596
rect 27960 20586 27988 21406
rect 26844 20580 26896 20586
rect 26844 20522 26896 20528
rect 27948 20580 28000 20586
rect 27948 20522 28000 20528
rect 27764 20104 27816 20110
rect 27764 20046 27816 20052
rect 27304 20036 27356 20042
rect 27304 19978 27356 19984
rect 27212 19084 27264 19090
rect 27212 19026 27264 19032
rect 27224 18342 27252 19026
rect 27316 19022 27344 19978
rect 27776 19362 27804 20046
rect 27948 19900 28000 19906
rect 27948 19842 28000 19848
rect 27960 19430 27988 19842
rect 27948 19424 28000 19430
rect 27948 19366 28000 19372
rect 27764 19356 27816 19362
rect 27764 19298 27816 19304
rect 27304 19016 27356 19022
rect 27304 18958 27356 18964
rect 27316 18410 27344 18958
rect 27304 18404 27356 18410
rect 27304 18346 27356 18352
rect 27776 18342 27804 19298
rect 28040 18948 28092 18954
rect 28040 18890 28092 18896
rect 27212 18336 27264 18342
rect 27212 18278 27264 18284
rect 27764 18336 27816 18342
rect 27764 18278 27816 18284
rect 27776 17866 27804 18278
rect 28052 18002 28080 18890
rect 28040 17996 28092 18002
rect 28040 17938 28092 17944
rect 27764 17860 27816 17866
rect 27764 17802 27816 17808
rect 27212 13984 27264 13990
rect 27212 13926 27264 13932
rect 26304 13638 26608 13666
rect 25832 12896 25884 12902
rect 25832 12838 25884 12844
rect 25832 12760 25884 12766
rect 25832 12702 25884 12708
rect 25844 12426 25872 12702
rect 25832 12420 25884 12426
rect 25832 12362 25884 12368
rect 25556 11740 25608 11746
rect 25556 11682 25608 11688
rect 25568 11474 25596 11682
rect 25556 11468 25608 11474
rect 25556 11410 25608 11416
rect 25372 11400 25424 11406
rect 25372 11342 25424 11348
rect 24116 11028 24412 11048
rect 24172 11026 24196 11028
rect 24252 11026 24276 11028
rect 24332 11026 24356 11028
rect 24194 10974 24196 11026
rect 24258 10974 24270 11026
rect 24332 10974 24334 11026
rect 24172 10972 24196 10974
rect 24252 10972 24276 10974
rect 24332 10972 24356 10974
rect 24116 10952 24412 10972
rect 24004 10510 24124 10538
rect 24096 9624 24124 10510
rect 26304 9624 26332 13638
rect 27224 13582 27252 13926
rect 28328 13666 28356 21610
rect 28420 17934 28448 26302
rect 28512 23442 28540 27390
rect 28972 26910 29000 28070
rect 29512 27992 29564 27998
rect 29512 27934 29564 27940
rect 29116 27892 29412 27912
rect 29172 27890 29196 27892
rect 29252 27890 29276 27892
rect 29332 27890 29356 27892
rect 29194 27838 29196 27890
rect 29258 27838 29270 27890
rect 29332 27838 29334 27890
rect 29172 27836 29196 27838
rect 29252 27836 29276 27838
rect 29332 27836 29356 27838
rect 29116 27816 29412 27836
rect 29524 26978 29552 27934
rect 29800 27114 29828 31266
rect 29972 30916 30024 30922
rect 29972 30858 30024 30864
rect 29984 29834 30012 30858
rect 30628 30446 30656 33034
rect 30800 30848 30852 30854
rect 30800 30790 30852 30796
rect 30616 30440 30668 30446
rect 30616 30382 30668 30388
rect 30812 30310 30840 30790
rect 30800 30304 30852 30310
rect 30800 30246 30852 30252
rect 29972 29828 30024 29834
rect 29972 29770 30024 29776
rect 29984 28746 30012 29770
rect 30892 29760 30944 29766
rect 30892 29702 30944 29708
rect 29972 28740 30024 28746
rect 29972 28682 30024 28688
rect 30904 27794 30932 29702
rect 31088 28202 31116 33879
rect 31456 33234 31484 35809
rect 33664 33642 33692 35809
rect 33652 33636 33704 33642
rect 33652 33578 33704 33584
rect 31444 33228 31496 33234
rect 31444 33170 31496 33176
rect 31260 31324 31312 31330
rect 31260 31266 31312 31272
rect 31272 30922 31300 31266
rect 31260 30916 31312 30922
rect 31260 30858 31312 30864
rect 31272 30446 31300 30858
rect 32640 30848 32692 30854
rect 32640 30790 32692 30796
rect 31810 30680 31866 30689
rect 31810 30615 31866 30624
rect 31260 30440 31312 30446
rect 31260 30382 31312 30388
rect 31444 30304 31496 30310
rect 31444 30246 31496 30252
rect 31168 29896 31220 29902
rect 31168 29838 31220 29844
rect 31180 29766 31208 29838
rect 31168 29760 31220 29766
rect 31168 29702 31220 29708
rect 31180 29222 31208 29702
rect 31168 29216 31220 29222
rect 31168 29158 31220 29164
rect 31456 29154 31484 30246
rect 31824 29970 31852 30615
rect 32652 30514 32680 30790
rect 32640 30508 32692 30514
rect 32640 30450 32692 30456
rect 31904 30168 31956 30174
rect 31904 30110 31956 30116
rect 32824 30168 32876 30174
rect 32824 30110 32876 30116
rect 31812 29964 31864 29970
rect 31812 29906 31864 29912
rect 31916 29902 31944 30110
rect 31904 29896 31956 29902
rect 31904 29838 31956 29844
rect 32836 29698 32864 30110
rect 32824 29692 32876 29698
rect 32824 29634 32876 29640
rect 32836 29222 32864 29634
rect 32824 29216 32876 29222
rect 32824 29158 32876 29164
rect 31444 29148 31496 29154
rect 31444 29090 31496 29096
rect 31456 28882 31484 29090
rect 31444 28876 31496 28882
rect 31444 28818 31496 28824
rect 31352 28740 31404 28746
rect 31352 28682 31404 28688
rect 31076 28196 31128 28202
rect 31076 28138 31128 28144
rect 30892 27788 30944 27794
rect 30892 27730 30944 27736
rect 30340 27584 30392 27590
rect 30340 27526 30392 27532
rect 30352 27114 30380 27526
rect 31258 27416 31314 27425
rect 31258 27351 31314 27360
rect 31272 27114 31300 27351
rect 29788 27108 29840 27114
rect 29788 27050 29840 27056
rect 30340 27108 30392 27114
rect 30340 27050 30392 27056
rect 31260 27108 31312 27114
rect 31260 27050 31312 27056
rect 29604 27040 29656 27046
rect 29604 26982 29656 26988
rect 29512 26972 29564 26978
rect 29512 26914 29564 26920
rect 28960 26904 29012 26910
rect 28960 26846 29012 26852
rect 28972 25482 29000 26846
rect 29116 26804 29412 26824
rect 29172 26802 29196 26804
rect 29252 26802 29276 26804
rect 29332 26802 29356 26804
rect 29194 26750 29196 26802
rect 29258 26750 29270 26802
rect 29332 26750 29334 26802
rect 29172 26748 29196 26750
rect 29252 26748 29276 26750
rect 29332 26748 29356 26750
rect 29116 26728 29412 26748
rect 29524 26570 29552 26914
rect 29616 26570 29644 26982
rect 29788 26972 29840 26978
rect 29788 26914 29840 26920
rect 29880 26972 29932 26978
rect 29880 26914 29932 26920
rect 29800 26638 29828 26914
rect 29788 26632 29840 26638
rect 29788 26574 29840 26580
rect 29512 26564 29564 26570
rect 29512 26506 29564 26512
rect 29604 26564 29656 26570
rect 29604 26506 29656 26512
rect 29616 25890 29644 26506
rect 29604 25884 29656 25890
rect 29604 25826 29656 25832
rect 29116 25716 29412 25736
rect 29172 25714 29196 25716
rect 29252 25714 29276 25716
rect 29332 25714 29356 25716
rect 29194 25662 29196 25714
rect 29258 25662 29270 25714
rect 29332 25662 29334 25714
rect 29172 25660 29196 25662
rect 29252 25660 29276 25662
rect 29332 25660 29356 25662
rect 29116 25640 29412 25660
rect 29512 25612 29564 25618
rect 29512 25554 29564 25560
rect 28960 25476 29012 25482
rect 28960 25418 29012 25424
rect 28592 25408 28644 25414
rect 28592 25350 28644 25356
rect 28604 24394 28632 25350
rect 28868 24456 28920 24462
rect 28868 24398 28920 24404
rect 28592 24388 28644 24394
rect 28592 24330 28644 24336
rect 28880 23782 28908 24398
rect 28972 24326 29000 25418
rect 29116 24628 29412 24648
rect 29172 24626 29196 24628
rect 29252 24626 29276 24628
rect 29332 24626 29356 24628
rect 29194 24574 29196 24626
rect 29258 24574 29270 24626
rect 29332 24574 29334 24626
rect 29172 24572 29196 24574
rect 29252 24572 29276 24574
rect 29332 24572 29356 24574
rect 29116 24552 29412 24572
rect 28960 24320 29012 24326
rect 28960 24262 29012 24268
rect 28868 23776 28920 23782
rect 28868 23718 28920 23724
rect 29116 23540 29412 23560
rect 29172 23538 29196 23540
rect 29252 23538 29276 23540
rect 29332 23538 29356 23540
rect 29194 23486 29196 23538
rect 29258 23486 29270 23538
rect 29332 23486 29334 23538
rect 29172 23484 29196 23486
rect 29252 23484 29276 23486
rect 29332 23484 29356 23486
rect 29116 23464 29412 23484
rect 28500 23436 28552 23442
rect 28500 23378 28552 23384
rect 28776 22756 28828 22762
rect 28776 22698 28828 22704
rect 28788 21826 28816 22698
rect 29116 22452 29412 22472
rect 29172 22450 29196 22452
rect 29252 22450 29276 22452
rect 29332 22450 29356 22452
rect 29194 22398 29196 22450
rect 29258 22398 29270 22450
rect 29332 22398 29334 22450
rect 29172 22396 29196 22398
rect 29252 22396 29276 22398
rect 29332 22396 29356 22398
rect 29116 22376 29412 22396
rect 29524 22354 29552 25554
rect 29800 25550 29828 26574
rect 29788 25544 29840 25550
rect 29788 25486 29840 25492
rect 29892 24870 29920 26914
rect 30248 26360 30300 26366
rect 30248 26302 30300 26308
rect 30260 26026 30288 26302
rect 30248 26020 30300 26026
rect 30248 25962 30300 25968
rect 30524 25952 30576 25958
rect 30524 25894 30576 25900
rect 30536 25550 30564 25894
rect 30524 25544 30576 25550
rect 30524 25486 30576 25492
rect 29880 24864 29932 24870
rect 29880 24806 29932 24812
rect 30340 24864 30392 24870
rect 30340 24806 30392 24812
rect 30248 24796 30300 24802
rect 30248 24738 30300 24744
rect 29788 24388 29840 24394
rect 29788 24330 29840 24336
rect 29800 23714 29828 24330
rect 29972 24320 30024 24326
rect 29972 24262 30024 24268
rect 29788 23708 29840 23714
rect 29788 23650 29840 23656
rect 29800 23442 29828 23650
rect 29788 23436 29840 23442
rect 29788 23378 29840 23384
rect 29604 23096 29656 23102
rect 29604 23038 29656 23044
rect 29512 22348 29564 22354
rect 29512 22290 29564 22296
rect 29512 22212 29564 22218
rect 29512 22154 29564 22160
rect 29328 22008 29380 22014
rect 29328 21950 29380 21956
rect 28788 21810 28908 21826
rect 28788 21804 28920 21810
rect 28788 21798 28868 21804
rect 28500 21532 28552 21538
rect 28500 21474 28552 21480
rect 28512 21266 28540 21474
rect 28500 21260 28552 21266
rect 28500 21202 28552 21208
rect 28500 19900 28552 19906
rect 28500 19842 28552 19848
rect 28512 19090 28540 19842
rect 28500 19084 28552 19090
rect 28500 19026 28552 19032
rect 28788 18954 28816 21798
rect 28868 21746 28920 21752
rect 29340 21606 29368 21950
rect 29328 21600 29380 21606
rect 29328 21542 29380 21548
rect 29524 21538 29552 22154
rect 29616 21606 29644 23038
rect 29880 22076 29932 22082
rect 29880 22018 29932 22024
rect 29892 21606 29920 22018
rect 29604 21600 29656 21606
rect 29604 21542 29656 21548
rect 29880 21600 29932 21606
rect 29880 21542 29932 21548
rect 29512 21532 29564 21538
rect 29512 21474 29564 21480
rect 29116 21364 29412 21384
rect 29172 21362 29196 21364
rect 29252 21362 29276 21364
rect 29332 21362 29356 21364
rect 29194 21310 29196 21362
rect 29258 21310 29270 21362
rect 29332 21310 29334 21362
rect 29172 21308 29196 21310
rect 29252 21308 29276 21310
rect 29332 21308 29356 21310
rect 29116 21288 29412 21308
rect 29524 21130 29552 21474
rect 29512 21124 29564 21130
rect 29512 21066 29564 21072
rect 29604 20444 29656 20450
rect 29604 20386 29656 20392
rect 29116 20276 29412 20296
rect 29172 20274 29196 20276
rect 29252 20274 29276 20276
rect 29332 20274 29356 20276
rect 29194 20222 29196 20274
rect 29258 20222 29270 20274
rect 29332 20222 29334 20274
rect 29172 20220 29196 20222
rect 29252 20220 29276 20222
rect 29332 20220 29356 20222
rect 29116 20200 29412 20220
rect 29616 20042 29644 20386
rect 29604 20036 29656 20042
rect 29604 19978 29656 19984
rect 29616 19566 29644 19978
rect 29696 19832 29748 19838
rect 29696 19774 29748 19780
rect 29604 19560 29656 19566
rect 29604 19502 29656 19508
rect 29116 19188 29412 19208
rect 29172 19186 29196 19188
rect 29252 19186 29276 19188
rect 29332 19186 29356 19188
rect 29194 19134 29196 19186
rect 29258 19134 29270 19186
rect 29332 19134 29334 19186
rect 29172 19132 29196 19134
rect 29252 19132 29276 19134
rect 29332 19132 29356 19134
rect 29116 19112 29412 19132
rect 28776 18948 28828 18954
rect 28776 18890 28828 18896
rect 29512 18744 29564 18750
rect 29512 18686 29564 18692
rect 29524 18410 29552 18686
rect 29616 18478 29644 19502
rect 29708 19430 29736 19774
rect 29696 19424 29748 19430
rect 29696 19366 29748 19372
rect 29604 18472 29656 18478
rect 29604 18414 29656 18420
rect 29512 18404 29564 18410
rect 29512 18346 29564 18352
rect 29116 18100 29412 18120
rect 29172 18098 29196 18100
rect 29252 18098 29276 18100
rect 29332 18098 29356 18100
rect 29194 18046 29196 18098
rect 29258 18046 29270 18098
rect 29332 18046 29334 18098
rect 29172 18044 29196 18046
rect 29252 18044 29276 18046
rect 29332 18044 29356 18046
rect 29116 18024 29412 18044
rect 28408 17928 28460 17934
rect 28408 17870 28460 17876
rect 28960 17792 29012 17798
rect 28960 17734 29012 17740
rect 28972 17118 29000 17734
rect 28960 17112 29012 17118
rect 28960 17054 29012 17060
rect 29116 17012 29412 17032
rect 29172 17010 29196 17012
rect 29252 17010 29276 17012
rect 29332 17010 29356 17012
rect 29194 16958 29196 17010
rect 29258 16958 29270 17010
rect 29332 16958 29334 17010
rect 29172 16956 29196 16958
rect 29252 16956 29276 16958
rect 29332 16956 29356 16958
rect 29116 16936 29412 16956
rect 29116 15924 29412 15944
rect 29172 15922 29196 15924
rect 29252 15922 29276 15924
rect 29332 15922 29356 15924
rect 29194 15870 29196 15922
rect 29258 15870 29270 15922
rect 29332 15870 29334 15922
rect 29172 15868 29196 15870
rect 29252 15868 29276 15870
rect 29332 15868 29356 15870
rect 29116 15848 29412 15868
rect 29116 14836 29412 14856
rect 29172 14834 29196 14836
rect 29252 14834 29276 14836
rect 29332 14834 29356 14836
rect 29194 14782 29196 14834
rect 29258 14782 29270 14834
rect 29332 14782 29334 14834
rect 29172 14780 29196 14782
rect 29252 14780 29276 14782
rect 29332 14780 29356 14782
rect 29116 14760 29412 14780
rect 29116 13748 29412 13768
rect 29172 13746 29196 13748
rect 29252 13746 29276 13748
rect 29332 13746 29356 13748
rect 29194 13694 29196 13746
rect 29258 13694 29270 13746
rect 29332 13694 29334 13746
rect 29172 13692 29196 13694
rect 29252 13692 29276 13694
rect 29332 13692 29356 13694
rect 29116 13672 29412 13692
rect 28328 13638 28724 13666
rect 27212 13576 27264 13582
rect 27212 13518 27264 13524
rect 26844 13440 26896 13446
rect 26844 13382 26896 13388
rect 26856 11882 26884 13382
rect 26844 11876 26896 11882
rect 26844 11818 26896 11824
rect 28696 9624 28724 13638
rect 29984 12834 30012 24262
rect 30260 23782 30288 24738
rect 30352 24394 30380 24806
rect 30536 24462 30564 25486
rect 30616 25476 30668 25482
rect 30616 25418 30668 25424
rect 30524 24456 30576 24462
rect 30524 24398 30576 24404
rect 30340 24388 30392 24394
rect 30340 24330 30392 24336
rect 30628 23889 30656 25418
rect 31364 25006 31392 28682
rect 31444 26564 31496 26570
rect 31444 26506 31496 26512
rect 31456 26094 31484 26506
rect 31444 26088 31496 26094
rect 31444 26030 31496 26036
rect 31536 25952 31588 25958
rect 31536 25894 31588 25900
rect 31548 25550 31576 25894
rect 32180 25884 32232 25890
rect 32180 25826 32232 25832
rect 31904 25816 31956 25822
rect 31904 25758 31956 25764
rect 31536 25544 31588 25550
rect 31536 25486 31588 25492
rect 30708 25000 30760 25006
rect 30708 24942 30760 24948
rect 31352 25000 31404 25006
rect 31352 24942 31404 24948
rect 30720 24394 30748 24942
rect 31168 24864 31220 24870
rect 31168 24806 31220 24812
rect 30708 24388 30760 24394
rect 30708 24330 30760 24336
rect 30720 23918 30748 24330
rect 31180 24326 31208 24806
rect 31364 24462 31392 24942
rect 31916 24462 31944 25758
rect 32192 25618 32220 25826
rect 32180 25612 32232 25618
rect 32180 25554 32232 25560
rect 32364 25476 32416 25482
rect 32364 25418 32416 25424
rect 32376 24870 32404 25418
rect 32364 24864 32416 24870
rect 32364 24806 32416 24812
rect 32376 24462 32404 24806
rect 31352 24456 31404 24462
rect 31352 24398 31404 24404
rect 31904 24456 31956 24462
rect 31904 24398 31956 24404
rect 32364 24456 32416 24462
rect 32364 24398 32416 24404
rect 31168 24320 31220 24326
rect 31168 24262 31220 24268
rect 30708 23912 30760 23918
rect 30614 23880 30670 23889
rect 30708 23854 30760 23860
rect 30614 23815 30670 23824
rect 30248 23776 30300 23782
rect 30248 23718 30300 23724
rect 30892 23300 30944 23306
rect 30892 23242 30944 23248
rect 30904 22762 30932 23242
rect 30892 22756 30944 22762
rect 30892 22698 30944 22704
rect 30248 22688 30300 22694
rect 30248 22630 30300 22636
rect 30800 22688 30852 22694
rect 30800 22630 30852 22636
rect 30260 22218 30288 22630
rect 30812 22218 30840 22630
rect 30248 22212 30300 22218
rect 30248 22154 30300 22160
rect 30800 22212 30852 22218
rect 30800 22154 30852 22160
rect 30064 22144 30116 22150
rect 30064 22086 30116 22092
rect 30076 21130 30104 22086
rect 30260 22014 30288 22154
rect 30248 22008 30300 22014
rect 30248 21950 30300 21956
rect 30156 21464 30208 21470
rect 30156 21406 30208 21412
rect 30168 21198 30196 21406
rect 30156 21192 30208 21198
rect 30156 21134 30208 21140
rect 30064 21124 30116 21130
rect 30064 21066 30116 21072
rect 30260 20654 30288 21950
rect 31180 21606 31208 24262
rect 31812 24184 31864 24190
rect 31812 24126 31864 24132
rect 31824 23850 31852 24126
rect 31812 23844 31864 23850
rect 31812 23786 31864 23792
rect 31260 22756 31312 22762
rect 31260 22698 31312 22704
rect 31272 22218 31300 22698
rect 31260 22212 31312 22218
rect 31260 22154 31312 22160
rect 31996 21736 32048 21742
rect 31996 21678 32048 21684
rect 32008 21606 32036 21678
rect 32180 21668 32232 21674
rect 32180 21610 32232 21616
rect 31168 21600 31220 21606
rect 31168 21542 31220 21548
rect 31996 21600 32048 21606
rect 31996 21542 32048 21548
rect 32088 21600 32140 21606
rect 32088 21542 32140 21548
rect 30248 20648 30300 20654
rect 32100 20625 32128 21542
rect 30248 20590 30300 20596
rect 32086 20616 32142 20625
rect 32086 20551 32142 20560
rect 30708 18880 30760 18886
rect 30708 18822 30760 18828
rect 30616 17112 30668 17118
rect 30614 17080 30616 17089
rect 30668 17080 30670 17089
rect 30614 17015 30670 17024
rect 30720 13825 30748 18822
rect 30706 13816 30762 13825
rect 30706 13751 30762 13760
rect 30616 13304 30668 13310
rect 30616 13246 30668 13252
rect 29972 12828 30024 12834
rect 29972 12770 30024 12776
rect 29116 12660 29412 12680
rect 29172 12658 29196 12660
rect 29252 12658 29276 12660
rect 29332 12658 29356 12660
rect 29194 12606 29196 12658
rect 29258 12606 29270 12658
rect 29332 12606 29334 12658
rect 29172 12604 29196 12606
rect 29252 12604 29276 12606
rect 29332 12604 29356 12606
rect 29116 12584 29412 12604
rect 29116 11572 29412 11592
rect 29172 11570 29196 11572
rect 29252 11570 29276 11572
rect 29332 11570 29356 11572
rect 29194 11518 29196 11570
rect 29258 11518 29270 11570
rect 29332 11518 29334 11570
rect 29172 11516 29196 11518
rect 29252 11516 29276 11518
rect 29332 11516 29356 11518
rect 29116 11496 29412 11516
rect 30628 10561 30656 13246
rect 32192 12306 32220 21610
rect 32192 12278 33140 12306
rect 30892 11332 30944 11338
rect 30892 11274 30944 11280
rect 30614 10552 30670 10561
rect 30614 10487 30670 10496
rect 30904 9624 30932 11274
rect 33112 9624 33140 12278
rect 10466 8824 10522 9624
rect 12674 8824 12730 9624
rect 14882 8824 14938 9624
rect 17274 8824 17330 9624
rect 19482 8824 19538 9624
rect 21690 8824 21746 9624
rect 24082 8824 24138 9624
rect 26290 8824 26346 9624
rect 28682 8824 28738 9624
rect 30890 8824 30946 9624
rect 33098 8824 33154 9624
<< via2 >>
rect 14116 33874 14172 33876
rect 14196 33874 14252 33876
rect 14276 33874 14332 33876
rect 14356 33874 14412 33876
rect 14116 33822 14142 33874
rect 14142 33822 14172 33874
rect 14196 33822 14206 33874
rect 14206 33822 14252 33874
rect 14276 33822 14322 33874
rect 14322 33822 14332 33874
rect 14356 33822 14386 33874
rect 14386 33822 14412 33874
rect 14116 33820 14172 33822
rect 14196 33820 14252 33822
rect 14276 33820 14332 33822
rect 14356 33820 14412 33822
rect 13962 33072 14018 33128
rect 14116 32786 14172 32788
rect 14196 32786 14252 32788
rect 14276 32786 14332 32788
rect 14356 32786 14412 32788
rect 14116 32734 14142 32786
rect 14142 32734 14172 32786
rect 14196 32734 14206 32786
rect 14206 32734 14252 32786
rect 14276 32734 14322 32786
rect 14322 32734 14332 32786
rect 14356 32734 14386 32786
rect 14386 32734 14412 32786
rect 14116 32732 14172 32734
rect 14196 32732 14252 32734
rect 14276 32732 14332 32734
rect 14356 32732 14412 32734
rect 14116 31698 14172 31700
rect 14196 31698 14252 31700
rect 14276 31698 14332 31700
rect 14356 31698 14412 31700
rect 14116 31646 14142 31698
rect 14142 31646 14172 31698
rect 14196 31646 14206 31698
rect 14206 31646 14252 31698
rect 14276 31646 14322 31698
rect 14322 31646 14332 31698
rect 14356 31646 14386 31698
rect 14386 31646 14412 31698
rect 14116 31644 14172 31646
rect 14196 31644 14252 31646
rect 14276 31644 14332 31646
rect 14356 31644 14412 31646
rect 14116 30610 14172 30612
rect 14196 30610 14252 30612
rect 14276 30610 14332 30612
rect 14356 30610 14412 30612
rect 14116 30558 14142 30610
rect 14142 30558 14172 30610
rect 14196 30558 14206 30610
rect 14206 30558 14252 30610
rect 14276 30558 14322 30610
rect 14322 30558 14332 30610
rect 14356 30558 14386 30610
rect 14386 30558 14412 30610
rect 14116 30556 14172 30558
rect 14196 30556 14252 30558
rect 14276 30556 14332 30558
rect 14356 30556 14412 30558
rect 13962 29808 14018 29864
rect 14116 29522 14172 29524
rect 14196 29522 14252 29524
rect 14276 29522 14332 29524
rect 14356 29522 14412 29524
rect 14116 29470 14142 29522
rect 14142 29470 14172 29522
rect 14196 29470 14206 29522
rect 14206 29470 14252 29522
rect 14276 29470 14322 29522
rect 14322 29470 14332 29522
rect 14356 29470 14386 29522
rect 14386 29470 14412 29522
rect 14116 29468 14172 29470
rect 14196 29468 14252 29470
rect 14276 29468 14332 29470
rect 14356 29468 14412 29470
rect 14116 28434 14172 28436
rect 14196 28434 14252 28436
rect 14276 28434 14332 28436
rect 14356 28434 14412 28436
rect 14116 28382 14142 28434
rect 14142 28382 14172 28434
rect 14196 28382 14206 28434
rect 14206 28382 14252 28434
rect 14276 28382 14322 28434
rect 14322 28382 14332 28434
rect 14356 28382 14386 28434
rect 14386 28382 14412 28434
rect 14116 28380 14172 28382
rect 14196 28380 14252 28382
rect 14276 28380 14332 28382
rect 14356 28380 14412 28382
rect 11938 26272 11994 26328
rect 14116 27346 14172 27348
rect 14196 27346 14252 27348
rect 14276 27346 14332 27348
rect 14356 27346 14412 27348
rect 14116 27294 14142 27346
rect 14142 27294 14172 27346
rect 14196 27294 14206 27346
rect 14206 27294 14252 27346
rect 14276 27294 14322 27346
rect 14322 27294 14332 27346
rect 14356 27294 14386 27346
rect 14386 27294 14412 27346
rect 14116 27292 14172 27294
rect 14196 27292 14252 27294
rect 14276 27292 14332 27294
rect 14356 27292 14412 27294
rect 14116 26258 14172 26260
rect 14196 26258 14252 26260
rect 14276 26258 14332 26260
rect 14356 26258 14412 26260
rect 14116 26206 14142 26258
rect 14142 26206 14172 26258
rect 14196 26206 14206 26258
rect 14206 26206 14252 26258
rect 14276 26206 14322 26258
rect 14322 26206 14332 26258
rect 14356 26206 14386 26258
rect 14386 26206 14412 26258
rect 14116 26204 14172 26206
rect 14196 26204 14252 26206
rect 14276 26204 14332 26206
rect 14356 26204 14412 26206
rect 13134 23008 13190 23064
rect 14116 25170 14172 25172
rect 14196 25170 14252 25172
rect 14276 25170 14332 25172
rect 14356 25170 14412 25172
rect 14116 25118 14142 25170
rect 14142 25118 14172 25170
rect 14196 25118 14206 25170
rect 14206 25118 14252 25170
rect 14276 25118 14322 25170
rect 14322 25118 14332 25170
rect 14356 25118 14386 25170
rect 14386 25118 14412 25170
rect 14116 25116 14172 25118
rect 14196 25116 14252 25118
rect 14276 25116 14332 25118
rect 14356 25116 14412 25118
rect 14116 24082 14172 24084
rect 14196 24082 14252 24084
rect 14276 24082 14332 24084
rect 14356 24082 14412 24084
rect 14116 24030 14142 24082
rect 14142 24030 14172 24082
rect 14196 24030 14206 24082
rect 14206 24030 14252 24082
rect 14276 24030 14322 24082
rect 14322 24030 14332 24082
rect 14356 24030 14386 24082
rect 14386 24030 14412 24082
rect 14116 24028 14172 24030
rect 14196 24028 14252 24030
rect 14276 24028 14332 24030
rect 14356 24028 14412 24030
rect 14116 22994 14172 22996
rect 14196 22994 14252 22996
rect 14276 22994 14332 22996
rect 14356 22994 14412 22996
rect 14116 22942 14142 22994
rect 14142 22942 14172 22994
rect 14196 22942 14206 22994
rect 14206 22942 14252 22994
rect 14276 22942 14322 22994
rect 14322 22942 14332 22994
rect 14356 22942 14386 22994
rect 14386 22942 14412 22994
rect 14116 22940 14172 22942
rect 14196 22940 14252 22942
rect 14276 22940 14332 22942
rect 14356 22940 14412 22942
rect 14116 21906 14172 21908
rect 14196 21906 14252 21908
rect 14276 21906 14332 21908
rect 14356 21906 14412 21908
rect 14116 21854 14142 21906
rect 14142 21854 14172 21906
rect 14196 21854 14206 21906
rect 14206 21854 14252 21906
rect 14276 21854 14322 21906
rect 14322 21854 14332 21906
rect 14356 21854 14386 21906
rect 14386 21854 14412 21906
rect 14116 21852 14172 21854
rect 14196 21852 14252 21854
rect 14276 21852 14332 21854
rect 14356 21852 14412 21854
rect 14116 20818 14172 20820
rect 14196 20818 14252 20820
rect 14276 20818 14332 20820
rect 14356 20818 14412 20820
rect 14116 20766 14142 20818
rect 14142 20766 14172 20818
rect 14196 20766 14206 20818
rect 14206 20766 14252 20818
rect 14276 20766 14322 20818
rect 14322 20766 14332 20818
rect 14356 20766 14386 20818
rect 14386 20766 14412 20818
rect 14116 20764 14172 20766
rect 14196 20764 14252 20766
rect 14276 20764 14332 20766
rect 14356 20764 14412 20766
rect 12674 19744 12730 19800
rect 14116 19730 14172 19732
rect 14196 19730 14252 19732
rect 14276 19730 14332 19732
rect 14356 19730 14412 19732
rect 14116 19678 14142 19730
rect 14142 19678 14172 19730
rect 14196 19678 14206 19730
rect 14206 19678 14252 19730
rect 14276 19678 14322 19730
rect 14322 19678 14332 19730
rect 14356 19678 14386 19730
rect 14386 19678 14412 19730
rect 14116 19676 14172 19678
rect 14196 19676 14252 19678
rect 14276 19676 14332 19678
rect 14356 19676 14412 19678
rect 19116 34418 19172 34420
rect 19196 34418 19252 34420
rect 19276 34418 19332 34420
rect 19356 34418 19412 34420
rect 19116 34366 19142 34418
rect 19142 34366 19172 34418
rect 19196 34366 19206 34418
rect 19206 34366 19252 34418
rect 19276 34366 19322 34418
rect 19322 34366 19332 34418
rect 19356 34366 19386 34418
rect 19386 34366 19412 34418
rect 19116 34364 19172 34366
rect 19196 34364 19252 34366
rect 19276 34364 19332 34366
rect 19356 34364 19412 34366
rect 19116 33330 19172 33332
rect 19196 33330 19252 33332
rect 19276 33330 19332 33332
rect 19356 33330 19412 33332
rect 19116 33278 19142 33330
rect 19142 33278 19172 33330
rect 19196 33278 19206 33330
rect 19206 33278 19252 33330
rect 19276 33278 19322 33330
rect 19322 33278 19332 33330
rect 19356 33278 19386 33330
rect 19386 33278 19412 33330
rect 19116 33276 19172 33278
rect 19196 33276 19252 33278
rect 19276 33276 19332 33278
rect 19356 33276 19412 33278
rect 19116 32242 19172 32244
rect 19196 32242 19252 32244
rect 19276 32242 19332 32244
rect 19356 32242 19412 32244
rect 19116 32190 19142 32242
rect 19142 32190 19172 32242
rect 19196 32190 19206 32242
rect 19206 32190 19252 32242
rect 19276 32190 19322 32242
rect 19322 32190 19332 32242
rect 19356 32190 19386 32242
rect 19386 32190 19412 32242
rect 19116 32188 19172 32190
rect 19196 32188 19252 32190
rect 19276 32188 19332 32190
rect 19356 32188 19412 32190
rect 19116 31154 19172 31156
rect 19196 31154 19252 31156
rect 19276 31154 19332 31156
rect 19356 31154 19412 31156
rect 19116 31102 19142 31154
rect 19142 31102 19172 31154
rect 19196 31102 19206 31154
rect 19206 31102 19252 31154
rect 19276 31102 19322 31154
rect 19322 31102 19332 31154
rect 19356 31102 19386 31154
rect 19386 31102 19412 31154
rect 19116 31100 19172 31102
rect 19196 31100 19252 31102
rect 19276 31100 19332 31102
rect 19356 31100 19412 31102
rect 19116 30066 19172 30068
rect 19196 30066 19252 30068
rect 19276 30066 19332 30068
rect 19356 30066 19412 30068
rect 19116 30014 19142 30066
rect 19142 30014 19172 30066
rect 19196 30014 19206 30066
rect 19206 30014 19252 30066
rect 19276 30014 19322 30066
rect 19322 30014 19332 30066
rect 19356 30014 19386 30066
rect 19386 30014 19412 30066
rect 19116 30012 19172 30014
rect 19196 30012 19252 30014
rect 19276 30012 19332 30014
rect 19356 30012 19412 30014
rect 19116 28978 19172 28980
rect 19196 28978 19252 28980
rect 19276 28978 19332 28980
rect 19356 28978 19412 28980
rect 19116 28926 19142 28978
rect 19142 28926 19172 28978
rect 19196 28926 19206 28978
rect 19206 28926 19252 28978
rect 19276 28926 19322 28978
rect 19322 28926 19332 28978
rect 19356 28926 19386 28978
rect 19386 28926 19412 28978
rect 19116 28924 19172 28926
rect 19196 28924 19252 28926
rect 19276 28924 19332 28926
rect 19356 28924 19412 28926
rect 19116 27890 19172 27892
rect 19196 27890 19252 27892
rect 19276 27890 19332 27892
rect 19356 27890 19412 27892
rect 19116 27838 19142 27890
rect 19142 27838 19172 27890
rect 19196 27838 19206 27890
rect 19206 27838 19252 27890
rect 19276 27838 19322 27890
rect 19322 27838 19332 27890
rect 19356 27838 19386 27890
rect 19386 27838 19412 27890
rect 19116 27836 19172 27838
rect 19196 27836 19252 27838
rect 19276 27836 19332 27838
rect 19356 27836 19412 27838
rect 19116 26802 19172 26804
rect 19196 26802 19252 26804
rect 19276 26802 19332 26804
rect 19356 26802 19412 26804
rect 19116 26750 19142 26802
rect 19142 26750 19172 26802
rect 19196 26750 19206 26802
rect 19206 26750 19252 26802
rect 19276 26750 19322 26802
rect 19322 26750 19332 26802
rect 19356 26750 19386 26802
rect 19386 26750 19412 26802
rect 19116 26748 19172 26750
rect 19196 26748 19252 26750
rect 19276 26748 19332 26750
rect 19356 26748 19412 26750
rect 19116 25714 19172 25716
rect 19196 25714 19252 25716
rect 19276 25714 19332 25716
rect 19356 25714 19412 25716
rect 19116 25662 19142 25714
rect 19142 25662 19172 25714
rect 19196 25662 19206 25714
rect 19206 25662 19252 25714
rect 19276 25662 19322 25714
rect 19322 25662 19332 25714
rect 19356 25662 19386 25714
rect 19386 25662 19412 25714
rect 19116 25660 19172 25662
rect 19196 25660 19252 25662
rect 19276 25660 19332 25662
rect 19356 25660 19412 25662
rect 18470 23144 18526 23200
rect 19116 24626 19172 24628
rect 19196 24626 19252 24628
rect 19276 24626 19332 24628
rect 19356 24626 19412 24628
rect 19116 24574 19142 24626
rect 19142 24574 19172 24626
rect 19196 24574 19206 24626
rect 19206 24574 19252 24626
rect 19276 24574 19322 24626
rect 19322 24574 19332 24626
rect 19356 24574 19386 24626
rect 19386 24574 19412 24626
rect 19116 24572 19172 24574
rect 19196 24572 19252 24574
rect 19276 24572 19332 24574
rect 19356 24572 19412 24574
rect 14116 18642 14172 18644
rect 14196 18642 14252 18644
rect 14276 18642 14332 18644
rect 14356 18642 14412 18644
rect 14116 18590 14142 18642
rect 14142 18590 14172 18642
rect 14196 18590 14206 18642
rect 14206 18590 14252 18642
rect 14276 18590 14322 18642
rect 14322 18590 14332 18642
rect 14356 18590 14386 18642
rect 14386 18590 14412 18642
rect 14116 18588 14172 18590
rect 14196 18588 14252 18590
rect 14276 18588 14332 18590
rect 14356 18588 14412 18590
rect 14116 17554 14172 17556
rect 14196 17554 14252 17556
rect 14276 17554 14332 17556
rect 14356 17554 14412 17556
rect 14116 17502 14142 17554
rect 14142 17502 14172 17554
rect 14196 17502 14206 17554
rect 14206 17502 14252 17554
rect 14276 17502 14322 17554
rect 14322 17502 14332 17554
rect 14356 17502 14386 17554
rect 14386 17502 14412 17554
rect 14116 17500 14172 17502
rect 14196 17500 14252 17502
rect 14276 17500 14332 17502
rect 14356 17500 14412 17502
rect 14116 16466 14172 16468
rect 14196 16466 14252 16468
rect 14276 16466 14332 16468
rect 14356 16466 14412 16468
rect 14116 16414 14142 16466
rect 14142 16414 14172 16466
rect 14196 16414 14206 16466
rect 14206 16414 14252 16466
rect 14276 16414 14322 16466
rect 14322 16414 14332 16466
rect 14356 16414 14386 16466
rect 14386 16414 14412 16466
rect 14116 16412 14172 16414
rect 14196 16412 14252 16414
rect 14276 16412 14332 16414
rect 14356 16412 14412 16414
rect 13962 16208 14018 16264
rect 14116 15378 14172 15380
rect 14196 15378 14252 15380
rect 14276 15378 14332 15380
rect 14356 15378 14412 15380
rect 14116 15326 14142 15378
rect 14142 15326 14172 15378
rect 14196 15326 14206 15378
rect 14206 15326 14252 15378
rect 14276 15326 14322 15378
rect 14322 15326 14332 15378
rect 14356 15326 14386 15378
rect 14386 15326 14412 15378
rect 14116 15324 14172 15326
rect 14196 15324 14252 15326
rect 14276 15324 14332 15326
rect 14356 15324 14412 15326
rect 12674 12964 12730 13000
rect 12674 12944 12676 12964
rect 12676 12944 12728 12964
rect 12728 12944 12730 12964
rect 14116 14290 14172 14292
rect 14196 14290 14252 14292
rect 14276 14290 14332 14292
rect 14356 14290 14412 14292
rect 14116 14238 14142 14290
rect 14142 14238 14172 14290
rect 14196 14238 14206 14290
rect 14206 14238 14252 14290
rect 14276 14238 14322 14290
rect 14322 14238 14332 14290
rect 14356 14238 14386 14290
rect 14386 14238 14412 14290
rect 14116 14236 14172 14238
rect 14196 14236 14252 14238
rect 14276 14236 14332 14238
rect 14356 14236 14412 14238
rect 19116 23538 19172 23540
rect 19196 23538 19252 23540
rect 19276 23538 19332 23540
rect 19356 23538 19412 23540
rect 19116 23486 19142 23538
rect 19142 23486 19172 23538
rect 19196 23486 19206 23538
rect 19206 23486 19252 23538
rect 19276 23486 19322 23538
rect 19322 23486 19332 23538
rect 19356 23486 19386 23538
rect 19386 23486 19412 23538
rect 19116 23484 19172 23486
rect 19196 23484 19252 23486
rect 19276 23484 19332 23486
rect 19356 23484 19412 23486
rect 19482 23180 19484 23200
rect 19484 23180 19536 23200
rect 19536 23180 19538 23200
rect 19482 23144 19538 23180
rect 19574 22736 19630 22792
rect 19116 22450 19172 22452
rect 19196 22450 19252 22452
rect 19276 22450 19332 22452
rect 19356 22450 19412 22452
rect 19116 22398 19142 22450
rect 19142 22398 19172 22450
rect 19196 22398 19206 22450
rect 19206 22398 19252 22450
rect 19276 22398 19322 22450
rect 19322 22398 19332 22450
rect 19356 22398 19386 22450
rect 19386 22398 19412 22450
rect 19116 22396 19172 22398
rect 19196 22396 19252 22398
rect 19276 22396 19332 22398
rect 19356 22396 19412 22398
rect 19116 21362 19172 21364
rect 19196 21362 19252 21364
rect 19276 21362 19332 21364
rect 19356 21362 19412 21364
rect 19116 21310 19142 21362
rect 19142 21310 19172 21362
rect 19196 21310 19206 21362
rect 19206 21310 19252 21362
rect 19276 21310 19322 21362
rect 19322 21310 19332 21362
rect 19356 21310 19386 21362
rect 19386 21310 19412 21362
rect 19116 21308 19172 21310
rect 19196 21308 19252 21310
rect 19276 21308 19332 21310
rect 19356 21308 19412 21310
rect 19116 20274 19172 20276
rect 19196 20274 19252 20276
rect 19276 20274 19332 20276
rect 19356 20274 19412 20276
rect 19116 20222 19142 20274
rect 19142 20222 19172 20274
rect 19196 20222 19206 20274
rect 19206 20222 19252 20274
rect 19276 20222 19322 20274
rect 19322 20222 19332 20274
rect 19356 20222 19386 20274
rect 19386 20222 19412 20274
rect 19116 20220 19172 20222
rect 19196 20220 19252 20222
rect 19276 20220 19332 20222
rect 19356 20220 19412 20222
rect 19116 19186 19172 19188
rect 19196 19186 19252 19188
rect 19276 19186 19332 19188
rect 19356 19186 19412 19188
rect 19116 19134 19142 19186
rect 19142 19134 19172 19186
rect 19196 19134 19206 19186
rect 19206 19134 19252 19186
rect 19276 19134 19322 19186
rect 19322 19134 19332 19186
rect 19356 19134 19386 19186
rect 19386 19134 19412 19186
rect 19116 19132 19172 19134
rect 19196 19132 19252 19134
rect 19276 19132 19332 19134
rect 19356 19132 19412 19134
rect 14116 13202 14172 13204
rect 14196 13202 14252 13204
rect 14276 13202 14332 13204
rect 14356 13202 14412 13204
rect 14116 13150 14142 13202
rect 14142 13150 14172 13202
rect 14196 13150 14206 13202
rect 14206 13150 14252 13202
rect 14276 13150 14322 13202
rect 14322 13150 14332 13202
rect 14356 13150 14386 13202
rect 14386 13150 14412 13202
rect 14116 13148 14172 13150
rect 14196 13148 14252 13150
rect 14276 13148 14332 13150
rect 14356 13148 14412 13150
rect 14116 12114 14172 12116
rect 14196 12114 14252 12116
rect 14276 12114 14332 12116
rect 14356 12114 14412 12116
rect 14116 12062 14142 12114
rect 14142 12062 14172 12114
rect 14196 12062 14206 12114
rect 14206 12062 14252 12114
rect 14276 12062 14322 12114
rect 14322 12062 14332 12114
rect 14356 12062 14386 12114
rect 14386 12062 14412 12114
rect 14116 12060 14172 12062
rect 14196 12060 14252 12062
rect 14276 12060 14332 12062
rect 14356 12060 14412 12062
rect 14116 11026 14172 11028
rect 14196 11026 14252 11028
rect 14276 11026 14332 11028
rect 14356 11026 14412 11028
rect 14116 10974 14142 11026
rect 14142 10974 14172 11026
rect 14196 10974 14206 11026
rect 14206 10974 14252 11026
rect 14276 10974 14322 11026
rect 14322 10974 14332 11026
rect 14356 10974 14386 11026
rect 14386 10974 14412 11026
rect 14116 10972 14172 10974
rect 14196 10972 14252 10974
rect 14276 10972 14332 10974
rect 14356 10972 14412 10974
rect 19116 18098 19172 18100
rect 19196 18098 19252 18100
rect 19276 18098 19332 18100
rect 19356 18098 19412 18100
rect 19116 18046 19142 18098
rect 19142 18046 19172 18098
rect 19196 18046 19206 18098
rect 19206 18046 19252 18098
rect 19276 18046 19322 18098
rect 19322 18046 19332 18098
rect 19356 18046 19386 18098
rect 19386 18046 19412 18098
rect 19116 18044 19172 18046
rect 19196 18044 19252 18046
rect 19276 18044 19332 18046
rect 19356 18044 19412 18046
rect 19116 17010 19172 17012
rect 19196 17010 19252 17012
rect 19276 17010 19332 17012
rect 19356 17010 19412 17012
rect 19116 16958 19142 17010
rect 19142 16958 19172 17010
rect 19196 16958 19206 17010
rect 19206 16958 19252 17010
rect 19276 16958 19322 17010
rect 19322 16958 19332 17010
rect 19356 16958 19386 17010
rect 19386 16958 19412 17010
rect 19116 16956 19172 16958
rect 19196 16956 19252 16958
rect 19276 16956 19332 16958
rect 19356 16956 19412 16958
rect 19116 15922 19172 15924
rect 19196 15922 19252 15924
rect 19276 15922 19332 15924
rect 19356 15922 19412 15924
rect 19116 15870 19142 15922
rect 19142 15870 19172 15922
rect 19196 15870 19206 15922
rect 19206 15870 19252 15922
rect 19276 15870 19322 15922
rect 19322 15870 19332 15922
rect 19356 15870 19386 15922
rect 19386 15870 19412 15922
rect 19116 15868 19172 15870
rect 19196 15868 19252 15870
rect 19276 15868 19332 15870
rect 19356 15868 19412 15870
rect 24116 33874 24172 33876
rect 24196 33874 24252 33876
rect 24276 33874 24332 33876
rect 24356 33874 24412 33876
rect 24116 33822 24142 33874
rect 24142 33822 24172 33874
rect 24196 33822 24206 33874
rect 24206 33822 24252 33874
rect 24276 33822 24322 33874
rect 24322 33822 24332 33874
rect 24356 33822 24386 33874
rect 24386 33822 24412 33874
rect 24116 33820 24172 33822
rect 24196 33820 24252 33822
rect 24276 33820 24332 33822
rect 24356 33820 24412 33822
rect 24116 32786 24172 32788
rect 24196 32786 24252 32788
rect 24276 32786 24332 32788
rect 24356 32786 24412 32788
rect 24116 32734 24142 32786
rect 24142 32734 24172 32786
rect 24196 32734 24206 32786
rect 24206 32734 24252 32786
rect 24276 32734 24322 32786
rect 24322 32734 24332 32786
rect 24356 32734 24386 32786
rect 24386 32734 24412 32786
rect 24116 32732 24172 32734
rect 24196 32732 24252 32734
rect 24276 32732 24332 32734
rect 24356 32732 24412 32734
rect 24116 31698 24172 31700
rect 24196 31698 24252 31700
rect 24276 31698 24332 31700
rect 24356 31698 24412 31700
rect 24116 31646 24142 31698
rect 24142 31646 24172 31698
rect 24196 31646 24206 31698
rect 24206 31646 24252 31698
rect 24276 31646 24322 31698
rect 24322 31646 24332 31698
rect 24356 31646 24386 31698
rect 24386 31646 24412 31698
rect 24116 31644 24172 31646
rect 24196 31644 24252 31646
rect 24276 31644 24332 31646
rect 24356 31644 24412 31646
rect 22518 24776 22574 24832
rect 24116 30610 24172 30612
rect 24196 30610 24252 30612
rect 24276 30610 24332 30612
rect 24356 30610 24412 30612
rect 24116 30558 24142 30610
rect 24142 30558 24172 30610
rect 24196 30558 24206 30610
rect 24206 30558 24252 30610
rect 24276 30558 24322 30610
rect 24322 30558 24332 30610
rect 24356 30558 24386 30610
rect 24386 30558 24412 30610
rect 24116 30556 24172 30558
rect 24196 30556 24252 30558
rect 24276 30556 24332 30558
rect 24356 30556 24412 30558
rect 24116 29522 24172 29524
rect 24196 29522 24252 29524
rect 24276 29522 24332 29524
rect 24356 29522 24412 29524
rect 24116 29470 24142 29522
rect 24142 29470 24172 29522
rect 24196 29470 24206 29522
rect 24206 29470 24252 29522
rect 24276 29470 24322 29522
rect 24322 29470 24332 29522
rect 24356 29470 24386 29522
rect 24386 29470 24412 29522
rect 24116 29468 24172 29470
rect 24196 29468 24252 29470
rect 24276 29468 24332 29470
rect 24356 29468 24412 29470
rect 24116 28434 24172 28436
rect 24196 28434 24252 28436
rect 24276 28434 24332 28436
rect 24356 28434 24412 28436
rect 24116 28382 24142 28434
rect 24142 28382 24172 28434
rect 24196 28382 24206 28434
rect 24206 28382 24252 28434
rect 24276 28382 24322 28434
rect 24322 28382 24332 28434
rect 24356 28382 24386 28434
rect 24386 28382 24412 28434
rect 24116 28380 24172 28382
rect 24196 28380 24252 28382
rect 24276 28380 24332 28382
rect 24356 28380 24412 28382
rect 24116 27346 24172 27348
rect 24196 27346 24252 27348
rect 24276 27346 24332 27348
rect 24356 27346 24412 27348
rect 24116 27294 24142 27346
rect 24142 27294 24172 27346
rect 24196 27294 24206 27346
rect 24206 27294 24252 27346
rect 24276 27294 24322 27346
rect 24322 27294 24332 27346
rect 24356 27294 24386 27346
rect 24386 27294 24412 27346
rect 24116 27292 24172 27294
rect 24196 27292 24252 27294
rect 24276 27292 24332 27294
rect 24356 27292 24412 27294
rect 24116 26258 24172 26260
rect 24196 26258 24252 26260
rect 24276 26258 24332 26260
rect 24356 26258 24412 26260
rect 24116 26206 24142 26258
rect 24142 26206 24172 26258
rect 24196 26206 24206 26258
rect 24206 26206 24252 26258
rect 24276 26206 24322 26258
rect 24322 26206 24332 26258
rect 24356 26206 24386 26258
rect 24386 26206 24412 26258
rect 24116 26204 24172 26206
rect 24196 26204 24252 26206
rect 24276 26204 24332 26206
rect 24356 26204 24412 26206
rect 24116 25170 24172 25172
rect 24196 25170 24252 25172
rect 24276 25170 24332 25172
rect 24356 25170 24412 25172
rect 24116 25118 24142 25170
rect 24142 25118 24172 25170
rect 24196 25118 24206 25170
rect 24206 25118 24252 25170
rect 24276 25118 24322 25170
rect 24322 25118 24332 25170
rect 24356 25118 24386 25170
rect 24386 25118 24412 25170
rect 24116 25116 24172 25118
rect 24196 25116 24252 25118
rect 24276 25116 24332 25118
rect 24356 25116 24412 25118
rect 24116 24082 24172 24084
rect 24196 24082 24252 24084
rect 24276 24082 24332 24084
rect 24356 24082 24412 24084
rect 24116 24030 24142 24082
rect 24142 24030 24172 24082
rect 24196 24030 24206 24082
rect 24206 24030 24252 24082
rect 24276 24030 24322 24082
rect 24322 24030 24332 24082
rect 24356 24030 24386 24082
rect 24386 24030 24412 24082
rect 24116 24028 24172 24030
rect 24196 24028 24252 24030
rect 24276 24028 24332 24030
rect 24356 24028 24412 24030
rect 24116 22994 24172 22996
rect 24196 22994 24252 22996
rect 24276 22994 24332 22996
rect 24356 22994 24412 22996
rect 24116 22942 24142 22994
rect 24142 22942 24172 22994
rect 24196 22942 24206 22994
rect 24206 22942 24252 22994
rect 24276 22942 24322 22994
rect 24322 22942 24332 22994
rect 24356 22942 24386 22994
rect 24386 22942 24412 22994
rect 24116 22940 24172 22942
rect 24196 22940 24252 22942
rect 24276 22940 24332 22942
rect 24356 22940 24412 22942
rect 24116 21906 24172 21908
rect 24196 21906 24252 21908
rect 24276 21906 24332 21908
rect 24356 21906 24412 21908
rect 24116 21854 24142 21906
rect 24142 21854 24172 21906
rect 24196 21854 24206 21906
rect 24206 21854 24252 21906
rect 24276 21854 24322 21906
rect 24322 21854 24332 21906
rect 24356 21854 24386 21906
rect 24386 21854 24412 21906
rect 24116 21852 24172 21854
rect 24196 21852 24252 21854
rect 24276 21852 24332 21854
rect 24356 21852 24412 21854
rect 24116 20818 24172 20820
rect 24196 20818 24252 20820
rect 24276 20818 24332 20820
rect 24356 20818 24412 20820
rect 24116 20766 24142 20818
rect 24142 20766 24172 20818
rect 24196 20766 24206 20818
rect 24206 20766 24252 20818
rect 24276 20766 24322 20818
rect 24322 20766 24332 20818
rect 24356 20766 24386 20818
rect 24386 20766 24412 20818
rect 24116 20764 24172 20766
rect 24196 20764 24252 20766
rect 24276 20764 24332 20766
rect 24356 20764 24412 20766
rect 19116 14834 19172 14836
rect 19196 14834 19252 14836
rect 19276 14834 19332 14836
rect 19356 14834 19412 14836
rect 19116 14782 19142 14834
rect 19142 14782 19172 14834
rect 19196 14782 19206 14834
rect 19206 14782 19252 14834
rect 19276 14782 19322 14834
rect 19322 14782 19332 14834
rect 19356 14782 19386 14834
rect 19386 14782 19412 14834
rect 19116 14780 19172 14782
rect 19196 14780 19252 14782
rect 19276 14780 19332 14782
rect 19356 14780 19412 14782
rect 19116 13746 19172 13748
rect 19196 13746 19252 13748
rect 19276 13746 19332 13748
rect 19356 13746 19412 13748
rect 19116 13694 19142 13746
rect 19142 13694 19172 13746
rect 19196 13694 19206 13746
rect 19206 13694 19252 13746
rect 19276 13694 19322 13746
rect 19322 13694 19332 13746
rect 19356 13694 19386 13746
rect 19386 13694 19412 13746
rect 19116 13692 19172 13694
rect 19196 13692 19252 13694
rect 19276 13692 19332 13694
rect 19356 13692 19412 13694
rect 19116 12658 19172 12660
rect 19196 12658 19252 12660
rect 19276 12658 19332 12660
rect 19356 12658 19412 12660
rect 19116 12606 19142 12658
rect 19142 12606 19172 12658
rect 19196 12606 19206 12658
rect 19206 12606 19252 12658
rect 19276 12606 19322 12658
rect 19322 12606 19332 12658
rect 19356 12606 19386 12658
rect 19386 12606 19412 12658
rect 19116 12604 19172 12606
rect 19196 12604 19252 12606
rect 19276 12604 19332 12606
rect 19356 12604 19412 12606
rect 19116 11570 19172 11572
rect 19196 11570 19252 11572
rect 19276 11570 19332 11572
rect 19356 11570 19412 11572
rect 19116 11518 19142 11570
rect 19142 11518 19172 11570
rect 19196 11518 19206 11570
rect 19206 11518 19252 11570
rect 19276 11518 19322 11570
rect 19322 11518 19332 11570
rect 19356 11518 19386 11570
rect 19386 11518 19412 11570
rect 19116 11516 19172 11518
rect 19196 11516 19252 11518
rect 19276 11516 19332 11518
rect 19356 11516 19412 11518
rect 24116 19730 24172 19732
rect 24196 19730 24252 19732
rect 24276 19730 24332 19732
rect 24356 19730 24412 19732
rect 24116 19678 24142 19730
rect 24142 19678 24172 19730
rect 24196 19678 24206 19730
rect 24206 19678 24252 19730
rect 24276 19678 24322 19730
rect 24322 19678 24332 19730
rect 24356 19678 24386 19730
rect 24386 19678 24412 19730
rect 24116 19676 24172 19678
rect 24196 19676 24252 19678
rect 24276 19676 24332 19678
rect 24356 19676 24412 19678
rect 24116 18642 24172 18644
rect 24196 18642 24252 18644
rect 24276 18642 24332 18644
rect 24356 18642 24412 18644
rect 24116 18590 24142 18642
rect 24142 18590 24172 18642
rect 24196 18590 24206 18642
rect 24206 18590 24252 18642
rect 24276 18590 24322 18642
rect 24322 18590 24332 18642
rect 24356 18590 24386 18642
rect 24386 18590 24412 18642
rect 24116 18588 24172 18590
rect 24196 18588 24252 18590
rect 24276 18588 24332 18590
rect 24356 18588 24412 18590
rect 24116 17554 24172 17556
rect 24196 17554 24252 17556
rect 24276 17554 24332 17556
rect 24356 17554 24412 17556
rect 24116 17502 24142 17554
rect 24142 17502 24172 17554
rect 24196 17502 24206 17554
rect 24206 17502 24252 17554
rect 24276 17502 24322 17554
rect 24322 17502 24332 17554
rect 24356 17502 24386 17554
rect 24386 17502 24412 17554
rect 24116 17500 24172 17502
rect 24196 17500 24252 17502
rect 24276 17500 24332 17502
rect 24356 17500 24412 17502
rect 24116 16466 24172 16468
rect 24196 16466 24252 16468
rect 24276 16466 24332 16468
rect 24356 16466 24412 16468
rect 24116 16414 24142 16466
rect 24142 16414 24172 16466
rect 24196 16414 24206 16466
rect 24206 16414 24252 16466
rect 24276 16414 24322 16466
rect 24322 16414 24332 16466
rect 24356 16414 24386 16466
rect 24386 16414 24412 16466
rect 24116 16412 24172 16414
rect 24196 16412 24252 16414
rect 24276 16412 24332 16414
rect 24356 16412 24412 16414
rect 24116 15378 24172 15380
rect 24196 15378 24252 15380
rect 24276 15378 24332 15380
rect 24356 15378 24412 15380
rect 24116 15326 24142 15378
rect 24142 15326 24172 15378
rect 24196 15326 24206 15378
rect 24206 15326 24252 15378
rect 24276 15326 24322 15378
rect 24322 15326 24332 15378
rect 24356 15326 24386 15378
rect 24386 15326 24412 15378
rect 24116 15324 24172 15326
rect 24196 15324 24252 15326
rect 24276 15324 24332 15326
rect 24356 15324 24412 15326
rect 24116 14290 24172 14292
rect 24196 14290 24252 14292
rect 24276 14290 24332 14292
rect 24356 14290 24412 14292
rect 24116 14238 24142 14290
rect 24142 14238 24172 14290
rect 24196 14238 24206 14290
rect 24206 14238 24252 14290
rect 24276 14238 24322 14290
rect 24322 14238 24332 14290
rect 24356 14238 24386 14290
rect 24386 14238 24412 14290
rect 24116 14236 24172 14238
rect 24196 14236 24252 14238
rect 24276 14236 24332 14238
rect 24356 14236 24412 14238
rect 24116 13202 24172 13204
rect 24196 13202 24252 13204
rect 24276 13202 24332 13204
rect 24356 13202 24412 13204
rect 24116 13150 24142 13202
rect 24142 13150 24172 13202
rect 24196 13150 24206 13202
rect 24206 13150 24252 13202
rect 24276 13150 24322 13202
rect 24322 13150 24332 13202
rect 24356 13150 24386 13202
rect 24386 13150 24412 13202
rect 24116 13148 24172 13150
rect 24196 13148 24252 13150
rect 24276 13148 24332 13150
rect 24356 13148 24412 13150
rect 24116 12114 24172 12116
rect 24196 12114 24252 12116
rect 24276 12114 24332 12116
rect 24356 12114 24412 12116
rect 24116 12062 24142 12114
rect 24142 12062 24172 12114
rect 24196 12062 24206 12114
rect 24206 12062 24252 12114
rect 24276 12062 24322 12114
rect 24322 12062 24332 12114
rect 24356 12062 24386 12114
rect 24386 12062 24412 12114
rect 24116 12060 24172 12062
rect 24196 12060 24252 12062
rect 24276 12060 24332 12062
rect 24356 12060 24412 12062
rect 25922 22756 25978 22792
rect 25922 22736 25924 22756
rect 25924 22736 25976 22756
rect 25976 22736 25978 22756
rect 29116 34418 29172 34420
rect 29196 34418 29252 34420
rect 29276 34418 29332 34420
rect 29356 34418 29412 34420
rect 29116 34366 29142 34418
rect 29142 34366 29172 34418
rect 29196 34366 29206 34418
rect 29206 34366 29252 34418
rect 29276 34366 29322 34418
rect 29322 34366 29332 34418
rect 29356 34366 29386 34418
rect 29386 34366 29412 34418
rect 29116 34364 29172 34366
rect 29196 34364 29252 34366
rect 29276 34364 29332 34366
rect 29356 34364 29412 34366
rect 26474 24776 26530 24832
rect 31074 33888 31130 33944
rect 29116 33330 29172 33332
rect 29196 33330 29252 33332
rect 29276 33330 29332 33332
rect 29356 33330 29412 33332
rect 29116 33278 29142 33330
rect 29142 33278 29172 33330
rect 29196 33278 29206 33330
rect 29206 33278 29252 33330
rect 29276 33278 29322 33330
rect 29322 33278 29332 33330
rect 29356 33278 29386 33330
rect 29386 33278 29412 33330
rect 29116 33276 29172 33278
rect 29196 33276 29252 33278
rect 29276 33276 29332 33278
rect 29356 33276 29412 33278
rect 29116 32242 29172 32244
rect 29196 32242 29252 32244
rect 29276 32242 29332 32244
rect 29356 32242 29412 32244
rect 29116 32190 29142 32242
rect 29142 32190 29172 32242
rect 29196 32190 29206 32242
rect 29206 32190 29252 32242
rect 29276 32190 29322 32242
rect 29322 32190 29332 32242
rect 29356 32190 29386 32242
rect 29386 32190 29412 32242
rect 29116 32188 29172 32190
rect 29196 32188 29252 32190
rect 29276 32188 29332 32190
rect 29356 32188 29412 32190
rect 29116 31154 29172 31156
rect 29196 31154 29252 31156
rect 29276 31154 29332 31156
rect 29356 31154 29412 31156
rect 29116 31102 29142 31154
rect 29142 31102 29172 31154
rect 29196 31102 29206 31154
rect 29206 31102 29252 31154
rect 29276 31102 29322 31154
rect 29322 31102 29332 31154
rect 29356 31102 29386 31154
rect 29386 31102 29412 31154
rect 29116 31100 29172 31102
rect 29196 31100 29252 31102
rect 29276 31100 29332 31102
rect 29356 31100 29412 31102
rect 29116 30066 29172 30068
rect 29196 30066 29252 30068
rect 29276 30066 29332 30068
rect 29356 30066 29412 30068
rect 29116 30014 29142 30066
rect 29142 30014 29172 30066
rect 29196 30014 29206 30066
rect 29206 30014 29252 30066
rect 29276 30014 29322 30066
rect 29322 30014 29332 30066
rect 29356 30014 29386 30066
rect 29386 30014 29412 30066
rect 29116 30012 29172 30014
rect 29196 30012 29252 30014
rect 29276 30012 29332 30014
rect 29356 30012 29412 30014
rect 29116 28978 29172 28980
rect 29196 28978 29252 28980
rect 29276 28978 29332 28980
rect 29356 28978 29412 28980
rect 29116 28926 29142 28978
rect 29142 28926 29172 28978
rect 29196 28926 29206 28978
rect 29206 28926 29252 28978
rect 29276 28926 29322 28978
rect 29322 28926 29332 28978
rect 29356 28926 29386 28978
rect 29386 28926 29412 28978
rect 29116 28924 29172 28926
rect 29196 28924 29252 28926
rect 29276 28924 29332 28926
rect 29356 28924 29412 28926
rect 27946 24796 28002 24832
rect 27946 24776 27948 24796
rect 27948 24776 28000 24796
rect 28000 24776 28002 24796
rect 24116 11026 24172 11028
rect 24196 11026 24252 11028
rect 24276 11026 24332 11028
rect 24356 11026 24412 11028
rect 24116 10974 24142 11026
rect 24142 10974 24172 11026
rect 24196 10974 24206 11026
rect 24206 10974 24252 11026
rect 24276 10974 24322 11026
rect 24322 10974 24332 11026
rect 24356 10974 24386 11026
rect 24386 10974 24412 11026
rect 24116 10972 24172 10974
rect 24196 10972 24252 10974
rect 24276 10972 24332 10974
rect 24356 10972 24412 10974
rect 29116 27890 29172 27892
rect 29196 27890 29252 27892
rect 29276 27890 29332 27892
rect 29356 27890 29412 27892
rect 29116 27838 29142 27890
rect 29142 27838 29172 27890
rect 29196 27838 29206 27890
rect 29206 27838 29252 27890
rect 29276 27838 29322 27890
rect 29322 27838 29332 27890
rect 29356 27838 29386 27890
rect 29386 27838 29412 27890
rect 29116 27836 29172 27838
rect 29196 27836 29252 27838
rect 29276 27836 29332 27838
rect 29356 27836 29412 27838
rect 31810 30624 31866 30680
rect 31258 27360 31314 27416
rect 29116 26802 29172 26804
rect 29196 26802 29252 26804
rect 29276 26802 29332 26804
rect 29356 26802 29412 26804
rect 29116 26750 29142 26802
rect 29142 26750 29172 26802
rect 29196 26750 29206 26802
rect 29206 26750 29252 26802
rect 29276 26750 29322 26802
rect 29322 26750 29332 26802
rect 29356 26750 29386 26802
rect 29386 26750 29412 26802
rect 29116 26748 29172 26750
rect 29196 26748 29252 26750
rect 29276 26748 29332 26750
rect 29356 26748 29412 26750
rect 29116 25714 29172 25716
rect 29196 25714 29252 25716
rect 29276 25714 29332 25716
rect 29356 25714 29412 25716
rect 29116 25662 29142 25714
rect 29142 25662 29172 25714
rect 29196 25662 29206 25714
rect 29206 25662 29252 25714
rect 29276 25662 29322 25714
rect 29322 25662 29332 25714
rect 29356 25662 29386 25714
rect 29386 25662 29412 25714
rect 29116 25660 29172 25662
rect 29196 25660 29252 25662
rect 29276 25660 29332 25662
rect 29356 25660 29412 25662
rect 29116 24626 29172 24628
rect 29196 24626 29252 24628
rect 29276 24626 29332 24628
rect 29356 24626 29412 24628
rect 29116 24574 29142 24626
rect 29142 24574 29172 24626
rect 29196 24574 29206 24626
rect 29206 24574 29252 24626
rect 29276 24574 29322 24626
rect 29322 24574 29332 24626
rect 29356 24574 29386 24626
rect 29386 24574 29412 24626
rect 29116 24572 29172 24574
rect 29196 24572 29252 24574
rect 29276 24572 29332 24574
rect 29356 24572 29412 24574
rect 29116 23538 29172 23540
rect 29196 23538 29252 23540
rect 29276 23538 29332 23540
rect 29356 23538 29412 23540
rect 29116 23486 29142 23538
rect 29142 23486 29172 23538
rect 29196 23486 29206 23538
rect 29206 23486 29252 23538
rect 29276 23486 29322 23538
rect 29322 23486 29332 23538
rect 29356 23486 29386 23538
rect 29386 23486 29412 23538
rect 29116 23484 29172 23486
rect 29196 23484 29252 23486
rect 29276 23484 29332 23486
rect 29356 23484 29412 23486
rect 29116 22450 29172 22452
rect 29196 22450 29252 22452
rect 29276 22450 29332 22452
rect 29356 22450 29412 22452
rect 29116 22398 29142 22450
rect 29142 22398 29172 22450
rect 29196 22398 29206 22450
rect 29206 22398 29252 22450
rect 29276 22398 29322 22450
rect 29322 22398 29332 22450
rect 29356 22398 29386 22450
rect 29386 22398 29412 22450
rect 29116 22396 29172 22398
rect 29196 22396 29252 22398
rect 29276 22396 29332 22398
rect 29356 22396 29412 22398
rect 29116 21362 29172 21364
rect 29196 21362 29252 21364
rect 29276 21362 29332 21364
rect 29356 21362 29412 21364
rect 29116 21310 29142 21362
rect 29142 21310 29172 21362
rect 29196 21310 29206 21362
rect 29206 21310 29252 21362
rect 29276 21310 29322 21362
rect 29322 21310 29332 21362
rect 29356 21310 29386 21362
rect 29386 21310 29412 21362
rect 29116 21308 29172 21310
rect 29196 21308 29252 21310
rect 29276 21308 29332 21310
rect 29356 21308 29412 21310
rect 29116 20274 29172 20276
rect 29196 20274 29252 20276
rect 29276 20274 29332 20276
rect 29356 20274 29412 20276
rect 29116 20222 29142 20274
rect 29142 20222 29172 20274
rect 29196 20222 29206 20274
rect 29206 20222 29252 20274
rect 29276 20222 29322 20274
rect 29322 20222 29332 20274
rect 29356 20222 29386 20274
rect 29386 20222 29412 20274
rect 29116 20220 29172 20222
rect 29196 20220 29252 20222
rect 29276 20220 29332 20222
rect 29356 20220 29412 20222
rect 29116 19186 29172 19188
rect 29196 19186 29252 19188
rect 29276 19186 29332 19188
rect 29356 19186 29412 19188
rect 29116 19134 29142 19186
rect 29142 19134 29172 19186
rect 29196 19134 29206 19186
rect 29206 19134 29252 19186
rect 29276 19134 29322 19186
rect 29322 19134 29332 19186
rect 29356 19134 29386 19186
rect 29386 19134 29412 19186
rect 29116 19132 29172 19134
rect 29196 19132 29252 19134
rect 29276 19132 29332 19134
rect 29356 19132 29412 19134
rect 29116 18098 29172 18100
rect 29196 18098 29252 18100
rect 29276 18098 29332 18100
rect 29356 18098 29412 18100
rect 29116 18046 29142 18098
rect 29142 18046 29172 18098
rect 29196 18046 29206 18098
rect 29206 18046 29252 18098
rect 29276 18046 29322 18098
rect 29322 18046 29332 18098
rect 29356 18046 29386 18098
rect 29386 18046 29412 18098
rect 29116 18044 29172 18046
rect 29196 18044 29252 18046
rect 29276 18044 29332 18046
rect 29356 18044 29412 18046
rect 29116 17010 29172 17012
rect 29196 17010 29252 17012
rect 29276 17010 29332 17012
rect 29356 17010 29412 17012
rect 29116 16958 29142 17010
rect 29142 16958 29172 17010
rect 29196 16958 29206 17010
rect 29206 16958 29252 17010
rect 29276 16958 29322 17010
rect 29322 16958 29332 17010
rect 29356 16958 29386 17010
rect 29386 16958 29412 17010
rect 29116 16956 29172 16958
rect 29196 16956 29252 16958
rect 29276 16956 29332 16958
rect 29356 16956 29412 16958
rect 29116 15922 29172 15924
rect 29196 15922 29252 15924
rect 29276 15922 29332 15924
rect 29356 15922 29412 15924
rect 29116 15870 29142 15922
rect 29142 15870 29172 15922
rect 29196 15870 29206 15922
rect 29206 15870 29252 15922
rect 29276 15870 29322 15922
rect 29322 15870 29332 15922
rect 29356 15870 29386 15922
rect 29386 15870 29412 15922
rect 29116 15868 29172 15870
rect 29196 15868 29252 15870
rect 29276 15868 29332 15870
rect 29356 15868 29412 15870
rect 29116 14834 29172 14836
rect 29196 14834 29252 14836
rect 29276 14834 29332 14836
rect 29356 14834 29412 14836
rect 29116 14782 29142 14834
rect 29142 14782 29172 14834
rect 29196 14782 29206 14834
rect 29206 14782 29252 14834
rect 29276 14782 29322 14834
rect 29322 14782 29332 14834
rect 29356 14782 29386 14834
rect 29386 14782 29412 14834
rect 29116 14780 29172 14782
rect 29196 14780 29252 14782
rect 29276 14780 29332 14782
rect 29356 14780 29412 14782
rect 29116 13746 29172 13748
rect 29196 13746 29252 13748
rect 29276 13746 29332 13748
rect 29356 13746 29412 13748
rect 29116 13694 29142 13746
rect 29142 13694 29172 13746
rect 29196 13694 29206 13746
rect 29206 13694 29252 13746
rect 29276 13694 29322 13746
rect 29322 13694 29332 13746
rect 29356 13694 29386 13746
rect 29386 13694 29412 13746
rect 29116 13692 29172 13694
rect 29196 13692 29252 13694
rect 29276 13692 29332 13694
rect 29356 13692 29412 13694
rect 30614 23824 30670 23880
rect 32086 20560 32142 20616
rect 30614 17060 30616 17080
rect 30616 17060 30668 17080
rect 30668 17060 30670 17080
rect 30614 17024 30670 17060
rect 30706 13760 30762 13816
rect 29116 12658 29172 12660
rect 29196 12658 29252 12660
rect 29276 12658 29332 12660
rect 29356 12658 29412 12660
rect 29116 12606 29142 12658
rect 29142 12606 29172 12658
rect 29196 12606 29206 12658
rect 29206 12606 29252 12658
rect 29276 12606 29322 12658
rect 29322 12606 29332 12658
rect 29356 12606 29386 12658
rect 29386 12606 29412 12658
rect 29116 12604 29172 12606
rect 29196 12604 29252 12606
rect 29276 12604 29332 12606
rect 29356 12604 29412 12606
rect 29116 11570 29172 11572
rect 29196 11570 29252 11572
rect 29276 11570 29332 11572
rect 29356 11570 29412 11572
rect 29116 11518 29142 11570
rect 29142 11518 29172 11570
rect 29196 11518 29206 11570
rect 29206 11518 29252 11570
rect 29276 11518 29322 11570
rect 29322 11518 29332 11570
rect 29356 11518 29386 11570
rect 29386 11518 29412 11570
rect 29116 11516 29172 11518
rect 29196 11516 29252 11518
rect 29276 11516 29332 11518
rect 29356 11516 29412 11518
rect 30614 10496 30670 10552
<< metal3 >>
rect 0 45384 45368 45392
rect 0 45320 8 45384
rect 72 45320 88 45384
rect 152 45320 168 45384
rect 232 45320 248 45384
rect 312 45320 328 45384
rect 392 45320 408 45384
rect 472 45320 488 45384
rect 552 45320 568 45384
rect 632 45320 648 45384
rect 712 45320 728 45384
rect 792 45320 808 45384
rect 872 45320 888 45384
rect 952 45320 968 45384
rect 1032 45320 1048 45384
rect 1112 45320 1128 45384
rect 1192 45320 1208 45384
rect 1272 45320 1288 45384
rect 1352 45320 1368 45384
rect 1432 45320 1448 45384
rect 1512 45320 1528 45384
rect 1592 45320 1608 45384
rect 1672 45320 1688 45384
rect 1752 45320 1768 45384
rect 1832 45320 1848 45384
rect 1912 45320 1928 45384
rect 1992 45320 2008 45384
rect 2072 45320 2088 45384
rect 2152 45320 2168 45384
rect 2232 45320 2248 45384
rect 2312 45320 2328 45384
rect 2392 45320 2408 45384
rect 2472 45320 2488 45384
rect 2552 45320 2568 45384
rect 2632 45320 2648 45384
rect 2712 45320 2728 45384
rect 2792 45320 2808 45384
rect 2872 45320 2888 45384
rect 2952 45320 2968 45384
rect 3032 45320 3048 45384
rect 3112 45320 3128 45384
rect 3192 45320 3208 45384
rect 3272 45320 3288 45384
rect 3352 45320 3368 45384
rect 3432 45320 3448 45384
rect 3512 45320 3528 45384
rect 3592 45320 3608 45384
rect 3672 45320 3688 45384
rect 3752 45320 3768 45384
rect 3832 45320 3848 45384
rect 3912 45320 3928 45384
rect 3992 45320 19112 45384
rect 19176 45320 19192 45384
rect 19256 45320 19272 45384
rect 19336 45320 19352 45384
rect 19416 45320 29112 45384
rect 29176 45320 29192 45384
rect 29256 45320 29272 45384
rect 29336 45320 29352 45384
rect 29416 45320 41376 45384
rect 41440 45320 41456 45384
rect 41520 45320 41536 45384
rect 41600 45320 41616 45384
rect 41680 45320 41696 45384
rect 41760 45320 41776 45384
rect 41840 45320 41856 45384
rect 41920 45320 41936 45384
rect 42000 45320 42016 45384
rect 42080 45320 42096 45384
rect 42160 45320 42176 45384
rect 42240 45320 42256 45384
rect 42320 45320 42336 45384
rect 42400 45320 42416 45384
rect 42480 45320 42496 45384
rect 42560 45320 42576 45384
rect 42640 45320 42656 45384
rect 42720 45320 42736 45384
rect 42800 45320 42816 45384
rect 42880 45320 42896 45384
rect 42960 45320 42976 45384
rect 43040 45320 43056 45384
rect 43120 45320 43136 45384
rect 43200 45320 43216 45384
rect 43280 45320 43296 45384
rect 43360 45320 43376 45384
rect 43440 45320 43456 45384
rect 43520 45320 43536 45384
rect 43600 45320 43616 45384
rect 43680 45320 43696 45384
rect 43760 45320 43776 45384
rect 43840 45320 43856 45384
rect 43920 45320 43936 45384
rect 44000 45320 44016 45384
rect 44080 45320 44096 45384
rect 44160 45320 44176 45384
rect 44240 45320 44256 45384
rect 44320 45320 44336 45384
rect 44400 45320 44416 45384
rect 44480 45320 44496 45384
rect 44560 45320 44576 45384
rect 44640 45320 44656 45384
rect 44720 45320 44736 45384
rect 44800 45320 44816 45384
rect 44880 45320 44896 45384
rect 44960 45320 44976 45384
rect 45040 45320 45056 45384
rect 45120 45320 45136 45384
rect 45200 45320 45216 45384
rect 45280 45320 45296 45384
rect 45360 45320 45368 45384
rect 0 45304 45368 45320
rect 0 45240 8 45304
rect 72 45240 88 45304
rect 152 45240 168 45304
rect 232 45240 248 45304
rect 312 45240 328 45304
rect 392 45240 408 45304
rect 472 45240 488 45304
rect 552 45240 568 45304
rect 632 45240 648 45304
rect 712 45240 728 45304
rect 792 45240 808 45304
rect 872 45240 888 45304
rect 952 45240 968 45304
rect 1032 45240 1048 45304
rect 1112 45240 1128 45304
rect 1192 45240 1208 45304
rect 1272 45240 1288 45304
rect 1352 45240 1368 45304
rect 1432 45240 1448 45304
rect 1512 45240 1528 45304
rect 1592 45240 1608 45304
rect 1672 45240 1688 45304
rect 1752 45240 1768 45304
rect 1832 45240 1848 45304
rect 1912 45240 1928 45304
rect 1992 45240 2008 45304
rect 2072 45240 2088 45304
rect 2152 45240 2168 45304
rect 2232 45240 2248 45304
rect 2312 45240 2328 45304
rect 2392 45240 2408 45304
rect 2472 45240 2488 45304
rect 2552 45240 2568 45304
rect 2632 45240 2648 45304
rect 2712 45240 2728 45304
rect 2792 45240 2808 45304
rect 2872 45240 2888 45304
rect 2952 45240 2968 45304
rect 3032 45240 3048 45304
rect 3112 45240 3128 45304
rect 3192 45240 3208 45304
rect 3272 45240 3288 45304
rect 3352 45240 3368 45304
rect 3432 45240 3448 45304
rect 3512 45240 3528 45304
rect 3592 45240 3608 45304
rect 3672 45240 3688 45304
rect 3752 45240 3768 45304
rect 3832 45240 3848 45304
rect 3912 45240 3928 45304
rect 3992 45240 19112 45304
rect 19176 45240 19192 45304
rect 19256 45240 19272 45304
rect 19336 45240 19352 45304
rect 19416 45240 29112 45304
rect 29176 45240 29192 45304
rect 29256 45240 29272 45304
rect 29336 45240 29352 45304
rect 29416 45240 41376 45304
rect 41440 45240 41456 45304
rect 41520 45240 41536 45304
rect 41600 45240 41616 45304
rect 41680 45240 41696 45304
rect 41760 45240 41776 45304
rect 41840 45240 41856 45304
rect 41920 45240 41936 45304
rect 42000 45240 42016 45304
rect 42080 45240 42096 45304
rect 42160 45240 42176 45304
rect 42240 45240 42256 45304
rect 42320 45240 42336 45304
rect 42400 45240 42416 45304
rect 42480 45240 42496 45304
rect 42560 45240 42576 45304
rect 42640 45240 42656 45304
rect 42720 45240 42736 45304
rect 42800 45240 42816 45304
rect 42880 45240 42896 45304
rect 42960 45240 42976 45304
rect 43040 45240 43056 45304
rect 43120 45240 43136 45304
rect 43200 45240 43216 45304
rect 43280 45240 43296 45304
rect 43360 45240 43376 45304
rect 43440 45240 43456 45304
rect 43520 45240 43536 45304
rect 43600 45240 43616 45304
rect 43680 45240 43696 45304
rect 43760 45240 43776 45304
rect 43840 45240 43856 45304
rect 43920 45240 43936 45304
rect 44000 45240 44016 45304
rect 44080 45240 44096 45304
rect 44160 45240 44176 45304
rect 44240 45240 44256 45304
rect 44320 45240 44336 45304
rect 44400 45240 44416 45304
rect 44480 45240 44496 45304
rect 44560 45240 44576 45304
rect 44640 45240 44656 45304
rect 44720 45240 44736 45304
rect 44800 45240 44816 45304
rect 44880 45240 44896 45304
rect 44960 45240 44976 45304
rect 45040 45240 45056 45304
rect 45120 45240 45136 45304
rect 45200 45240 45216 45304
rect 45280 45240 45296 45304
rect 45360 45240 45368 45304
rect 0 45224 45368 45240
rect 0 45160 8 45224
rect 72 45160 88 45224
rect 152 45160 168 45224
rect 232 45160 248 45224
rect 312 45160 328 45224
rect 392 45160 408 45224
rect 472 45160 488 45224
rect 552 45160 568 45224
rect 632 45160 648 45224
rect 712 45160 728 45224
rect 792 45160 808 45224
rect 872 45160 888 45224
rect 952 45160 968 45224
rect 1032 45160 1048 45224
rect 1112 45160 1128 45224
rect 1192 45160 1208 45224
rect 1272 45160 1288 45224
rect 1352 45160 1368 45224
rect 1432 45160 1448 45224
rect 1512 45160 1528 45224
rect 1592 45160 1608 45224
rect 1672 45160 1688 45224
rect 1752 45160 1768 45224
rect 1832 45160 1848 45224
rect 1912 45160 1928 45224
rect 1992 45160 2008 45224
rect 2072 45160 2088 45224
rect 2152 45160 2168 45224
rect 2232 45160 2248 45224
rect 2312 45160 2328 45224
rect 2392 45160 2408 45224
rect 2472 45160 2488 45224
rect 2552 45160 2568 45224
rect 2632 45160 2648 45224
rect 2712 45160 2728 45224
rect 2792 45160 2808 45224
rect 2872 45160 2888 45224
rect 2952 45160 2968 45224
rect 3032 45160 3048 45224
rect 3112 45160 3128 45224
rect 3192 45160 3208 45224
rect 3272 45160 3288 45224
rect 3352 45160 3368 45224
rect 3432 45160 3448 45224
rect 3512 45160 3528 45224
rect 3592 45160 3608 45224
rect 3672 45160 3688 45224
rect 3752 45160 3768 45224
rect 3832 45160 3848 45224
rect 3912 45160 3928 45224
rect 3992 45160 19112 45224
rect 19176 45160 19192 45224
rect 19256 45160 19272 45224
rect 19336 45160 19352 45224
rect 19416 45160 29112 45224
rect 29176 45160 29192 45224
rect 29256 45160 29272 45224
rect 29336 45160 29352 45224
rect 29416 45160 41376 45224
rect 41440 45160 41456 45224
rect 41520 45160 41536 45224
rect 41600 45160 41616 45224
rect 41680 45160 41696 45224
rect 41760 45160 41776 45224
rect 41840 45160 41856 45224
rect 41920 45160 41936 45224
rect 42000 45160 42016 45224
rect 42080 45160 42096 45224
rect 42160 45160 42176 45224
rect 42240 45160 42256 45224
rect 42320 45160 42336 45224
rect 42400 45160 42416 45224
rect 42480 45160 42496 45224
rect 42560 45160 42576 45224
rect 42640 45160 42656 45224
rect 42720 45160 42736 45224
rect 42800 45160 42816 45224
rect 42880 45160 42896 45224
rect 42960 45160 42976 45224
rect 43040 45160 43056 45224
rect 43120 45160 43136 45224
rect 43200 45160 43216 45224
rect 43280 45160 43296 45224
rect 43360 45160 43376 45224
rect 43440 45160 43456 45224
rect 43520 45160 43536 45224
rect 43600 45160 43616 45224
rect 43680 45160 43696 45224
rect 43760 45160 43776 45224
rect 43840 45160 43856 45224
rect 43920 45160 43936 45224
rect 44000 45160 44016 45224
rect 44080 45160 44096 45224
rect 44160 45160 44176 45224
rect 44240 45160 44256 45224
rect 44320 45160 44336 45224
rect 44400 45160 44416 45224
rect 44480 45160 44496 45224
rect 44560 45160 44576 45224
rect 44640 45160 44656 45224
rect 44720 45160 44736 45224
rect 44800 45160 44816 45224
rect 44880 45160 44896 45224
rect 44960 45160 44976 45224
rect 45040 45160 45056 45224
rect 45120 45160 45136 45224
rect 45200 45160 45216 45224
rect 45280 45160 45296 45224
rect 45360 45160 45368 45224
rect 0 45144 45368 45160
rect 0 45080 8 45144
rect 72 45080 88 45144
rect 152 45080 168 45144
rect 232 45080 248 45144
rect 312 45080 328 45144
rect 392 45080 408 45144
rect 472 45080 488 45144
rect 552 45080 568 45144
rect 632 45080 648 45144
rect 712 45080 728 45144
rect 792 45080 808 45144
rect 872 45080 888 45144
rect 952 45080 968 45144
rect 1032 45080 1048 45144
rect 1112 45080 1128 45144
rect 1192 45080 1208 45144
rect 1272 45080 1288 45144
rect 1352 45080 1368 45144
rect 1432 45080 1448 45144
rect 1512 45080 1528 45144
rect 1592 45080 1608 45144
rect 1672 45080 1688 45144
rect 1752 45080 1768 45144
rect 1832 45080 1848 45144
rect 1912 45080 1928 45144
rect 1992 45080 2008 45144
rect 2072 45080 2088 45144
rect 2152 45080 2168 45144
rect 2232 45080 2248 45144
rect 2312 45080 2328 45144
rect 2392 45080 2408 45144
rect 2472 45080 2488 45144
rect 2552 45080 2568 45144
rect 2632 45080 2648 45144
rect 2712 45080 2728 45144
rect 2792 45080 2808 45144
rect 2872 45080 2888 45144
rect 2952 45080 2968 45144
rect 3032 45080 3048 45144
rect 3112 45080 3128 45144
rect 3192 45080 3208 45144
rect 3272 45080 3288 45144
rect 3352 45080 3368 45144
rect 3432 45080 3448 45144
rect 3512 45080 3528 45144
rect 3592 45080 3608 45144
rect 3672 45080 3688 45144
rect 3752 45080 3768 45144
rect 3832 45080 3848 45144
rect 3912 45080 3928 45144
rect 3992 45080 19112 45144
rect 19176 45080 19192 45144
rect 19256 45080 19272 45144
rect 19336 45080 19352 45144
rect 19416 45080 29112 45144
rect 29176 45080 29192 45144
rect 29256 45080 29272 45144
rect 29336 45080 29352 45144
rect 29416 45080 41376 45144
rect 41440 45080 41456 45144
rect 41520 45080 41536 45144
rect 41600 45080 41616 45144
rect 41680 45080 41696 45144
rect 41760 45080 41776 45144
rect 41840 45080 41856 45144
rect 41920 45080 41936 45144
rect 42000 45080 42016 45144
rect 42080 45080 42096 45144
rect 42160 45080 42176 45144
rect 42240 45080 42256 45144
rect 42320 45080 42336 45144
rect 42400 45080 42416 45144
rect 42480 45080 42496 45144
rect 42560 45080 42576 45144
rect 42640 45080 42656 45144
rect 42720 45080 42736 45144
rect 42800 45080 42816 45144
rect 42880 45080 42896 45144
rect 42960 45080 42976 45144
rect 43040 45080 43056 45144
rect 43120 45080 43136 45144
rect 43200 45080 43216 45144
rect 43280 45080 43296 45144
rect 43360 45080 43376 45144
rect 43440 45080 43456 45144
rect 43520 45080 43536 45144
rect 43600 45080 43616 45144
rect 43680 45080 43696 45144
rect 43760 45080 43776 45144
rect 43840 45080 43856 45144
rect 43920 45080 43936 45144
rect 44000 45080 44016 45144
rect 44080 45080 44096 45144
rect 44160 45080 44176 45144
rect 44240 45080 44256 45144
rect 44320 45080 44336 45144
rect 44400 45080 44416 45144
rect 44480 45080 44496 45144
rect 44560 45080 44576 45144
rect 44640 45080 44656 45144
rect 44720 45080 44736 45144
rect 44800 45080 44816 45144
rect 44880 45080 44896 45144
rect 44960 45080 44976 45144
rect 45040 45080 45056 45144
rect 45120 45080 45136 45144
rect 45200 45080 45216 45144
rect 45280 45080 45296 45144
rect 45360 45080 45368 45144
rect 0 45064 45368 45080
rect 0 45000 8 45064
rect 72 45000 88 45064
rect 152 45000 168 45064
rect 232 45000 248 45064
rect 312 45000 328 45064
rect 392 45000 408 45064
rect 472 45000 488 45064
rect 552 45000 568 45064
rect 632 45000 648 45064
rect 712 45000 728 45064
rect 792 45000 808 45064
rect 872 45000 888 45064
rect 952 45000 968 45064
rect 1032 45000 1048 45064
rect 1112 45000 1128 45064
rect 1192 45000 1208 45064
rect 1272 45000 1288 45064
rect 1352 45000 1368 45064
rect 1432 45000 1448 45064
rect 1512 45000 1528 45064
rect 1592 45000 1608 45064
rect 1672 45000 1688 45064
rect 1752 45000 1768 45064
rect 1832 45000 1848 45064
rect 1912 45000 1928 45064
rect 1992 45000 2008 45064
rect 2072 45000 2088 45064
rect 2152 45000 2168 45064
rect 2232 45000 2248 45064
rect 2312 45000 2328 45064
rect 2392 45000 2408 45064
rect 2472 45000 2488 45064
rect 2552 45000 2568 45064
rect 2632 45000 2648 45064
rect 2712 45000 2728 45064
rect 2792 45000 2808 45064
rect 2872 45000 2888 45064
rect 2952 45000 2968 45064
rect 3032 45000 3048 45064
rect 3112 45000 3128 45064
rect 3192 45000 3208 45064
rect 3272 45000 3288 45064
rect 3352 45000 3368 45064
rect 3432 45000 3448 45064
rect 3512 45000 3528 45064
rect 3592 45000 3608 45064
rect 3672 45000 3688 45064
rect 3752 45000 3768 45064
rect 3832 45000 3848 45064
rect 3912 45000 3928 45064
rect 3992 45000 19112 45064
rect 19176 45000 19192 45064
rect 19256 45000 19272 45064
rect 19336 45000 19352 45064
rect 19416 45000 29112 45064
rect 29176 45000 29192 45064
rect 29256 45000 29272 45064
rect 29336 45000 29352 45064
rect 29416 45000 41376 45064
rect 41440 45000 41456 45064
rect 41520 45000 41536 45064
rect 41600 45000 41616 45064
rect 41680 45000 41696 45064
rect 41760 45000 41776 45064
rect 41840 45000 41856 45064
rect 41920 45000 41936 45064
rect 42000 45000 42016 45064
rect 42080 45000 42096 45064
rect 42160 45000 42176 45064
rect 42240 45000 42256 45064
rect 42320 45000 42336 45064
rect 42400 45000 42416 45064
rect 42480 45000 42496 45064
rect 42560 45000 42576 45064
rect 42640 45000 42656 45064
rect 42720 45000 42736 45064
rect 42800 45000 42816 45064
rect 42880 45000 42896 45064
rect 42960 45000 42976 45064
rect 43040 45000 43056 45064
rect 43120 45000 43136 45064
rect 43200 45000 43216 45064
rect 43280 45000 43296 45064
rect 43360 45000 43376 45064
rect 43440 45000 43456 45064
rect 43520 45000 43536 45064
rect 43600 45000 43616 45064
rect 43680 45000 43696 45064
rect 43760 45000 43776 45064
rect 43840 45000 43856 45064
rect 43920 45000 43936 45064
rect 44000 45000 44016 45064
rect 44080 45000 44096 45064
rect 44160 45000 44176 45064
rect 44240 45000 44256 45064
rect 44320 45000 44336 45064
rect 44400 45000 44416 45064
rect 44480 45000 44496 45064
rect 44560 45000 44576 45064
rect 44640 45000 44656 45064
rect 44720 45000 44736 45064
rect 44800 45000 44816 45064
rect 44880 45000 44896 45064
rect 44960 45000 44976 45064
rect 45040 45000 45056 45064
rect 45120 45000 45136 45064
rect 45200 45000 45216 45064
rect 45280 45000 45296 45064
rect 45360 45000 45368 45064
rect 0 44984 45368 45000
rect 0 44920 8 44984
rect 72 44920 88 44984
rect 152 44920 168 44984
rect 232 44920 248 44984
rect 312 44920 328 44984
rect 392 44920 408 44984
rect 472 44920 488 44984
rect 552 44920 568 44984
rect 632 44920 648 44984
rect 712 44920 728 44984
rect 792 44920 808 44984
rect 872 44920 888 44984
rect 952 44920 968 44984
rect 1032 44920 1048 44984
rect 1112 44920 1128 44984
rect 1192 44920 1208 44984
rect 1272 44920 1288 44984
rect 1352 44920 1368 44984
rect 1432 44920 1448 44984
rect 1512 44920 1528 44984
rect 1592 44920 1608 44984
rect 1672 44920 1688 44984
rect 1752 44920 1768 44984
rect 1832 44920 1848 44984
rect 1912 44920 1928 44984
rect 1992 44920 2008 44984
rect 2072 44920 2088 44984
rect 2152 44920 2168 44984
rect 2232 44920 2248 44984
rect 2312 44920 2328 44984
rect 2392 44920 2408 44984
rect 2472 44920 2488 44984
rect 2552 44920 2568 44984
rect 2632 44920 2648 44984
rect 2712 44920 2728 44984
rect 2792 44920 2808 44984
rect 2872 44920 2888 44984
rect 2952 44920 2968 44984
rect 3032 44920 3048 44984
rect 3112 44920 3128 44984
rect 3192 44920 3208 44984
rect 3272 44920 3288 44984
rect 3352 44920 3368 44984
rect 3432 44920 3448 44984
rect 3512 44920 3528 44984
rect 3592 44920 3608 44984
rect 3672 44920 3688 44984
rect 3752 44920 3768 44984
rect 3832 44920 3848 44984
rect 3912 44920 3928 44984
rect 3992 44920 19112 44984
rect 19176 44920 19192 44984
rect 19256 44920 19272 44984
rect 19336 44920 19352 44984
rect 19416 44920 29112 44984
rect 29176 44920 29192 44984
rect 29256 44920 29272 44984
rect 29336 44920 29352 44984
rect 29416 44920 41376 44984
rect 41440 44920 41456 44984
rect 41520 44920 41536 44984
rect 41600 44920 41616 44984
rect 41680 44920 41696 44984
rect 41760 44920 41776 44984
rect 41840 44920 41856 44984
rect 41920 44920 41936 44984
rect 42000 44920 42016 44984
rect 42080 44920 42096 44984
rect 42160 44920 42176 44984
rect 42240 44920 42256 44984
rect 42320 44920 42336 44984
rect 42400 44920 42416 44984
rect 42480 44920 42496 44984
rect 42560 44920 42576 44984
rect 42640 44920 42656 44984
rect 42720 44920 42736 44984
rect 42800 44920 42816 44984
rect 42880 44920 42896 44984
rect 42960 44920 42976 44984
rect 43040 44920 43056 44984
rect 43120 44920 43136 44984
rect 43200 44920 43216 44984
rect 43280 44920 43296 44984
rect 43360 44920 43376 44984
rect 43440 44920 43456 44984
rect 43520 44920 43536 44984
rect 43600 44920 43616 44984
rect 43680 44920 43696 44984
rect 43760 44920 43776 44984
rect 43840 44920 43856 44984
rect 43920 44920 43936 44984
rect 44000 44920 44016 44984
rect 44080 44920 44096 44984
rect 44160 44920 44176 44984
rect 44240 44920 44256 44984
rect 44320 44920 44336 44984
rect 44400 44920 44416 44984
rect 44480 44920 44496 44984
rect 44560 44920 44576 44984
rect 44640 44920 44656 44984
rect 44720 44920 44736 44984
rect 44800 44920 44816 44984
rect 44880 44920 44896 44984
rect 44960 44920 44976 44984
rect 45040 44920 45056 44984
rect 45120 44920 45136 44984
rect 45200 44920 45216 44984
rect 45280 44920 45296 44984
rect 45360 44920 45368 44984
rect 0 44904 45368 44920
rect 0 44840 8 44904
rect 72 44840 88 44904
rect 152 44840 168 44904
rect 232 44840 248 44904
rect 312 44840 328 44904
rect 392 44840 408 44904
rect 472 44840 488 44904
rect 552 44840 568 44904
rect 632 44840 648 44904
rect 712 44840 728 44904
rect 792 44840 808 44904
rect 872 44840 888 44904
rect 952 44840 968 44904
rect 1032 44840 1048 44904
rect 1112 44840 1128 44904
rect 1192 44840 1208 44904
rect 1272 44840 1288 44904
rect 1352 44840 1368 44904
rect 1432 44840 1448 44904
rect 1512 44840 1528 44904
rect 1592 44840 1608 44904
rect 1672 44840 1688 44904
rect 1752 44840 1768 44904
rect 1832 44840 1848 44904
rect 1912 44840 1928 44904
rect 1992 44840 2008 44904
rect 2072 44840 2088 44904
rect 2152 44840 2168 44904
rect 2232 44840 2248 44904
rect 2312 44840 2328 44904
rect 2392 44840 2408 44904
rect 2472 44840 2488 44904
rect 2552 44840 2568 44904
rect 2632 44840 2648 44904
rect 2712 44840 2728 44904
rect 2792 44840 2808 44904
rect 2872 44840 2888 44904
rect 2952 44840 2968 44904
rect 3032 44840 3048 44904
rect 3112 44840 3128 44904
rect 3192 44840 3208 44904
rect 3272 44840 3288 44904
rect 3352 44840 3368 44904
rect 3432 44840 3448 44904
rect 3512 44840 3528 44904
rect 3592 44840 3608 44904
rect 3672 44840 3688 44904
rect 3752 44840 3768 44904
rect 3832 44840 3848 44904
rect 3912 44840 3928 44904
rect 3992 44840 19112 44904
rect 19176 44840 19192 44904
rect 19256 44840 19272 44904
rect 19336 44840 19352 44904
rect 19416 44840 29112 44904
rect 29176 44840 29192 44904
rect 29256 44840 29272 44904
rect 29336 44840 29352 44904
rect 29416 44840 41376 44904
rect 41440 44840 41456 44904
rect 41520 44840 41536 44904
rect 41600 44840 41616 44904
rect 41680 44840 41696 44904
rect 41760 44840 41776 44904
rect 41840 44840 41856 44904
rect 41920 44840 41936 44904
rect 42000 44840 42016 44904
rect 42080 44840 42096 44904
rect 42160 44840 42176 44904
rect 42240 44840 42256 44904
rect 42320 44840 42336 44904
rect 42400 44840 42416 44904
rect 42480 44840 42496 44904
rect 42560 44840 42576 44904
rect 42640 44840 42656 44904
rect 42720 44840 42736 44904
rect 42800 44840 42816 44904
rect 42880 44840 42896 44904
rect 42960 44840 42976 44904
rect 43040 44840 43056 44904
rect 43120 44840 43136 44904
rect 43200 44840 43216 44904
rect 43280 44840 43296 44904
rect 43360 44840 43376 44904
rect 43440 44840 43456 44904
rect 43520 44840 43536 44904
rect 43600 44840 43616 44904
rect 43680 44840 43696 44904
rect 43760 44840 43776 44904
rect 43840 44840 43856 44904
rect 43920 44840 43936 44904
rect 44000 44840 44016 44904
rect 44080 44840 44096 44904
rect 44160 44840 44176 44904
rect 44240 44840 44256 44904
rect 44320 44840 44336 44904
rect 44400 44840 44416 44904
rect 44480 44840 44496 44904
rect 44560 44840 44576 44904
rect 44640 44840 44656 44904
rect 44720 44840 44736 44904
rect 44800 44840 44816 44904
rect 44880 44840 44896 44904
rect 44960 44840 44976 44904
rect 45040 44840 45056 44904
rect 45120 44840 45136 44904
rect 45200 44840 45216 44904
rect 45280 44840 45296 44904
rect 45360 44840 45368 44904
rect 0 44824 45368 44840
rect 0 44760 8 44824
rect 72 44760 88 44824
rect 152 44760 168 44824
rect 232 44760 248 44824
rect 312 44760 328 44824
rect 392 44760 408 44824
rect 472 44760 488 44824
rect 552 44760 568 44824
rect 632 44760 648 44824
rect 712 44760 728 44824
rect 792 44760 808 44824
rect 872 44760 888 44824
rect 952 44760 968 44824
rect 1032 44760 1048 44824
rect 1112 44760 1128 44824
rect 1192 44760 1208 44824
rect 1272 44760 1288 44824
rect 1352 44760 1368 44824
rect 1432 44760 1448 44824
rect 1512 44760 1528 44824
rect 1592 44760 1608 44824
rect 1672 44760 1688 44824
rect 1752 44760 1768 44824
rect 1832 44760 1848 44824
rect 1912 44760 1928 44824
rect 1992 44760 2008 44824
rect 2072 44760 2088 44824
rect 2152 44760 2168 44824
rect 2232 44760 2248 44824
rect 2312 44760 2328 44824
rect 2392 44760 2408 44824
rect 2472 44760 2488 44824
rect 2552 44760 2568 44824
rect 2632 44760 2648 44824
rect 2712 44760 2728 44824
rect 2792 44760 2808 44824
rect 2872 44760 2888 44824
rect 2952 44760 2968 44824
rect 3032 44760 3048 44824
rect 3112 44760 3128 44824
rect 3192 44760 3208 44824
rect 3272 44760 3288 44824
rect 3352 44760 3368 44824
rect 3432 44760 3448 44824
rect 3512 44760 3528 44824
rect 3592 44760 3608 44824
rect 3672 44760 3688 44824
rect 3752 44760 3768 44824
rect 3832 44760 3848 44824
rect 3912 44760 3928 44824
rect 3992 44760 19112 44824
rect 19176 44760 19192 44824
rect 19256 44760 19272 44824
rect 19336 44760 19352 44824
rect 19416 44760 29112 44824
rect 29176 44760 29192 44824
rect 29256 44760 29272 44824
rect 29336 44760 29352 44824
rect 29416 44760 41376 44824
rect 41440 44760 41456 44824
rect 41520 44760 41536 44824
rect 41600 44760 41616 44824
rect 41680 44760 41696 44824
rect 41760 44760 41776 44824
rect 41840 44760 41856 44824
rect 41920 44760 41936 44824
rect 42000 44760 42016 44824
rect 42080 44760 42096 44824
rect 42160 44760 42176 44824
rect 42240 44760 42256 44824
rect 42320 44760 42336 44824
rect 42400 44760 42416 44824
rect 42480 44760 42496 44824
rect 42560 44760 42576 44824
rect 42640 44760 42656 44824
rect 42720 44760 42736 44824
rect 42800 44760 42816 44824
rect 42880 44760 42896 44824
rect 42960 44760 42976 44824
rect 43040 44760 43056 44824
rect 43120 44760 43136 44824
rect 43200 44760 43216 44824
rect 43280 44760 43296 44824
rect 43360 44760 43376 44824
rect 43440 44760 43456 44824
rect 43520 44760 43536 44824
rect 43600 44760 43616 44824
rect 43680 44760 43696 44824
rect 43760 44760 43776 44824
rect 43840 44760 43856 44824
rect 43920 44760 43936 44824
rect 44000 44760 44016 44824
rect 44080 44760 44096 44824
rect 44160 44760 44176 44824
rect 44240 44760 44256 44824
rect 44320 44760 44336 44824
rect 44400 44760 44416 44824
rect 44480 44760 44496 44824
rect 44560 44760 44576 44824
rect 44640 44760 44656 44824
rect 44720 44760 44736 44824
rect 44800 44760 44816 44824
rect 44880 44760 44896 44824
rect 44960 44760 44976 44824
rect 45040 44760 45056 44824
rect 45120 44760 45136 44824
rect 45200 44760 45216 44824
rect 45280 44760 45296 44824
rect 45360 44760 45368 44824
rect 0 44744 45368 44760
rect 0 44680 8 44744
rect 72 44680 88 44744
rect 152 44680 168 44744
rect 232 44680 248 44744
rect 312 44680 328 44744
rect 392 44680 408 44744
rect 472 44680 488 44744
rect 552 44680 568 44744
rect 632 44680 648 44744
rect 712 44680 728 44744
rect 792 44680 808 44744
rect 872 44680 888 44744
rect 952 44680 968 44744
rect 1032 44680 1048 44744
rect 1112 44680 1128 44744
rect 1192 44680 1208 44744
rect 1272 44680 1288 44744
rect 1352 44680 1368 44744
rect 1432 44680 1448 44744
rect 1512 44680 1528 44744
rect 1592 44680 1608 44744
rect 1672 44680 1688 44744
rect 1752 44680 1768 44744
rect 1832 44680 1848 44744
rect 1912 44680 1928 44744
rect 1992 44680 2008 44744
rect 2072 44680 2088 44744
rect 2152 44680 2168 44744
rect 2232 44680 2248 44744
rect 2312 44680 2328 44744
rect 2392 44680 2408 44744
rect 2472 44680 2488 44744
rect 2552 44680 2568 44744
rect 2632 44680 2648 44744
rect 2712 44680 2728 44744
rect 2792 44680 2808 44744
rect 2872 44680 2888 44744
rect 2952 44680 2968 44744
rect 3032 44680 3048 44744
rect 3112 44680 3128 44744
rect 3192 44680 3208 44744
rect 3272 44680 3288 44744
rect 3352 44680 3368 44744
rect 3432 44680 3448 44744
rect 3512 44680 3528 44744
rect 3592 44680 3608 44744
rect 3672 44680 3688 44744
rect 3752 44680 3768 44744
rect 3832 44680 3848 44744
rect 3912 44680 3928 44744
rect 3992 44680 19112 44744
rect 19176 44680 19192 44744
rect 19256 44680 19272 44744
rect 19336 44680 19352 44744
rect 19416 44680 29112 44744
rect 29176 44680 29192 44744
rect 29256 44680 29272 44744
rect 29336 44680 29352 44744
rect 29416 44680 41376 44744
rect 41440 44680 41456 44744
rect 41520 44680 41536 44744
rect 41600 44680 41616 44744
rect 41680 44680 41696 44744
rect 41760 44680 41776 44744
rect 41840 44680 41856 44744
rect 41920 44680 41936 44744
rect 42000 44680 42016 44744
rect 42080 44680 42096 44744
rect 42160 44680 42176 44744
rect 42240 44680 42256 44744
rect 42320 44680 42336 44744
rect 42400 44680 42416 44744
rect 42480 44680 42496 44744
rect 42560 44680 42576 44744
rect 42640 44680 42656 44744
rect 42720 44680 42736 44744
rect 42800 44680 42816 44744
rect 42880 44680 42896 44744
rect 42960 44680 42976 44744
rect 43040 44680 43056 44744
rect 43120 44680 43136 44744
rect 43200 44680 43216 44744
rect 43280 44680 43296 44744
rect 43360 44680 43376 44744
rect 43440 44680 43456 44744
rect 43520 44680 43536 44744
rect 43600 44680 43616 44744
rect 43680 44680 43696 44744
rect 43760 44680 43776 44744
rect 43840 44680 43856 44744
rect 43920 44680 43936 44744
rect 44000 44680 44016 44744
rect 44080 44680 44096 44744
rect 44160 44680 44176 44744
rect 44240 44680 44256 44744
rect 44320 44680 44336 44744
rect 44400 44680 44416 44744
rect 44480 44680 44496 44744
rect 44560 44680 44576 44744
rect 44640 44680 44656 44744
rect 44720 44680 44736 44744
rect 44800 44680 44816 44744
rect 44880 44680 44896 44744
rect 44960 44680 44976 44744
rect 45040 44680 45056 44744
rect 45120 44680 45136 44744
rect 45200 44680 45216 44744
rect 45280 44680 45296 44744
rect 45360 44680 45368 44744
rect 0 44664 45368 44680
rect 0 44600 8 44664
rect 72 44600 88 44664
rect 152 44600 168 44664
rect 232 44600 248 44664
rect 312 44600 328 44664
rect 392 44600 408 44664
rect 472 44600 488 44664
rect 552 44600 568 44664
rect 632 44600 648 44664
rect 712 44600 728 44664
rect 792 44600 808 44664
rect 872 44600 888 44664
rect 952 44600 968 44664
rect 1032 44600 1048 44664
rect 1112 44600 1128 44664
rect 1192 44600 1208 44664
rect 1272 44600 1288 44664
rect 1352 44600 1368 44664
rect 1432 44600 1448 44664
rect 1512 44600 1528 44664
rect 1592 44600 1608 44664
rect 1672 44600 1688 44664
rect 1752 44600 1768 44664
rect 1832 44600 1848 44664
rect 1912 44600 1928 44664
rect 1992 44600 2008 44664
rect 2072 44600 2088 44664
rect 2152 44600 2168 44664
rect 2232 44600 2248 44664
rect 2312 44600 2328 44664
rect 2392 44600 2408 44664
rect 2472 44600 2488 44664
rect 2552 44600 2568 44664
rect 2632 44600 2648 44664
rect 2712 44600 2728 44664
rect 2792 44600 2808 44664
rect 2872 44600 2888 44664
rect 2952 44600 2968 44664
rect 3032 44600 3048 44664
rect 3112 44600 3128 44664
rect 3192 44600 3208 44664
rect 3272 44600 3288 44664
rect 3352 44600 3368 44664
rect 3432 44600 3448 44664
rect 3512 44600 3528 44664
rect 3592 44600 3608 44664
rect 3672 44600 3688 44664
rect 3752 44600 3768 44664
rect 3832 44600 3848 44664
rect 3912 44600 3928 44664
rect 3992 44600 19112 44664
rect 19176 44600 19192 44664
rect 19256 44600 19272 44664
rect 19336 44600 19352 44664
rect 19416 44600 29112 44664
rect 29176 44600 29192 44664
rect 29256 44600 29272 44664
rect 29336 44600 29352 44664
rect 29416 44600 41376 44664
rect 41440 44600 41456 44664
rect 41520 44600 41536 44664
rect 41600 44600 41616 44664
rect 41680 44600 41696 44664
rect 41760 44600 41776 44664
rect 41840 44600 41856 44664
rect 41920 44600 41936 44664
rect 42000 44600 42016 44664
rect 42080 44600 42096 44664
rect 42160 44600 42176 44664
rect 42240 44600 42256 44664
rect 42320 44600 42336 44664
rect 42400 44600 42416 44664
rect 42480 44600 42496 44664
rect 42560 44600 42576 44664
rect 42640 44600 42656 44664
rect 42720 44600 42736 44664
rect 42800 44600 42816 44664
rect 42880 44600 42896 44664
rect 42960 44600 42976 44664
rect 43040 44600 43056 44664
rect 43120 44600 43136 44664
rect 43200 44600 43216 44664
rect 43280 44600 43296 44664
rect 43360 44600 43376 44664
rect 43440 44600 43456 44664
rect 43520 44600 43536 44664
rect 43600 44600 43616 44664
rect 43680 44600 43696 44664
rect 43760 44600 43776 44664
rect 43840 44600 43856 44664
rect 43920 44600 43936 44664
rect 44000 44600 44016 44664
rect 44080 44600 44096 44664
rect 44160 44600 44176 44664
rect 44240 44600 44256 44664
rect 44320 44600 44336 44664
rect 44400 44600 44416 44664
rect 44480 44600 44496 44664
rect 44560 44600 44576 44664
rect 44640 44600 44656 44664
rect 44720 44600 44736 44664
rect 44800 44600 44816 44664
rect 44880 44600 44896 44664
rect 44960 44600 44976 44664
rect 45040 44600 45056 44664
rect 45120 44600 45136 44664
rect 45200 44600 45216 44664
rect 45280 44600 45296 44664
rect 45360 44600 45368 44664
rect 0 44584 45368 44600
rect 0 44520 8 44584
rect 72 44520 88 44584
rect 152 44520 168 44584
rect 232 44520 248 44584
rect 312 44520 328 44584
rect 392 44520 408 44584
rect 472 44520 488 44584
rect 552 44520 568 44584
rect 632 44520 648 44584
rect 712 44520 728 44584
rect 792 44520 808 44584
rect 872 44520 888 44584
rect 952 44520 968 44584
rect 1032 44520 1048 44584
rect 1112 44520 1128 44584
rect 1192 44520 1208 44584
rect 1272 44520 1288 44584
rect 1352 44520 1368 44584
rect 1432 44520 1448 44584
rect 1512 44520 1528 44584
rect 1592 44520 1608 44584
rect 1672 44520 1688 44584
rect 1752 44520 1768 44584
rect 1832 44520 1848 44584
rect 1912 44520 1928 44584
rect 1992 44520 2008 44584
rect 2072 44520 2088 44584
rect 2152 44520 2168 44584
rect 2232 44520 2248 44584
rect 2312 44520 2328 44584
rect 2392 44520 2408 44584
rect 2472 44520 2488 44584
rect 2552 44520 2568 44584
rect 2632 44520 2648 44584
rect 2712 44520 2728 44584
rect 2792 44520 2808 44584
rect 2872 44520 2888 44584
rect 2952 44520 2968 44584
rect 3032 44520 3048 44584
rect 3112 44520 3128 44584
rect 3192 44520 3208 44584
rect 3272 44520 3288 44584
rect 3352 44520 3368 44584
rect 3432 44520 3448 44584
rect 3512 44520 3528 44584
rect 3592 44520 3608 44584
rect 3672 44520 3688 44584
rect 3752 44520 3768 44584
rect 3832 44520 3848 44584
rect 3912 44520 3928 44584
rect 3992 44520 19112 44584
rect 19176 44520 19192 44584
rect 19256 44520 19272 44584
rect 19336 44520 19352 44584
rect 19416 44520 29112 44584
rect 29176 44520 29192 44584
rect 29256 44520 29272 44584
rect 29336 44520 29352 44584
rect 29416 44520 41376 44584
rect 41440 44520 41456 44584
rect 41520 44520 41536 44584
rect 41600 44520 41616 44584
rect 41680 44520 41696 44584
rect 41760 44520 41776 44584
rect 41840 44520 41856 44584
rect 41920 44520 41936 44584
rect 42000 44520 42016 44584
rect 42080 44520 42096 44584
rect 42160 44520 42176 44584
rect 42240 44520 42256 44584
rect 42320 44520 42336 44584
rect 42400 44520 42416 44584
rect 42480 44520 42496 44584
rect 42560 44520 42576 44584
rect 42640 44520 42656 44584
rect 42720 44520 42736 44584
rect 42800 44520 42816 44584
rect 42880 44520 42896 44584
rect 42960 44520 42976 44584
rect 43040 44520 43056 44584
rect 43120 44520 43136 44584
rect 43200 44520 43216 44584
rect 43280 44520 43296 44584
rect 43360 44520 43376 44584
rect 43440 44520 43456 44584
rect 43520 44520 43536 44584
rect 43600 44520 43616 44584
rect 43680 44520 43696 44584
rect 43760 44520 43776 44584
rect 43840 44520 43856 44584
rect 43920 44520 43936 44584
rect 44000 44520 44016 44584
rect 44080 44520 44096 44584
rect 44160 44520 44176 44584
rect 44240 44520 44256 44584
rect 44320 44520 44336 44584
rect 44400 44520 44416 44584
rect 44480 44520 44496 44584
rect 44560 44520 44576 44584
rect 44640 44520 44656 44584
rect 44720 44520 44736 44584
rect 44800 44520 44816 44584
rect 44880 44520 44896 44584
rect 44960 44520 44976 44584
rect 45040 44520 45056 44584
rect 45120 44520 45136 44584
rect 45200 44520 45216 44584
rect 45280 44520 45296 44584
rect 45360 44520 45368 44584
rect 0 44504 45368 44520
rect 0 44440 8 44504
rect 72 44440 88 44504
rect 152 44440 168 44504
rect 232 44440 248 44504
rect 312 44440 328 44504
rect 392 44440 408 44504
rect 472 44440 488 44504
rect 552 44440 568 44504
rect 632 44440 648 44504
rect 712 44440 728 44504
rect 792 44440 808 44504
rect 872 44440 888 44504
rect 952 44440 968 44504
rect 1032 44440 1048 44504
rect 1112 44440 1128 44504
rect 1192 44440 1208 44504
rect 1272 44440 1288 44504
rect 1352 44440 1368 44504
rect 1432 44440 1448 44504
rect 1512 44440 1528 44504
rect 1592 44440 1608 44504
rect 1672 44440 1688 44504
rect 1752 44440 1768 44504
rect 1832 44440 1848 44504
rect 1912 44440 1928 44504
rect 1992 44440 2008 44504
rect 2072 44440 2088 44504
rect 2152 44440 2168 44504
rect 2232 44440 2248 44504
rect 2312 44440 2328 44504
rect 2392 44440 2408 44504
rect 2472 44440 2488 44504
rect 2552 44440 2568 44504
rect 2632 44440 2648 44504
rect 2712 44440 2728 44504
rect 2792 44440 2808 44504
rect 2872 44440 2888 44504
rect 2952 44440 2968 44504
rect 3032 44440 3048 44504
rect 3112 44440 3128 44504
rect 3192 44440 3208 44504
rect 3272 44440 3288 44504
rect 3352 44440 3368 44504
rect 3432 44440 3448 44504
rect 3512 44440 3528 44504
rect 3592 44440 3608 44504
rect 3672 44440 3688 44504
rect 3752 44440 3768 44504
rect 3832 44440 3848 44504
rect 3912 44440 3928 44504
rect 3992 44440 19112 44504
rect 19176 44440 19192 44504
rect 19256 44440 19272 44504
rect 19336 44440 19352 44504
rect 19416 44440 29112 44504
rect 29176 44440 29192 44504
rect 29256 44440 29272 44504
rect 29336 44440 29352 44504
rect 29416 44440 41376 44504
rect 41440 44440 41456 44504
rect 41520 44440 41536 44504
rect 41600 44440 41616 44504
rect 41680 44440 41696 44504
rect 41760 44440 41776 44504
rect 41840 44440 41856 44504
rect 41920 44440 41936 44504
rect 42000 44440 42016 44504
rect 42080 44440 42096 44504
rect 42160 44440 42176 44504
rect 42240 44440 42256 44504
rect 42320 44440 42336 44504
rect 42400 44440 42416 44504
rect 42480 44440 42496 44504
rect 42560 44440 42576 44504
rect 42640 44440 42656 44504
rect 42720 44440 42736 44504
rect 42800 44440 42816 44504
rect 42880 44440 42896 44504
rect 42960 44440 42976 44504
rect 43040 44440 43056 44504
rect 43120 44440 43136 44504
rect 43200 44440 43216 44504
rect 43280 44440 43296 44504
rect 43360 44440 43376 44504
rect 43440 44440 43456 44504
rect 43520 44440 43536 44504
rect 43600 44440 43616 44504
rect 43680 44440 43696 44504
rect 43760 44440 43776 44504
rect 43840 44440 43856 44504
rect 43920 44440 43936 44504
rect 44000 44440 44016 44504
rect 44080 44440 44096 44504
rect 44160 44440 44176 44504
rect 44240 44440 44256 44504
rect 44320 44440 44336 44504
rect 44400 44440 44416 44504
rect 44480 44440 44496 44504
rect 44560 44440 44576 44504
rect 44640 44440 44656 44504
rect 44720 44440 44736 44504
rect 44800 44440 44816 44504
rect 44880 44440 44896 44504
rect 44960 44440 44976 44504
rect 45040 44440 45056 44504
rect 45120 44440 45136 44504
rect 45200 44440 45216 44504
rect 45280 44440 45296 44504
rect 45360 44440 45368 44504
rect 0 44424 45368 44440
rect 0 44360 8 44424
rect 72 44360 88 44424
rect 152 44360 168 44424
rect 232 44360 248 44424
rect 312 44360 328 44424
rect 392 44360 408 44424
rect 472 44360 488 44424
rect 552 44360 568 44424
rect 632 44360 648 44424
rect 712 44360 728 44424
rect 792 44360 808 44424
rect 872 44360 888 44424
rect 952 44360 968 44424
rect 1032 44360 1048 44424
rect 1112 44360 1128 44424
rect 1192 44360 1208 44424
rect 1272 44360 1288 44424
rect 1352 44360 1368 44424
rect 1432 44360 1448 44424
rect 1512 44360 1528 44424
rect 1592 44360 1608 44424
rect 1672 44360 1688 44424
rect 1752 44360 1768 44424
rect 1832 44360 1848 44424
rect 1912 44360 1928 44424
rect 1992 44360 2008 44424
rect 2072 44360 2088 44424
rect 2152 44360 2168 44424
rect 2232 44360 2248 44424
rect 2312 44360 2328 44424
rect 2392 44360 2408 44424
rect 2472 44360 2488 44424
rect 2552 44360 2568 44424
rect 2632 44360 2648 44424
rect 2712 44360 2728 44424
rect 2792 44360 2808 44424
rect 2872 44360 2888 44424
rect 2952 44360 2968 44424
rect 3032 44360 3048 44424
rect 3112 44360 3128 44424
rect 3192 44360 3208 44424
rect 3272 44360 3288 44424
rect 3352 44360 3368 44424
rect 3432 44360 3448 44424
rect 3512 44360 3528 44424
rect 3592 44360 3608 44424
rect 3672 44360 3688 44424
rect 3752 44360 3768 44424
rect 3832 44360 3848 44424
rect 3912 44360 3928 44424
rect 3992 44360 19112 44424
rect 19176 44360 19192 44424
rect 19256 44360 19272 44424
rect 19336 44360 19352 44424
rect 19416 44360 29112 44424
rect 29176 44360 29192 44424
rect 29256 44360 29272 44424
rect 29336 44360 29352 44424
rect 29416 44360 41376 44424
rect 41440 44360 41456 44424
rect 41520 44360 41536 44424
rect 41600 44360 41616 44424
rect 41680 44360 41696 44424
rect 41760 44360 41776 44424
rect 41840 44360 41856 44424
rect 41920 44360 41936 44424
rect 42000 44360 42016 44424
rect 42080 44360 42096 44424
rect 42160 44360 42176 44424
rect 42240 44360 42256 44424
rect 42320 44360 42336 44424
rect 42400 44360 42416 44424
rect 42480 44360 42496 44424
rect 42560 44360 42576 44424
rect 42640 44360 42656 44424
rect 42720 44360 42736 44424
rect 42800 44360 42816 44424
rect 42880 44360 42896 44424
rect 42960 44360 42976 44424
rect 43040 44360 43056 44424
rect 43120 44360 43136 44424
rect 43200 44360 43216 44424
rect 43280 44360 43296 44424
rect 43360 44360 43376 44424
rect 43440 44360 43456 44424
rect 43520 44360 43536 44424
rect 43600 44360 43616 44424
rect 43680 44360 43696 44424
rect 43760 44360 43776 44424
rect 43840 44360 43856 44424
rect 43920 44360 43936 44424
rect 44000 44360 44016 44424
rect 44080 44360 44096 44424
rect 44160 44360 44176 44424
rect 44240 44360 44256 44424
rect 44320 44360 44336 44424
rect 44400 44360 44416 44424
rect 44480 44360 44496 44424
rect 44560 44360 44576 44424
rect 44640 44360 44656 44424
rect 44720 44360 44736 44424
rect 44800 44360 44816 44424
rect 44880 44360 44896 44424
rect 44960 44360 44976 44424
rect 45040 44360 45056 44424
rect 45120 44360 45136 44424
rect 45200 44360 45216 44424
rect 45280 44360 45296 44424
rect 45360 44360 45368 44424
rect 0 44344 45368 44360
rect 0 44280 8 44344
rect 72 44280 88 44344
rect 152 44280 168 44344
rect 232 44280 248 44344
rect 312 44280 328 44344
rect 392 44280 408 44344
rect 472 44280 488 44344
rect 552 44280 568 44344
rect 632 44280 648 44344
rect 712 44280 728 44344
rect 792 44280 808 44344
rect 872 44280 888 44344
rect 952 44280 968 44344
rect 1032 44280 1048 44344
rect 1112 44280 1128 44344
rect 1192 44280 1208 44344
rect 1272 44280 1288 44344
rect 1352 44280 1368 44344
rect 1432 44280 1448 44344
rect 1512 44280 1528 44344
rect 1592 44280 1608 44344
rect 1672 44280 1688 44344
rect 1752 44280 1768 44344
rect 1832 44280 1848 44344
rect 1912 44280 1928 44344
rect 1992 44280 2008 44344
rect 2072 44280 2088 44344
rect 2152 44280 2168 44344
rect 2232 44280 2248 44344
rect 2312 44280 2328 44344
rect 2392 44280 2408 44344
rect 2472 44280 2488 44344
rect 2552 44280 2568 44344
rect 2632 44280 2648 44344
rect 2712 44280 2728 44344
rect 2792 44280 2808 44344
rect 2872 44280 2888 44344
rect 2952 44280 2968 44344
rect 3032 44280 3048 44344
rect 3112 44280 3128 44344
rect 3192 44280 3208 44344
rect 3272 44280 3288 44344
rect 3352 44280 3368 44344
rect 3432 44280 3448 44344
rect 3512 44280 3528 44344
rect 3592 44280 3608 44344
rect 3672 44280 3688 44344
rect 3752 44280 3768 44344
rect 3832 44280 3848 44344
rect 3912 44280 3928 44344
rect 3992 44280 19112 44344
rect 19176 44280 19192 44344
rect 19256 44280 19272 44344
rect 19336 44280 19352 44344
rect 19416 44280 29112 44344
rect 29176 44280 29192 44344
rect 29256 44280 29272 44344
rect 29336 44280 29352 44344
rect 29416 44280 41376 44344
rect 41440 44280 41456 44344
rect 41520 44280 41536 44344
rect 41600 44280 41616 44344
rect 41680 44280 41696 44344
rect 41760 44280 41776 44344
rect 41840 44280 41856 44344
rect 41920 44280 41936 44344
rect 42000 44280 42016 44344
rect 42080 44280 42096 44344
rect 42160 44280 42176 44344
rect 42240 44280 42256 44344
rect 42320 44280 42336 44344
rect 42400 44280 42416 44344
rect 42480 44280 42496 44344
rect 42560 44280 42576 44344
rect 42640 44280 42656 44344
rect 42720 44280 42736 44344
rect 42800 44280 42816 44344
rect 42880 44280 42896 44344
rect 42960 44280 42976 44344
rect 43040 44280 43056 44344
rect 43120 44280 43136 44344
rect 43200 44280 43216 44344
rect 43280 44280 43296 44344
rect 43360 44280 43376 44344
rect 43440 44280 43456 44344
rect 43520 44280 43536 44344
rect 43600 44280 43616 44344
rect 43680 44280 43696 44344
rect 43760 44280 43776 44344
rect 43840 44280 43856 44344
rect 43920 44280 43936 44344
rect 44000 44280 44016 44344
rect 44080 44280 44096 44344
rect 44160 44280 44176 44344
rect 44240 44280 44256 44344
rect 44320 44280 44336 44344
rect 44400 44280 44416 44344
rect 44480 44280 44496 44344
rect 44560 44280 44576 44344
rect 44640 44280 44656 44344
rect 44720 44280 44736 44344
rect 44800 44280 44816 44344
rect 44880 44280 44896 44344
rect 44960 44280 44976 44344
rect 45040 44280 45056 44344
rect 45120 44280 45136 44344
rect 45200 44280 45216 44344
rect 45280 44280 45296 44344
rect 45360 44280 45368 44344
rect 0 44264 45368 44280
rect 0 44200 8 44264
rect 72 44200 88 44264
rect 152 44200 168 44264
rect 232 44200 248 44264
rect 312 44200 328 44264
rect 392 44200 408 44264
rect 472 44200 488 44264
rect 552 44200 568 44264
rect 632 44200 648 44264
rect 712 44200 728 44264
rect 792 44200 808 44264
rect 872 44200 888 44264
rect 952 44200 968 44264
rect 1032 44200 1048 44264
rect 1112 44200 1128 44264
rect 1192 44200 1208 44264
rect 1272 44200 1288 44264
rect 1352 44200 1368 44264
rect 1432 44200 1448 44264
rect 1512 44200 1528 44264
rect 1592 44200 1608 44264
rect 1672 44200 1688 44264
rect 1752 44200 1768 44264
rect 1832 44200 1848 44264
rect 1912 44200 1928 44264
rect 1992 44200 2008 44264
rect 2072 44200 2088 44264
rect 2152 44200 2168 44264
rect 2232 44200 2248 44264
rect 2312 44200 2328 44264
rect 2392 44200 2408 44264
rect 2472 44200 2488 44264
rect 2552 44200 2568 44264
rect 2632 44200 2648 44264
rect 2712 44200 2728 44264
rect 2792 44200 2808 44264
rect 2872 44200 2888 44264
rect 2952 44200 2968 44264
rect 3032 44200 3048 44264
rect 3112 44200 3128 44264
rect 3192 44200 3208 44264
rect 3272 44200 3288 44264
rect 3352 44200 3368 44264
rect 3432 44200 3448 44264
rect 3512 44200 3528 44264
rect 3592 44200 3608 44264
rect 3672 44200 3688 44264
rect 3752 44200 3768 44264
rect 3832 44200 3848 44264
rect 3912 44200 3928 44264
rect 3992 44200 19112 44264
rect 19176 44200 19192 44264
rect 19256 44200 19272 44264
rect 19336 44200 19352 44264
rect 19416 44200 29112 44264
rect 29176 44200 29192 44264
rect 29256 44200 29272 44264
rect 29336 44200 29352 44264
rect 29416 44200 41376 44264
rect 41440 44200 41456 44264
rect 41520 44200 41536 44264
rect 41600 44200 41616 44264
rect 41680 44200 41696 44264
rect 41760 44200 41776 44264
rect 41840 44200 41856 44264
rect 41920 44200 41936 44264
rect 42000 44200 42016 44264
rect 42080 44200 42096 44264
rect 42160 44200 42176 44264
rect 42240 44200 42256 44264
rect 42320 44200 42336 44264
rect 42400 44200 42416 44264
rect 42480 44200 42496 44264
rect 42560 44200 42576 44264
rect 42640 44200 42656 44264
rect 42720 44200 42736 44264
rect 42800 44200 42816 44264
rect 42880 44200 42896 44264
rect 42960 44200 42976 44264
rect 43040 44200 43056 44264
rect 43120 44200 43136 44264
rect 43200 44200 43216 44264
rect 43280 44200 43296 44264
rect 43360 44200 43376 44264
rect 43440 44200 43456 44264
rect 43520 44200 43536 44264
rect 43600 44200 43616 44264
rect 43680 44200 43696 44264
rect 43760 44200 43776 44264
rect 43840 44200 43856 44264
rect 43920 44200 43936 44264
rect 44000 44200 44016 44264
rect 44080 44200 44096 44264
rect 44160 44200 44176 44264
rect 44240 44200 44256 44264
rect 44320 44200 44336 44264
rect 44400 44200 44416 44264
rect 44480 44200 44496 44264
rect 44560 44200 44576 44264
rect 44640 44200 44656 44264
rect 44720 44200 44736 44264
rect 44800 44200 44816 44264
rect 44880 44200 44896 44264
rect 44960 44200 44976 44264
rect 45040 44200 45056 44264
rect 45120 44200 45136 44264
rect 45200 44200 45216 44264
rect 45280 44200 45296 44264
rect 45360 44200 45368 44264
rect 0 44184 45368 44200
rect 0 44120 8 44184
rect 72 44120 88 44184
rect 152 44120 168 44184
rect 232 44120 248 44184
rect 312 44120 328 44184
rect 392 44120 408 44184
rect 472 44120 488 44184
rect 552 44120 568 44184
rect 632 44120 648 44184
rect 712 44120 728 44184
rect 792 44120 808 44184
rect 872 44120 888 44184
rect 952 44120 968 44184
rect 1032 44120 1048 44184
rect 1112 44120 1128 44184
rect 1192 44120 1208 44184
rect 1272 44120 1288 44184
rect 1352 44120 1368 44184
rect 1432 44120 1448 44184
rect 1512 44120 1528 44184
rect 1592 44120 1608 44184
rect 1672 44120 1688 44184
rect 1752 44120 1768 44184
rect 1832 44120 1848 44184
rect 1912 44120 1928 44184
rect 1992 44120 2008 44184
rect 2072 44120 2088 44184
rect 2152 44120 2168 44184
rect 2232 44120 2248 44184
rect 2312 44120 2328 44184
rect 2392 44120 2408 44184
rect 2472 44120 2488 44184
rect 2552 44120 2568 44184
rect 2632 44120 2648 44184
rect 2712 44120 2728 44184
rect 2792 44120 2808 44184
rect 2872 44120 2888 44184
rect 2952 44120 2968 44184
rect 3032 44120 3048 44184
rect 3112 44120 3128 44184
rect 3192 44120 3208 44184
rect 3272 44120 3288 44184
rect 3352 44120 3368 44184
rect 3432 44120 3448 44184
rect 3512 44120 3528 44184
rect 3592 44120 3608 44184
rect 3672 44120 3688 44184
rect 3752 44120 3768 44184
rect 3832 44120 3848 44184
rect 3912 44120 3928 44184
rect 3992 44120 19112 44184
rect 19176 44120 19192 44184
rect 19256 44120 19272 44184
rect 19336 44120 19352 44184
rect 19416 44120 29112 44184
rect 29176 44120 29192 44184
rect 29256 44120 29272 44184
rect 29336 44120 29352 44184
rect 29416 44120 41376 44184
rect 41440 44120 41456 44184
rect 41520 44120 41536 44184
rect 41600 44120 41616 44184
rect 41680 44120 41696 44184
rect 41760 44120 41776 44184
rect 41840 44120 41856 44184
rect 41920 44120 41936 44184
rect 42000 44120 42016 44184
rect 42080 44120 42096 44184
rect 42160 44120 42176 44184
rect 42240 44120 42256 44184
rect 42320 44120 42336 44184
rect 42400 44120 42416 44184
rect 42480 44120 42496 44184
rect 42560 44120 42576 44184
rect 42640 44120 42656 44184
rect 42720 44120 42736 44184
rect 42800 44120 42816 44184
rect 42880 44120 42896 44184
rect 42960 44120 42976 44184
rect 43040 44120 43056 44184
rect 43120 44120 43136 44184
rect 43200 44120 43216 44184
rect 43280 44120 43296 44184
rect 43360 44120 43376 44184
rect 43440 44120 43456 44184
rect 43520 44120 43536 44184
rect 43600 44120 43616 44184
rect 43680 44120 43696 44184
rect 43760 44120 43776 44184
rect 43840 44120 43856 44184
rect 43920 44120 43936 44184
rect 44000 44120 44016 44184
rect 44080 44120 44096 44184
rect 44160 44120 44176 44184
rect 44240 44120 44256 44184
rect 44320 44120 44336 44184
rect 44400 44120 44416 44184
rect 44480 44120 44496 44184
rect 44560 44120 44576 44184
rect 44640 44120 44656 44184
rect 44720 44120 44736 44184
rect 44800 44120 44816 44184
rect 44880 44120 44896 44184
rect 44960 44120 44976 44184
rect 45040 44120 45056 44184
rect 45120 44120 45136 44184
rect 45200 44120 45216 44184
rect 45280 44120 45296 44184
rect 45360 44120 45368 44184
rect 0 44104 45368 44120
rect 0 44040 8 44104
rect 72 44040 88 44104
rect 152 44040 168 44104
rect 232 44040 248 44104
rect 312 44040 328 44104
rect 392 44040 408 44104
rect 472 44040 488 44104
rect 552 44040 568 44104
rect 632 44040 648 44104
rect 712 44040 728 44104
rect 792 44040 808 44104
rect 872 44040 888 44104
rect 952 44040 968 44104
rect 1032 44040 1048 44104
rect 1112 44040 1128 44104
rect 1192 44040 1208 44104
rect 1272 44040 1288 44104
rect 1352 44040 1368 44104
rect 1432 44040 1448 44104
rect 1512 44040 1528 44104
rect 1592 44040 1608 44104
rect 1672 44040 1688 44104
rect 1752 44040 1768 44104
rect 1832 44040 1848 44104
rect 1912 44040 1928 44104
rect 1992 44040 2008 44104
rect 2072 44040 2088 44104
rect 2152 44040 2168 44104
rect 2232 44040 2248 44104
rect 2312 44040 2328 44104
rect 2392 44040 2408 44104
rect 2472 44040 2488 44104
rect 2552 44040 2568 44104
rect 2632 44040 2648 44104
rect 2712 44040 2728 44104
rect 2792 44040 2808 44104
rect 2872 44040 2888 44104
rect 2952 44040 2968 44104
rect 3032 44040 3048 44104
rect 3112 44040 3128 44104
rect 3192 44040 3208 44104
rect 3272 44040 3288 44104
rect 3352 44040 3368 44104
rect 3432 44040 3448 44104
rect 3512 44040 3528 44104
rect 3592 44040 3608 44104
rect 3672 44040 3688 44104
rect 3752 44040 3768 44104
rect 3832 44040 3848 44104
rect 3912 44040 3928 44104
rect 3992 44040 19112 44104
rect 19176 44040 19192 44104
rect 19256 44040 19272 44104
rect 19336 44040 19352 44104
rect 19416 44040 29112 44104
rect 29176 44040 29192 44104
rect 29256 44040 29272 44104
rect 29336 44040 29352 44104
rect 29416 44040 41376 44104
rect 41440 44040 41456 44104
rect 41520 44040 41536 44104
rect 41600 44040 41616 44104
rect 41680 44040 41696 44104
rect 41760 44040 41776 44104
rect 41840 44040 41856 44104
rect 41920 44040 41936 44104
rect 42000 44040 42016 44104
rect 42080 44040 42096 44104
rect 42160 44040 42176 44104
rect 42240 44040 42256 44104
rect 42320 44040 42336 44104
rect 42400 44040 42416 44104
rect 42480 44040 42496 44104
rect 42560 44040 42576 44104
rect 42640 44040 42656 44104
rect 42720 44040 42736 44104
rect 42800 44040 42816 44104
rect 42880 44040 42896 44104
rect 42960 44040 42976 44104
rect 43040 44040 43056 44104
rect 43120 44040 43136 44104
rect 43200 44040 43216 44104
rect 43280 44040 43296 44104
rect 43360 44040 43376 44104
rect 43440 44040 43456 44104
rect 43520 44040 43536 44104
rect 43600 44040 43616 44104
rect 43680 44040 43696 44104
rect 43760 44040 43776 44104
rect 43840 44040 43856 44104
rect 43920 44040 43936 44104
rect 44000 44040 44016 44104
rect 44080 44040 44096 44104
rect 44160 44040 44176 44104
rect 44240 44040 44256 44104
rect 44320 44040 44336 44104
rect 44400 44040 44416 44104
rect 44480 44040 44496 44104
rect 44560 44040 44576 44104
rect 44640 44040 44656 44104
rect 44720 44040 44736 44104
rect 44800 44040 44816 44104
rect 44880 44040 44896 44104
rect 44960 44040 44976 44104
rect 45040 44040 45056 44104
rect 45120 44040 45136 44104
rect 45200 44040 45216 44104
rect 45280 44040 45296 44104
rect 45360 44040 45368 44104
rect 0 44024 45368 44040
rect 0 43960 8 44024
rect 72 43960 88 44024
rect 152 43960 168 44024
rect 232 43960 248 44024
rect 312 43960 328 44024
rect 392 43960 408 44024
rect 472 43960 488 44024
rect 552 43960 568 44024
rect 632 43960 648 44024
rect 712 43960 728 44024
rect 792 43960 808 44024
rect 872 43960 888 44024
rect 952 43960 968 44024
rect 1032 43960 1048 44024
rect 1112 43960 1128 44024
rect 1192 43960 1208 44024
rect 1272 43960 1288 44024
rect 1352 43960 1368 44024
rect 1432 43960 1448 44024
rect 1512 43960 1528 44024
rect 1592 43960 1608 44024
rect 1672 43960 1688 44024
rect 1752 43960 1768 44024
rect 1832 43960 1848 44024
rect 1912 43960 1928 44024
rect 1992 43960 2008 44024
rect 2072 43960 2088 44024
rect 2152 43960 2168 44024
rect 2232 43960 2248 44024
rect 2312 43960 2328 44024
rect 2392 43960 2408 44024
rect 2472 43960 2488 44024
rect 2552 43960 2568 44024
rect 2632 43960 2648 44024
rect 2712 43960 2728 44024
rect 2792 43960 2808 44024
rect 2872 43960 2888 44024
rect 2952 43960 2968 44024
rect 3032 43960 3048 44024
rect 3112 43960 3128 44024
rect 3192 43960 3208 44024
rect 3272 43960 3288 44024
rect 3352 43960 3368 44024
rect 3432 43960 3448 44024
rect 3512 43960 3528 44024
rect 3592 43960 3608 44024
rect 3672 43960 3688 44024
rect 3752 43960 3768 44024
rect 3832 43960 3848 44024
rect 3912 43960 3928 44024
rect 3992 43960 19112 44024
rect 19176 43960 19192 44024
rect 19256 43960 19272 44024
rect 19336 43960 19352 44024
rect 19416 43960 29112 44024
rect 29176 43960 29192 44024
rect 29256 43960 29272 44024
rect 29336 43960 29352 44024
rect 29416 43960 41376 44024
rect 41440 43960 41456 44024
rect 41520 43960 41536 44024
rect 41600 43960 41616 44024
rect 41680 43960 41696 44024
rect 41760 43960 41776 44024
rect 41840 43960 41856 44024
rect 41920 43960 41936 44024
rect 42000 43960 42016 44024
rect 42080 43960 42096 44024
rect 42160 43960 42176 44024
rect 42240 43960 42256 44024
rect 42320 43960 42336 44024
rect 42400 43960 42416 44024
rect 42480 43960 42496 44024
rect 42560 43960 42576 44024
rect 42640 43960 42656 44024
rect 42720 43960 42736 44024
rect 42800 43960 42816 44024
rect 42880 43960 42896 44024
rect 42960 43960 42976 44024
rect 43040 43960 43056 44024
rect 43120 43960 43136 44024
rect 43200 43960 43216 44024
rect 43280 43960 43296 44024
rect 43360 43960 43376 44024
rect 43440 43960 43456 44024
rect 43520 43960 43536 44024
rect 43600 43960 43616 44024
rect 43680 43960 43696 44024
rect 43760 43960 43776 44024
rect 43840 43960 43856 44024
rect 43920 43960 43936 44024
rect 44000 43960 44016 44024
rect 44080 43960 44096 44024
rect 44160 43960 44176 44024
rect 44240 43960 44256 44024
rect 44320 43960 44336 44024
rect 44400 43960 44416 44024
rect 44480 43960 44496 44024
rect 44560 43960 44576 44024
rect 44640 43960 44656 44024
rect 44720 43960 44736 44024
rect 44800 43960 44816 44024
rect 44880 43960 44896 44024
rect 44960 43960 44976 44024
rect 45040 43960 45056 44024
rect 45120 43960 45136 44024
rect 45200 43960 45216 44024
rect 45280 43960 45296 44024
rect 45360 43960 45368 44024
rect 0 43944 45368 43960
rect 0 43880 8 43944
rect 72 43880 88 43944
rect 152 43880 168 43944
rect 232 43880 248 43944
rect 312 43880 328 43944
rect 392 43880 408 43944
rect 472 43880 488 43944
rect 552 43880 568 43944
rect 632 43880 648 43944
rect 712 43880 728 43944
rect 792 43880 808 43944
rect 872 43880 888 43944
rect 952 43880 968 43944
rect 1032 43880 1048 43944
rect 1112 43880 1128 43944
rect 1192 43880 1208 43944
rect 1272 43880 1288 43944
rect 1352 43880 1368 43944
rect 1432 43880 1448 43944
rect 1512 43880 1528 43944
rect 1592 43880 1608 43944
rect 1672 43880 1688 43944
rect 1752 43880 1768 43944
rect 1832 43880 1848 43944
rect 1912 43880 1928 43944
rect 1992 43880 2008 43944
rect 2072 43880 2088 43944
rect 2152 43880 2168 43944
rect 2232 43880 2248 43944
rect 2312 43880 2328 43944
rect 2392 43880 2408 43944
rect 2472 43880 2488 43944
rect 2552 43880 2568 43944
rect 2632 43880 2648 43944
rect 2712 43880 2728 43944
rect 2792 43880 2808 43944
rect 2872 43880 2888 43944
rect 2952 43880 2968 43944
rect 3032 43880 3048 43944
rect 3112 43880 3128 43944
rect 3192 43880 3208 43944
rect 3272 43880 3288 43944
rect 3352 43880 3368 43944
rect 3432 43880 3448 43944
rect 3512 43880 3528 43944
rect 3592 43880 3608 43944
rect 3672 43880 3688 43944
rect 3752 43880 3768 43944
rect 3832 43880 3848 43944
rect 3912 43880 3928 43944
rect 3992 43880 19112 43944
rect 19176 43880 19192 43944
rect 19256 43880 19272 43944
rect 19336 43880 19352 43944
rect 19416 43880 29112 43944
rect 29176 43880 29192 43944
rect 29256 43880 29272 43944
rect 29336 43880 29352 43944
rect 29416 43880 41376 43944
rect 41440 43880 41456 43944
rect 41520 43880 41536 43944
rect 41600 43880 41616 43944
rect 41680 43880 41696 43944
rect 41760 43880 41776 43944
rect 41840 43880 41856 43944
rect 41920 43880 41936 43944
rect 42000 43880 42016 43944
rect 42080 43880 42096 43944
rect 42160 43880 42176 43944
rect 42240 43880 42256 43944
rect 42320 43880 42336 43944
rect 42400 43880 42416 43944
rect 42480 43880 42496 43944
rect 42560 43880 42576 43944
rect 42640 43880 42656 43944
rect 42720 43880 42736 43944
rect 42800 43880 42816 43944
rect 42880 43880 42896 43944
rect 42960 43880 42976 43944
rect 43040 43880 43056 43944
rect 43120 43880 43136 43944
rect 43200 43880 43216 43944
rect 43280 43880 43296 43944
rect 43360 43880 43376 43944
rect 43440 43880 43456 43944
rect 43520 43880 43536 43944
rect 43600 43880 43616 43944
rect 43680 43880 43696 43944
rect 43760 43880 43776 43944
rect 43840 43880 43856 43944
rect 43920 43880 43936 43944
rect 44000 43880 44016 43944
rect 44080 43880 44096 43944
rect 44160 43880 44176 43944
rect 44240 43880 44256 43944
rect 44320 43880 44336 43944
rect 44400 43880 44416 43944
rect 44480 43880 44496 43944
rect 44560 43880 44576 43944
rect 44640 43880 44656 43944
rect 44720 43880 44736 43944
rect 44800 43880 44816 43944
rect 44880 43880 44896 43944
rect 44960 43880 44976 43944
rect 45040 43880 45056 43944
rect 45120 43880 45136 43944
rect 45200 43880 45216 43944
rect 45280 43880 45296 43944
rect 45360 43880 45368 43944
rect 0 43864 45368 43880
rect 0 43800 8 43864
rect 72 43800 88 43864
rect 152 43800 168 43864
rect 232 43800 248 43864
rect 312 43800 328 43864
rect 392 43800 408 43864
rect 472 43800 488 43864
rect 552 43800 568 43864
rect 632 43800 648 43864
rect 712 43800 728 43864
rect 792 43800 808 43864
rect 872 43800 888 43864
rect 952 43800 968 43864
rect 1032 43800 1048 43864
rect 1112 43800 1128 43864
rect 1192 43800 1208 43864
rect 1272 43800 1288 43864
rect 1352 43800 1368 43864
rect 1432 43800 1448 43864
rect 1512 43800 1528 43864
rect 1592 43800 1608 43864
rect 1672 43800 1688 43864
rect 1752 43800 1768 43864
rect 1832 43800 1848 43864
rect 1912 43800 1928 43864
rect 1992 43800 2008 43864
rect 2072 43800 2088 43864
rect 2152 43800 2168 43864
rect 2232 43800 2248 43864
rect 2312 43800 2328 43864
rect 2392 43800 2408 43864
rect 2472 43800 2488 43864
rect 2552 43800 2568 43864
rect 2632 43800 2648 43864
rect 2712 43800 2728 43864
rect 2792 43800 2808 43864
rect 2872 43800 2888 43864
rect 2952 43800 2968 43864
rect 3032 43800 3048 43864
rect 3112 43800 3128 43864
rect 3192 43800 3208 43864
rect 3272 43800 3288 43864
rect 3352 43800 3368 43864
rect 3432 43800 3448 43864
rect 3512 43800 3528 43864
rect 3592 43800 3608 43864
rect 3672 43800 3688 43864
rect 3752 43800 3768 43864
rect 3832 43800 3848 43864
rect 3912 43800 3928 43864
rect 3992 43800 19112 43864
rect 19176 43800 19192 43864
rect 19256 43800 19272 43864
rect 19336 43800 19352 43864
rect 19416 43800 29112 43864
rect 29176 43800 29192 43864
rect 29256 43800 29272 43864
rect 29336 43800 29352 43864
rect 29416 43800 41376 43864
rect 41440 43800 41456 43864
rect 41520 43800 41536 43864
rect 41600 43800 41616 43864
rect 41680 43800 41696 43864
rect 41760 43800 41776 43864
rect 41840 43800 41856 43864
rect 41920 43800 41936 43864
rect 42000 43800 42016 43864
rect 42080 43800 42096 43864
rect 42160 43800 42176 43864
rect 42240 43800 42256 43864
rect 42320 43800 42336 43864
rect 42400 43800 42416 43864
rect 42480 43800 42496 43864
rect 42560 43800 42576 43864
rect 42640 43800 42656 43864
rect 42720 43800 42736 43864
rect 42800 43800 42816 43864
rect 42880 43800 42896 43864
rect 42960 43800 42976 43864
rect 43040 43800 43056 43864
rect 43120 43800 43136 43864
rect 43200 43800 43216 43864
rect 43280 43800 43296 43864
rect 43360 43800 43376 43864
rect 43440 43800 43456 43864
rect 43520 43800 43536 43864
rect 43600 43800 43616 43864
rect 43680 43800 43696 43864
rect 43760 43800 43776 43864
rect 43840 43800 43856 43864
rect 43920 43800 43936 43864
rect 44000 43800 44016 43864
rect 44080 43800 44096 43864
rect 44160 43800 44176 43864
rect 44240 43800 44256 43864
rect 44320 43800 44336 43864
rect 44400 43800 44416 43864
rect 44480 43800 44496 43864
rect 44560 43800 44576 43864
rect 44640 43800 44656 43864
rect 44720 43800 44736 43864
rect 44800 43800 44816 43864
rect 44880 43800 44896 43864
rect 44960 43800 44976 43864
rect 45040 43800 45056 43864
rect 45120 43800 45136 43864
rect 45200 43800 45216 43864
rect 45280 43800 45296 43864
rect 45360 43800 45368 43864
rect 0 43784 45368 43800
rect 0 43720 8 43784
rect 72 43720 88 43784
rect 152 43720 168 43784
rect 232 43720 248 43784
rect 312 43720 328 43784
rect 392 43720 408 43784
rect 472 43720 488 43784
rect 552 43720 568 43784
rect 632 43720 648 43784
rect 712 43720 728 43784
rect 792 43720 808 43784
rect 872 43720 888 43784
rect 952 43720 968 43784
rect 1032 43720 1048 43784
rect 1112 43720 1128 43784
rect 1192 43720 1208 43784
rect 1272 43720 1288 43784
rect 1352 43720 1368 43784
rect 1432 43720 1448 43784
rect 1512 43720 1528 43784
rect 1592 43720 1608 43784
rect 1672 43720 1688 43784
rect 1752 43720 1768 43784
rect 1832 43720 1848 43784
rect 1912 43720 1928 43784
rect 1992 43720 2008 43784
rect 2072 43720 2088 43784
rect 2152 43720 2168 43784
rect 2232 43720 2248 43784
rect 2312 43720 2328 43784
rect 2392 43720 2408 43784
rect 2472 43720 2488 43784
rect 2552 43720 2568 43784
rect 2632 43720 2648 43784
rect 2712 43720 2728 43784
rect 2792 43720 2808 43784
rect 2872 43720 2888 43784
rect 2952 43720 2968 43784
rect 3032 43720 3048 43784
rect 3112 43720 3128 43784
rect 3192 43720 3208 43784
rect 3272 43720 3288 43784
rect 3352 43720 3368 43784
rect 3432 43720 3448 43784
rect 3512 43720 3528 43784
rect 3592 43720 3608 43784
rect 3672 43720 3688 43784
rect 3752 43720 3768 43784
rect 3832 43720 3848 43784
rect 3912 43720 3928 43784
rect 3992 43720 19112 43784
rect 19176 43720 19192 43784
rect 19256 43720 19272 43784
rect 19336 43720 19352 43784
rect 19416 43720 29112 43784
rect 29176 43720 29192 43784
rect 29256 43720 29272 43784
rect 29336 43720 29352 43784
rect 29416 43720 41376 43784
rect 41440 43720 41456 43784
rect 41520 43720 41536 43784
rect 41600 43720 41616 43784
rect 41680 43720 41696 43784
rect 41760 43720 41776 43784
rect 41840 43720 41856 43784
rect 41920 43720 41936 43784
rect 42000 43720 42016 43784
rect 42080 43720 42096 43784
rect 42160 43720 42176 43784
rect 42240 43720 42256 43784
rect 42320 43720 42336 43784
rect 42400 43720 42416 43784
rect 42480 43720 42496 43784
rect 42560 43720 42576 43784
rect 42640 43720 42656 43784
rect 42720 43720 42736 43784
rect 42800 43720 42816 43784
rect 42880 43720 42896 43784
rect 42960 43720 42976 43784
rect 43040 43720 43056 43784
rect 43120 43720 43136 43784
rect 43200 43720 43216 43784
rect 43280 43720 43296 43784
rect 43360 43720 43376 43784
rect 43440 43720 43456 43784
rect 43520 43720 43536 43784
rect 43600 43720 43616 43784
rect 43680 43720 43696 43784
rect 43760 43720 43776 43784
rect 43840 43720 43856 43784
rect 43920 43720 43936 43784
rect 44000 43720 44016 43784
rect 44080 43720 44096 43784
rect 44160 43720 44176 43784
rect 44240 43720 44256 43784
rect 44320 43720 44336 43784
rect 44400 43720 44416 43784
rect 44480 43720 44496 43784
rect 44560 43720 44576 43784
rect 44640 43720 44656 43784
rect 44720 43720 44736 43784
rect 44800 43720 44816 43784
rect 44880 43720 44896 43784
rect 44960 43720 44976 43784
rect 45040 43720 45056 43784
rect 45120 43720 45136 43784
rect 45200 43720 45216 43784
rect 45280 43720 45296 43784
rect 45360 43720 45368 43784
rect 0 43704 45368 43720
rect 0 43640 8 43704
rect 72 43640 88 43704
rect 152 43640 168 43704
rect 232 43640 248 43704
rect 312 43640 328 43704
rect 392 43640 408 43704
rect 472 43640 488 43704
rect 552 43640 568 43704
rect 632 43640 648 43704
rect 712 43640 728 43704
rect 792 43640 808 43704
rect 872 43640 888 43704
rect 952 43640 968 43704
rect 1032 43640 1048 43704
rect 1112 43640 1128 43704
rect 1192 43640 1208 43704
rect 1272 43640 1288 43704
rect 1352 43640 1368 43704
rect 1432 43640 1448 43704
rect 1512 43640 1528 43704
rect 1592 43640 1608 43704
rect 1672 43640 1688 43704
rect 1752 43640 1768 43704
rect 1832 43640 1848 43704
rect 1912 43640 1928 43704
rect 1992 43640 2008 43704
rect 2072 43640 2088 43704
rect 2152 43640 2168 43704
rect 2232 43640 2248 43704
rect 2312 43640 2328 43704
rect 2392 43640 2408 43704
rect 2472 43640 2488 43704
rect 2552 43640 2568 43704
rect 2632 43640 2648 43704
rect 2712 43640 2728 43704
rect 2792 43640 2808 43704
rect 2872 43640 2888 43704
rect 2952 43640 2968 43704
rect 3032 43640 3048 43704
rect 3112 43640 3128 43704
rect 3192 43640 3208 43704
rect 3272 43640 3288 43704
rect 3352 43640 3368 43704
rect 3432 43640 3448 43704
rect 3512 43640 3528 43704
rect 3592 43640 3608 43704
rect 3672 43640 3688 43704
rect 3752 43640 3768 43704
rect 3832 43640 3848 43704
rect 3912 43640 3928 43704
rect 3992 43640 19112 43704
rect 19176 43640 19192 43704
rect 19256 43640 19272 43704
rect 19336 43640 19352 43704
rect 19416 43640 29112 43704
rect 29176 43640 29192 43704
rect 29256 43640 29272 43704
rect 29336 43640 29352 43704
rect 29416 43640 41376 43704
rect 41440 43640 41456 43704
rect 41520 43640 41536 43704
rect 41600 43640 41616 43704
rect 41680 43640 41696 43704
rect 41760 43640 41776 43704
rect 41840 43640 41856 43704
rect 41920 43640 41936 43704
rect 42000 43640 42016 43704
rect 42080 43640 42096 43704
rect 42160 43640 42176 43704
rect 42240 43640 42256 43704
rect 42320 43640 42336 43704
rect 42400 43640 42416 43704
rect 42480 43640 42496 43704
rect 42560 43640 42576 43704
rect 42640 43640 42656 43704
rect 42720 43640 42736 43704
rect 42800 43640 42816 43704
rect 42880 43640 42896 43704
rect 42960 43640 42976 43704
rect 43040 43640 43056 43704
rect 43120 43640 43136 43704
rect 43200 43640 43216 43704
rect 43280 43640 43296 43704
rect 43360 43640 43376 43704
rect 43440 43640 43456 43704
rect 43520 43640 43536 43704
rect 43600 43640 43616 43704
rect 43680 43640 43696 43704
rect 43760 43640 43776 43704
rect 43840 43640 43856 43704
rect 43920 43640 43936 43704
rect 44000 43640 44016 43704
rect 44080 43640 44096 43704
rect 44160 43640 44176 43704
rect 44240 43640 44256 43704
rect 44320 43640 44336 43704
rect 44400 43640 44416 43704
rect 44480 43640 44496 43704
rect 44560 43640 44576 43704
rect 44640 43640 44656 43704
rect 44720 43640 44736 43704
rect 44800 43640 44816 43704
rect 44880 43640 44896 43704
rect 44960 43640 44976 43704
rect 45040 43640 45056 43704
rect 45120 43640 45136 43704
rect 45200 43640 45216 43704
rect 45280 43640 45296 43704
rect 45360 43640 45368 43704
rect 0 43624 45368 43640
rect 0 43560 8 43624
rect 72 43560 88 43624
rect 152 43560 168 43624
rect 232 43560 248 43624
rect 312 43560 328 43624
rect 392 43560 408 43624
rect 472 43560 488 43624
rect 552 43560 568 43624
rect 632 43560 648 43624
rect 712 43560 728 43624
rect 792 43560 808 43624
rect 872 43560 888 43624
rect 952 43560 968 43624
rect 1032 43560 1048 43624
rect 1112 43560 1128 43624
rect 1192 43560 1208 43624
rect 1272 43560 1288 43624
rect 1352 43560 1368 43624
rect 1432 43560 1448 43624
rect 1512 43560 1528 43624
rect 1592 43560 1608 43624
rect 1672 43560 1688 43624
rect 1752 43560 1768 43624
rect 1832 43560 1848 43624
rect 1912 43560 1928 43624
rect 1992 43560 2008 43624
rect 2072 43560 2088 43624
rect 2152 43560 2168 43624
rect 2232 43560 2248 43624
rect 2312 43560 2328 43624
rect 2392 43560 2408 43624
rect 2472 43560 2488 43624
rect 2552 43560 2568 43624
rect 2632 43560 2648 43624
rect 2712 43560 2728 43624
rect 2792 43560 2808 43624
rect 2872 43560 2888 43624
rect 2952 43560 2968 43624
rect 3032 43560 3048 43624
rect 3112 43560 3128 43624
rect 3192 43560 3208 43624
rect 3272 43560 3288 43624
rect 3352 43560 3368 43624
rect 3432 43560 3448 43624
rect 3512 43560 3528 43624
rect 3592 43560 3608 43624
rect 3672 43560 3688 43624
rect 3752 43560 3768 43624
rect 3832 43560 3848 43624
rect 3912 43560 3928 43624
rect 3992 43560 19112 43624
rect 19176 43560 19192 43624
rect 19256 43560 19272 43624
rect 19336 43560 19352 43624
rect 19416 43560 29112 43624
rect 29176 43560 29192 43624
rect 29256 43560 29272 43624
rect 29336 43560 29352 43624
rect 29416 43560 41376 43624
rect 41440 43560 41456 43624
rect 41520 43560 41536 43624
rect 41600 43560 41616 43624
rect 41680 43560 41696 43624
rect 41760 43560 41776 43624
rect 41840 43560 41856 43624
rect 41920 43560 41936 43624
rect 42000 43560 42016 43624
rect 42080 43560 42096 43624
rect 42160 43560 42176 43624
rect 42240 43560 42256 43624
rect 42320 43560 42336 43624
rect 42400 43560 42416 43624
rect 42480 43560 42496 43624
rect 42560 43560 42576 43624
rect 42640 43560 42656 43624
rect 42720 43560 42736 43624
rect 42800 43560 42816 43624
rect 42880 43560 42896 43624
rect 42960 43560 42976 43624
rect 43040 43560 43056 43624
rect 43120 43560 43136 43624
rect 43200 43560 43216 43624
rect 43280 43560 43296 43624
rect 43360 43560 43376 43624
rect 43440 43560 43456 43624
rect 43520 43560 43536 43624
rect 43600 43560 43616 43624
rect 43680 43560 43696 43624
rect 43760 43560 43776 43624
rect 43840 43560 43856 43624
rect 43920 43560 43936 43624
rect 44000 43560 44016 43624
rect 44080 43560 44096 43624
rect 44160 43560 44176 43624
rect 44240 43560 44256 43624
rect 44320 43560 44336 43624
rect 44400 43560 44416 43624
rect 44480 43560 44496 43624
rect 44560 43560 44576 43624
rect 44640 43560 44656 43624
rect 44720 43560 44736 43624
rect 44800 43560 44816 43624
rect 44880 43560 44896 43624
rect 44960 43560 44976 43624
rect 45040 43560 45056 43624
rect 45120 43560 45136 43624
rect 45200 43560 45216 43624
rect 45280 43560 45296 43624
rect 45360 43560 45368 43624
rect 0 43544 45368 43560
rect 0 43480 8 43544
rect 72 43480 88 43544
rect 152 43480 168 43544
rect 232 43480 248 43544
rect 312 43480 328 43544
rect 392 43480 408 43544
rect 472 43480 488 43544
rect 552 43480 568 43544
rect 632 43480 648 43544
rect 712 43480 728 43544
rect 792 43480 808 43544
rect 872 43480 888 43544
rect 952 43480 968 43544
rect 1032 43480 1048 43544
rect 1112 43480 1128 43544
rect 1192 43480 1208 43544
rect 1272 43480 1288 43544
rect 1352 43480 1368 43544
rect 1432 43480 1448 43544
rect 1512 43480 1528 43544
rect 1592 43480 1608 43544
rect 1672 43480 1688 43544
rect 1752 43480 1768 43544
rect 1832 43480 1848 43544
rect 1912 43480 1928 43544
rect 1992 43480 2008 43544
rect 2072 43480 2088 43544
rect 2152 43480 2168 43544
rect 2232 43480 2248 43544
rect 2312 43480 2328 43544
rect 2392 43480 2408 43544
rect 2472 43480 2488 43544
rect 2552 43480 2568 43544
rect 2632 43480 2648 43544
rect 2712 43480 2728 43544
rect 2792 43480 2808 43544
rect 2872 43480 2888 43544
rect 2952 43480 2968 43544
rect 3032 43480 3048 43544
rect 3112 43480 3128 43544
rect 3192 43480 3208 43544
rect 3272 43480 3288 43544
rect 3352 43480 3368 43544
rect 3432 43480 3448 43544
rect 3512 43480 3528 43544
rect 3592 43480 3608 43544
rect 3672 43480 3688 43544
rect 3752 43480 3768 43544
rect 3832 43480 3848 43544
rect 3912 43480 3928 43544
rect 3992 43480 19112 43544
rect 19176 43480 19192 43544
rect 19256 43480 19272 43544
rect 19336 43480 19352 43544
rect 19416 43480 29112 43544
rect 29176 43480 29192 43544
rect 29256 43480 29272 43544
rect 29336 43480 29352 43544
rect 29416 43480 41376 43544
rect 41440 43480 41456 43544
rect 41520 43480 41536 43544
rect 41600 43480 41616 43544
rect 41680 43480 41696 43544
rect 41760 43480 41776 43544
rect 41840 43480 41856 43544
rect 41920 43480 41936 43544
rect 42000 43480 42016 43544
rect 42080 43480 42096 43544
rect 42160 43480 42176 43544
rect 42240 43480 42256 43544
rect 42320 43480 42336 43544
rect 42400 43480 42416 43544
rect 42480 43480 42496 43544
rect 42560 43480 42576 43544
rect 42640 43480 42656 43544
rect 42720 43480 42736 43544
rect 42800 43480 42816 43544
rect 42880 43480 42896 43544
rect 42960 43480 42976 43544
rect 43040 43480 43056 43544
rect 43120 43480 43136 43544
rect 43200 43480 43216 43544
rect 43280 43480 43296 43544
rect 43360 43480 43376 43544
rect 43440 43480 43456 43544
rect 43520 43480 43536 43544
rect 43600 43480 43616 43544
rect 43680 43480 43696 43544
rect 43760 43480 43776 43544
rect 43840 43480 43856 43544
rect 43920 43480 43936 43544
rect 44000 43480 44016 43544
rect 44080 43480 44096 43544
rect 44160 43480 44176 43544
rect 44240 43480 44256 43544
rect 44320 43480 44336 43544
rect 44400 43480 44416 43544
rect 44480 43480 44496 43544
rect 44560 43480 44576 43544
rect 44640 43480 44656 43544
rect 44720 43480 44736 43544
rect 44800 43480 44816 43544
rect 44880 43480 44896 43544
rect 44960 43480 44976 43544
rect 45040 43480 45056 43544
rect 45120 43480 45136 43544
rect 45200 43480 45216 43544
rect 45280 43480 45296 43544
rect 45360 43480 45368 43544
rect 0 43464 45368 43480
rect 0 43400 8 43464
rect 72 43400 88 43464
rect 152 43400 168 43464
rect 232 43400 248 43464
rect 312 43400 328 43464
rect 392 43400 408 43464
rect 472 43400 488 43464
rect 552 43400 568 43464
rect 632 43400 648 43464
rect 712 43400 728 43464
rect 792 43400 808 43464
rect 872 43400 888 43464
rect 952 43400 968 43464
rect 1032 43400 1048 43464
rect 1112 43400 1128 43464
rect 1192 43400 1208 43464
rect 1272 43400 1288 43464
rect 1352 43400 1368 43464
rect 1432 43400 1448 43464
rect 1512 43400 1528 43464
rect 1592 43400 1608 43464
rect 1672 43400 1688 43464
rect 1752 43400 1768 43464
rect 1832 43400 1848 43464
rect 1912 43400 1928 43464
rect 1992 43400 2008 43464
rect 2072 43400 2088 43464
rect 2152 43400 2168 43464
rect 2232 43400 2248 43464
rect 2312 43400 2328 43464
rect 2392 43400 2408 43464
rect 2472 43400 2488 43464
rect 2552 43400 2568 43464
rect 2632 43400 2648 43464
rect 2712 43400 2728 43464
rect 2792 43400 2808 43464
rect 2872 43400 2888 43464
rect 2952 43400 2968 43464
rect 3032 43400 3048 43464
rect 3112 43400 3128 43464
rect 3192 43400 3208 43464
rect 3272 43400 3288 43464
rect 3352 43400 3368 43464
rect 3432 43400 3448 43464
rect 3512 43400 3528 43464
rect 3592 43400 3608 43464
rect 3672 43400 3688 43464
rect 3752 43400 3768 43464
rect 3832 43400 3848 43464
rect 3912 43400 3928 43464
rect 3992 43400 19112 43464
rect 19176 43400 19192 43464
rect 19256 43400 19272 43464
rect 19336 43400 19352 43464
rect 19416 43400 29112 43464
rect 29176 43400 29192 43464
rect 29256 43400 29272 43464
rect 29336 43400 29352 43464
rect 29416 43400 41376 43464
rect 41440 43400 41456 43464
rect 41520 43400 41536 43464
rect 41600 43400 41616 43464
rect 41680 43400 41696 43464
rect 41760 43400 41776 43464
rect 41840 43400 41856 43464
rect 41920 43400 41936 43464
rect 42000 43400 42016 43464
rect 42080 43400 42096 43464
rect 42160 43400 42176 43464
rect 42240 43400 42256 43464
rect 42320 43400 42336 43464
rect 42400 43400 42416 43464
rect 42480 43400 42496 43464
rect 42560 43400 42576 43464
rect 42640 43400 42656 43464
rect 42720 43400 42736 43464
rect 42800 43400 42816 43464
rect 42880 43400 42896 43464
rect 42960 43400 42976 43464
rect 43040 43400 43056 43464
rect 43120 43400 43136 43464
rect 43200 43400 43216 43464
rect 43280 43400 43296 43464
rect 43360 43400 43376 43464
rect 43440 43400 43456 43464
rect 43520 43400 43536 43464
rect 43600 43400 43616 43464
rect 43680 43400 43696 43464
rect 43760 43400 43776 43464
rect 43840 43400 43856 43464
rect 43920 43400 43936 43464
rect 44000 43400 44016 43464
rect 44080 43400 44096 43464
rect 44160 43400 44176 43464
rect 44240 43400 44256 43464
rect 44320 43400 44336 43464
rect 44400 43400 44416 43464
rect 44480 43400 44496 43464
rect 44560 43400 44576 43464
rect 44640 43400 44656 43464
rect 44720 43400 44736 43464
rect 44800 43400 44816 43464
rect 44880 43400 44896 43464
rect 44960 43400 44976 43464
rect 45040 43400 45056 43464
rect 45120 43400 45136 43464
rect 45200 43400 45216 43464
rect 45280 43400 45296 43464
rect 45360 43400 45368 43464
rect 0 43384 45368 43400
rect 0 43320 8 43384
rect 72 43320 88 43384
rect 152 43320 168 43384
rect 232 43320 248 43384
rect 312 43320 328 43384
rect 392 43320 408 43384
rect 472 43320 488 43384
rect 552 43320 568 43384
rect 632 43320 648 43384
rect 712 43320 728 43384
rect 792 43320 808 43384
rect 872 43320 888 43384
rect 952 43320 968 43384
rect 1032 43320 1048 43384
rect 1112 43320 1128 43384
rect 1192 43320 1208 43384
rect 1272 43320 1288 43384
rect 1352 43320 1368 43384
rect 1432 43320 1448 43384
rect 1512 43320 1528 43384
rect 1592 43320 1608 43384
rect 1672 43320 1688 43384
rect 1752 43320 1768 43384
rect 1832 43320 1848 43384
rect 1912 43320 1928 43384
rect 1992 43320 2008 43384
rect 2072 43320 2088 43384
rect 2152 43320 2168 43384
rect 2232 43320 2248 43384
rect 2312 43320 2328 43384
rect 2392 43320 2408 43384
rect 2472 43320 2488 43384
rect 2552 43320 2568 43384
rect 2632 43320 2648 43384
rect 2712 43320 2728 43384
rect 2792 43320 2808 43384
rect 2872 43320 2888 43384
rect 2952 43320 2968 43384
rect 3032 43320 3048 43384
rect 3112 43320 3128 43384
rect 3192 43320 3208 43384
rect 3272 43320 3288 43384
rect 3352 43320 3368 43384
rect 3432 43320 3448 43384
rect 3512 43320 3528 43384
rect 3592 43320 3608 43384
rect 3672 43320 3688 43384
rect 3752 43320 3768 43384
rect 3832 43320 3848 43384
rect 3912 43320 3928 43384
rect 3992 43320 19112 43384
rect 19176 43320 19192 43384
rect 19256 43320 19272 43384
rect 19336 43320 19352 43384
rect 19416 43320 29112 43384
rect 29176 43320 29192 43384
rect 29256 43320 29272 43384
rect 29336 43320 29352 43384
rect 29416 43320 41376 43384
rect 41440 43320 41456 43384
rect 41520 43320 41536 43384
rect 41600 43320 41616 43384
rect 41680 43320 41696 43384
rect 41760 43320 41776 43384
rect 41840 43320 41856 43384
rect 41920 43320 41936 43384
rect 42000 43320 42016 43384
rect 42080 43320 42096 43384
rect 42160 43320 42176 43384
rect 42240 43320 42256 43384
rect 42320 43320 42336 43384
rect 42400 43320 42416 43384
rect 42480 43320 42496 43384
rect 42560 43320 42576 43384
rect 42640 43320 42656 43384
rect 42720 43320 42736 43384
rect 42800 43320 42816 43384
rect 42880 43320 42896 43384
rect 42960 43320 42976 43384
rect 43040 43320 43056 43384
rect 43120 43320 43136 43384
rect 43200 43320 43216 43384
rect 43280 43320 43296 43384
rect 43360 43320 43376 43384
rect 43440 43320 43456 43384
rect 43520 43320 43536 43384
rect 43600 43320 43616 43384
rect 43680 43320 43696 43384
rect 43760 43320 43776 43384
rect 43840 43320 43856 43384
rect 43920 43320 43936 43384
rect 44000 43320 44016 43384
rect 44080 43320 44096 43384
rect 44160 43320 44176 43384
rect 44240 43320 44256 43384
rect 44320 43320 44336 43384
rect 44400 43320 44416 43384
rect 44480 43320 44496 43384
rect 44560 43320 44576 43384
rect 44640 43320 44656 43384
rect 44720 43320 44736 43384
rect 44800 43320 44816 43384
rect 44880 43320 44896 43384
rect 44960 43320 44976 43384
rect 45040 43320 45056 43384
rect 45120 43320 45136 43384
rect 45200 43320 45216 43384
rect 45280 43320 45296 43384
rect 45360 43320 45368 43384
rect 0 43304 45368 43320
rect 0 43240 8 43304
rect 72 43240 88 43304
rect 152 43240 168 43304
rect 232 43240 248 43304
rect 312 43240 328 43304
rect 392 43240 408 43304
rect 472 43240 488 43304
rect 552 43240 568 43304
rect 632 43240 648 43304
rect 712 43240 728 43304
rect 792 43240 808 43304
rect 872 43240 888 43304
rect 952 43240 968 43304
rect 1032 43240 1048 43304
rect 1112 43240 1128 43304
rect 1192 43240 1208 43304
rect 1272 43240 1288 43304
rect 1352 43240 1368 43304
rect 1432 43240 1448 43304
rect 1512 43240 1528 43304
rect 1592 43240 1608 43304
rect 1672 43240 1688 43304
rect 1752 43240 1768 43304
rect 1832 43240 1848 43304
rect 1912 43240 1928 43304
rect 1992 43240 2008 43304
rect 2072 43240 2088 43304
rect 2152 43240 2168 43304
rect 2232 43240 2248 43304
rect 2312 43240 2328 43304
rect 2392 43240 2408 43304
rect 2472 43240 2488 43304
rect 2552 43240 2568 43304
rect 2632 43240 2648 43304
rect 2712 43240 2728 43304
rect 2792 43240 2808 43304
rect 2872 43240 2888 43304
rect 2952 43240 2968 43304
rect 3032 43240 3048 43304
rect 3112 43240 3128 43304
rect 3192 43240 3208 43304
rect 3272 43240 3288 43304
rect 3352 43240 3368 43304
rect 3432 43240 3448 43304
rect 3512 43240 3528 43304
rect 3592 43240 3608 43304
rect 3672 43240 3688 43304
rect 3752 43240 3768 43304
rect 3832 43240 3848 43304
rect 3912 43240 3928 43304
rect 3992 43240 19112 43304
rect 19176 43240 19192 43304
rect 19256 43240 19272 43304
rect 19336 43240 19352 43304
rect 19416 43240 29112 43304
rect 29176 43240 29192 43304
rect 29256 43240 29272 43304
rect 29336 43240 29352 43304
rect 29416 43240 41376 43304
rect 41440 43240 41456 43304
rect 41520 43240 41536 43304
rect 41600 43240 41616 43304
rect 41680 43240 41696 43304
rect 41760 43240 41776 43304
rect 41840 43240 41856 43304
rect 41920 43240 41936 43304
rect 42000 43240 42016 43304
rect 42080 43240 42096 43304
rect 42160 43240 42176 43304
rect 42240 43240 42256 43304
rect 42320 43240 42336 43304
rect 42400 43240 42416 43304
rect 42480 43240 42496 43304
rect 42560 43240 42576 43304
rect 42640 43240 42656 43304
rect 42720 43240 42736 43304
rect 42800 43240 42816 43304
rect 42880 43240 42896 43304
rect 42960 43240 42976 43304
rect 43040 43240 43056 43304
rect 43120 43240 43136 43304
rect 43200 43240 43216 43304
rect 43280 43240 43296 43304
rect 43360 43240 43376 43304
rect 43440 43240 43456 43304
rect 43520 43240 43536 43304
rect 43600 43240 43616 43304
rect 43680 43240 43696 43304
rect 43760 43240 43776 43304
rect 43840 43240 43856 43304
rect 43920 43240 43936 43304
rect 44000 43240 44016 43304
rect 44080 43240 44096 43304
rect 44160 43240 44176 43304
rect 44240 43240 44256 43304
rect 44320 43240 44336 43304
rect 44400 43240 44416 43304
rect 44480 43240 44496 43304
rect 44560 43240 44576 43304
rect 44640 43240 44656 43304
rect 44720 43240 44736 43304
rect 44800 43240 44816 43304
rect 44880 43240 44896 43304
rect 44960 43240 44976 43304
rect 45040 43240 45056 43304
rect 45120 43240 45136 43304
rect 45200 43240 45216 43304
rect 45280 43240 45296 43304
rect 45360 43240 45368 43304
rect 0 43224 45368 43240
rect 0 43160 8 43224
rect 72 43160 88 43224
rect 152 43160 168 43224
rect 232 43160 248 43224
rect 312 43160 328 43224
rect 392 43160 408 43224
rect 472 43160 488 43224
rect 552 43160 568 43224
rect 632 43160 648 43224
rect 712 43160 728 43224
rect 792 43160 808 43224
rect 872 43160 888 43224
rect 952 43160 968 43224
rect 1032 43160 1048 43224
rect 1112 43160 1128 43224
rect 1192 43160 1208 43224
rect 1272 43160 1288 43224
rect 1352 43160 1368 43224
rect 1432 43160 1448 43224
rect 1512 43160 1528 43224
rect 1592 43160 1608 43224
rect 1672 43160 1688 43224
rect 1752 43160 1768 43224
rect 1832 43160 1848 43224
rect 1912 43160 1928 43224
rect 1992 43160 2008 43224
rect 2072 43160 2088 43224
rect 2152 43160 2168 43224
rect 2232 43160 2248 43224
rect 2312 43160 2328 43224
rect 2392 43160 2408 43224
rect 2472 43160 2488 43224
rect 2552 43160 2568 43224
rect 2632 43160 2648 43224
rect 2712 43160 2728 43224
rect 2792 43160 2808 43224
rect 2872 43160 2888 43224
rect 2952 43160 2968 43224
rect 3032 43160 3048 43224
rect 3112 43160 3128 43224
rect 3192 43160 3208 43224
rect 3272 43160 3288 43224
rect 3352 43160 3368 43224
rect 3432 43160 3448 43224
rect 3512 43160 3528 43224
rect 3592 43160 3608 43224
rect 3672 43160 3688 43224
rect 3752 43160 3768 43224
rect 3832 43160 3848 43224
rect 3912 43160 3928 43224
rect 3992 43160 19112 43224
rect 19176 43160 19192 43224
rect 19256 43160 19272 43224
rect 19336 43160 19352 43224
rect 19416 43160 29112 43224
rect 29176 43160 29192 43224
rect 29256 43160 29272 43224
rect 29336 43160 29352 43224
rect 29416 43160 41376 43224
rect 41440 43160 41456 43224
rect 41520 43160 41536 43224
rect 41600 43160 41616 43224
rect 41680 43160 41696 43224
rect 41760 43160 41776 43224
rect 41840 43160 41856 43224
rect 41920 43160 41936 43224
rect 42000 43160 42016 43224
rect 42080 43160 42096 43224
rect 42160 43160 42176 43224
rect 42240 43160 42256 43224
rect 42320 43160 42336 43224
rect 42400 43160 42416 43224
rect 42480 43160 42496 43224
rect 42560 43160 42576 43224
rect 42640 43160 42656 43224
rect 42720 43160 42736 43224
rect 42800 43160 42816 43224
rect 42880 43160 42896 43224
rect 42960 43160 42976 43224
rect 43040 43160 43056 43224
rect 43120 43160 43136 43224
rect 43200 43160 43216 43224
rect 43280 43160 43296 43224
rect 43360 43160 43376 43224
rect 43440 43160 43456 43224
rect 43520 43160 43536 43224
rect 43600 43160 43616 43224
rect 43680 43160 43696 43224
rect 43760 43160 43776 43224
rect 43840 43160 43856 43224
rect 43920 43160 43936 43224
rect 44000 43160 44016 43224
rect 44080 43160 44096 43224
rect 44160 43160 44176 43224
rect 44240 43160 44256 43224
rect 44320 43160 44336 43224
rect 44400 43160 44416 43224
rect 44480 43160 44496 43224
rect 44560 43160 44576 43224
rect 44640 43160 44656 43224
rect 44720 43160 44736 43224
rect 44800 43160 44816 43224
rect 44880 43160 44896 43224
rect 44960 43160 44976 43224
rect 45040 43160 45056 43224
rect 45120 43160 45136 43224
rect 45200 43160 45216 43224
rect 45280 43160 45296 43224
rect 45360 43160 45368 43224
rect 0 43144 45368 43160
rect 0 43080 8 43144
rect 72 43080 88 43144
rect 152 43080 168 43144
rect 232 43080 248 43144
rect 312 43080 328 43144
rect 392 43080 408 43144
rect 472 43080 488 43144
rect 552 43080 568 43144
rect 632 43080 648 43144
rect 712 43080 728 43144
rect 792 43080 808 43144
rect 872 43080 888 43144
rect 952 43080 968 43144
rect 1032 43080 1048 43144
rect 1112 43080 1128 43144
rect 1192 43080 1208 43144
rect 1272 43080 1288 43144
rect 1352 43080 1368 43144
rect 1432 43080 1448 43144
rect 1512 43080 1528 43144
rect 1592 43080 1608 43144
rect 1672 43080 1688 43144
rect 1752 43080 1768 43144
rect 1832 43080 1848 43144
rect 1912 43080 1928 43144
rect 1992 43080 2008 43144
rect 2072 43080 2088 43144
rect 2152 43080 2168 43144
rect 2232 43080 2248 43144
rect 2312 43080 2328 43144
rect 2392 43080 2408 43144
rect 2472 43080 2488 43144
rect 2552 43080 2568 43144
rect 2632 43080 2648 43144
rect 2712 43080 2728 43144
rect 2792 43080 2808 43144
rect 2872 43080 2888 43144
rect 2952 43080 2968 43144
rect 3032 43080 3048 43144
rect 3112 43080 3128 43144
rect 3192 43080 3208 43144
rect 3272 43080 3288 43144
rect 3352 43080 3368 43144
rect 3432 43080 3448 43144
rect 3512 43080 3528 43144
rect 3592 43080 3608 43144
rect 3672 43080 3688 43144
rect 3752 43080 3768 43144
rect 3832 43080 3848 43144
rect 3912 43080 3928 43144
rect 3992 43080 19112 43144
rect 19176 43080 19192 43144
rect 19256 43080 19272 43144
rect 19336 43080 19352 43144
rect 19416 43080 29112 43144
rect 29176 43080 29192 43144
rect 29256 43080 29272 43144
rect 29336 43080 29352 43144
rect 29416 43080 41376 43144
rect 41440 43080 41456 43144
rect 41520 43080 41536 43144
rect 41600 43080 41616 43144
rect 41680 43080 41696 43144
rect 41760 43080 41776 43144
rect 41840 43080 41856 43144
rect 41920 43080 41936 43144
rect 42000 43080 42016 43144
rect 42080 43080 42096 43144
rect 42160 43080 42176 43144
rect 42240 43080 42256 43144
rect 42320 43080 42336 43144
rect 42400 43080 42416 43144
rect 42480 43080 42496 43144
rect 42560 43080 42576 43144
rect 42640 43080 42656 43144
rect 42720 43080 42736 43144
rect 42800 43080 42816 43144
rect 42880 43080 42896 43144
rect 42960 43080 42976 43144
rect 43040 43080 43056 43144
rect 43120 43080 43136 43144
rect 43200 43080 43216 43144
rect 43280 43080 43296 43144
rect 43360 43080 43376 43144
rect 43440 43080 43456 43144
rect 43520 43080 43536 43144
rect 43600 43080 43616 43144
rect 43680 43080 43696 43144
rect 43760 43080 43776 43144
rect 43840 43080 43856 43144
rect 43920 43080 43936 43144
rect 44000 43080 44016 43144
rect 44080 43080 44096 43144
rect 44160 43080 44176 43144
rect 44240 43080 44256 43144
rect 44320 43080 44336 43144
rect 44400 43080 44416 43144
rect 44480 43080 44496 43144
rect 44560 43080 44576 43144
rect 44640 43080 44656 43144
rect 44720 43080 44736 43144
rect 44800 43080 44816 43144
rect 44880 43080 44896 43144
rect 44960 43080 44976 43144
rect 45040 43080 45056 43144
rect 45120 43080 45136 43144
rect 45200 43080 45216 43144
rect 45280 43080 45296 43144
rect 45360 43080 45368 43144
rect 0 43064 45368 43080
rect 0 43000 8 43064
rect 72 43000 88 43064
rect 152 43000 168 43064
rect 232 43000 248 43064
rect 312 43000 328 43064
rect 392 43000 408 43064
rect 472 43000 488 43064
rect 552 43000 568 43064
rect 632 43000 648 43064
rect 712 43000 728 43064
rect 792 43000 808 43064
rect 872 43000 888 43064
rect 952 43000 968 43064
rect 1032 43000 1048 43064
rect 1112 43000 1128 43064
rect 1192 43000 1208 43064
rect 1272 43000 1288 43064
rect 1352 43000 1368 43064
rect 1432 43000 1448 43064
rect 1512 43000 1528 43064
rect 1592 43000 1608 43064
rect 1672 43000 1688 43064
rect 1752 43000 1768 43064
rect 1832 43000 1848 43064
rect 1912 43000 1928 43064
rect 1992 43000 2008 43064
rect 2072 43000 2088 43064
rect 2152 43000 2168 43064
rect 2232 43000 2248 43064
rect 2312 43000 2328 43064
rect 2392 43000 2408 43064
rect 2472 43000 2488 43064
rect 2552 43000 2568 43064
rect 2632 43000 2648 43064
rect 2712 43000 2728 43064
rect 2792 43000 2808 43064
rect 2872 43000 2888 43064
rect 2952 43000 2968 43064
rect 3032 43000 3048 43064
rect 3112 43000 3128 43064
rect 3192 43000 3208 43064
rect 3272 43000 3288 43064
rect 3352 43000 3368 43064
rect 3432 43000 3448 43064
rect 3512 43000 3528 43064
rect 3592 43000 3608 43064
rect 3672 43000 3688 43064
rect 3752 43000 3768 43064
rect 3832 43000 3848 43064
rect 3912 43000 3928 43064
rect 3992 43000 19112 43064
rect 19176 43000 19192 43064
rect 19256 43000 19272 43064
rect 19336 43000 19352 43064
rect 19416 43000 29112 43064
rect 29176 43000 29192 43064
rect 29256 43000 29272 43064
rect 29336 43000 29352 43064
rect 29416 43000 41376 43064
rect 41440 43000 41456 43064
rect 41520 43000 41536 43064
rect 41600 43000 41616 43064
rect 41680 43000 41696 43064
rect 41760 43000 41776 43064
rect 41840 43000 41856 43064
rect 41920 43000 41936 43064
rect 42000 43000 42016 43064
rect 42080 43000 42096 43064
rect 42160 43000 42176 43064
rect 42240 43000 42256 43064
rect 42320 43000 42336 43064
rect 42400 43000 42416 43064
rect 42480 43000 42496 43064
rect 42560 43000 42576 43064
rect 42640 43000 42656 43064
rect 42720 43000 42736 43064
rect 42800 43000 42816 43064
rect 42880 43000 42896 43064
rect 42960 43000 42976 43064
rect 43040 43000 43056 43064
rect 43120 43000 43136 43064
rect 43200 43000 43216 43064
rect 43280 43000 43296 43064
rect 43360 43000 43376 43064
rect 43440 43000 43456 43064
rect 43520 43000 43536 43064
rect 43600 43000 43616 43064
rect 43680 43000 43696 43064
rect 43760 43000 43776 43064
rect 43840 43000 43856 43064
rect 43920 43000 43936 43064
rect 44000 43000 44016 43064
rect 44080 43000 44096 43064
rect 44160 43000 44176 43064
rect 44240 43000 44256 43064
rect 44320 43000 44336 43064
rect 44400 43000 44416 43064
rect 44480 43000 44496 43064
rect 44560 43000 44576 43064
rect 44640 43000 44656 43064
rect 44720 43000 44736 43064
rect 44800 43000 44816 43064
rect 44880 43000 44896 43064
rect 44960 43000 44976 43064
rect 45040 43000 45056 43064
rect 45120 43000 45136 43064
rect 45200 43000 45216 43064
rect 45280 43000 45296 43064
rect 45360 43000 45368 43064
rect 0 42984 45368 43000
rect 0 42920 8 42984
rect 72 42920 88 42984
rect 152 42920 168 42984
rect 232 42920 248 42984
rect 312 42920 328 42984
rect 392 42920 408 42984
rect 472 42920 488 42984
rect 552 42920 568 42984
rect 632 42920 648 42984
rect 712 42920 728 42984
rect 792 42920 808 42984
rect 872 42920 888 42984
rect 952 42920 968 42984
rect 1032 42920 1048 42984
rect 1112 42920 1128 42984
rect 1192 42920 1208 42984
rect 1272 42920 1288 42984
rect 1352 42920 1368 42984
rect 1432 42920 1448 42984
rect 1512 42920 1528 42984
rect 1592 42920 1608 42984
rect 1672 42920 1688 42984
rect 1752 42920 1768 42984
rect 1832 42920 1848 42984
rect 1912 42920 1928 42984
rect 1992 42920 2008 42984
rect 2072 42920 2088 42984
rect 2152 42920 2168 42984
rect 2232 42920 2248 42984
rect 2312 42920 2328 42984
rect 2392 42920 2408 42984
rect 2472 42920 2488 42984
rect 2552 42920 2568 42984
rect 2632 42920 2648 42984
rect 2712 42920 2728 42984
rect 2792 42920 2808 42984
rect 2872 42920 2888 42984
rect 2952 42920 2968 42984
rect 3032 42920 3048 42984
rect 3112 42920 3128 42984
rect 3192 42920 3208 42984
rect 3272 42920 3288 42984
rect 3352 42920 3368 42984
rect 3432 42920 3448 42984
rect 3512 42920 3528 42984
rect 3592 42920 3608 42984
rect 3672 42920 3688 42984
rect 3752 42920 3768 42984
rect 3832 42920 3848 42984
rect 3912 42920 3928 42984
rect 3992 42920 19112 42984
rect 19176 42920 19192 42984
rect 19256 42920 19272 42984
rect 19336 42920 19352 42984
rect 19416 42920 29112 42984
rect 29176 42920 29192 42984
rect 29256 42920 29272 42984
rect 29336 42920 29352 42984
rect 29416 42920 41376 42984
rect 41440 42920 41456 42984
rect 41520 42920 41536 42984
rect 41600 42920 41616 42984
rect 41680 42920 41696 42984
rect 41760 42920 41776 42984
rect 41840 42920 41856 42984
rect 41920 42920 41936 42984
rect 42000 42920 42016 42984
rect 42080 42920 42096 42984
rect 42160 42920 42176 42984
rect 42240 42920 42256 42984
rect 42320 42920 42336 42984
rect 42400 42920 42416 42984
rect 42480 42920 42496 42984
rect 42560 42920 42576 42984
rect 42640 42920 42656 42984
rect 42720 42920 42736 42984
rect 42800 42920 42816 42984
rect 42880 42920 42896 42984
rect 42960 42920 42976 42984
rect 43040 42920 43056 42984
rect 43120 42920 43136 42984
rect 43200 42920 43216 42984
rect 43280 42920 43296 42984
rect 43360 42920 43376 42984
rect 43440 42920 43456 42984
rect 43520 42920 43536 42984
rect 43600 42920 43616 42984
rect 43680 42920 43696 42984
rect 43760 42920 43776 42984
rect 43840 42920 43856 42984
rect 43920 42920 43936 42984
rect 44000 42920 44016 42984
rect 44080 42920 44096 42984
rect 44160 42920 44176 42984
rect 44240 42920 44256 42984
rect 44320 42920 44336 42984
rect 44400 42920 44416 42984
rect 44480 42920 44496 42984
rect 44560 42920 44576 42984
rect 44640 42920 44656 42984
rect 44720 42920 44736 42984
rect 44800 42920 44816 42984
rect 44880 42920 44896 42984
rect 44960 42920 44976 42984
rect 45040 42920 45056 42984
rect 45120 42920 45136 42984
rect 45200 42920 45216 42984
rect 45280 42920 45296 42984
rect 45360 42920 45368 42984
rect 0 42904 45368 42920
rect 0 42840 8 42904
rect 72 42840 88 42904
rect 152 42840 168 42904
rect 232 42840 248 42904
rect 312 42840 328 42904
rect 392 42840 408 42904
rect 472 42840 488 42904
rect 552 42840 568 42904
rect 632 42840 648 42904
rect 712 42840 728 42904
rect 792 42840 808 42904
rect 872 42840 888 42904
rect 952 42840 968 42904
rect 1032 42840 1048 42904
rect 1112 42840 1128 42904
rect 1192 42840 1208 42904
rect 1272 42840 1288 42904
rect 1352 42840 1368 42904
rect 1432 42840 1448 42904
rect 1512 42840 1528 42904
rect 1592 42840 1608 42904
rect 1672 42840 1688 42904
rect 1752 42840 1768 42904
rect 1832 42840 1848 42904
rect 1912 42840 1928 42904
rect 1992 42840 2008 42904
rect 2072 42840 2088 42904
rect 2152 42840 2168 42904
rect 2232 42840 2248 42904
rect 2312 42840 2328 42904
rect 2392 42840 2408 42904
rect 2472 42840 2488 42904
rect 2552 42840 2568 42904
rect 2632 42840 2648 42904
rect 2712 42840 2728 42904
rect 2792 42840 2808 42904
rect 2872 42840 2888 42904
rect 2952 42840 2968 42904
rect 3032 42840 3048 42904
rect 3112 42840 3128 42904
rect 3192 42840 3208 42904
rect 3272 42840 3288 42904
rect 3352 42840 3368 42904
rect 3432 42840 3448 42904
rect 3512 42840 3528 42904
rect 3592 42840 3608 42904
rect 3672 42840 3688 42904
rect 3752 42840 3768 42904
rect 3832 42840 3848 42904
rect 3912 42840 3928 42904
rect 3992 42840 19112 42904
rect 19176 42840 19192 42904
rect 19256 42840 19272 42904
rect 19336 42840 19352 42904
rect 19416 42840 29112 42904
rect 29176 42840 29192 42904
rect 29256 42840 29272 42904
rect 29336 42840 29352 42904
rect 29416 42840 41376 42904
rect 41440 42840 41456 42904
rect 41520 42840 41536 42904
rect 41600 42840 41616 42904
rect 41680 42840 41696 42904
rect 41760 42840 41776 42904
rect 41840 42840 41856 42904
rect 41920 42840 41936 42904
rect 42000 42840 42016 42904
rect 42080 42840 42096 42904
rect 42160 42840 42176 42904
rect 42240 42840 42256 42904
rect 42320 42840 42336 42904
rect 42400 42840 42416 42904
rect 42480 42840 42496 42904
rect 42560 42840 42576 42904
rect 42640 42840 42656 42904
rect 42720 42840 42736 42904
rect 42800 42840 42816 42904
rect 42880 42840 42896 42904
rect 42960 42840 42976 42904
rect 43040 42840 43056 42904
rect 43120 42840 43136 42904
rect 43200 42840 43216 42904
rect 43280 42840 43296 42904
rect 43360 42840 43376 42904
rect 43440 42840 43456 42904
rect 43520 42840 43536 42904
rect 43600 42840 43616 42904
rect 43680 42840 43696 42904
rect 43760 42840 43776 42904
rect 43840 42840 43856 42904
rect 43920 42840 43936 42904
rect 44000 42840 44016 42904
rect 44080 42840 44096 42904
rect 44160 42840 44176 42904
rect 44240 42840 44256 42904
rect 44320 42840 44336 42904
rect 44400 42840 44416 42904
rect 44480 42840 44496 42904
rect 44560 42840 44576 42904
rect 44640 42840 44656 42904
rect 44720 42840 44736 42904
rect 44800 42840 44816 42904
rect 44880 42840 44896 42904
rect 44960 42840 44976 42904
rect 45040 42840 45056 42904
rect 45120 42840 45136 42904
rect 45200 42840 45216 42904
rect 45280 42840 45296 42904
rect 45360 42840 45368 42904
rect 0 42824 45368 42840
rect 0 42760 8 42824
rect 72 42760 88 42824
rect 152 42760 168 42824
rect 232 42760 248 42824
rect 312 42760 328 42824
rect 392 42760 408 42824
rect 472 42760 488 42824
rect 552 42760 568 42824
rect 632 42760 648 42824
rect 712 42760 728 42824
rect 792 42760 808 42824
rect 872 42760 888 42824
rect 952 42760 968 42824
rect 1032 42760 1048 42824
rect 1112 42760 1128 42824
rect 1192 42760 1208 42824
rect 1272 42760 1288 42824
rect 1352 42760 1368 42824
rect 1432 42760 1448 42824
rect 1512 42760 1528 42824
rect 1592 42760 1608 42824
rect 1672 42760 1688 42824
rect 1752 42760 1768 42824
rect 1832 42760 1848 42824
rect 1912 42760 1928 42824
rect 1992 42760 2008 42824
rect 2072 42760 2088 42824
rect 2152 42760 2168 42824
rect 2232 42760 2248 42824
rect 2312 42760 2328 42824
rect 2392 42760 2408 42824
rect 2472 42760 2488 42824
rect 2552 42760 2568 42824
rect 2632 42760 2648 42824
rect 2712 42760 2728 42824
rect 2792 42760 2808 42824
rect 2872 42760 2888 42824
rect 2952 42760 2968 42824
rect 3032 42760 3048 42824
rect 3112 42760 3128 42824
rect 3192 42760 3208 42824
rect 3272 42760 3288 42824
rect 3352 42760 3368 42824
rect 3432 42760 3448 42824
rect 3512 42760 3528 42824
rect 3592 42760 3608 42824
rect 3672 42760 3688 42824
rect 3752 42760 3768 42824
rect 3832 42760 3848 42824
rect 3912 42760 3928 42824
rect 3992 42760 19112 42824
rect 19176 42760 19192 42824
rect 19256 42760 19272 42824
rect 19336 42760 19352 42824
rect 19416 42760 29112 42824
rect 29176 42760 29192 42824
rect 29256 42760 29272 42824
rect 29336 42760 29352 42824
rect 29416 42760 41376 42824
rect 41440 42760 41456 42824
rect 41520 42760 41536 42824
rect 41600 42760 41616 42824
rect 41680 42760 41696 42824
rect 41760 42760 41776 42824
rect 41840 42760 41856 42824
rect 41920 42760 41936 42824
rect 42000 42760 42016 42824
rect 42080 42760 42096 42824
rect 42160 42760 42176 42824
rect 42240 42760 42256 42824
rect 42320 42760 42336 42824
rect 42400 42760 42416 42824
rect 42480 42760 42496 42824
rect 42560 42760 42576 42824
rect 42640 42760 42656 42824
rect 42720 42760 42736 42824
rect 42800 42760 42816 42824
rect 42880 42760 42896 42824
rect 42960 42760 42976 42824
rect 43040 42760 43056 42824
rect 43120 42760 43136 42824
rect 43200 42760 43216 42824
rect 43280 42760 43296 42824
rect 43360 42760 43376 42824
rect 43440 42760 43456 42824
rect 43520 42760 43536 42824
rect 43600 42760 43616 42824
rect 43680 42760 43696 42824
rect 43760 42760 43776 42824
rect 43840 42760 43856 42824
rect 43920 42760 43936 42824
rect 44000 42760 44016 42824
rect 44080 42760 44096 42824
rect 44160 42760 44176 42824
rect 44240 42760 44256 42824
rect 44320 42760 44336 42824
rect 44400 42760 44416 42824
rect 44480 42760 44496 42824
rect 44560 42760 44576 42824
rect 44640 42760 44656 42824
rect 44720 42760 44736 42824
rect 44800 42760 44816 42824
rect 44880 42760 44896 42824
rect 44960 42760 44976 42824
rect 45040 42760 45056 42824
rect 45120 42760 45136 42824
rect 45200 42760 45216 42824
rect 45280 42760 45296 42824
rect 45360 42760 45368 42824
rect 0 42744 45368 42760
rect 0 42680 8 42744
rect 72 42680 88 42744
rect 152 42680 168 42744
rect 232 42680 248 42744
rect 312 42680 328 42744
rect 392 42680 408 42744
rect 472 42680 488 42744
rect 552 42680 568 42744
rect 632 42680 648 42744
rect 712 42680 728 42744
rect 792 42680 808 42744
rect 872 42680 888 42744
rect 952 42680 968 42744
rect 1032 42680 1048 42744
rect 1112 42680 1128 42744
rect 1192 42680 1208 42744
rect 1272 42680 1288 42744
rect 1352 42680 1368 42744
rect 1432 42680 1448 42744
rect 1512 42680 1528 42744
rect 1592 42680 1608 42744
rect 1672 42680 1688 42744
rect 1752 42680 1768 42744
rect 1832 42680 1848 42744
rect 1912 42680 1928 42744
rect 1992 42680 2008 42744
rect 2072 42680 2088 42744
rect 2152 42680 2168 42744
rect 2232 42680 2248 42744
rect 2312 42680 2328 42744
rect 2392 42680 2408 42744
rect 2472 42680 2488 42744
rect 2552 42680 2568 42744
rect 2632 42680 2648 42744
rect 2712 42680 2728 42744
rect 2792 42680 2808 42744
rect 2872 42680 2888 42744
rect 2952 42680 2968 42744
rect 3032 42680 3048 42744
rect 3112 42680 3128 42744
rect 3192 42680 3208 42744
rect 3272 42680 3288 42744
rect 3352 42680 3368 42744
rect 3432 42680 3448 42744
rect 3512 42680 3528 42744
rect 3592 42680 3608 42744
rect 3672 42680 3688 42744
rect 3752 42680 3768 42744
rect 3832 42680 3848 42744
rect 3912 42680 3928 42744
rect 3992 42680 19112 42744
rect 19176 42680 19192 42744
rect 19256 42680 19272 42744
rect 19336 42680 19352 42744
rect 19416 42680 29112 42744
rect 29176 42680 29192 42744
rect 29256 42680 29272 42744
rect 29336 42680 29352 42744
rect 29416 42680 41376 42744
rect 41440 42680 41456 42744
rect 41520 42680 41536 42744
rect 41600 42680 41616 42744
rect 41680 42680 41696 42744
rect 41760 42680 41776 42744
rect 41840 42680 41856 42744
rect 41920 42680 41936 42744
rect 42000 42680 42016 42744
rect 42080 42680 42096 42744
rect 42160 42680 42176 42744
rect 42240 42680 42256 42744
rect 42320 42680 42336 42744
rect 42400 42680 42416 42744
rect 42480 42680 42496 42744
rect 42560 42680 42576 42744
rect 42640 42680 42656 42744
rect 42720 42680 42736 42744
rect 42800 42680 42816 42744
rect 42880 42680 42896 42744
rect 42960 42680 42976 42744
rect 43040 42680 43056 42744
rect 43120 42680 43136 42744
rect 43200 42680 43216 42744
rect 43280 42680 43296 42744
rect 43360 42680 43376 42744
rect 43440 42680 43456 42744
rect 43520 42680 43536 42744
rect 43600 42680 43616 42744
rect 43680 42680 43696 42744
rect 43760 42680 43776 42744
rect 43840 42680 43856 42744
rect 43920 42680 43936 42744
rect 44000 42680 44016 42744
rect 44080 42680 44096 42744
rect 44160 42680 44176 42744
rect 44240 42680 44256 42744
rect 44320 42680 44336 42744
rect 44400 42680 44416 42744
rect 44480 42680 44496 42744
rect 44560 42680 44576 42744
rect 44640 42680 44656 42744
rect 44720 42680 44736 42744
rect 44800 42680 44816 42744
rect 44880 42680 44896 42744
rect 44960 42680 44976 42744
rect 45040 42680 45056 42744
rect 45120 42680 45136 42744
rect 45200 42680 45216 42744
rect 45280 42680 45296 42744
rect 45360 42680 45368 42744
rect 0 42664 45368 42680
rect 0 42600 8 42664
rect 72 42600 88 42664
rect 152 42600 168 42664
rect 232 42600 248 42664
rect 312 42600 328 42664
rect 392 42600 408 42664
rect 472 42600 488 42664
rect 552 42600 568 42664
rect 632 42600 648 42664
rect 712 42600 728 42664
rect 792 42600 808 42664
rect 872 42600 888 42664
rect 952 42600 968 42664
rect 1032 42600 1048 42664
rect 1112 42600 1128 42664
rect 1192 42600 1208 42664
rect 1272 42600 1288 42664
rect 1352 42600 1368 42664
rect 1432 42600 1448 42664
rect 1512 42600 1528 42664
rect 1592 42600 1608 42664
rect 1672 42600 1688 42664
rect 1752 42600 1768 42664
rect 1832 42600 1848 42664
rect 1912 42600 1928 42664
rect 1992 42600 2008 42664
rect 2072 42600 2088 42664
rect 2152 42600 2168 42664
rect 2232 42600 2248 42664
rect 2312 42600 2328 42664
rect 2392 42600 2408 42664
rect 2472 42600 2488 42664
rect 2552 42600 2568 42664
rect 2632 42600 2648 42664
rect 2712 42600 2728 42664
rect 2792 42600 2808 42664
rect 2872 42600 2888 42664
rect 2952 42600 2968 42664
rect 3032 42600 3048 42664
rect 3112 42600 3128 42664
rect 3192 42600 3208 42664
rect 3272 42600 3288 42664
rect 3352 42600 3368 42664
rect 3432 42600 3448 42664
rect 3512 42600 3528 42664
rect 3592 42600 3608 42664
rect 3672 42600 3688 42664
rect 3752 42600 3768 42664
rect 3832 42600 3848 42664
rect 3912 42600 3928 42664
rect 3992 42600 19112 42664
rect 19176 42600 19192 42664
rect 19256 42600 19272 42664
rect 19336 42600 19352 42664
rect 19416 42600 29112 42664
rect 29176 42600 29192 42664
rect 29256 42600 29272 42664
rect 29336 42600 29352 42664
rect 29416 42600 41376 42664
rect 41440 42600 41456 42664
rect 41520 42600 41536 42664
rect 41600 42600 41616 42664
rect 41680 42600 41696 42664
rect 41760 42600 41776 42664
rect 41840 42600 41856 42664
rect 41920 42600 41936 42664
rect 42000 42600 42016 42664
rect 42080 42600 42096 42664
rect 42160 42600 42176 42664
rect 42240 42600 42256 42664
rect 42320 42600 42336 42664
rect 42400 42600 42416 42664
rect 42480 42600 42496 42664
rect 42560 42600 42576 42664
rect 42640 42600 42656 42664
rect 42720 42600 42736 42664
rect 42800 42600 42816 42664
rect 42880 42600 42896 42664
rect 42960 42600 42976 42664
rect 43040 42600 43056 42664
rect 43120 42600 43136 42664
rect 43200 42600 43216 42664
rect 43280 42600 43296 42664
rect 43360 42600 43376 42664
rect 43440 42600 43456 42664
rect 43520 42600 43536 42664
rect 43600 42600 43616 42664
rect 43680 42600 43696 42664
rect 43760 42600 43776 42664
rect 43840 42600 43856 42664
rect 43920 42600 43936 42664
rect 44000 42600 44016 42664
rect 44080 42600 44096 42664
rect 44160 42600 44176 42664
rect 44240 42600 44256 42664
rect 44320 42600 44336 42664
rect 44400 42600 44416 42664
rect 44480 42600 44496 42664
rect 44560 42600 44576 42664
rect 44640 42600 44656 42664
rect 44720 42600 44736 42664
rect 44800 42600 44816 42664
rect 44880 42600 44896 42664
rect 44960 42600 44976 42664
rect 45040 42600 45056 42664
rect 45120 42600 45136 42664
rect 45200 42600 45216 42664
rect 45280 42600 45296 42664
rect 45360 42600 45368 42664
rect 0 42584 45368 42600
rect 0 42520 8 42584
rect 72 42520 88 42584
rect 152 42520 168 42584
rect 232 42520 248 42584
rect 312 42520 328 42584
rect 392 42520 408 42584
rect 472 42520 488 42584
rect 552 42520 568 42584
rect 632 42520 648 42584
rect 712 42520 728 42584
rect 792 42520 808 42584
rect 872 42520 888 42584
rect 952 42520 968 42584
rect 1032 42520 1048 42584
rect 1112 42520 1128 42584
rect 1192 42520 1208 42584
rect 1272 42520 1288 42584
rect 1352 42520 1368 42584
rect 1432 42520 1448 42584
rect 1512 42520 1528 42584
rect 1592 42520 1608 42584
rect 1672 42520 1688 42584
rect 1752 42520 1768 42584
rect 1832 42520 1848 42584
rect 1912 42520 1928 42584
rect 1992 42520 2008 42584
rect 2072 42520 2088 42584
rect 2152 42520 2168 42584
rect 2232 42520 2248 42584
rect 2312 42520 2328 42584
rect 2392 42520 2408 42584
rect 2472 42520 2488 42584
rect 2552 42520 2568 42584
rect 2632 42520 2648 42584
rect 2712 42520 2728 42584
rect 2792 42520 2808 42584
rect 2872 42520 2888 42584
rect 2952 42520 2968 42584
rect 3032 42520 3048 42584
rect 3112 42520 3128 42584
rect 3192 42520 3208 42584
rect 3272 42520 3288 42584
rect 3352 42520 3368 42584
rect 3432 42520 3448 42584
rect 3512 42520 3528 42584
rect 3592 42520 3608 42584
rect 3672 42520 3688 42584
rect 3752 42520 3768 42584
rect 3832 42520 3848 42584
rect 3912 42520 3928 42584
rect 3992 42520 19112 42584
rect 19176 42520 19192 42584
rect 19256 42520 19272 42584
rect 19336 42520 19352 42584
rect 19416 42520 29112 42584
rect 29176 42520 29192 42584
rect 29256 42520 29272 42584
rect 29336 42520 29352 42584
rect 29416 42520 41376 42584
rect 41440 42520 41456 42584
rect 41520 42520 41536 42584
rect 41600 42520 41616 42584
rect 41680 42520 41696 42584
rect 41760 42520 41776 42584
rect 41840 42520 41856 42584
rect 41920 42520 41936 42584
rect 42000 42520 42016 42584
rect 42080 42520 42096 42584
rect 42160 42520 42176 42584
rect 42240 42520 42256 42584
rect 42320 42520 42336 42584
rect 42400 42520 42416 42584
rect 42480 42520 42496 42584
rect 42560 42520 42576 42584
rect 42640 42520 42656 42584
rect 42720 42520 42736 42584
rect 42800 42520 42816 42584
rect 42880 42520 42896 42584
rect 42960 42520 42976 42584
rect 43040 42520 43056 42584
rect 43120 42520 43136 42584
rect 43200 42520 43216 42584
rect 43280 42520 43296 42584
rect 43360 42520 43376 42584
rect 43440 42520 43456 42584
rect 43520 42520 43536 42584
rect 43600 42520 43616 42584
rect 43680 42520 43696 42584
rect 43760 42520 43776 42584
rect 43840 42520 43856 42584
rect 43920 42520 43936 42584
rect 44000 42520 44016 42584
rect 44080 42520 44096 42584
rect 44160 42520 44176 42584
rect 44240 42520 44256 42584
rect 44320 42520 44336 42584
rect 44400 42520 44416 42584
rect 44480 42520 44496 42584
rect 44560 42520 44576 42584
rect 44640 42520 44656 42584
rect 44720 42520 44736 42584
rect 44800 42520 44816 42584
rect 44880 42520 44896 42584
rect 44960 42520 44976 42584
rect 45040 42520 45056 42584
rect 45120 42520 45136 42584
rect 45200 42520 45216 42584
rect 45280 42520 45296 42584
rect 45360 42520 45368 42584
rect 0 42504 45368 42520
rect 0 42440 8 42504
rect 72 42440 88 42504
rect 152 42440 168 42504
rect 232 42440 248 42504
rect 312 42440 328 42504
rect 392 42440 408 42504
rect 472 42440 488 42504
rect 552 42440 568 42504
rect 632 42440 648 42504
rect 712 42440 728 42504
rect 792 42440 808 42504
rect 872 42440 888 42504
rect 952 42440 968 42504
rect 1032 42440 1048 42504
rect 1112 42440 1128 42504
rect 1192 42440 1208 42504
rect 1272 42440 1288 42504
rect 1352 42440 1368 42504
rect 1432 42440 1448 42504
rect 1512 42440 1528 42504
rect 1592 42440 1608 42504
rect 1672 42440 1688 42504
rect 1752 42440 1768 42504
rect 1832 42440 1848 42504
rect 1912 42440 1928 42504
rect 1992 42440 2008 42504
rect 2072 42440 2088 42504
rect 2152 42440 2168 42504
rect 2232 42440 2248 42504
rect 2312 42440 2328 42504
rect 2392 42440 2408 42504
rect 2472 42440 2488 42504
rect 2552 42440 2568 42504
rect 2632 42440 2648 42504
rect 2712 42440 2728 42504
rect 2792 42440 2808 42504
rect 2872 42440 2888 42504
rect 2952 42440 2968 42504
rect 3032 42440 3048 42504
rect 3112 42440 3128 42504
rect 3192 42440 3208 42504
rect 3272 42440 3288 42504
rect 3352 42440 3368 42504
rect 3432 42440 3448 42504
rect 3512 42440 3528 42504
rect 3592 42440 3608 42504
rect 3672 42440 3688 42504
rect 3752 42440 3768 42504
rect 3832 42440 3848 42504
rect 3912 42440 3928 42504
rect 3992 42440 19112 42504
rect 19176 42440 19192 42504
rect 19256 42440 19272 42504
rect 19336 42440 19352 42504
rect 19416 42440 29112 42504
rect 29176 42440 29192 42504
rect 29256 42440 29272 42504
rect 29336 42440 29352 42504
rect 29416 42440 41376 42504
rect 41440 42440 41456 42504
rect 41520 42440 41536 42504
rect 41600 42440 41616 42504
rect 41680 42440 41696 42504
rect 41760 42440 41776 42504
rect 41840 42440 41856 42504
rect 41920 42440 41936 42504
rect 42000 42440 42016 42504
rect 42080 42440 42096 42504
rect 42160 42440 42176 42504
rect 42240 42440 42256 42504
rect 42320 42440 42336 42504
rect 42400 42440 42416 42504
rect 42480 42440 42496 42504
rect 42560 42440 42576 42504
rect 42640 42440 42656 42504
rect 42720 42440 42736 42504
rect 42800 42440 42816 42504
rect 42880 42440 42896 42504
rect 42960 42440 42976 42504
rect 43040 42440 43056 42504
rect 43120 42440 43136 42504
rect 43200 42440 43216 42504
rect 43280 42440 43296 42504
rect 43360 42440 43376 42504
rect 43440 42440 43456 42504
rect 43520 42440 43536 42504
rect 43600 42440 43616 42504
rect 43680 42440 43696 42504
rect 43760 42440 43776 42504
rect 43840 42440 43856 42504
rect 43920 42440 43936 42504
rect 44000 42440 44016 42504
rect 44080 42440 44096 42504
rect 44160 42440 44176 42504
rect 44240 42440 44256 42504
rect 44320 42440 44336 42504
rect 44400 42440 44416 42504
rect 44480 42440 44496 42504
rect 44560 42440 44576 42504
rect 44640 42440 44656 42504
rect 44720 42440 44736 42504
rect 44800 42440 44816 42504
rect 44880 42440 44896 42504
rect 44960 42440 44976 42504
rect 45040 42440 45056 42504
rect 45120 42440 45136 42504
rect 45200 42440 45216 42504
rect 45280 42440 45296 42504
rect 45360 42440 45368 42504
rect 0 42424 45368 42440
rect 0 42360 8 42424
rect 72 42360 88 42424
rect 152 42360 168 42424
rect 232 42360 248 42424
rect 312 42360 328 42424
rect 392 42360 408 42424
rect 472 42360 488 42424
rect 552 42360 568 42424
rect 632 42360 648 42424
rect 712 42360 728 42424
rect 792 42360 808 42424
rect 872 42360 888 42424
rect 952 42360 968 42424
rect 1032 42360 1048 42424
rect 1112 42360 1128 42424
rect 1192 42360 1208 42424
rect 1272 42360 1288 42424
rect 1352 42360 1368 42424
rect 1432 42360 1448 42424
rect 1512 42360 1528 42424
rect 1592 42360 1608 42424
rect 1672 42360 1688 42424
rect 1752 42360 1768 42424
rect 1832 42360 1848 42424
rect 1912 42360 1928 42424
rect 1992 42360 2008 42424
rect 2072 42360 2088 42424
rect 2152 42360 2168 42424
rect 2232 42360 2248 42424
rect 2312 42360 2328 42424
rect 2392 42360 2408 42424
rect 2472 42360 2488 42424
rect 2552 42360 2568 42424
rect 2632 42360 2648 42424
rect 2712 42360 2728 42424
rect 2792 42360 2808 42424
rect 2872 42360 2888 42424
rect 2952 42360 2968 42424
rect 3032 42360 3048 42424
rect 3112 42360 3128 42424
rect 3192 42360 3208 42424
rect 3272 42360 3288 42424
rect 3352 42360 3368 42424
rect 3432 42360 3448 42424
rect 3512 42360 3528 42424
rect 3592 42360 3608 42424
rect 3672 42360 3688 42424
rect 3752 42360 3768 42424
rect 3832 42360 3848 42424
rect 3912 42360 3928 42424
rect 3992 42360 19112 42424
rect 19176 42360 19192 42424
rect 19256 42360 19272 42424
rect 19336 42360 19352 42424
rect 19416 42360 29112 42424
rect 29176 42360 29192 42424
rect 29256 42360 29272 42424
rect 29336 42360 29352 42424
rect 29416 42360 41376 42424
rect 41440 42360 41456 42424
rect 41520 42360 41536 42424
rect 41600 42360 41616 42424
rect 41680 42360 41696 42424
rect 41760 42360 41776 42424
rect 41840 42360 41856 42424
rect 41920 42360 41936 42424
rect 42000 42360 42016 42424
rect 42080 42360 42096 42424
rect 42160 42360 42176 42424
rect 42240 42360 42256 42424
rect 42320 42360 42336 42424
rect 42400 42360 42416 42424
rect 42480 42360 42496 42424
rect 42560 42360 42576 42424
rect 42640 42360 42656 42424
rect 42720 42360 42736 42424
rect 42800 42360 42816 42424
rect 42880 42360 42896 42424
rect 42960 42360 42976 42424
rect 43040 42360 43056 42424
rect 43120 42360 43136 42424
rect 43200 42360 43216 42424
rect 43280 42360 43296 42424
rect 43360 42360 43376 42424
rect 43440 42360 43456 42424
rect 43520 42360 43536 42424
rect 43600 42360 43616 42424
rect 43680 42360 43696 42424
rect 43760 42360 43776 42424
rect 43840 42360 43856 42424
rect 43920 42360 43936 42424
rect 44000 42360 44016 42424
rect 44080 42360 44096 42424
rect 44160 42360 44176 42424
rect 44240 42360 44256 42424
rect 44320 42360 44336 42424
rect 44400 42360 44416 42424
rect 44480 42360 44496 42424
rect 44560 42360 44576 42424
rect 44640 42360 44656 42424
rect 44720 42360 44736 42424
rect 44800 42360 44816 42424
rect 44880 42360 44896 42424
rect 44960 42360 44976 42424
rect 45040 42360 45056 42424
rect 45120 42360 45136 42424
rect 45200 42360 45216 42424
rect 45280 42360 45296 42424
rect 45360 42360 45368 42424
rect 0 42344 45368 42360
rect 0 42280 8 42344
rect 72 42280 88 42344
rect 152 42280 168 42344
rect 232 42280 248 42344
rect 312 42280 328 42344
rect 392 42280 408 42344
rect 472 42280 488 42344
rect 552 42280 568 42344
rect 632 42280 648 42344
rect 712 42280 728 42344
rect 792 42280 808 42344
rect 872 42280 888 42344
rect 952 42280 968 42344
rect 1032 42280 1048 42344
rect 1112 42280 1128 42344
rect 1192 42280 1208 42344
rect 1272 42280 1288 42344
rect 1352 42280 1368 42344
rect 1432 42280 1448 42344
rect 1512 42280 1528 42344
rect 1592 42280 1608 42344
rect 1672 42280 1688 42344
rect 1752 42280 1768 42344
rect 1832 42280 1848 42344
rect 1912 42280 1928 42344
rect 1992 42280 2008 42344
rect 2072 42280 2088 42344
rect 2152 42280 2168 42344
rect 2232 42280 2248 42344
rect 2312 42280 2328 42344
rect 2392 42280 2408 42344
rect 2472 42280 2488 42344
rect 2552 42280 2568 42344
rect 2632 42280 2648 42344
rect 2712 42280 2728 42344
rect 2792 42280 2808 42344
rect 2872 42280 2888 42344
rect 2952 42280 2968 42344
rect 3032 42280 3048 42344
rect 3112 42280 3128 42344
rect 3192 42280 3208 42344
rect 3272 42280 3288 42344
rect 3352 42280 3368 42344
rect 3432 42280 3448 42344
rect 3512 42280 3528 42344
rect 3592 42280 3608 42344
rect 3672 42280 3688 42344
rect 3752 42280 3768 42344
rect 3832 42280 3848 42344
rect 3912 42280 3928 42344
rect 3992 42280 19112 42344
rect 19176 42280 19192 42344
rect 19256 42280 19272 42344
rect 19336 42280 19352 42344
rect 19416 42280 29112 42344
rect 29176 42280 29192 42344
rect 29256 42280 29272 42344
rect 29336 42280 29352 42344
rect 29416 42280 41376 42344
rect 41440 42280 41456 42344
rect 41520 42280 41536 42344
rect 41600 42280 41616 42344
rect 41680 42280 41696 42344
rect 41760 42280 41776 42344
rect 41840 42280 41856 42344
rect 41920 42280 41936 42344
rect 42000 42280 42016 42344
rect 42080 42280 42096 42344
rect 42160 42280 42176 42344
rect 42240 42280 42256 42344
rect 42320 42280 42336 42344
rect 42400 42280 42416 42344
rect 42480 42280 42496 42344
rect 42560 42280 42576 42344
rect 42640 42280 42656 42344
rect 42720 42280 42736 42344
rect 42800 42280 42816 42344
rect 42880 42280 42896 42344
rect 42960 42280 42976 42344
rect 43040 42280 43056 42344
rect 43120 42280 43136 42344
rect 43200 42280 43216 42344
rect 43280 42280 43296 42344
rect 43360 42280 43376 42344
rect 43440 42280 43456 42344
rect 43520 42280 43536 42344
rect 43600 42280 43616 42344
rect 43680 42280 43696 42344
rect 43760 42280 43776 42344
rect 43840 42280 43856 42344
rect 43920 42280 43936 42344
rect 44000 42280 44016 42344
rect 44080 42280 44096 42344
rect 44160 42280 44176 42344
rect 44240 42280 44256 42344
rect 44320 42280 44336 42344
rect 44400 42280 44416 42344
rect 44480 42280 44496 42344
rect 44560 42280 44576 42344
rect 44640 42280 44656 42344
rect 44720 42280 44736 42344
rect 44800 42280 44816 42344
rect 44880 42280 44896 42344
rect 44960 42280 44976 42344
rect 45040 42280 45056 42344
rect 45120 42280 45136 42344
rect 45200 42280 45216 42344
rect 45280 42280 45296 42344
rect 45360 42280 45368 42344
rect 0 42264 45368 42280
rect 0 42200 8 42264
rect 72 42200 88 42264
rect 152 42200 168 42264
rect 232 42200 248 42264
rect 312 42200 328 42264
rect 392 42200 408 42264
rect 472 42200 488 42264
rect 552 42200 568 42264
rect 632 42200 648 42264
rect 712 42200 728 42264
rect 792 42200 808 42264
rect 872 42200 888 42264
rect 952 42200 968 42264
rect 1032 42200 1048 42264
rect 1112 42200 1128 42264
rect 1192 42200 1208 42264
rect 1272 42200 1288 42264
rect 1352 42200 1368 42264
rect 1432 42200 1448 42264
rect 1512 42200 1528 42264
rect 1592 42200 1608 42264
rect 1672 42200 1688 42264
rect 1752 42200 1768 42264
rect 1832 42200 1848 42264
rect 1912 42200 1928 42264
rect 1992 42200 2008 42264
rect 2072 42200 2088 42264
rect 2152 42200 2168 42264
rect 2232 42200 2248 42264
rect 2312 42200 2328 42264
rect 2392 42200 2408 42264
rect 2472 42200 2488 42264
rect 2552 42200 2568 42264
rect 2632 42200 2648 42264
rect 2712 42200 2728 42264
rect 2792 42200 2808 42264
rect 2872 42200 2888 42264
rect 2952 42200 2968 42264
rect 3032 42200 3048 42264
rect 3112 42200 3128 42264
rect 3192 42200 3208 42264
rect 3272 42200 3288 42264
rect 3352 42200 3368 42264
rect 3432 42200 3448 42264
rect 3512 42200 3528 42264
rect 3592 42200 3608 42264
rect 3672 42200 3688 42264
rect 3752 42200 3768 42264
rect 3832 42200 3848 42264
rect 3912 42200 3928 42264
rect 3992 42200 19112 42264
rect 19176 42200 19192 42264
rect 19256 42200 19272 42264
rect 19336 42200 19352 42264
rect 19416 42200 29112 42264
rect 29176 42200 29192 42264
rect 29256 42200 29272 42264
rect 29336 42200 29352 42264
rect 29416 42200 41376 42264
rect 41440 42200 41456 42264
rect 41520 42200 41536 42264
rect 41600 42200 41616 42264
rect 41680 42200 41696 42264
rect 41760 42200 41776 42264
rect 41840 42200 41856 42264
rect 41920 42200 41936 42264
rect 42000 42200 42016 42264
rect 42080 42200 42096 42264
rect 42160 42200 42176 42264
rect 42240 42200 42256 42264
rect 42320 42200 42336 42264
rect 42400 42200 42416 42264
rect 42480 42200 42496 42264
rect 42560 42200 42576 42264
rect 42640 42200 42656 42264
rect 42720 42200 42736 42264
rect 42800 42200 42816 42264
rect 42880 42200 42896 42264
rect 42960 42200 42976 42264
rect 43040 42200 43056 42264
rect 43120 42200 43136 42264
rect 43200 42200 43216 42264
rect 43280 42200 43296 42264
rect 43360 42200 43376 42264
rect 43440 42200 43456 42264
rect 43520 42200 43536 42264
rect 43600 42200 43616 42264
rect 43680 42200 43696 42264
rect 43760 42200 43776 42264
rect 43840 42200 43856 42264
rect 43920 42200 43936 42264
rect 44000 42200 44016 42264
rect 44080 42200 44096 42264
rect 44160 42200 44176 42264
rect 44240 42200 44256 42264
rect 44320 42200 44336 42264
rect 44400 42200 44416 42264
rect 44480 42200 44496 42264
rect 44560 42200 44576 42264
rect 44640 42200 44656 42264
rect 44720 42200 44736 42264
rect 44800 42200 44816 42264
rect 44880 42200 44896 42264
rect 44960 42200 44976 42264
rect 45040 42200 45056 42264
rect 45120 42200 45136 42264
rect 45200 42200 45216 42264
rect 45280 42200 45296 42264
rect 45360 42200 45368 42264
rect 0 42184 45368 42200
rect 0 42120 8 42184
rect 72 42120 88 42184
rect 152 42120 168 42184
rect 232 42120 248 42184
rect 312 42120 328 42184
rect 392 42120 408 42184
rect 472 42120 488 42184
rect 552 42120 568 42184
rect 632 42120 648 42184
rect 712 42120 728 42184
rect 792 42120 808 42184
rect 872 42120 888 42184
rect 952 42120 968 42184
rect 1032 42120 1048 42184
rect 1112 42120 1128 42184
rect 1192 42120 1208 42184
rect 1272 42120 1288 42184
rect 1352 42120 1368 42184
rect 1432 42120 1448 42184
rect 1512 42120 1528 42184
rect 1592 42120 1608 42184
rect 1672 42120 1688 42184
rect 1752 42120 1768 42184
rect 1832 42120 1848 42184
rect 1912 42120 1928 42184
rect 1992 42120 2008 42184
rect 2072 42120 2088 42184
rect 2152 42120 2168 42184
rect 2232 42120 2248 42184
rect 2312 42120 2328 42184
rect 2392 42120 2408 42184
rect 2472 42120 2488 42184
rect 2552 42120 2568 42184
rect 2632 42120 2648 42184
rect 2712 42120 2728 42184
rect 2792 42120 2808 42184
rect 2872 42120 2888 42184
rect 2952 42120 2968 42184
rect 3032 42120 3048 42184
rect 3112 42120 3128 42184
rect 3192 42120 3208 42184
rect 3272 42120 3288 42184
rect 3352 42120 3368 42184
rect 3432 42120 3448 42184
rect 3512 42120 3528 42184
rect 3592 42120 3608 42184
rect 3672 42120 3688 42184
rect 3752 42120 3768 42184
rect 3832 42120 3848 42184
rect 3912 42120 3928 42184
rect 3992 42120 19112 42184
rect 19176 42120 19192 42184
rect 19256 42120 19272 42184
rect 19336 42120 19352 42184
rect 19416 42120 29112 42184
rect 29176 42120 29192 42184
rect 29256 42120 29272 42184
rect 29336 42120 29352 42184
rect 29416 42120 41376 42184
rect 41440 42120 41456 42184
rect 41520 42120 41536 42184
rect 41600 42120 41616 42184
rect 41680 42120 41696 42184
rect 41760 42120 41776 42184
rect 41840 42120 41856 42184
rect 41920 42120 41936 42184
rect 42000 42120 42016 42184
rect 42080 42120 42096 42184
rect 42160 42120 42176 42184
rect 42240 42120 42256 42184
rect 42320 42120 42336 42184
rect 42400 42120 42416 42184
rect 42480 42120 42496 42184
rect 42560 42120 42576 42184
rect 42640 42120 42656 42184
rect 42720 42120 42736 42184
rect 42800 42120 42816 42184
rect 42880 42120 42896 42184
rect 42960 42120 42976 42184
rect 43040 42120 43056 42184
rect 43120 42120 43136 42184
rect 43200 42120 43216 42184
rect 43280 42120 43296 42184
rect 43360 42120 43376 42184
rect 43440 42120 43456 42184
rect 43520 42120 43536 42184
rect 43600 42120 43616 42184
rect 43680 42120 43696 42184
rect 43760 42120 43776 42184
rect 43840 42120 43856 42184
rect 43920 42120 43936 42184
rect 44000 42120 44016 42184
rect 44080 42120 44096 42184
rect 44160 42120 44176 42184
rect 44240 42120 44256 42184
rect 44320 42120 44336 42184
rect 44400 42120 44416 42184
rect 44480 42120 44496 42184
rect 44560 42120 44576 42184
rect 44640 42120 44656 42184
rect 44720 42120 44736 42184
rect 44800 42120 44816 42184
rect 44880 42120 44896 42184
rect 44960 42120 44976 42184
rect 45040 42120 45056 42184
rect 45120 42120 45136 42184
rect 45200 42120 45216 42184
rect 45280 42120 45296 42184
rect 45360 42120 45368 42184
rect 0 42104 45368 42120
rect 0 42040 8 42104
rect 72 42040 88 42104
rect 152 42040 168 42104
rect 232 42040 248 42104
rect 312 42040 328 42104
rect 392 42040 408 42104
rect 472 42040 488 42104
rect 552 42040 568 42104
rect 632 42040 648 42104
rect 712 42040 728 42104
rect 792 42040 808 42104
rect 872 42040 888 42104
rect 952 42040 968 42104
rect 1032 42040 1048 42104
rect 1112 42040 1128 42104
rect 1192 42040 1208 42104
rect 1272 42040 1288 42104
rect 1352 42040 1368 42104
rect 1432 42040 1448 42104
rect 1512 42040 1528 42104
rect 1592 42040 1608 42104
rect 1672 42040 1688 42104
rect 1752 42040 1768 42104
rect 1832 42040 1848 42104
rect 1912 42040 1928 42104
rect 1992 42040 2008 42104
rect 2072 42040 2088 42104
rect 2152 42040 2168 42104
rect 2232 42040 2248 42104
rect 2312 42040 2328 42104
rect 2392 42040 2408 42104
rect 2472 42040 2488 42104
rect 2552 42040 2568 42104
rect 2632 42040 2648 42104
rect 2712 42040 2728 42104
rect 2792 42040 2808 42104
rect 2872 42040 2888 42104
rect 2952 42040 2968 42104
rect 3032 42040 3048 42104
rect 3112 42040 3128 42104
rect 3192 42040 3208 42104
rect 3272 42040 3288 42104
rect 3352 42040 3368 42104
rect 3432 42040 3448 42104
rect 3512 42040 3528 42104
rect 3592 42040 3608 42104
rect 3672 42040 3688 42104
rect 3752 42040 3768 42104
rect 3832 42040 3848 42104
rect 3912 42040 3928 42104
rect 3992 42040 19112 42104
rect 19176 42040 19192 42104
rect 19256 42040 19272 42104
rect 19336 42040 19352 42104
rect 19416 42040 29112 42104
rect 29176 42040 29192 42104
rect 29256 42040 29272 42104
rect 29336 42040 29352 42104
rect 29416 42040 41376 42104
rect 41440 42040 41456 42104
rect 41520 42040 41536 42104
rect 41600 42040 41616 42104
rect 41680 42040 41696 42104
rect 41760 42040 41776 42104
rect 41840 42040 41856 42104
rect 41920 42040 41936 42104
rect 42000 42040 42016 42104
rect 42080 42040 42096 42104
rect 42160 42040 42176 42104
rect 42240 42040 42256 42104
rect 42320 42040 42336 42104
rect 42400 42040 42416 42104
rect 42480 42040 42496 42104
rect 42560 42040 42576 42104
rect 42640 42040 42656 42104
rect 42720 42040 42736 42104
rect 42800 42040 42816 42104
rect 42880 42040 42896 42104
rect 42960 42040 42976 42104
rect 43040 42040 43056 42104
rect 43120 42040 43136 42104
rect 43200 42040 43216 42104
rect 43280 42040 43296 42104
rect 43360 42040 43376 42104
rect 43440 42040 43456 42104
rect 43520 42040 43536 42104
rect 43600 42040 43616 42104
rect 43680 42040 43696 42104
rect 43760 42040 43776 42104
rect 43840 42040 43856 42104
rect 43920 42040 43936 42104
rect 44000 42040 44016 42104
rect 44080 42040 44096 42104
rect 44160 42040 44176 42104
rect 44240 42040 44256 42104
rect 44320 42040 44336 42104
rect 44400 42040 44416 42104
rect 44480 42040 44496 42104
rect 44560 42040 44576 42104
rect 44640 42040 44656 42104
rect 44720 42040 44736 42104
rect 44800 42040 44816 42104
rect 44880 42040 44896 42104
rect 44960 42040 44976 42104
rect 45040 42040 45056 42104
rect 45120 42040 45136 42104
rect 45200 42040 45216 42104
rect 45280 42040 45296 42104
rect 45360 42040 45368 42104
rect 0 42024 45368 42040
rect 0 41960 8 42024
rect 72 41960 88 42024
rect 152 41960 168 42024
rect 232 41960 248 42024
rect 312 41960 328 42024
rect 392 41960 408 42024
rect 472 41960 488 42024
rect 552 41960 568 42024
rect 632 41960 648 42024
rect 712 41960 728 42024
rect 792 41960 808 42024
rect 872 41960 888 42024
rect 952 41960 968 42024
rect 1032 41960 1048 42024
rect 1112 41960 1128 42024
rect 1192 41960 1208 42024
rect 1272 41960 1288 42024
rect 1352 41960 1368 42024
rect 1432 41960 1448 42024
rect 1512 41960 1528 42024
rect 1592 41960 1608 42024
rect 1672 41960 1688 42024
rect 1752 41960 1768 42024
rect 1832 41960 1848 42024
rect 1912 41960 1928 42024
rect 1992 41960 2008 42024
rect 2072 41960 2088 42024
rect 2152 41960 2168 42024
rect 2232 41960 2248 42024
rect 2312 41960 2328 42024
rect 2392 41960 2408 42024
rect 2472 41960 2488 42024
rect 2552 41960 2568 42024
rect 2632 41960 2648 42024
rect 2712 41960 2728 42024
rect 2792 41960 2808 42024
rect 2872 41960 2888 42024
rect 2952 41960 2968 42024
rect 3032 41960 3048 42024
rect 3112 41960 3128 42024
rect 3192 41960 3208 42024
rect 3272 41960 3288 42024
rect 3352 41960 3368 42024
rect 3432 41960 3448 42024
rect 3512 41960 3528 42024
rect 3592 41960 3608 42024
rect 3672 41960 3688 42024
rect 3752 41960 3768 42024
rect 3832 41960 3848 42024
rect 3912 41960 3928 42024
rect 3992 41960 19112 42024
rect 19176 41960 19192 42024
rect 19256 41960 19272 42024
rect 19336 41960 19352 42024
rect 19416 41960 29112 42024
rect 29176 41960 29192 42024
rect 29256 41960 29272 42024
rect 29336 41960 29352 42024
rect 29416 41960 41376 42024
rect 41440 41960 41456 42024
rect 41520 41960 41536 42024
rect 41600 41960 41616 42024
rect 41680 41960 41696 42024
rect 41760 41960 41776 42024
rect 41840 41960 41856 42024
rect 41920 41960 41936 42024
rect 42000 41960 42016 42024
rect 42080 41960 42096 42024
rect 42160 41960 42176 42024
rect 42240 41960 42256 42024
rect 42320 41960 42336 42024
rect 42400 41960 42416 42024
rect 42480 41960 42496 42024
rect 42560 41960 42576 42024
rect 42640 41960 42656 42024
rect 42720 41960 42736 42024
rect 42800 41960 42816 42024
rect 42880 41960 42896 42024
rect 42960 41960 42976 42024
rect 43040 41960 43056 42024
rect 43120 41960 43136 42024
rect 43200 41960 43216 42024
rect 43280 41960 43296 42024
rect 43360 41960 43376 42024
rect 43440 41960 43456 42024
rect 43520 41960 43536 42024
rect 43600 41960 43616 42024
rect 43680 41960 43696 42024
rect 43760 41960 43776 42024
rect 43840 41960 43856 42024
rect 43920 41960 43936 42024
rect 44000 41960 44016 42024
rect 44080 41960 44096 42024
rect 44160 41960 44176 42024
rect 44240 41960 44256 42024
rect 44320 41960 44336 42024
rect 44400 41960 44416 42024
rect 44480 41960 44496 42024
rect 44560 41960 44576 42024
rect 44640 41960 44656 42024
rect 44720 41960 44736 42024
rect 44800 41960 44816 42024
rect 44880 41960 44896 42024
rect 44960 41960 44976 42024
rect 45040 41960 45056 42024
rect 45120 41960 45136 42024
rect 45200 41960 45216 42024
rect 45280 41960 45296 42024
rect 45360 41960 45368 42024
rect 0 41944 45368 41960
rect 0 41880 8 41944
rect 72 41880 88 41944
rect 152 41880 168 41944
rect 232 41880 248 41944
rect 312 41880 328 41944
rect 392 41880 408 41944
rect 472 41880 488 41944
rect 552 41880 568 41944
rect 632 41880 648 41944
rect 712 41880 728 41944
rect 792 41880 808 41944
rect 872 41880 888 41944
rect 952 41880 968 41944
rect 1032 41880 1048 41944
rect 1112 41880 1128 41944
rect 1192 41880 1208 41944
rect 1272 41880 1288 41944
rect 1352 41880 1368 41944
rect 1432 41880 1448 41944
rect 1512 41880 1528 41944
rect 1592 41880 1608 41944
rect 1672 41880 1688 41944
rect 1752 41880 1768 41944
rect 1832 41880 1848 41944
rect 1912 41880 1928 41944
rect 1992 41880 2008 41944
rect 2072 41880 2088 41944
rect 2152 41880 2168 41944
rect 2232 41880 2248 41944
rect 2312 41880 2328 41944
rect 2392 41880 2408 41944
rect 2472 41880 2488 41944
rect 2552 41880 2568 41944
rect 2632 41880 2648 41944
rect 2712 41880 2728 41944
rect 2792 41880 2808 41944
rect 2872 41880 2888 41944
rect 2952 41880 2968 41944
rect 3032 41880 3048 41944
rect 3112 41880 3128 41944
rect 3192 41880 3208 41944
rect 3272 41880 3288 41944
rect 3352 41880 3368 41944
rect 3432 41880 3448 41944
rect 3512 41880 3528 41944
rect 3592 41880 3608 41944
rect 3672 41880 3688 41944
rect 3752 41880 3768 41944
rect 3832 41880 3848 41944
rect 3912 41880 3928 41944
rect 3992 41880 19112 41944
rect 19176 41880 19192 41944
rect 19256 41880 19272 41944
rect 19336 41880 19352 41944
rect 19416 41880 29112 41944
rect 29176 41880 29192 41944
rect 29256 41880 29272 41944
rect 29336 41880 29352 41944
rect 29416 41880 41376 41944
rect 41440 41880 41456 41944
rect 41520 41880 41536 41944
rect 41600 41880 41616 41944
rect 41680 41880 41696 41944
rect 41760 41880 41776 41944
rect 41840 41880 41856 41944
rect 41920 41880 41936 41944
rect 42000 41880 42016 41944
rect 42080 41880 42096 41944
rect 42160 41880 42176 41944
rect 42240 41880 42256 41944
rect 42320 41880 42336 41944
rect 42400 41880 42416 41944
rect 42480 41880 42496 41944
rect 42560 41880 42576 41944
rect 42640 41880 42656 41944
rect 42720 41880 42736 41944
rect 42800 41880 42816 41944
rect 42880 41880 42896 41944
rect 42960 41880 42976 41944
rect 43040 41880 43056 41944
rect 43120 41880 43136 41944
rect 43200 41880 43216 41944
rect 43280 41880 43296 41944
rect 43360 41880 43376 41944
rect 43440 41880 43456 41944
rect 43520 41880 43536 41944
rect 43600 41880 43616 41944
rect 43680 41880 43696 41944
rect 43760 41880 43776 41944
rect 43840 41880 43856 41944
rect 43920 41880 43936 41944
rect 44000 41880 44016 41944
rect 44080 41880 44096 41944
rect 44160 41880 44176 41944
rect 44240 41880 44256 41944
rect 44320 41880 44336 41944
rect 44400 41880 44416 41944
rect 44480 41880 44496 41944
rect 44560 41880 44576 41944
rect 44640 41880 44656 41944
rect 44720 41880 44736 41944
rect 44800 41880 44816 41944
rect 44880 41880 44896 41944
rect 44960 41880 44976 41944
rect 45040 41880 45056 41944
rect 45120 41880 45136 41944
rect 45200 41880 45216 41944
rect 45280 41880 45296 41944
rect 45360 41880 45368 41944
rect 0 41864 45368 41880
rect 0 41800 8 41864
rect 72 41800 88 41864
rect 152 41800 168 41864
rect 232 41800 248 41864
rect 312 41800 328 41864
rect 392 41800 408 41864
rect 472 41800 488 41864
rect 552 41800 568 41864
rect 632 41800 648 41864
rect 712 41800 728 41864
rect 792 41800 808 41864
rect 872 41800 888 41864
rect 952 41800 968 41864
rect 1032 41800 1048 41864
rect 1112 41800 1128 41864
rect 1192 41800 1208 41864
rect 1272 41800 1288 41864
rect 1352 41800 1368 41864
rect 1432 41800 1448 41864
rect 1512 41800 1528 41864
rect 1592 41800 1608 41864
rect 1672 41800 1688 41864
rect 1752 41800 1768 41864
rect 1832 41800 1848 41864
rect 1912 41800 1928 41864
rect 1992 41800 2008 41864
rect 2072 41800 2088 41864
rect 2152 41800 2168 41864
rect 2232 41800 2248 41864
rect 2312 41800 2328 41864
rect 2392 41800 2408 41864
rect 2472 41800 2488 41864
rect 2552 41800 2568 41864
rect 2632 41800 2648 41864
rect 2712 41800 2728 41864
rect 2792 41800 2808 41864
rect 2872 41800 2888 41864
rect 2952 41800 2968 41864
rect 3032 41800 3048 41864
rect 3112 41800 3128 41864
rect 3192 41800 3208 41864
rect 3272 41800 3288 41864
rect 3352 41800 3368 41864
rect 3432 41800 3448 41864
rect 3512 41800 3528 41864
rect 3592 41800 3608 41864
rect 3672 41800 3688 41864
rect 3752 41800 3768 41864
rect 3832 41800 3848 41864
rect 3912 41800 3928 41864
rect 3992 41800 19112 41864
rect 19176 41800 19192 41864
rect 19256 41800 19272 41864
rect 19336 41800 19352 41864
rect 19416 41800 29112 41864
rect 29176 41800 29192 41864
rect 29256 41800 29272 41864
rect 29336 41800 29352 41864
rect 29416 41800 41376 41864
rect 41440 41800 41456 41864
rect 41520 41800 41536 41864
rect 41600 41800 41616 41864
rect 41680 41800 41696 41864
rect 41760 41800 41776 41864
rect 41840 41800 41856 41864
rect 41920 41800 41936 41864
rect 42000 41800 42016 41864
rect 42080 41800 42096 41864
rect 42160 41800 42176 41864
rect 42240 41800 42256 41864
rect 42320 41800 42336 41864
rect 42400 41800 42416 41864
rect 42480 41800 42496 41864
rect 42560 41800 42576 41864
rect 42640 41800 42656 41864
rect 42720 41800 42736 41864
rect 42800 41800 42816 41864
rect 42880 41800 42896 41864
rect 42960 41800 42976 41864
rect 43040 41800 43056 41864
rect 43120 41800 43136 41864
rect 43200 41800 43216 41864
rect 43280 41800 43296 41864
rect 43360 41800 43376 41864
rect 43440 41800 43456 41864
rect 43520 41800 43536 41864
rect 43600 41800 43616 41864
rect 43680 41800 43696 41864
rect 43760 41800 43776 41864
rect 43840 41800 43856 41864
rect 43920 41800 43936 41864
rect 44000 41800 44016 41864
rect 44080 41800 44096 41864
rect 44160 41800 44176 41864
rect 44240 41800 44256 41864
rect 44320 41800 44336 41864
rect 44400 41800 44416 41864
rect 44480 41800 44496 41864
rect 44560 41800 44576 41864
rect 44640 41800 44656 41864
rect 44720 41800 44736 41864
rect 44800 41800 44816 41864
rect 44880 41800 44896 41864
rect 44960 41800 44976 41864
rect 45040 41800 45056 41864
rect 45120 41800 45136 41864
rect 45200 41800 45216 41864
rect 45280 41800 45296 41864
rect 45360 41800 45368 41864
rect 0 41784 45368 41800
rect 0 41720 8 41784
rect 72 41720 88 41784
rect 152 41720 168 41784
rect 232 41720 248 41784
rect 312 41720 328 41784
rect 392 41720 408 41784
rect 472 41720 488 41784
rect 552 41720 568 41784
rect 632 41720 648 41784
rect 712 41720 728 41784
rect 792 41720 808 41784
rect 872 41720 888 41784
rect 952 41720 968 41784
rect 1032 41720 1048 41784
rect 1112 41720 1128 41784
rect 1192 41720 1208 41784
rect 1272 41720 1288 41784
rect 1352 41720 1368 41784
rect 1432 41720 1448 41784
rect 1512 41720 1528 41784
rect 1592 41720 1608 41784
rect 1672 41720 1688 41784
rect 1752 41720 1768 41784
rect 1832 41720 1848 41784
rect 1912 41720 1928 41784
rect 1992 41720 2008 41784
rect 2072 41720 2088 41784
rect 2152 41720 2168 41784
rect 2232 41720 2248 41784
rect 2312 41720 2328 41784
rect 2392 41720 2408 41784
rect 2472 41720 2488 41784
rect 2552 41720 2568 41784
rect 2632 41720 2648 41784
rect 2712 41720 2728 41784
rect 2792 41720 2808 41784
rect 2872 41720 2888 41784
rect 2952 41720 2968 41784
rect 3032 41720 3048 41784
rect 3112 41720 3128 41784
rect 3192 41720 3208 41784
rect 3272 41720 3288 41784
rect 3352 41720 3368 41784
rect 3432 41720 3448 41784
rect 3512 41720 3528 41784
rect 3592 41720 3608 41784
rect 3672 41720 3688 41784
rect 3752 41720 3768 41784
rect 3832 41720 3848 41784
rect 3912 41720 3928 41784
rect 3992 41720 19112 41784
rect 19176 41720 19192 41784
rect 19256 41720 19272 41784
rect 19336 41720 19352 41784
rect 19416 41720 29112 41784
rect 29176 41720 29192 41784
rect 29256 41720 29272 41784
rect 29336 41720 29352 41784
rect 29416 41720 41376 41784
rect 41440 41720 41456 41784
rect 41520 41720 41536 41784
rect 41600 41720 41616 41784
rect 41680 41720 41696 41784
rect 41760 41720 41776 41784
rect 41840 41720 41856 41784
rect 41920 41720 41936 41784
rect 42000 41720 42016 41784
rect 42080 41720 42096 41784
rect 42160 41720 42176 41784
rect 42240 41720 42256 41784
rect 42320 41720 42336 41784
rect 42400 41720 42416 41784
rect 42480 41720 42496 41784
rect 42560 41720 42576 41784
rect 42640 41720 42656 41784
rect 42720 41720 42736 41784
rect 42800 41720 42816 41784
rect 42880 41720 42896 41784
rect 42960 41720 42976 41784
rect 43040 41720 43056 41784
rect 43120 41720 43136 41784
rect 43200 41720 43216 41784
rect 43280 41720 43296 41784
rect 43360 41720 43376 41784
rect 43440 41720 43456 41784
rect 43520 41720 43536 41784
rect 43600 41720 43616 41784
rect 43680 41720 43696 41784
rect 43760 41720 43776 41784
rect 43840 41720 43856 41784
rect 43920 41720 43936 41784
rect 44000 41720 44016 41784
rect 44080 41720 44096 41784
rect 44160 41720 44176 41784
rect 44240 41720 44256 41784
rect 44320 41720 44336 41784
rect 44400 41720 44416 41784
rect 44480 41720 44496 41784
rect 44560 41720 44576 41784
rect 44640 41720 44656 41784
rect 44720 41720 44736 41784
rect 44800 41720 44816 41784
rect 44880 41720 44896 41784
rect 44960 41720 44976 41784
rect 45040 41720 45056 41784
rect 45120 41720 45136 41784
rect 45200 41720 45216 41784
rect 45280 41720 45296 41784
rect 45360 41720 45368 41784
rect 0 41704 45368 41720
rect 0 41640 8 41704
rect 72 41640 88 41704
rect 152 41640 168 41704
rect 232 41640 248 41704
rect 312 41640 328 41704
rect 392 41640 408 41704
rect 472 41640 488 41704
rect 552 41640 568 41704
rect 632 41640 648 41704
rect 712 41640 728 41704
rect 792 41640 808 41704
rect 872 41640 888 41704
rect 952 41640 968 41704
rect 1032 41640 1048 41704
rect 1112 41640 1128 41704
rect 1192 41640 1208 41704
rect 1272 41640 1288 41704
rect 1352 41640 1368 41704
rect 1432 41640 1448 41704
rect 1512 41640 1528 41704
rect 1592 41640 1608 41704
rect 1672 41640 1688 41704
rect 1752 41640 1768 41704
rect 1832 41640 1848 41704
rect 1912 41640 1928 41704
rect 1992 41640 2008 41704
rect 2072 41640 2088 41704
rect 2152 41640 2168 41704
rect 2232 41640 2248 41704
rect 2312 41640 2328 41704
rect 2392 41640 2408 41704
rect 2472 41640 2488 41704
rect 2552 41640 2568 41704
rect 2632 41640 2648 41704
rect 2712 41640 2728 41704
rect 2792 41640 2808 41704
rect 2872 41640 2888 41704
rect 2952 41640 2968 41704
rect 3032 41640 3048 41704
rect 3112 41640 3128 41704
rect 3192 41640 3208 41704
rect 3272 41640 3288 41704
rect 3352 41640 3368 41704
rect 3432 41640 3448 41704
rect 3512 41640 3528 41704
rect 3592 41640 3608 41704
rect 3672 41640 3688 41704
rect 3752 41640 3768 41704
rect 3832 41640 3848 41704
rect 3912 41640 3928 41704
rect 3992 41640 19112 41704
rect 19176 41640 19192 41704
rect 19256 41640 19272 41704
rect 19336 41640 19352 41704
rect 19416 41640 29112 41704
rect 29176 41640 29192 41704
rect 29256 41640 29272 41704
rect 29336 41640 29352 41704
rect 29416 41640 41376 41704
rect 41440 41640 41456 41704
rect 41520 41640 41536 41704
rect 41600 41640 41616 41704
rect 41680 41640 41696 41704
rect 41760 41640 41776 41704
rect 41840 41640 41856 41704
rect 41920 41640 41936 41704
rect 42000 41640 42016 41704
rect 42080 41640 42096 41704
rect 42160 41640 42176 41704
rect 42240 41640 42256 41704
rect 42320 41640 42336 41704
rect 42400 41640 42416 41704
rect 42480 41640 42496 41704
rect 42560 41640 42576 41704
rect 42640 41640 42656 41704
rect 42720 41640 42736 41704
rect 42800 41640 42816 41704
rect 42880 41640 42896 41704
rect 42960 41640 42976 41704
rect 43040 41640 43056 41704
rect 43120 41640 43136 41704
rect 43200 41640 43216 41704
rect 43280 41640 43296 41704
rect 43360 41640 43376 41704
rect 43440 41640 43456 41704
rect 43520 41640 43536 41704
rect 43600 41640 43616 41704
rect 43680 41640 43696 41704
rect 43760 41640 43776 41704
rect 43840 41640 43856 41704
rect 43920 41640 43936 41704
rect 44000 41640 44016 41704
rect 44080 41640 44096 41704
rect 44160 41640 44176 41704
rect 44240 41640 44256 41704
rect 44320 41640 44336 41704
rect 44400 41640 44416 41704
rect 44480 41640 44496 41704
rect 44560 41640 44576 41704
rect 44640 41640 44656 41704
rect 44720 41640 44736 41704
rect 44800 41640 44816 41704
rect 44880 41640 44896 41704
rect 44960 41640 44976 41704
rect 45040 41640 45056 41704
rect 45120 41640 45136 41704
rect 45200 41640 45216 41704
rect 45280 41640 45296 41704
rect 45360 41640 45368 41704
rect 0 41624 45368 41640
rect 0 41560 8 41624
rect 72 41560 88 41624
rect 152 41560 168 41624
rect 232 41560 248 41624
rect 312 41560 328 41624
rect 392 41560 408 41624
rect 472 41560 488 41624
rect 552 41560 568 41624
rect 632 41560 648 41624
rect 712 41560 728 41624
rect 792 41560 808 41624
rect 872 41560 888 41624
rect 952 41560 968 41624
rect 1032 41560 1048 41624
rect 1112 41560 1128 41624
rect 1192 41560 1208 41624
rect 1272 41560 1288 41624
rect 1352 41560 1368 41624
rect 1432 41560 1448 41624
rect 1512 41560 1528 41624
rect 1592 41560 1608 41624
rect 1672 41560 1688 41624
rect 1752 41560 1768 41624
rect 1832 41560 1848 41624
rect 1912 41560 1928 41624
rect 1992 41560 2008 41624
rect 2072 41560 2088 41624
rect 2152 41560 2168 41624
rect 2232 41560 2248 41624
rect 2312 41560 2328 41624
rect 2392 41560 2408 41624
rect 2472 41560 2488 41624
rect 2552 41560 2568 41624
rect 2632 41560 2648 41624
rect 2712 41560 2728 41624
rect 2792 41560 2808 41624
rect 2872 41560 2888 41624
rect 2952 41560 2968 41624
rect 3032 41560 3048 41624
rect 3112 41560 3128 41624
rect 3192 41560 3208 41624
rect 3272 41560 3288 41624
rect 3352 41560 3368 41624
rect 3432 41560 3448 41624
rect 3512 41560 3528 41624
rect 3592 41560 3608 41624
rect 3672 41560 3688 41624
rect 3752 41560 3768 41624
rect 3832 41560 3848 41624
rect 3912 41560 3928 41624
rect 3992 41560 19112 41624
rect 19176 41560 19192 41624
rect 19256 41560 19272 41624
rect 19336 41560 19352 41624
rect 19416 41560 29112 41624
rect 29176 41560 29192 41624
rect 29256 41560 29272 41624
rect 29336 41560 29352 41624
rect 29416 41560 41376 41624
rect 41440 41560 41456 41624
rect 41520 41560 41536 41624
rect 41600 41560 41616 41624
rect 41680 41560 41696 41624
rect 41760 41560 41776 41624
rect 41840 41560 41856 41624
rect 41920 41560 41936 41624
rect 42000 41560 42016 41624
rect 42080 41560 42096 41624
rect 42160 41560 42176 41624
rect 42240 41560 42256 41624
rect 42320 41560 42336 41624
rect 42400 41560 42416 41624
rect 42480 41560 42496 41624
rect 42560 41560 42576 41624
rect 42640 41560 42656 41624
rect 42720 41560 42736 41624
rect 42800 41560 42816 41624
rect 42880 41560 42896 41624
rect 42960 41560 42976 41624
rect 43040 41560 43056 41624
rect 43120 41560 43136 41624
rect 43200 41560 43216 41624
rect 43280 41560 43296 41624
rect 43360 41560 43376 41624
rect 43440 41560 43456 41624
rect 43520 41560 43536 41624
rect 43600 41560 43616 41624
rect 43680 41560 43696 41624
rect 43760 41560 43776 41624
rect 43840 41560 43856 41624
rect 43920 41560 43936 41624
rect 44000 41560 44016 41624
rect 44080 41560 44096 41624
rect 44160 41560 44176 41624
rect 44240 41560 44256 41624
rect 44320 41560 44336 41624
rect 44400 41560 44416 41624
rect 44480 41560 44496 41624
rect 44560 41560 44576 41624
rect 44640 41560 44656 41624
rect 44720 41560 44736 41624
rect 44800 41560 44816 41624
rect 44880 41560 44896 41624
rect 44960 41560 44976 41624
rect 45040 41560 45056 41624
rect 45120 41560 45136 41624
rect 45200 41560 45216 41624
rect 45280 41560 45296 41624
rect 45360 41560 45368 41624
rect 0 41544 45368 41560
rect 0 41480 8 41544
rect 72 41480 88 41544
rect 152 41480 168 41544
rect 232 41480 248 41544
rect 312 41480 328 41544
rect 392 41480 408 41544
rect 472 41480 488 41544
rect 552 41480 568 41544
rect 632 41480 648 41544
rect 712 41480 728 41544
rect 792 41480 808 41544
rect 872 41480 888 41544
rect 952 41480 968 41544
rect 1032 41480 1048 41544
rect 1112 41480 1128 41544
rect 1192 41480 1208 41544
rect 1272 41480 1288 41544
rect 1352 41480 1368 41544
rect 1432 41480 1448 41544
rect 1512 41480 1528 41544
rect 1592 41480 1608 41544
rect 1672 41480 1688 41544
rect 1752 41480 1768 41544
rect 1832 41480 1848 41544
rect 1912 41480 1928 41544
rect 1992 41480 2008 41544
rect 2072 41480 2088 41544
rect 2152 41480 2168 41544
rect 2232 41480 2248 41544
rect 2312 41480 2328 41544
rect 2392 41480 2408 41544
rect 2472 41480 2488 41544
rect 2552 41480 2568 41544
rect 2632 41480 2648 41544
rect 2712 41480 2728 41544
rect 2792 41480 2808 41544
rect 2872 41480 2888 41544
rect 2952 41480 2968 41544
rect 3032 41480 3048 41544
rect 3112 41480 3128 41544
rect 3192 41480 3208 41544
rect 3272 41480 3288 41544
rect 3352 41480 3368 41544
rect 3432 41480 3448 41544
rect 3512 41480 3528 41544
rect 3592 41480 3608 41544
rect 3672 41480 3688 41544
rect 3752 41480 3768 41544
rect 3832 41480 3848 41544
rect 3912 41480 3928 41544
rect 3992 41480 19112 41544
rect 19176 41480 19192 41544
rect 19256 41480 19272 41544
rect 19336 41480 19352 41544
rect 19416 41480 29112 41544
rect 29176 41480 29192 41544
rect 29256 41480 29272 41544
rect 29336 41480 29352 41544
rect 29416 41480 41376 41544
rect 41440 41480 41456 41544
rect 41520 41480 41536 41544
rect 41600 41480 41616 41544
rect 41680 41480 41696 41544
rect 41760 41480 41776 41544
rect 41840 41480 41856 41544
rect 41920 41480 41936 41544
rect 42000 41480 42016 41544
rect 42080 41480 42096 41544
rect 42160 41480 42176 41544
rect 42240 41480 42256 41544
rect 42320 41480 42336 41544
rect 42400 41480 42416 41544
rect 42480 41480 42496 41544
rect 42560 41480 42576 41544
rect 42640 41480 42656 41544
rect 42720 41480 42736 41544
rect 42800 41480 42816 41544
rect 42880 41480 42896 41544
rect 42960 41480 42976 41544
rect 43040 41480 43056 41544
rect 43120 41480 43136 41544
rect 43200 41480 43216 41544
rect 43280 41480 43296 41544
rect 43360 41480 43376 41544
rect 43440 41480 43456 41544
rect 43520 41480 43536 41544
rect 43600 41480 43616 41544
rect 43680 41480 43696 41544
rect 43760 41480 43776 41544
rect 43840 41480 43856 41544
rect 43920 41480 43936 41544
rect 44000 41480 44016 41544
rect 44080 41480 44096 41544
rect 44160 41480 44176 41544
rect 44240 41480 44256 41544
rect 44320 41480 44336 41544
rect 44400 41480 44416 41544
rect 44480 41480 44496 41544
rect 44560 41480 44576 41544
rect 44640 41480 44656 41544
rect 44720 41480 44736 41544
rect 44800 41480 44816 41544
rect 44880 41480 44896 41544
rect 44960 41480 44976 41544
rect 45040 41480 45056 41544
rect 45120 41480 45136 41544
rect 45200 41480 45216 41544
rect 45280 41480 45296 41544
rect 45360 41480 45368 41544
rect 0 41464 45368 41480
rect 0 41400 8 41464
rect 72 41400 88 41464
rect 152 41400 168 41464
rect 232 41400 248 41464
rect 312 41400 328 41464
rect 392 41400 408 41464
rect 472 41400 488 41464
rect 552 41400 568 41464
rect 632 41400 648 41464
rect 712 41400 728 41464
rect 792 41400 808 41464
rect 872 41400 888 41464
rect 952 41400 968 41464
rect 1032 41400 1048 41464
rect 1112 41400 1128 41464
rect 1192 41400 1208 41464
rect 1272 41400 1288 41464
rect 1352 41400 1368 41464
rect 1432 41400 1448 41464
rect 1512 41400 1528 41464
rect 1592 41400 1608 41464
rect 1672 41400 1688 41464
rect 1752 41400 1768 41464
rect 1832 41400 1848 41464
rect 1912 41400 1928 41464
rect 1992 41400 2008 41464
rect 2072 41400 2088 41464
rect 2152 41400 2168 41464
rect 2232 41400 2248 41464
rect 2312 41400 2328 41464
rect 2392 41400 2408 41464
rect 2472 41400 2488 41464
rect 2552 41400 2568 41464
rect 2632 41400 2648 41464
rect 2712 41400 2728 41464
rect 2792 41400 2808 41464
rect 2872 41400 2888 41464
rect 2952 41400 2968 41464
rect 3032 41400 3048 41464
rect 3112 41400 3128 41464
rect 3192 41400 3208 41464
rect 3272 41400 3288 41464
rect 3352 41400 3368 41464
rect 3432 41400 3448 41464
rect 3512 41400 3528 41464
rect 3592 41400 3608 41464
rect 3672 41400 3688 41464
rect 3752 41400 3768 41464
rect 3832 41400 3848 41464
rect 3912 41400 3928 41464
rect 3992 41400 19112 41464
rect 19176 41400 19192 41464
rect 19256 41400 19272 41464
rect 19336 41400 19352 41464
rect 19416 41400 29112 41464
rect 29176 41400 29192 41464
rect 29256 41400 29272 41464
rect 29336 41400 29352 41464
rect 29416 41400 41376 41464
rect 41440 41400 41456 41464
rect 41520 41400 41536 41464
rect 41600 41400 41616 41464
rect 41680 41400 41696 41464
rect 41760 41400 41776 41464
rect 41840 41400 41856 41464
rect 41920 41400 41936 41464
rect 42000 41400 42016 41464
rect 42080 41400 42096 41464
rect 42160 41400 42176 41464
rect 42240 41400 42256 41464
rect 42320 41400 42336 41464
rect 42400 41400 42416 41464
rect 42480 41400 42496 41464
rect 42560 41400 42576 41464
rect 42640 41400 42656 41464
rect 42720 41400 42736 41464
rect 42800 41400 42816 41464
rect 42880 41400 42896 41464
rect 42960 41400 42976 41464
rect 43040 41400 43056 41464
rect 43120 41400 43136 41464
rect 43200 41400 43216 41464
rect 43280 41400 43296 41464
rect 43360 41400 43376 41464
rect 43440 41400 43456 41464
rect 43520 41400 43536 41464
rect 43600 41400 43616 41464
rect 43680 41400 43696 41464
rect 43760 41400 43776 41464
rect 43840 41400 43856 41464
rect 43920 41400 43936 41464
rect 44000 41400 44016 41464
rect 44080 41400 44096 41464
rect 44160 41400 44176 41464
rect 44240 41400 44256 41464
rect 44320 41400 44336 41464
rect 44400 41400 44416 41464
rect 44480 41400 44496 41464
rect 44560 41400 44576 41464
rect 44640 41400 44656 41464
rect 44720 41400 44736 41464
rect 44800 41400 44816 41464
rect 44880 41400 44896 41464
rect 44960 41400 44976 41464
rect 45040 41400 45056 41464
rect 45120 41400 45136 41464
rect 45200 41400 45216 41464
rect 45280 41400 45296 41464
rect 45360 41400 45368 41464
rect 0 41392 45368 41400
rect 5000 40384 40368 40392
rect 5000 40320 5008 40384
rect 5072 40320 5088 40384
rect 5152 40320 5168 40384
rect 5232 40320 5248 40384
rect 5312 40320 5328 40384
rect 5392 40320 5408 40384
rect 5472 40320 5488 40384
rect 5552 40320 5568 40384
rect 5632 40320 5648 40384
rect 5712 40320 5728 40384
rect 5792 40320 5808 40384
rect 5872 40320 5888 40384
rect 5952 40320 5968 40384
rect 6032 40320 6048 40384
rect 6112 40320 6128 40384
rect 6192 40320 6208 40384
rect 6272 40320 6288 40384
rect 6352 40320 6368 40384
rect 6432 40320 6448 40384
rect 6512 40320 6528 40384
rect 6592 40320 6608 40384
rect 6672 40320 6688 40384
rect 6752 40320 6768 40384
rect 6832 40320 6848 40384
rect 6912 40320 6928 40384
rect 6992 40320 7008 40384
rect 7072 40320 7088 40384
rect 7152 40320 7168 40384
rect 7232 40320 7248 40384
rect 7312 40320 7328 40384
rect 7392 40320 7408 40384
rect 7472 40320 7488 40384
rect 7552 40320 7568 40384
rect 7632 40320 7648 40384
rect 7712 40320 7728 40384
rect 7792 40320 7808 40384
rect 7872 40320 7888 40384
rect 7952 40320 7968 40384
rect 8032 40320 8048 40384
rect 8112 40320 8128 40384
rect 8192 40320 8208 40384
rect 8272 40320 8288 40384
rect 8352 40320 8368 40384
rect 8432 40320 8448 40384
rect 8512 40320 8528 40384
rect 8592 40320 8608 40384
rect 8672 40320 8688 40384
rect 8752 40320 8768 40384
rect 8832 40320 8848 40384
rect 8912 40320 8928 40384
rect 8992 40320 14112 40384
rect 14176 40320 14192 40384
rect 14256 40320 14272 40384
rect 14336 40320 14352 40384
rect 14416 40320 24112 40384
rect 24176 40320 24192 40384
rect 24256 40320 24272 40384
rect 24336 40320 24352 40384
rect 24416 40320 36376 40384
rect 36440 40320 36456 40384
rect 36520 40320 36536 40384
rect 36600 40320 36616 40384
rect 36680 40320 36696 40384
rect 36760 40320 36776 40384
rect 36840 40320 36856 40384
rect 36920 40320 36936 40384
rect 37000 40320 37016 40384
rect 37080 40320 37096 40384
rect 37160 40320 37176 40384
rect 37240 40320 37256 40384
rect 37320 40320 37336 40384
rect 37400 40320 37416 40384
rect 37480 40320 37496 40384
rect 37560 40320 37576 40384
rect 37640 40320 37656 40384
rect 37720 40320 37736 40384
rect 37800 40320 37816 40384
rect 37880 40320 37896 40384
rect 37960 40320 37976 40384
rect 38040 40320 38056 40384
rect 38120 40320 38136 40384
rect 38200 40320 38216 40384
rect 38280 40320 38296 40384
rect 38360 40320 38376 40384
rect 38440 40320 38456 40384
rect 38520 40320 38536 40384
rect 38600 40320 38616 40384
rect 38680 40320 38696 40384
rect 38760 40320 38776 40384
rect 38840 40320 38856 40384
rect 38920 40320 38936 40384
rect 39000 40320 39016 40384
rect 39080 40320 39096 40384
rect 39160 40320 39176 40384
rect 39240 40320 39256 40384
rect 39320 40320 39336 40384
rect 39400 40320 39416 40384
rect 39480 40320 39496 40384
rect 39560 40320 39576 40384
rect 39640 40320 39656 40384
rect 39720 40320 39736 40384
rect 39800 40320 39816 40384
rect 39880 40320 39896 40384
rect 39960 40320 39976 40384
rect 40040 40320 40056 40384
rect 40120 40320 40136 40384
rect 40200 40320 40216 40384
rect 40280 40320 40296 40384
rect 40360 40320 40368 40384
rect 5000 40304 40368 40320
rect 5000 40240 5008 40304
rect 5072 40240 5088 40304
rect 5152 40240 5168 40304
rect 5232 40240 5248 40304
rect 5312 40240 5328 40304
rect 5392 40240 5408 40304
rect 5472 40240 5488 40304
rect 5552 40240 5568 40304
rect 5632 40240 5648 40304
rect 5712 40240 5728 40304
rect 5792 40240 5808 40304
rect 5872 40240 5888 40304
rect 5952 40240 5968 40304
rect 6032 40240 6048 40304
rect 6112 40240 6128 40304
rect 6192 40240 6208 40304
rect 6272 40240 6288 40304
rect 6352 40240 6368 40304
rect 6432 40240 6448 40304
rect 6512 40240 6528 40304
rect 6592 40240 6608 40304
rect 6672 40240 6688 40304
rect 6752 40240 6768 40304
rect 6832 40240 6848 40304
rect 6912 40240 6928 40304
rect 6992 40240 7008 40304
rect 7072 40240 7088 40304
rect 7152 40240 7168 40304
rect 7232 40240 7248 40304
rect 7312 40240 7328 40304
rect 7392 40240 7408 40304
rect 7472 40240 7488 40304
rect 7552 40240 7568 40304
rect 7632 40240 7648 40304
rect 7712 40240 7728 40304
rect 7792 40240 7808 40304
rect 7872 40240 7888 40304
rect 7952 40240 7968 40304
rect 8032 40240 8048 40304
rect 8112 40240 8128 40304
rect 8192 40240 8208 40304
rect 8272 40240 8288 40304
rect 8352 40240 8368 40304
rect 8432 40240 8448 40304
rect 8512 40240 8528 40304
rect 8592 40240 8608 40304
rect 8672 40240 8688 40304
rect 8752 40240 8768 40304
rect 8832 40240 8848 40304
rect 8912 40240 8928 40304
rect 8992 40240 14112 40304
rect 14176 40240 14192 40304
rect 14256 40240 14272 40304
rect 14336 40240 14352 40304
rect 14416 40240 24112 40304
rect 24176 40240 24192 40304
rect 24256 40240 24272 40304
rect 24336 40240 24352 40304
rect 24416 40240 36376 40304
rect 36440 40240 36456 40304
rect 36520 40240 36536 40304
rect 36600 40240 36616 40304
rect 36680 40240 36696 40304
rect 36760 40240 36776 40304
rect 36840 40240 36856 40304
rect 36920 40240 36936 40304
rect 37000 40240 37016 40304
rect 37080 40240 37096 40304
rect 37160 40240 37176 40304
rect 37240 40240 37256 40304
rect 37320 40240 37336 40304
rect 37400 40240 37416 40304
rect 37480 40240 37496 40304
rect 37560 40240 37576 40304
rect 37640 40240 37656 40304
rect 37720 40240 37736 40304
rect 37800 40240 37816 40304
rect 37880 40240 37896 40304
rect 37960 40240 37976 40304
rect 38040 40240 38056 40304
rect 38120 40240 38136 40304
rect 38200 40240 38216 40304
rect 38280 40240 38296 40304
rect 38360 40240 38376 40304
rect 38440 40240 38456 40304
rect 38520 40240 38536 40304
rect 38600 40240 38616 40304
rect 38680 40240 38696 40304
rect 38760 40240 38776 40304
rect 38840 40240 38856 40304
rect 38920 40240 38936 40304
rect 39000 40240 39016 40304
rect 39080 40240 39096 40304
rect 39160 40240 39176 40304
rect 39240 40240 39256 40304
rect 39320 40240 39336 40304
rect 39400 40240 39416 40304
rect 39480 40240 39496 40304
rect 39560 40240 39576 40304
rect 39640 40240 39656 40304
rect 39720 40240 39736 40304
rect 39800 40240 39816 40304
rect 39880 40240 39896 40304
rect 39960 40240 39976 40304
rect 40040 40240 40056 40304
rect 40120 40240 40136 40304
rect 40200 40240 40216 40304
rect 40280 40240 40296 40304
rect 40360 40240 40368 40304
rect 5000 40224 40368 40240
rect 5000 40160 5008 40224
rect 5072 40160 5088 40224
rect 5152 40160 5168 40224
rect 5232 40160 5248 40224
rect 5312 40160 5328 40224
rect 5392 40160 5408 40224
rect 5472 40160 5488 40224
rect 5552 40160 5568 40224
rect 5632 40160 5648 40224
rect 5712 40160 5728 40224
rect 5792 40160 5808 40224
rect 5872 40160 5888 40224
rect 5952 40160 5968 40224
rect 6032 40160 6048 40224
rect 6112 40160 6128 40224
rect 6192 40160 6208 40224
rect 6272 40160 6288 40224
rect 6352 40160 6368 40224
rect 6432 40160 6448 40224
rect 6512 40160 6528 40224
rect 6592 40160 6608 40224
rect 6672 40160 6688 40224
rect 6752 40160 6768 40224
rect 6832 40160 6848 40224
rect 6912 40160 6928 40224
rect 6992 40160 7008 40224
rect 7072 40160 7088 40224
rect 7152 40160 7168 40224
rect 7232 40160 7248 40224
rect 7312 40160 7328 40224
rect 7392 40160 7408 40224
rect 7472 40160 7488 40224
rect 7552 40160 7568 40224
rect 7632 40160 7648 40224
rect 7712 40160 7728 40224
rect 7792 40160 7808 40224
rect 7872 40160 7888 40224
rect 7952 40160 7968 40224
rect 8032 40160 8048 40224
rect 8112 40160 8128 40224
rect 8192 40160 8208 40224
rect 8272 40160 8288 40224
rect 8352 40160 8368 40224
rect 8432 40160 8448 40224
rect 8512 40160 8528 40224
rect 8592 40160 8608 40224
rect 8672 40160 8688 40224
rect 8752 40160 8768 40224
rect 8832 40160 8848 40224
rect 8912 40160 8928 40224
rect 8992 40160 14112 40224
rect 14176 40160 14192 40224
rect 14256 40160 14272 40224
rect 14336 40160 14352 40224
rect 14416 40160 24112 40224
rect 24176 40160 24192 40224
rect 24256 40160 24272 40224
rect 24336 40160 24352 40224
rect 24416 40160 36376 40224
rect 36440 40160 36456 40224
rect 36520 40160 36536 40224
rect 36600 40160 36616 40224
rect 36680 40160 36696 40224
rect 36760 40160 36776 40224
rect 36840 40160 36856 40224
rect 36920 40160 36936 40224
rect 37000 40160 37016 40224
rect 37080 40160 37096 40224
rect 37160 40160 37176 40224
rect 37240 40160 37256 40224
rect 37320 40160 37336 40224
rect 37400 40160 37416 40224
rect 37480 40160 37496 40224
rect 37560 40160 37576 40224
rect 37640 40160 37656 40224
rect 37720 40160 37736 40224
rect 37800 40160 37816 40224
rect 37880 40160 37896 40224
rect 37960 40160 37976 40224
rect 38040 40160 38056 40224
rect 38120 40160 38136 40224
rect 38200 40160 38216 40224
rect 38280 40160 38296 40224
rect 38360 40160 38376 40224
rect 38440 40160 38456 40224
rect 38520 40160 38536 40224
rect 38600 40160 38616 40224
rect 38680 40160 38696 40224
rect 38760 40160 38776 40224
rect 38840 40160 38856 40224
rect 38920 40160 38936 40224
rect 39000 40160 39016 40224
rect 39080 40160 39096 40224
rect 39160 40160 39176 40224
rect 39240 40160 39256 40224
rect 39320 40160 39336 40224
rect 39400 40160 39416 40224
rect 39480 40160 39496 40224
rect 39560 40160 39576 40224
rect 39640 40160 39656 40224
rect 39720 40160 39736 40224
rect 39800 40160 39816 40224
rect 39880 40160 39896 40224
rect 39960 40160 39976 40224
rect 40040 40160 40056 40224
rect 40120 40160 40136 40224
rect 40200 40160 40216 40224
rect 40280 40160 40296 40224
rect 40360 40160 40368 40224
rect 5000 40144 40368 40160
rect 5000 40080 5008 40144
rect 5072 40080 5088 40144
rect 5152 40080 5168 40144
rect 5232 40080 5248 40144
rect 5312 40080 5328 40144
rect 5392 40080 5408 40144
rect 5472 40080 5488 40144
rect 5552 40080 5568 40144
rect 5632 40080 5648 40144
rect 5712 40080 5728 40144
rect 5792 40080 5808 40144
rect 5872 40080 5888 40144
rect 5952 40080 5968 40144
rect 6032 40080 6048 40144
rect 6112 40080 6128 40144
rect 6192 40080 6208 40144
rect 6272 40080 6288 40144
rect 6352 40080 6368 40144
rect 6432 40080 6448 40144
rect 6512 40080 6528 40144
rect 6592 40080 6608 40144
rect 6672 40080 6688 40144
rect 6752 40080 6768 40144
rect 6832 40080 6848 40144
rect 6912 40080 6928 40144
rect 6992 40080 7008 40144
rect 7072 40080 7088 40144
rect 7152 40080 7168 40144
rect 7232 40080 7248 40144
rect 7312 40080 7328 40144
rect 7392 40080 7408 40144
rect 7472 40080 7488 40144
rect 7552 40080 7568 40144
rect 7632 40080 7648 40144
rect 7712 40080 7728 40144
rect 7792 40080 7808 40144
rect 7872 40080 7888 40144
rect 7952 40080 7968 40144
rect 8032 40080 8048 40144
rect 8112 40080 8128 40144
rect 8192 40080 8208 40144
rect 8272 40080 8288 40144
rect 8352 40080 8368 40144
rect 8432 40080 8448 40144
rect 8512 40080 8528 40144
rect 8592 40080 8608 40144
rect 8672 40080 8688 40144
rect 8752 40080 8768 40144
rect 8832 40080 8848 40144
rect 8912 40080 8928 40144
rect 8992 40080 14112 40144
rect 14176 40080 14192 40144
rect 14256 40080 14272 40144
rect 14336 40080 14352 40144
rect 14416 40080 24112 40144
rect 24176 40080 24192 40144
rect 24256 40080 24272 40144
rect 24336 40080 24352 40144
rect 24416 40080 36376 40144
rect 36440 40080 36456 40144
rect 36520 40080 36536 40144
rect 36600 40080 36616 40144
rect 36680 40080 36696 40144
rect 36760 40080 36776 40144
rect 36840 40080 36856 40144
rect 36920 40080 36936 40144
rect 37000 40080 37016 40144
rect 37080 40080 37096 40144
rect 37160 40080 37176 40144
rect 37240 40080 37256 40144
rect 37320 40080 37336 40144
rect 37400 40080 37416 40144
rect 37480 40080 37496 40144
rect 37560 40080 37576 40144
rect 37640 40080 37656 40144
rect 37720 40080 37736 40144
rect 37800 40080 37816 40144
rect 37880 40080 37896 40144
rect 37960 40080 37976 40144
rect 38040 40080 38056 40144
rect 38120 40080 38136 40144
rect 38200 40080 38216 40144
rect 38280 40080 38296 40144
rect 38360 40080 38376 40144
rect 38440 40080 38456 40144
rect 38520 40080 38536 40144
rect 38600 40080 38616 40144
rect 38680 40080 38696 40144
rect 38760 40080 38776 40144
rect 38840 40080 38856 40144
rect 38920 40080 38936 40144
rect 39000 40080 39016 40144
rect 39080 40080 39096 40144
rect 39160 40080 39176 40144
rect 39240 40080 39256 40144
rect 39320 40080 39336 40144
rect 39400 40080 39416 40144
rect 39480 40080 39496 40144
rect 39560 40080 39576 40144
rect 39640 40080 39656 40144
rect 39720 40080 39736 40144
rect 39800 40080 39816 40144
rect 39880 40080 39896 40144
rect 39960 40080 39976 40144
rect 40040 40080 40056 40144
rect 40120 40080 40136 40144
rect 40200 40080 40216 40144
rect 40280 40080 40296 40144
rect 40360 40080 40368 40144
rect 5000 40064 40368 40080
rect 5000 40000 5008 40064
rect 5072 40000 5088 40064
rect 5152 40000 5168 40064
rect 5232 40000 5248 40064
rect 5312 40000 5328 40064
rect 5392 40000 5408 40064
rect 5472 40000 5488 40064
rect 5552 40000 5568 40064
rect 5632 40000 5648 40064
rect 5712 40000 5728 40064
rect 5792 40000 5808 40064
rect 5872 40000 5888 40064
rect 5952 40000 5968 40064
rect 6032 40000 6048 40064
rect 6112 40000 6128 40064
rect 6192 40000 6208 40064
rect 6272 40000 6288 40064
rect 6352 40000 6368 40064
rect 6432 40000 6448 40064
rect 6512 40000 6528 40064
rect 6592 40000 6608 40064
rect 6672 40000 6688 40064
rect 6752 40000 6768 40064
rect 6832 40000 6848 40064
rect 6912 40000 6928 40064
rect 6992 40000 7008 40064
rect 7072 40000 7088 40064
rect 7152 40000 7168 40064
rect 7232 40000 7248 40064
rect 7312 40000 7328 40064
rect 7392 40000 7408 40064
rect 7472 40000 7488 40064
rect 7552 40000 7568 40064
rect 7632 40000 7648 40064
rect 7712 40000 7728 40064
rect 7792 40000 7808 40064
rect 7872 40000 7888 40064
rect 7952 40000 7968 40064
rect 8032 40000 8048 40064
rect 8112 40000 8128 40064
rect 8192 40000 8208 40064
rect 8272 40000 8288 40064
rect 8352 40000 8368 40064
rect 8432 40000 8448 40064
rect 8512 40000 8528 40064
rect 8592 40000 8608 40064
rect 8672 40000 8688 40064
rect 8752 40000 8768 40064
rect 8832 40000 8848 40064
rect 8912 40000 8928 40064
rect 8992 40000 14112 40064
rect 14176 40000 14192 40064
rect 14256 40000 14272 40064
rect 14336 40000 14352 40064
rect 14416 40000 24112 40064
rect 24176 40000 24192 40064
rect 24256 40000 24272 40064
rect 24336 40000 24352 40064
rect 24416 40000 36376 40064
rect 36440 40000 36456 40064
rect 36520 40000 36536 40064
rect 36600 40000 36616 40064
rect 36680 40000 36696 40064
rect 36760 40000 36776 40064
rect 36840 40000 36856 40064
rect 36920 40000 36936 40064
rect 37000 40000 37016 40064
rect 37080 40000 37096 40064
rect 37160 40000 37176 40064
rect 37240 40000 37256 40064
rect 37320 40000 37336 40064
rect 37400 40000 37416 40064
rect 37480 40000 37496 40064
rect 37560 40000 37576 40064
rect 37640 40000 37656 40064
rect 37720 40000 37736 40064
rect 37800 40000 37816 40064
rect 37880 40000 37896 40064
rect 37960 40000 37976 40064
rect 38040 40000 38056 40064
rect 38120 40000 38136 40064
rect 38200 40000 38216 40064
rect 38280 40000 38296 40064
rect 38360 40000 38376 40064
rect 38440 40000 38456 40064
rect 38520 40000 38536 40064
rect 38600 40000 38616 40064
rect 38680 40000 38696 40064
rect 38760 40000 38776 40064
rect 38840 40000 38856 40064
rect 38920 40000 38936 40064
rect 39000 40000 39016 40064
rect 39080 40000 39096 40064
rect 39160 40000 39176 40064
rect 39240 40000 39256 40064
rect 39320 40000 39336 40064
rect 39400 40000 39416 40064
rect 39480 40000 39496 40064
rect 39560 40000 39576 40064
rect 39640 40000 39656 40064
rect 39720 40000 39736 40064
rect 39800 40000 39816 40064
rect 39880 40000 39896 40064
rect 39960 40000 39976 40064
rect 40040 40000 40056 40064
rect 40120 40000 40136 40064
rect 40200 40000 40216 40064
rect 40280 40000 40296 40064
rect 40360 40000 40368 40064
rect 5000 39984 40368 40000
rect 5000 39920 5008 39984
rect 5072 39920 5088 39984
rect 5152 39920 5168 39984
rect 5232 39920 5248 39984
rect 5312 39920 5328 39984
rect 5392 39920 5408 39984
rect 5472 39920 5488 39984
rect 5552 39920 5568 39984
rect 5632 39920 5648 39984
rect 5712 39920 5728 39984
rect 5792 39920 5808 39984
rect 5872 39920 5888 39984
rect 5952 39920 5968 39984
rect 6032 39920 6048 39984
rect 6112 39920 6128 39984
rect 6192 39920 6208 39984
rect 6272 39920 6288 39984
rect 6352 39920 6368 39984
rect 6432 39920 6448 39984
rect 6512 39920 6528 39984
rect 6592 39920 6608 39984
rect 6672 39920 6688 39984
rect 6752 39920 6768 39984
rect 6832 39920 6848 39984
rect 6912 39920 6928 39984
rect 6992 39920 7008 39984
rect 7072 39920 7088 39984
rect 7152 39920 7168 39984
rect 7232 39920 7248 39984
rect 7312 39920 7328 39984
rect 7392 39920 7408 39984
rect 7472 39920 7488 39984
rect 7552 39920 7568 39984
rect 7632 39920 7648 39984
rect 7712 39920 7728 39984
rect 7792 39920 7808 39984
rect 7872 39920 7888 39984
rect 7952 39920 7968 39984
rect 8032 39920 8048 39984
rect 8112 39920 8128 39984
rect 8192 39920 8208 39984
rect 8272 39920 8288 39984
rect 8352 39920 8368 39984
rect 8432 39920 8448 39984
rect 8512 39920 8528 39984
rect 8592 39920 8608 39984
rect 8672 39920 8688 39984
rect 8752 39920 8768 39984
rect 8832 39920 8848 39984
rect 8912 39920 8928 39984
rect 8992 39920 14112 39984
rect 14176 39920 14192 39984
rect 14256 39920 14272 39984
rect 14336 39920 14352 39984
rect 14416 39920 24112 39984
rect 24176 39920 24192 39984
rect 24256 39920 24272 39984
rect 24336 39920 24352 39984
rect 24416 39920 36376 39984
rect 36440 39920 36456 39984
rect 36520 39920 36536 39984
rect 36600 39920 36616 39984
rect 36680 39920 36696 39984
rect 36760 39920 36776 39984
rect 36840 39920 36856 39984
rect 36920 39920 36936 39984
rect 37000 39920 37016 39984
rect 37080 39920 37096 39984
rect 37160 39920 37176 39984
rect 37240 39920 37256 39984
rect 37320 39920 37336 39984
rect 37400 39920 37416 39984
rect 37480 39920 37496 39984
rect 37560 39920 37576 39984
rect 37640 39920 37656 39984
rect 37720 39920 37736 39984
rect 37800 39920 37816 39984
rect 37880 39920 37896 39984
rect 37960 39920 37976 39984
rect 38040 39920 38056 39984
rect 38120 39920 38136 39984
rect 38200 39920 38216 39984
rect 38280 39920 38296 39984
rect 38360 39920 38376 39984
rect 38440 39920 38456 39984
rect 38520 39920 38536 39984
rect 38600 39920 38616 39984
rect 38680 39920 38696 39984
rect 38760 39920 38776 39984
rect 38840 39920 38856 39984
rect 38920 39920 38936 39984
rect 39000 39920 39016 39984
rect 39080 39920 39096 39984
rect 39160 39920 39176 39984
rect 39240 39920 39256 39984
rect 39320 39920 39336 39984
rect 39400 39920 39416 39984
rect 39480 39920 39496 39984
rect 39560 39920 39576 39984
rect 39640 39920 39656 39984
rect 39720 39920 39736 39984
rect 39800 39920 39816 39984
rect 39880 39920 39896 39984
rect 39960 39920 39976 39984
rect 40040 39920 40056 39984
rect 40120 39920 40136 39984
rect 40200 39920 40216 39984
rect 40280 39920 40296 39984
rect 40360 39920 40368 39984
rect 5000 39904 40368 39920
rect 5000 39840 5008 39904
rect 5072 39840 5088 39904
rect 5152 39840 5168 39904
rect 5232 39840 5248 39904
rect 5312 39840 5328 39904
rect 5392 39840 5408 39904
rect 5472 39840 5488 39904
rect 5552 39840 5568 39904
rect 5632 39840 5648 39904
rect 5712 39840 5728 39904
rect 5792 39840 5808 39904
rect 5872 39840 5888 39904
rect 5952 39840 5968 39904
rect 6032 39840 6048 39904
rect 6112 39840 6128 39904
rect 6192 39840 6208 39904
rect 6272 39840 6288 39904
rect 6352 39840 6368 39904
rect 6432 39840 6448 39904
rect 6512 39840 6528 39904
rect 6592 39840 6608 39904
rect 6672 39840 6688 39904
rect 6752 39840 6768 39904
rect 6832 39840 6848 39904
rect 6912 39840 6928 39904
rect 6992 39840 7008 39904
rect 7072 39840 7088 39904
rect 7152 39840 7168 39904
rect 7232 39840 7248 39904
rect 7312 39840 7328 39904
rect 7392 39840 7408 39904
rect 7472 39840 7488 39904
rect 7552 39840 7568 39904
rect 7632 39840 7648 39904
rect 7712 39840 7728 39904
rect 7792 39840 7808 39904
rect 7872 39840 7888 39904
rect 7952 39840 7968 39904
rect 8032 39840 8048 39904
rect 8112 39840 8128 39904
rect 8192 39840 8208 39904
rect 8272 39840 8288 39904
rect 8352 39840 8368 39904
rect 8432 39840 8448 39904
rect 8512 39840 8528 39904
rect 8592 39840 8608 39904
rect 8672 39840 8688 39904
rect 8752 39840 8768 39904
rect 8832 39840 8848 39904
rect 8912 39840 8928 39904
rect 8992 39840 14112 39904
rect 14176 39840 14192 39904
rect 14256 39840 14272 39904
rect 14336 39840 14352 39904
rect 14416 39840 24112 39904
rect 24176 39840 24192 39904
rect 24256 39840 24272 39904
rect 24336 39840 24352 39904
rect 24416 39840 36376 39904
rect 36440 39840 36456 39904
rect 36520 39840 36536 39904
rect 36600 39840 36616 39904
rect 36680 39840 36696 39904
rect 36760 39840 36776 39904
rect 36840 39840 36856 39904
rect 36920 39840 36936 39904
rect 37000 39840 37016 39904
rect 37080 39840 37096 39904
rect 37160 39840 37176 39904
rect 37240 39840 37256 39904
rect 37320 39840 37336 39904
rect 37400 39840 37416 39904
rect 37480 39840 37496 39904
rect 37560 39840 37576 39904
rect 37640 39840 37656 39904
rect 37720 39840 37736 39904
rect 37800 39840 37816 39904
rect 37880 39840 37896 39904
rect 37960 39840 37976 39904
rect 38040 39840 38056 39904
rect 38120 39840 38136 39904
rect 38200 39840 38216 39904
rect 38280 39840 38296 39904
rect 38360 39840 38376 39904
rect 38440 39840 38456 39904
rect 38520 39840 38536 39904
rect 38600 39840 38616 39904
rect 38680 39840 38696 39904
rect 38760 39840 38776 39904
rect 38840 39840 38856 39904
rect 38920 39840 38936 39904
rect 39000 39840 39016 39904
rect 39080 39840 39096 39904
rect 39160 39840 39176 39904
rect 39240 39840 39256 39904
rect 39320 39840 39336 39904
rect 39400 39840 39416 39904
rect 39480 39840 39496 39904
rect 39560 39840 39576 39904
rect 39640 39840 39656 39904
rect 39720 39840 39736 39904
rect 39800 39840 39816 39904
rect 39880 39840 39896 39904
rect 39960 39840 39976 39904
rect 40040 39840 40056 39904
rect 40120 39840 40136 39904
rect 40200 39840 40216 39904
rect 40280 39840 40296 39904
rect 40360 39840 40368 39904
rect 5000 39824 40368 39840
rect 5000 39760 5008 39824
rect 5072 39760 5088 39824
rect 5152 39760 5168 39824
rect 5232 39760 5248 39824
rect 5312 39760 5328 39824
rect 5392 39760 5408 39824
rect 5472 39760 5488 39824
rect 5552 39760 5568 39824
rect 5632 39760 5648 39824
rect 5712 39760 5728 39824
rect 5792 39760 5808 39824
rect 5872 39760 5888 39824
rect 5952 39760 5968 39824
rect 6032 39760 6048 39824
rect 6112 39760 6128 39824
rect 6192 39760 6208 39824
rect 6272 39760 6288 39824
rect 6352 39760 6368 39824
rect 6432 39760 6448 39824
rect 6512 39760 6528 39824
rect 6592 39760 6608 39824
rect 6672 39760 6688 39824
rect 6752 39760 6768 39824
rect 6832 39760 6848 39824
rect 6912 39760 6928 39824
rect 6992 39760 7008 39824
rect 7072 39760 7088 39824
rect 7152 39760 7168 39824
rect 7232 39760 7248 39824
rect 7312 39760 7328 39824
rect 7392 39760 7408 39824
rect 7472 39760 7488 39824
rect 7552 39760 7568 39824
rect 7632 39760 7648 39824
rect 7712 39760 7728 39824
rect 7792 39760 7808 39824
rect 7872 39760 7888 39824
rect 7952 39760 7968 39824
rect 8032 39760 8048 39824
rect 8112 39760 8128 39824
rect 8192 39760 8208 39824
rect 8272 39760 8288 39824
rect 8352 39760 8368 39824
rect 8432 39760 8448 39824
rect 8512 39760 8528 39824
rect 8592 39760 8608 39824
rect 8672 39760 8688 39824
rect 8752 39760 8768 39824
rect 8832 39760 8848 39824
rect 8912 39760 8928 39824
rect 8992 39760 14112 39824
rect 14176 39760 14192 39824
rect 14256 39760 14272 39824
rect 14336 39760 14352 39824
rect 14416 39760 24112 39824
rect 24176 39760 24192 39824
rect 24256 39760 24272 39824
rect 24336 39760 24352 39824
rect 24416 39760 36376 39824
rect 36440 39760 36456 39824
rect 36520 39760 36536 39824
rect 36600 39760 36616 39824
rect 36680 39760 36696 39824
rect 36760 39760 36776 39824
rect 36840 39760 36856 39824
rect 36920 39760 36936 39824
rect 37000 39760 37016 39824
rect 37080 39760 37096 39824
rect 37160 39760 37176 39824
rect 37240 39760 37256 39824
rect 37320 39760 37336 39824
rect 37400 39760 37416 39824
rect 37480 39760 37496 39824
rect 37560 39760 37576 39824
rect 37640 39760 37656 39824
rect 37720 39760 37736 39824
rect 37800 39760 37816 39824
rect 37880 39760 37896 39824
rect 37960 39760 37976 39824
rect 38040 39760 38056 39824
rect 38120 39760 38136 39824
rect 38200 39760 38216 39824
rect 38280 39760 38296 39824
rect 38360 39760 38376 39824
rect 38440 39760 38456 39824
rect 38520 39760 38536 39824
rect 38600 39760 38616 39824
rect 38680 39760 38696 39824
rect 38760 39760 38776 39824
rect 38840 39760 38856 39824
rect 38920 39760 38936 39824
rect 39000 39760 39016 39824
rect 39080 39760 39096 39824
rect 39160 39760 39176 39824
rect 39240 39760 39256 39824
rect 39320 39760 39336 39824
rect 39400 39760 39416 39824
rect 39480 39760 39496 39824
rect 39560 39760 39576 39824
rect 39640 39760 39656 39824
rect 39720 39760 39736 39824
rect 39800 39760 39816 39824
rect 39880 39760 39896 39824
rect 39960 39760 39976 39824
rect 40040 39760 40056 39824
rect 40120 39760 40136 39824
rect 40200 39760 40216 39824
rect 40280 39760 40296 39824
rect 40360 39760 40368 39824
rect 5000 39744 40368 39760
rect 5000 39680 5008 39744
rect 5072 39680 5088 39744
rect 5152 39680 5168 39744
rect 5232 39680 5248 39744
rect 5312 39680 5328 39744
rect 5392 39680 5408 39744
rect 5472 39680 5488 39744
rect 5552 39680 5568 39744
rect 5632 39680 5648 39744
rect 5712 39680 5728 39744
rect 5792 39680 5808 39744
rect 5872 39680 5888 39744
rect 5952 39680 5968 39744
rect 6032 39680 6048 39744
rect 6112 39680 6128 39744
rect 6192 39680 6208 39744
rect 6272 39680 6288 39744
rect 6352 39680 6368 39744
rect 6432 39680 6448 39744
rect 6512 39680 6528 39744
rect 6592 39680 6608 39744
rect 6672 39680 6688 39744
rect 6752 39680 6768 39744
rect 6832 39680 6848 39744
rect 6912 39680 6928 39744
rect 6992 39680 7008 39744
rect 7072 39680 7088 39744
rect 7152 39680 7168 39744
rect 7232 39680 7248 39744
rect 7312 39680 7328 39744
rect 7392 39680 7408 39744
rect 7472 39680 7488 39744
rect 7552 39680 7568 39744
rect 7632 39680 7648 39744
rect 7712 39680 7728 39744
rect 7792 39680 7808 39744
rect 7872 39680 7888 39744
rect 7952 39680 7968 39744
rect 8032 39680 8048 39744
rect 8112 39680 8128 39744
rect 8192 39680 8208 39744
rect 8272 39680 8288 39744
rect 8352 39680 8368 39744
rect 8432 39680 8448 39744
rect 8512 39680 8528 39744
rect 8592 39680 8608 39744
rect 8672 39680 8688 39744
rect 8752 39680 8768 39744
rect 8832 39680 8848 39744
rect 8912 39680 8928 39744
rect 8992 39680 14112 39744
rect 14176 39680 14192 39744
rect 14256 39680 14272 39744
rect 14336 39680 14352 39744
rect 14416 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 36376 39744
rect 36440 39680 36456 39744
rect 36520 39680 36536 39744
rect 36600 39680 36616 39744
rect 36680 39680 36696 39744
rect 36760 39680 36776 39744
rect 36840 39680 36856 39744
rect 36920 39680 36936 39744
rect 37000 39680 37016 39744
rect 37080 39680 37096 39744
rect 37160 39680 37176 39744
rect 37240 39680 37256 39744
rect 37320 39680 37336 39744
rect 37400 39680 37416 39744
rect 37480 39680 37496 39744
rect 37560 39680 37576 39744
rect 37640 39680 37656 39744
rect 37720 39680 37736 39744
rect 37800 39680 37816 39744
rect 37880 39680 37896 39744
rect 37960 39680 37976 39744
rect 38040 39680 38056 39744
rect 38120 39680 38136 39744
rect 38200 39680 38216 39744
rect 38280 39680 38296 39744
rect 38360 39680 38376 39744
rect 38440 39680 38456 39744
rect 38520 39680 38536 39744
rect 38600 39680 38616 39744
rect 38680 39680 38696 39744
rect 38760 39680 38776 39744
rect 38840 39680 38856 39744
rect 38920 39680 38936 39744
rect 39000 39680 39016 39744
rect 39080 39680 39096 39744
rect 39160 39680 39176 39744
rect 39240 39680 39256 39744
rect 39320 39680 39336 39744
rect 39400 39680 39416 39744
rect 39480 39680 39496 39744
rect 39560 39680 39576 39744
rect 39640 39680 39656 39744
rect 39720 39680 39736 39744
rect 39800 39680 39816 39744
rect 39880 39680 39896 39744
rect 39960 39680 39976 39744
rect 40040 39680 40056 39744
rect 40120 39680 40136 39744
rect 40200 39680 40216 39744
rect 40280 39680 40296 39744
rect 40360 39680 40368 39744
rect 5000 39664 40368 39680
rect 5000 39600 5008 39664
rect 5072 39600 5088 39664
rect 5152 39600 5168 39664
rect 5232 39600 5248 39664
rect 5312 39600 5328 39664
rect 5392 39600 5408 39664
rect 5472 39600 5488 39664
rect 5552 39600 5568 39664
rect 5632 39600 5648 39664
rect 5712 39600 5728 39664
rect 5792 39600 5808 39664
rect 5872 39600 5888 39664
rect 5952 39600 5968 39664
rect 6032 39600 6048 39664
rect 6112 39600 6128 39664
rect 6192 39600 6208 39664
rect 6272 39600 6288 39664
rect 6352 39600 6368 39664
rect 6432 39600 6448 39664
rect 6512 39600 6528 39664
rect 6592 39600 6608 39664
rect 6672 39600 6688 39664
rect 6752 39600 6768 39664
rect 6832 39600 6848 39664
rect 6912 39600 6928 39664
rect 6992 39600 7008 39664
rect 7072 39600 7088 39664
rect 7152 39600 7168 39664
rect 7232 39600 7248 39664
rect 7312 39600 7328 39664
rect 7392 39600 7408 39664
rect 7472 39600 7488 39664
rect 7552 39600 7568 39664
rect 7632 39600 7648 39664
rect 7712 39600 7728 39664
rect 7792 39600 7808 39664
rect 7872 39600 7888 39664
rect 7952 39600 7968 39664
rect 8032 39600 8048 39664
rect 8112 39600 8128 39664
rect 8192 39600 8208 39664
rect 8272 39600 8288 39664
rect 8352 39600 8368 39664
rect 8432 39600 8448 39664
rect 8512 39600 8528 39664
rect 8592 39600 8608 39664
rect 8672 39600 8688 39664
rect 8752 39600 8768 39664
rect 8832 39600 8848 39664
rect 8912 39600 8928 39664
rect 8992 39600 14112 39664
rect 14176 39600 14192 39664
rect 14256 39600 14272 39664
rect 14336 39600 14352 39664
rect 14416 39600 24112 39664
rect 24176 39600 24192 39664
rect 24256 39600 24272 39664
rect 24336 39600 24352 39664
rect 24416 39600 36376 39664
rect 36440 39600 36456 39664
rect 36520 39600 36536 39664
rect 36600 39600 36616 39664
rect 36680 39600 36696 39664
rect 36760 39600 36776 39664
rect 36840 39600 36856 39664
rect 36920 39600 36936 39664
rect 37000 39600 37016 39664
rect 37080 39600 37096 39664
rect 37160 39600 37176 39664
rect 37240 39600 37256 39664
rect 37320 39600 37336 39664
rect 37400 39600 37416 39664
rect 37480 39600 37496 39664
rect 37560 39600 37576 39664
rect 37640 39600 37656 39664
rect 37720 39600 37736 39664
rect 37800 39600 37816 39664
rect 37880 39600 37896 39664
rect 37960 39600 37976 39664
rect 38040 39600 38056 39664
rect 38120 39600 38136 39664
rect 38200 39600 38216 39664
rect 38280 39600 38296 39664
rect 38360 39600 38376 39664
rect 38440 39600 38456 39664
rect 38520 39600 38536 39664
rect 38600 39600 38616 39664
rect 38680 39600 38696 39664
rect 38760 39600 38776 39664
rect 38840 39600 38856 39664
rect 38920 39600 38936 39664
rect 39000 39600 39016 39664
rect 39080 39600 39096 39664
rect 39160 39600 39176 39664
rect 39240 39600 39256 39664
rect 39320 39600 39336 39664
rect 39400 39600 39416 39664
rect 39480 39600 39496 39664
rect 39560 39600 39576 39664
rect 39640 39600 39656 39664
rect 39720 39600 39736 39664
rect 39800 39600 39816 39664
rect 39880 39600 39896 39664
rect 39960 39600 39976 39664
rect 40040 39600 40056 39664
rect 40120 39600 40136 39664
rect 40200 39600 40216 39664
rect 40280 39600 40296 39664
rect 40360 39600 40368 39664
rect 5000 39584 40368 39600
rect 5000 39520 5008 39584
rect 5072 39520 5088 39584
rect 5152 39520 5168 39584
rect 5232 39520 5248 39584
rect 5312 39520 5328 39584
rect 5392 39520 5408 39584
rect 5472 39520 5488 39584
rect 5552 39520 5568 39584
rect 5632 39520 5648 39584
rect 5712 39520 5728 39584
rect 5792 39520 5808 39584
rect 5872 39520 5888 39584
rect 5952 39520 5968 39584
rect 6032 39520 6048 39584
rect 6112 39520 6128 39584
rect 6192 39520 6208 39584
rect 6272 39520 6288 39584
rect 6352 39520 6368 39584
rect 6432 39520 6448 39584
rect 6512 39520 6528 39584
rect 6592 39520 6608 39584
rect 6672 39520 6688 39584
rect 6752 39520 6768 39584
rect 6832 39520 6848 39584
rect 6912 39520 6928 39584
rect 6992 39520 7008 39584
rect 7072 39520 7088 39584
rect 7152 39520 7168 39584
rect 7232 39520 7248 39584
rect 7312 39520 7328 39584
rect 7392 39520 7408 39584
rect 7472 39520 7488 39584
rect 7552 39520 7568 39584
rect 7632 39520 7648 39584
rect 7712 39520 7728 39584
rect 7792 39520 7808 39584
rect 7872 39520 7888 39584
rect 7952 39520 7968 39584
rect 8032 39520 8048 39584
rect 8112 39520 8128 39584
rect 8192 39520 8208 39584
rect 8272 39520 8288 39584
rect 8352 39520 8368 39584
rect 8432 39520 8448 39584
rect 8512 39520 8528 39584
rect 8592 39520 8608 39584
rect 8672 39520 8688 39584
rect 8752 39520 8768 39584
rect 8832 39520 8848 39584
rect 8912 39520 8928 39584
rect 8992 39520 14112 39584
rect 14176 39520 14192 39584
rect 14256 39520 14272 39584
rect 14336 39520 14352 39584
rect 14416 39520 24112 39584
rect 24176 39520 24192 39584
rect 24256 39520 24272 39584
rect 24336 39520 24352 39584
rect 24416 39520 36376 39584
rect 36440 39520 36456 39584
rect 36520 39520 36536 39584
rect 36600 39520 36616 39584
rect 36680 39520 36696 39584
rect 36760 39520 36776 39584
rect 36840 39520 36856 39584
rect 36920 39520 36936 39584
rect 37000 39520 37016 39584
rect 37080 39520 37096 39584
rect 37160 39520 37176 39584
rect 37240 39520 37256 39584
rect 37320 39520 37336 39584
rect 37400 39520 37416 39584
rect 37480 39520 37496 39584
rect 37560 39520 37576 39584
rect 37640 39520 37656 39584
rect 37720 39520 37736 39584
rect 37800 39520 37816 39584
rect 37880 39520 37896 39584
rect 37960 39520 37976 39584
rect 38040 39520 38056 39584
rect 38120 39520 38136 39584
rect 38200 39520 38216 39584
rect 38280 39520 38296 39584
rect 38360 39520 38376 39584
rect 38440 39520 38456 39584
rect 38520 39520 38536 39584
rect 38600 39520 38616 39584
rect 38680 39520 38696 39584
rect 38760 39520 38776 39584
rect 38840 39520 38856 39584
rect 38920 39520 38936 39584
rect 39000 39520 39016 39584
rect 39080 39520 39096 39584
rect 39160 39520 39176 39584
rect 39240 39520 39256 39584
rect 39320 39520 39336 39584
rect 39400 39520 39416 39584
rect 39480 39520 39496 39584
rect 39560 39520 39576 39584
rect 39640 39520 39656 39584
rect 39720 39520 39736 39584
rect 39800 39520 39816 39584
rect 39880 39520 39896 39584
rect 39960 39520 39976 39584
rect 40040 39520 40056 39584
rect 40120 39520 40136 39584
rect 40200 39520 40216 39584
rect 40280 39520 40296 39584
rect 40360 39520 40368 39584
rect 5000 39504 40368 39520
rect 5000 39440 5008 39504
rect 5072 39440 5088 39504
rect 5152 39440 5168 39504
rect 5232 39440 5248 39504
rect 5312 39440 5328 39504
rect 5392 39440 5408 39504
rect 5472 39440 5488 39504
rect 5552 39440 5568 39504
rect 5632 39440 5648 39504
rect 5712 39440 5728 39504
rect 5792 39440 5808 39504
rect 5872 39440 5888 39504
rect 5952 39440 5968 39504
rect 6032 39440 6048 39504
rect 6112 39440 6128 39504
rect 6192 39440 6208 39504
rect 6272 39440 6288 39504
rect 6352 39440 6368 39504
rect 6432 39440 6448 39504
rect 6512 39440 6528 39504
rect 6592 39440 6608 39504
rect 6672 39440 6688 39504
rect 6752 39440 6768 39504
rect 6832 39440 6848 39504
rect 6912 39440 6928 39504
rect 6992 39440 7008 39504
rect 7072 39440 7088 39504
rect 7152 39440 7168 39504
rect 7232 39440 7248 39504
rect 7312 39440 7328 39504
rect 7392 39440 7408 39504
rect 7472 39440 7488 39504
rect 7552 39440 7568 39504
rect 7632 39440 7648 39504
rect 7712 39440 7728 39504
rect 7792 39440 7808 39504
rect 7872 39440 7888 39504
rect 7952 39440 7968 39504
rect 8032 39440 8048 39504
rect 8112 39440 8128 39504
rect 8192 39440 8208 39504
rect 8272 39440 8288 39504
rect 8352 39440 8368 39504
rect 8432 39440 8448 39504
rect 8512 39440 8528 39504
rect 8592 39440 8608 39504
rect 8672 39440 8688 39504
rect 8752 39440 8768 39504
rect 8832 39440 8848 39504
rect 8912 39440 8928 39504
rect 8992 39440 14112 39504
rect 14176 39440 14192 39504
rect 14256 39440 14272 39504
rect 14336 39440 14352 39504
rect 14416 39440 24112 39504
rect 24176 39440 24192 39504
rect 24256 39440 24272 39504
rect 24336 39440 24352 39504
rect 24416 39440 36376 39504
rect 36440 39440 36456 39504
rect 36520 39440 36536 39504
rect 36600 39440 36616 39504
rect 36680 39440 36696 39504
rect 36760 39440 36776 39504
rect 36840 39440 36856 39504
rect 36920 39440 36936 39504
rect 37000 39440 37016 39504
rect 37080 39440 37096 39504
rect 37160 39440 37176 39504
rect 37240 39440 37256 39504
rect 37320 39440 37336 39504
rect 37400 39440 37416 39504
rect 37480 39440 37496 39504
rect 37560 39440 37576 39504
rect 37640 39440 37656 39504
rect 37720 39440 37736 39504
rect 37800 39440 37816 39504
rect 37880 39440 37896 39504
rect 37960 39440 37976 39504
rect 38040 39440 38056 39504
rect 38120 39440 38136 39504
rect 38200 39440 38216 39504
rect 38280 39440 38296 39504
rect 38360 39440 38376 39504
rect 38440 39440 38456 39504
rect 38520 39440 38536 39504
rect 38600 39440 38616 39504
rect 38680 39440 38696 39504
rect 38760 39440 38776 39504
rect 38840 39440 38856 39504
rect 38920 39440 38936 39504
rect 39000 39440 39016 39504
rect 39080 39440 39096 39504
rect 39160 39440 39176 39504
rect 39240 39440 39256 39504
rect 39320 39440 39336 39504
rect 39400 39440 39416 39504
rect 39480 39440 39496 39504
rect 39560 39440 39576 39504
rect 39640 39440 39656 39504
rect 39720 39440 39736 39504
rect 39800 39440 39816 39504
rect 39880 39440 39896 39504
rect 39960 39440 39976 39504
rect 40040 39440 40056 39504
rect 40120 39440 40136 39504
rect 40200 39440 40216 39504
rect 40280 39440 40296 39504
rect 40360 39440 40368 39504
rect 5000 39424 40368 39440
rect 5000 39360 5008 39424
rect 5072 39360 5088 39424
rect 5152 39360 5168 39424
rect 5232 39360 5248 39424
rect 5312 39360 5328 39424
rect 5392 39360 5408 39424
rect 5472 39360 5488 39424
rect 5552 39360 5568 39424
rect 5632 39360 5648 39424
rect 5712 39360 5728 39424
rect 5792 39360 5808 39424
rect 5872 39360 5888 39424
rect 5952 39360 5968 39424
rect 6032 39360 6048 39424
rect 6112 39360 6128 39424
rect 6192 39360 6208 39424
rect 6272 39360 6288 39424
rect 6352 39360 6368 39424
rect 6432 39360 6448 39424
rect 6512 39360 6528 39424
rect 6592 39360 6608 39424
rect 6672 39360 6688 39424
rect 6752 39360 6768 39424
rect 6832 39360 6848 39424
rect 6912 39360 6928 39424
rect 6992 39360 7008 39424
rect 7072 39360 7088 39424
rect 7152 39360 7168 39424
rect 7232 39360 7248 39424
rect 7312 39360 7328 39424
rect 7392 39360 7408 39424
rect 7472 39360 7488 39424
rect 7552 39360 7568 39424
rect 7632 39360 7648 39424
rect 7712 39360 7728 39424
rect 7792 39360 7808 39424
rect 7872 39360 7888 39424
rect 7952 39360 7968 39424
rect 8032 39360 8048 39424
rect 8112 39360 8128 39424
rect 8192 39360 8208 39424
rect 8272 39360 8288 39424
rect 8352 39360 8368 39424
rect 8432 39360 8448 39424
rect 8512 39360 8528 39424
rect 8592 39360 8608 39424
rect 8672 39360 8688 39424
rect 8752 39360 8768 39424
rect 8832 39360 8848 39424
rect 8912 39360 8928 39424
rect 8992 39360 14112 39424
rect 14176 39360 14192 39424
rect 14256 39360 14272 39424
rect 14336 39360 14352 39424
rect 14416 39360 24112 39424
rect 24176 39360 24192 39424
rect 24256 39360 24272 39424
rect 24336 39360 24352 39424
rect 24416 39360 36376 39424
rect 36440 39360 36456 39424
rect 36520 39360 36536 39424
rect 36600 39360 36616 39424
rect 36680 39360 36696 39424
rect 36760 39360 36776 39424
rect 36840 39360 36856 39424
rect 36920 39360 36936 39424
rect 37000 39360 37016 39424
rect 37080 39360 37096 39424
rect 37160 39360 37176 39424
rect 37240 39360 37256 39424
rect 37320 39360 37336 39424
rect 37400 39360 37416 39424
rect 37480 39360 37496 39424
rect 37560 39360 37576 39424
rect 37640 39360 37656 39424
rect 37720 39360 37736 39424
rect 37800 39360 37816 39424
rect 37880 39360 37896 39424
rect 37960 39360 37976 39424
rect 38040 39360 38056 39424
rect 38120 39360 38136 39424
rect 38200 39360 38216 39424
rect 38280 39360 38296 39424
rect 38360 39360 38376 39424
rect 38440 39360 38456 39424
rect 38520 39360 38536 39424
rect 38600 39360 38616 39424
rect 38680 39360 38696 39424
rect 38760 39360 38776 39424
rect 38840 39360 38856 39424
rect 38920 39360 38936 39424
rect 39000 39360 39016 39424
rect 39080 39360 39096 39424
rect 39160 39360 39176 39424
rect 39240 39360 39256 39424
rect 39320 39360 39336 39424
rect 39400 39360 39416 39424
rect 39480 39360 39496 39424
rect 39560 39360 39576 39424
rect 39640 39360 39656 39424
rect 39720 39360 39736 39424
rect 39800 39360 39816 39424
rect 39880 39360 39896 39424
rect 39960 39360 39976 39424
rect 40040 39360 40056 39424
rect 40120 39360 40136 39424
rect 40200 39360 40216 39424
rect 40280 39360 40296 39424
rect 40360 39360 40368 39424
rect 5000 39344 40368 39360
rect 5000 39280 5008 39344
rect 5072 39280 5088 39344
rect 5152 39280 5168 39344
rect 5232 39280 5248 39344
rect 5312 39280 5328 39344
rect 5392 39280 5408 39344
rect 5472 39280 5488 39344
rect 5552 39280 5568 39344
rect 5632 39280 5648 39344
rect 5712 39280 5728 39344
rect 5792 39280 5808 39344
rect 5872 39280 5888 39344
rect 5952 39280 5968 39344
rect 6032 39280 6048 39344
rect 6112 39280 6128 39344
rect 6192 39280 6208 39344
rect 6272 39280 6288 39344
rect 6352 39280 6368 39344
rect 6432 39280 6448 39344
rect 6512 39280 6528 39344
rect 6592 39280 6608 39344
rect 6672 39280 6688 39344
rect 6752 39280 6768 39344
rect 6832 39280 6848 39344
rect 6912 39280 6928 39344
rect 6992 39280 7008 39344
rect 7072 39280 7088 39344
rect 7152 39280 7168 39344
rect 7232 39280 7248 39344
rect 7312 39280 7328 39344
rect 7392 39280 7408 39344
rect 7472 39280 7488 39344
rect 7552 39280 7568 39344
rect 7632 39280 7648 39344
rect 7712 39280 7728 39344
rect 7792 39280 7808 39344
rect 7872 39280 7888 39344
rect 7952 39280 7968 39344
rect 8032 39280 8048 39344
rect 8112 39280 8128 39344
rect 8192 39280 8208 39344
rect 8272 39280 8288 39344
rect 8352 39280 8368 39344
rect 8432 39280 8448 39344
rect 8512 39280 8528 39344
rect 8592 39280 8608 39344
rect 8672 39280 8688 39344
rect 8752 39280 8768 39344
rect 8832 39280 8848 39344
rect 8912 39280 8928 39344
rect 8992 39280 14112 39344
rect 14176 39280 14192 39344
rect 14256 39280 14272 39344
rect 14336 39280 14352 39344
rect 14416 39280 24112 39344
rect 24176 39280 24192 39344
rect 24256 39280 24272 39344
rect 24336 39280 24352 39344
rect 24416 39280 36376 39344
rect 36440 39280 36456 39344
rect 36520 39280 36536 39344
rect 36600 39280 36616 39344
rect 36680 39280 36696 39344
rect 36760 39280 36776 39344
rect 36840 39280 36856 39344
rect 36920 39280 36936 39344
rect 37000 39280 37016 39344
rect 37080 39280 37096 39344
rect 37160 39280 37176 39344
rect 37240 39280 37256 39344
rect 37320 39280 37336 39344
rect 37400 39280 37416 39344
rect 37480 39280 37496 39344
rect 37560 39280 37576 39344
rect 37640 39280 37656 39344
rect 37720 39280 37736 39344
rect 37800 39280 37816 39344
rect 37880 39280 37896 39344
rect 37960 39280 37976 39344
rect 38040 39280 38056 39344
rect 38120 39280 38136 39344
rect 38200 39280 38216 39344
rect 38280 39280 38296 39344
rect 38360 39280 38376 39344
rect 38440 39280 38456 39344
rect 38520 39280 38536 39344
rect 38600 39280 38616 39344
rect 38680 39280 38696 39344
rect 38760 39280 38776 39344
rect 38840 39280 38856 39344
rect 38920 39280 38936 39344
rect 39000 39280 39016 39344
rect 39080 39280 39096 39344
rect 39160 39280 39176 39344
rect 39240 39280 39256 39344
rect 39320 39280 39336 39344
rect 39400 39280 39416 39344
rect 39480 39280 39496 39344
rect 39560 39280 39576 39344
rect 39640 39280 39656 39344
rect 39720 39280 39736 39344
rect 39800 39280 39816 39344
rect 39880 39280 39896 39344
rect 39960 39280 39976 39344
rect 40040 39280 40056 39344
rect 40120 39280 40136 39344
rect 40200 39280 40216 39344
rect 40280 39280 40296 39344
rect 40360 39280 40368 39344
rect 5000 39264 40368 39280
rect 5000 39200 5008 39264
rect 5072 39200 5088 39264
rect 5152 39200 5168 39264
rect 5232 39200 5248 39264
rect 5312 39200 5328 39264
rect 5392 39200 5408 39264
rect 5472 39200 5488 39264
rect 5552 39200 5568 39264
rect 5632 39200 5648 39264
rect 5712 39200 5728 39264
rect 5792 39200 5808 39264
rect 5872 39200 5888 39264
rect 5952 39200 5968 39264
rect 6032 39200 6048 39264
rect 6112 39200 6128 39264
rect 6192 39200 6208 39264
rect 6272 39200 6288 39264
rect 6352 39200 6368 39264
rect 6432 39200 6448 39264
rect 6512 39200 6528 39264
rect 6592 39200 6608 39264
rect 6672 39200 6688 39264
rect 6752 39200 6768 39264
rect 6832 39200 6848 39264
rect 6912 39200 6928 39264
rect 6992 39200 7008 39264
rect 7072 39200 7088 39264
rect 7152 39200 7168 39264
rect 7232 39200 7248 39264
rect 7312 39200 7328 39264
rect 7392 39200 7408 39264
rect 7472 39200 7488 39264
rect 7552 39200 7568 39264
rect 7632 39200 7648 39264
rect 7712 39200 7728 39264
rect 7792 39200 7808 39264
rect 7872 39200 7888 39264
rect 7952 39200 7968 39264
rect 8032 39200 8048 39264
rect 8112 39200 8128 39264
rect 8192 39200 8208 39264
rect 8272 39200 8288 39264
rect 8352 39200 8368 39264
rect 8432 39200 8448 39264
rect 8512 39200 8528 39264
rect 8592 39200 8608 39264
rect 8672 39200 8688 39264
rect 8752 39200 8768 39264
rect 8832 39200 8848 39264
rect 8912 39200 8928 39264
rect 8992 39200 14112 39264
rect 14176 39200 14192 39264
rect 14256 39200 14272 39264
rect 14336 39200 14352 39264
rect 14416 39200 24112 39264
rect 24176 39200 24192 39264
rect 24256 39200 24272 39264
rect 24336 39200 24352 39264
rect 24416 39200 36376 39264
rect 36440 39200 36456 39264
rect 36520 39200 36536 39264
rect 36600 39200 36616 39264
rect 36680 39200 36696 39264
rect 36760 39200 36776 39264
rect 36840 39200 36856 39264
rect 36920 39200 36936 39264
rect 37000 39200 37016 39264
rect 37080 39200 37096 39264
rect 37160 39200 37176 39264
rect 37240 39200 37256 39264
rect 37320 39200 37336 39264
rect 37400 39200 37416 39264
rect 37480 39200 37496 39264
rect 37560 39200 37576 39264
rect 37640 39200 37656 39264
rect 37720 39200 37736 39264
rect 37800 39200 37816 39264
rect 37880 39200 37896 39264
rect 37960 39200 37976 39264
rect 38040 39200 38056 39264
rect 38120 39200 38136 39264
rect 38200 39200 38216 39264
rect 38280 39200 38296 39264
rect 38360 39200 38376 39264
rect 38440 39200 38456 39264
rect 38520 39200 38536 39264
rect 38600 39200 38616 39264
rect 38680 39200 38696 39264
rect 38760 39200 38776 39264
rect 38840 39200 38856 39264
rect 38920 39200 38936 39264
rect 39000 39200 39016 39264
rect 39080 39200 39096 39264
rect 39160 39200 39176 39264
rect 39240 39200 39256 39264
rect 39320 39200 39336 39264
rect 39400 39200 39416 39264
rect 39480 39200 39496 39264
rect 39560 39200 39576 39264
rect 39640 39200 39656 39264
rect 39720 39200 39736 39264
rect 39800 39200 39816 39264
rect 39880 39200 39896 39264
rect 39960 39200 39976 39264
rect 40040 39200 40056 39264
rect 40120 39200 40136 39264
rect 40200 39200 40216 39264
rect 40280 39200 40296 39264
rect 40360 39200 40368 39264
rect 5000 39184 40368 39200
rect 5000 39120 5008 39184
rect 5072 39120 5088 39184
rect 5152 39120 5168 39184
rect 5232 39120 5248 39184
rect 5312 39120 5328 39184
rect 5392 39120 5408 39184
rect 5472 39120 5488 39184
rect 5552 39120 5568 39184
rect 5632 39120 5648 39184
rect 5712 39120 5728 39184
rect 5792 39120 5808 39184
rect 5872 39120 5888 39184
rect 5952 39120 5968 39184
rect 6032 39120 6048 39184
rect 6112 39120 6128 39184
rect 6192 39120 6208 39184
rect 6272 39120 6288 39184
rect 6352 39120 6368 39184
rect 6432 39120 6448 39184
rect 6512 39120 6528 39184
rect 6592 39120 6608 39184
rect 6672 39120 6688 39184
rect 6752 39120 6768 39184
rect 6832 39120 6848 39184
rect 6912 39120 6928 39184
rect 6992 39120 7008 39184
rect 7072 39120 7088 39184
rect 7152 39120 7168 39184
rect 7232 39120 7248 39184
rect 7312 39120 7328 39184
rect 7392 39120 7408 39184
rect 7472 39120 7488 39184
rect 7552 39120 7568 39184
rect 7632 39120 7648 39184
rect 7712 39120 7728 39184
rect 7792 39120 7808 39184
rect 7872 39120 7888 39184
rect 7952 39120 7968 39184
rect 8032 39120 8048 39184
rect 8112 39120 8128 39184
rect 8192 39120 8208 39184
rect 8272 39120 8288 39184
rect 8352 39120 8368 39184
rect 8432 39120 8448 39184
rect 8512 39120 8528 39184
rect 8592 39120 8608 39184
rect 8672 39120 8688 39184
rect 8752 39120 8768 39184
rect 8832 39120 8848 39184
rect 8912 39120 8928 39184
rect 8992 39120 14112 39184
rect 14176 39120 14192 39184
rect 14256 39120 14272 39184
rect 14336 39120 14352 39184
rect 14416 39120 24112 39184
rect 24176 39120 24192 39184
rect 24256 39120 24272 39184
rect 24336 39120 24352 39184
rect 24416 39120 36376 39184
rect 36440 39120 36456 39184
rect 36520 39120 36536 39184
rect 36600 39120 36616 39184
rect 36680 39120 36696 39184
rect 36760 39120 36776 39184
rect 36840 39120 36856 39184
rect 36920 39120 36936 39184
rect 37000 39120 37016 39184
rect 37080 39120 37096 39184
rect 37160 39120 37176 39184
rect 37240 39120 37256 39184
rect 37320 39120 37336 39184
rect 37400 39120 37416 39184
rect 37480 39120 37496 39184
rect 37560 39120 37576 39184
rect 37640 39120 37656 39184
rect 37720 39120 37736 39184
rect 37800 39120 37816 39184
rect 37880 39120 37896 39184
rect 37960 39120 37976 39184
rect 38040 39120 38056 39184
rect 38120 39120 38136 39184
rect 38200 39120 38216 39184
rect 38280 39120 38296 39184
rect 38360 39120 38376 39184
rect 38440 39120 38456 39184
rect 38520 39120 38536 39184
rect 38600 39120 38616 39184
rect 38680 39120 38696 39184
rect 38760 39120 38776 39184
rect 38840 39120 38856 39184
rect 38920 39120 38936 39184
rect 39000 39120 39016 39184
rect 39080 39120 39096 39184
rect 39160 39120 39176 39184
rect 39240 39120 39256 39184
rect 39320 39120 39336 39184
rect 39400 39120 39416 39184
rect 39480 39120 39496 39184
rect 39560 39120 39576 39184
rect 39640 39120 39656 39184
rect 39720 39120 39736 39184
rect 39800 39120 39816 39184
rect 39880 39120 39896 39184
rect 39960 39120 39976 39184
rect 40040 39120 40056 39184
rect 40120 39120 40136 39184
rect 40200 39120 40216 39184
rect 40280 39120 40296 39184
rect 40360 39120 40368 39184
rect 5000 39104 40368 39120
rect 5000 39040 5008 39104
rect 5072 39040 5088 39104
rect 5152 39040 5168 39104
rect 5232 39040 5248 39104
rect 5312 39040 5328 39104
rect 5392 39040 5408 39104
rect 5472 39040 5488 39104
rect 5552 39040 5568 39104
rect 5632 39040 5648 39104
rect 5712 39040 5728 39104
rect 5792 39040 5808 39104
rect 5872 39040 5888 39104
rect 5952 39040 5968 39104
rect 6032 39040 6048 39104
rect 6112 39040 6128 39104
rect 6192 39040 6208 39104
rect 6272 39040 6288 39104
rect 6352 39040 6368 39104
rect 6432 39040 6448 39104
rect 6512 39040 6528 39104
rect 6592 39040 6608 39104
rect 6672 39040 6688 39104
rect 6752 39040 6768 39104
rect 6832 39040 6848 39104
rect 6912 39040 6928 39104
rect 6992 39040 7008 39104
rect 7072 39040 7088 39104
rect 7152 39040 7168 39104
rect 7232 39040 7248 39104
rect 7312 39040 7328 39104
rect 7392 39040 7408 39104
rect 7472 39040 7488 39104
rect 7552 39040 7568 39104
rect 7632 39040 7648 39104
rect 7712 39040 7728 39104
rect 7792 39040 7808 39104
rect 7872 39040 7888 39104
rect 7952 39040 7968 39104
rect 8032 39040 8048 39104
rect 8112 39040 8128 39104
rect 8192 39040 8208 39104
rect 8272 39040 8288 39104
rect 8352 39040 8368 39104
rect 8432 39040 8448 39104
rect 8512 39040 8528 39104
rect 8592 39040 8608 39104
rect 8672 39040 8688 39104
rect 8752 39040 8768 39104
rect 8832 39040 8848 39104
rect 8912 39040 8928 39104
rect 8992 39040 14112 39104
rect 14176 39040 14192 39104
rect 14256 39040 14272 39104
rect 14336 39040 14352 39104
rect 14416 39040 24112 39104
rect 24176 39040 24192 39104
rect 24256 39040 24272 39104
rect 24336 39040 24352 39104
rect 24416 39040 36376 39104
rect 36440 39040 36456 39104
rect 36520 39040 36536 39104
rect 36600 39040 36616 39104
rect 36680 39040 36696 39104
rect 36760 39040 36776 39104
rect 36840 39040 36856 39104
rect 36920 39040 36936 39104
rect 37000 39040 37016 39104
rect 37080 39040 37096 39104
rect 37160 39040 37176 39104
rect 37240 39040 37256 39104
rect 37320 39040 37336 39104
rect 37400 39040 37416 39104
rect 37480 39040 37496 39104
rect 37560 39040 37576 39104
rect 37640 39040 37656 39104
rect 37720 39040 37736 39104
rect 37800 39040 37816 39104
rect 37880 39040 37896 39104
rect 37960 39040 37976 39104
rect 38040 39040 38056 39104
rect 38120 39040 38136 39104
rect 38200 39040 38216 39104
rect 38280 39040 38296 39104
rect 38360 39040 38376 39104
rect 38440 39040 38456 39104
rect 38520 39040 38536 39104
rect 38600 39040 38616 39104
rect 38680 39040 38696 39104
rect 38760 39040 38776 39104
rect 38840 39040 38856 39104
rect 38920 39040 38936 39104
rect 39000 39040 39016 39104
rect 39080 39040 39096 39104
rect 39160 39040 39176 39104
rect 39240 39040 39256 39104
rect 39320 39040 39336 39104
rect 39400 39040 39416 39104
rect 39480 39040 39496 39104
rect 39560 39040 39576 39104
rect 39640 39040 39656 39104
rect 39720 39040 39736 39104
rect 39800 39040 39816 39104
rect 39880 39040 39896 39104
rect 39960 39040 39976 39104
rect 40040 39040 40056 39104
rect 40120 39040 40136 39104
rect 40200 39040 40216 39104
rect 40280 39040 40296 39104
rect 40360 39040 40368 39104
rect 5000 39024 40368 39040
rect 5000 38960 5008 39024
rect 5072 38960 5088 39024
rect 5152 38960 5168 39024
rect 5232 38960 5248 39024
rect 5312 38960 5328 39024
rect 5392 38960 5408 39024
rect 5472 38960 5488 39024
rect 5552 38960 5568 39024
rect 5632 38960 5648 39024
rect 5712 38960 5728 39024
rect 5792 38960 5808 39024
rect 5872 38960 5888 39024
rect 5952 38960 5968 39024
rect 6032 38960 6048 39024
rect 6112 38960 6128 39024
rect 6192 38960 6208 39024
rect 6272 38960 6288 39024
rect 6352 38960 6368 39024
rect 6432 38960 6448 39024
rect 6512 38960 6528 39024
rect 6592 38960 6608 39024
rect 6672 38960 6688 39024
rect 6752 38960 6768 39024
rect 6832 38960 6848 39024
rect 6912 38960 6928 39024
rect 6992 38960 7008 39024
rect 7072 38960 7088 39024
rect 7152 38960 7168 39024
rect 7232 38960 7248 39024
rect 7312 38960 7328 39024
rect 7392 38960 7408 39024
rect 7472 38960 7488 39024
rect 7552 38960 7568 39024
rect 7632 38960 7648 39024
rect 7712 38960 7728 39024
rect 7792 38960 7808 39024
rect 7872 38960 7888 39024
rect 7952 38960 7968 39024
rect 8032 38960 8048 39024
rect 8112 38960 8128 39024
rect 8192 38960 8208 39024
rect 8272 38960 8288 39024
rect 8352 38960 8368 39024
rect 8432 38960 8448 39024
rect 8512 38960 8528 39024
rect 8592 38960 8608 39024
rect 8672 38960 8688 39024
rect 8752 38960 8768 39024
rect 8832 38960 8848 39024
rect 8912 38960 8928 39024
rect 8992 38960 14112 39024
rect 14176 38960 14192 39024
rect 14256 38960 14272 39024
rect 14336 38960 14352 39024
rect 14416 38960 24112 39024
rect 24176 38960 24192 39024
rect 24256 38960 24272 39024
rect 24336 38960 24352 39024
rect 24416 38960 36376 39024
rect 36440 38960 36456 39024
rect 36520 38960 36536 39024
rect 36600 38960 36616 39024
rect 36680 38960 36696 39024
rect 36760 38960 36776 39024
rect 36840 38960 36856 39024
rect 36920 38960 36936 39024
rect 37000 38960 37016 39024
rect 37080 38960 37096 39024
rect 37160 38960 37176 39024
rect 37240 38960 37256 39024
rect 37320 38960 37336 39024
rect 37400 38960 37416 39024
rect 37480 38960 37496 39024
rect 37560 38960 37576 39024
rect 37640 38960 37656 39024
rect 37720 38960 37736 39024
rect 37800 38960 37816 39024
rect 37880 38960 37896 39024
rect 37960 38960 37976 39024
rect 38040 38960 38056 39024
rect 38120 38960 38136 39024
rect 38200 38960 38216 39024
rect 38280 38960 38296 39024
rect 38360 38960 38376 39024
rect 38440 38960 38456 39024
rect 38520 38960 38536 39024
rect 38600 38960 38616 39024
rect 38680 38960 38696 39024
rect 38760 38960 38776 39024
rect 38840 38960 38856 39024
rect 38920 38960 38936 39024
rect 39000 38960 39016 39024
rect 39080 38960 39096 39024
rect 39160 38960 39176 39024
rect 39240 38960 39256 39024
rect 39320 38960 39336 39024
rect 39400 38960 39416 39024
rect 39480 38960 39496 39024
rect 39560 38960 39576 39024
rect 39640 38960 39656 39024
rect 39720 38960 39736 39024
rect 39800 38960 39816 39024
rect 39880 38960 39896 39024
rect 39960 38960 39976 39024
rect 40040 38960 40056 39024
rect 40120 38960 40136 39024
rect 40200 38960 40216 39024
rect 40280 38960 40296 39024
rect 40360 38960 40368 39024
rect 5000 38944 40368 38960
rect 5000 38880 5008 38944
rect 5072 38880 5088 38944
rect 5152 38880 5168 38944
rect 5232 38880 5248 38944
rect 5312 38880 5328 38944
rect 5392 38880 5408 38944
rect 5472 38880 5488 38944
rect 5552 38880 5568 38944
rect 5632 38880 5648 38944
rect 5712 38880 5728 38944
rect 5792 38880 5808 38944
rect 5872 38880 5888 38944
rect 5952 38880 5968 38944
rect 6032 38880 6048 38944
rect 6112 38880 6128 38944
rect 6192 38880 6208 38944
rect 6272 38880 6288 38944
rect 6352 38880 6368 38944
rect 6432 38880 6448 38944
rect 6512 38880 6528 38944
rect 6592 38880 6608 38944
rect 6672 38880 6688 38944
rect 6752 38880 6768 38944
rect 6832 38880 6848 38944
rect 6912 38880 6928 38944
rect 6992 38880 7008 38944
rect 7072 38880 7088 38944
rect 7152 38880 7168 38944
rect 7232 38880 7248 38944
rect 7312 38880 7328 38944
rect 7392 38880 7408 38944
rect 7472 38880 7488 38944
rect 7552 38880 7568 38944
rect 7632 38880 7648 38944
rect 7712 38880 7728 38944
rect 7792 38880 7808 38944
rect 7872 38880 7888 38944
rect 7952 38880 7968 38944
rect 8032 38880 8048 38944
rect 8112 38880 8128 38944
rect 8192 38880 8208 38944
rect 8272 38880 8288 38944
rect 8352 38880 8368 38944
rect 8432 38880 8448 38944
rect 8512 38880 8528 38944
rect 8592 38880 8608 38944
rect 8672 38880 8688 38944
rect 8752 38880 8768 38944
rect 8832 38880 8848 38944
rect 8912 38880 8928 38944
rect 8992 38880 14112 38944
rect 14176 38880 14192 38944
rect 14256 38880 14272 38944
rect 14336 38880 14352 38944
rect 14416 38880 24112 38944
rect 24176 38880 24192 38944
rect 24256 38880 24272 38944
rect 24336 38880 24352 38944
rect 24416 38880 36376 38944
rect 36440 38880 36456 38944
rect 36520 38880 36536 38944
rect 36600 38880 36616 38944
rect 36680 38880 36696 38944
rect 36760 38880 36776 38944
rect 36840 38880 36856 38944
rect 36920 38880 36936 38944
rect 37000 38880 37016 38944
rect 37080 38880 37096 38944
rect 37160 38880 37176 38944
rect 37240 38880 37256 38944
rect 37320 38880 37336 38944
rect 37400 38880 37416 38944
rect 37480 38880 37496 38944
rect 37560 38880 37576 38944
rect 37640 38880 37656 38944
rect 37720 38880 37736 38944
rect 37800 38880 37816 38944
rect 37880 38880 37896 38944
rect 37960 38880 37976 38944
rect 38040 38880 38056 38944
rect 38120 38880 38136 38944
rect 38200 38880 38216 38944
rect 38280 38880 38296 38944
rect 38360 38880 38376 38944
rect 38440 38880 38456 38944
rect 38520 38880 38536 38944
rect 38600 38880 38616 38944
rect 38680 38880 38696 38944
rect 38760 38880 38776 38944
rect 38840 38880 38856 38944
rect 38920 38880 38936 38944
rect 39000 38880 39016 38944
rect 39080 38880 39096 38944
rect 39160 38880 39176 38944
rect 39240 38880 39256 38944
rect 39320 38880 39336 38944
rect 39400 38880 39416 38944
rect 39480 38880 39496 38944
rect 39560 38880 39576 38944
rect 39640 38880 39656 38944
rect 39720 38880 39736 38944
rect 39800 38880 39816 38944
rect 39880 38880 39896 38944
rect 39960 38880 39976 38944
rect 40040 38880 40056 38944
rect 40120 38880 40136 38944
rect 40200 38880 40216 38944
rect 40280 38880 40296 38944
rect 40360 38880 40368 38944
rect 5000 38864 40368 38880
rect 5000 38800 5008 38864
rect 5072 38800 5088 38864
rect 5152 38800 5168 38864
rect 5232 38800 5248 38864
rect 5312 38800 5328 38864
rect 5392 38800 5408 38864
rect 5472 38800 5488 38864
rect 5552 38800 5568 38864
rect 5632 38800 5648 38864
rect 5712 38800 5728 38864
rect 5792 38800 5808 38864
rect 5872 38800 5888 38864
rect 5952 38800 5968 38864
rect 6032 38800 6048 38864
rect 6112 38800 6128 38864
rect 6192 38800 6208 38864
rect 6272 38800 6288 38864
rect 6352 38800 6368 38864
rect 6432 38800 6448 38864
rect 6512 38800 6528 38864
rect 6592 38800 6608 38864
rect 6672 38800 6688 38864
rect 6752 38800 6768 38864
rect 6832 38800 6848 38864
rect 6912 38800 6928 38864
rect 6992 38800 7008 38864
rect 7072 38800 7088 38864
rect 7152 38800 7168 38864
rect 7232 38800 7248 38864
rect 7312 38800 7328 38864
rect 7392 38800 7408 38864
rect 7472 38800 7488 38864
rect 7552 38800 7568 38864
rect 7632 38800 7648 38864
rect 7712 38800 7728 38864
rect 7792 38800 7808 38864
rect 7872 38800 7888 38864
rect 7952 38800 7968 38864
rect 8032 38800 8048 38864
rect 8112 38800 8128 38864
rect 8192 38800 8208 38864
rect 8272 38800 8288 38864
rect 8352 38800 8368 38864
rect 8432 38800 8448 38864
rect 8512 38800 8528 38864
rect 8592 38800 8608 38864
rect 8672 38800 8688 38864
rect 8752 38800 8768 38864
rect 8832 38800 8848 38864
rect 8912 38800 8928 38864
rect 8992 38800 14112 38864
rect 14176 38800 14192 38864
rect 14256 38800 14272 38864
rect 14336 38800 14352 38864
rect 14416 38800 24112 38864
rect 24176 38800 24192 38864
rect 24256 38800 24272 38864
rect 24336 38800 24352 38864
rect 24416 38800 36376 38864
rect 36440 38800 36456 38864
rect 36520 38800 36536 38864
rect 36600 38800 36616 38864
rect 36680 38800 36696 38864
rect 36760 38800 36776 38864
rect 36840 38800 36856 38864
rect 36920 38800 36936 38864
rect 37000 38800 37016 38864
rect 37080 38800 37096 38864
rect 37160 38800 37176 38864
rect 37240 38800 37256 38864
rect 37320 38800 37336 38864
rect 37400 38800 37416 38864
rect 37480 38800 37496 38864
rect 37560 38800 37576 38864
rect 37640 38800 37656 38864
rect 37720 38800 37736 38864
rect 37800 38800 37816 38864
rect 37880 38800 37896 38864
rect 37960 38800 37976 38864
rect 38040 38800 38056 38864
rect 38120 38800 38136 38864
rect 38200 38800 38216 38864
rect 38280 38800 38296 38864
rect 38360 38800 38376 38864
rect 38440 38800 38456 38864
rect 38520 38800 38536 38864
rect 38600 38800 38616 38864
rect 38680 38800 38696 38864
rect 38760 38800 38776 38864
rect 38840 38800 38856 38864
rect 38920 38800 38936 38864
rect 39000 38800 39016 38864
rect 39080 38800 39096 38864
rect 39160 38800 39176 38864
rect 39240 38800 39256 38864
rect 39320 38800 39336 38864
rect 39400 38800 39416 38864
rect 39480 38800 39496 38864
rect 39560 38800 39576 38864
rect 39640 38800 39656 38864
rect 39720 38800 39736 38864
rect 39800 38800 39816 38864
rect 39880 38800 39896 38864
rect 39960 38800 39976 38864
rect 40040 38800 40056 38864
rect 40120 38800 40136 38864
rect 40200 38800 40216 38864
rect 40280 38800 40296 38864
rect 40360 38800 40368 38864
rect 5000 38784 40368 38800
rect 5000 38720 5008 38784
rect 5072 38720 5088 38784
rect 5152 38720 5168 38784
rect 5232 38720 5248 38784
rect 5312 38720 5328 38784
rect 5392 38720 5408 38784
rect 5472 38720 5488 38784
rect 5552 38720 5568 38784
rect 5632 38720 5648 38784
rect 5712 38720 5728 38784
rect 5792 38720 5808 38784
rect 5872 38720 5888 38784
rect 5952 38720 5968 38784
rect 6032 38720 6048 38784
rect 6112 38720 6128 38784
rect 6192 38720 6208 38784
rect 6272 38720 6288 38784
rect 6352 38720 6368 38784
rect 6432 38720 6448 38784
rect 6512 38720 6528 38784
rect 6592 38720 6608 38784
rect 6672 38720 6688 38784
rect 6752 38720 6768 38784
rect 6832 38720 6848 38784
rect 6912 38720 6928 38784
rect 6992 38720 7008 38784
rect 7072 38720 7088 38784
rect 7152 38720 7168 38784
rect 7232 38720 7248 38784
rect 7312 38720 7328 38784
rect 7392 38720 7408 38784
rect 7472 38720 7488 38784
rect 7552 38720 7568 38784
rect 7632 38720 7648 38784
rect 7712 38720 7728 38784
rect 7792 38720 7808 38784
rect 7872 38720 7888 38784
rect 7952 38720 7968 38784
rect 8032 38720 8048 38784
rect 8112 38720 8128 38784
rect 8192 38720 8208 38784
rect 8272 38720 8288 38784
rect 8352 38720 8368 38784
rect 8432 38720 8448 38784
rect 8512 38720 8528 38784
rect 8592 38720 8608 38784
rect 8672 38720 8688 38784
rect 8752 38720 8768 38784
rect 8832 38720 8848 38784
rect 8912 38720 8928 38784
rect 8992 38720 14112 38784
rect 14176 38720 14192 38784
rect 14256 38720 14272 38784
rect 14336 38720 14352 38784
rect 14416 38720 24112 38784
rect 24176 38720 24192 38784
rect 24256 38720 24272 38784
rect 24336 38720 24352 38784
rect 24416 38720 36376 38784
rect 36440 38720 36456 38784
rect 36520 38720 36536 38784
rect 36600 38720 36616 38784
rect 36680 38720 36696 38784
rect 36760 38720 36776 38784
rect 36840 38720 36856 38784
rect 36920 38720 36936 38784
rect 37000 38720 37016 38784
rect 37080 38720 37096 38784
rect 37160 38720 37176 38784
rect 37240 38720 37256 38784
rect 37320 38720 37336 38784
rect 37400 38720 37416 38784
rect 37480 38720 37496 38784
rect 37560 38720 37576 38784
rect 37640 38720 37656 38784
rect 37720 38720 37736 38784
rect 37800 38720 37816 38784
rect 37880 38720 37896 38784
rect 37960 38720 37976 38784
rect 38040 38720 38056 38784
rect 38120 38720 38136 38784
rect 38200 38720 38216 38784
rect 38280 38720 38296 38784
rect 38360 38720 38376 38784
rect 38440 38720 38456 38784
rect 38520 38720 38536 38784
rect 38600 38720 38616 38784
rect 38680 38720 38696 38784
rect 38760 38720 38776 38784
rect 38840 38720 38856 38784
rect 38920 38720 38936 38784
rect 39000 38720 39016 38784
rect 39080 38720 39096 38784
rect 39160 38720 39176 38784
rect 39240 38720 39256 38784
rect 39320 38720 39336 38784
rect 39400 38720 39416 38784
rect 39480 38720 39496 38784
rect 39560 38720 39576 38784
rect 39640 38720 39656 38784
rect 39720 38720 39736 38784
rect 39800 38720 39816 38784
rect 39880 38720 39896 38784
rect 39960 38720 39976 38784
rect 40040 38720 40056 38784
rect 40120 38720 40136 38784
rect 40200 38720 40216 38784
rect 40280 38720 40296 38784
rect 40360 38720 40368 38784
rect 5000 38704 40368 38720
rect 5000 38640 5008 38704
rect 5072 38640 5088 38704
rect 5152 38640 5168 38704
rect 5232 38640 5248 38704
rect 5312 38640 5328 38704
rect 5392 38640 5408 38704
rect 5472 38640 5488 38704
rect 5552 38640 5568 38704
rect 5632 38640 5648 38704
rect 5712 38640 5728 38704
rect 5792 38640 5808 38704
rect 5872 38640 5888 38704
rect 5952 38640 5968 38704
rect 6032 38640 6048 38704
rect 6112 38640 6128 38704
rect 6192 38640 6208 38704
rect 6272 38640 6288 38704
rect 6352 38640 6368 38704
rect 6432 38640 6448 38704
rect 6512 38640 6528 38704
rect 6592 38640 6608 38704
rect 6672 38640 6688 38704
rect 6752 38640 6768 38704
rect 6832 38640 6848 38704
rect 6912 38640 6928 38704
rect 6992 38640 7008 38704
rect 7072 38640 7088 38704
rect 7152 38640 7168 38704
rect 7232 38640 7248 38704
rect 7312 38640 7328 38704
rect 7392 38640 7408 38704
rect 7472 38640 7488 38704
rect 7552 38640 7568 38704
rect 7632 38640 7648 38704
rect 7712 38640 7728 38704
rect 7792 38640 7808 38704
rect 7872 38640 7888 38704
rect 7952 38640 7968 38704
rect 8032 38640 8048 38704
rect 8112 38640 8128 38704
rect 8192 38640 8208 38704
rect 8272 38640 8288 38704
rect 8352 38640 8368 38704
rect 8432 38640 8448 38704
rect 8512 38640 8528 38704
rect 8592 38640 8608 38704
rect 8672 38640 8688 38704
rect 8752 38640 8768 38704
rect 8832 38640 8848 38704
rect 8912 38640 8928 38704
rect 8992 38640 14112 38704
rect 14176 38640 14192 38704
rect 14256 38640 14272 38704
rect 14336 38640 14352 38704
rect 14416 38640 24112 38704
rect 24176 38640 24192 38704
rect 24256 38640 24272 38704
rect 24336 38640 24352 38704
rect 24416 38640 36376 38704
rect 36440 38640 36456 38704
rect 36520 38640 36536 38704
rect 36600 38640 36616 38704
rect 36680 38640 36696 38704
rect 36760 38640 36776 38704
rect 36840 38640 36856 38704
rect 36920 38640 36936 38704
rect 37000 38640 37016 38704
rect 37080 38640 37096 38704
rect 37160 38640 37176 38704
rect 37240 38640 37256 38704
rect 37320 38640 37336 38704
rect 37400 38640 37416 38704
rect 37480 38640 37496 38704
rect 37560 38640 37576 38704
rect 37640 38640 37656 38704
rect 37720 38640 37736 38704
rect 37800 38640 37816 38704
rect 37880 38640 37896 38704
rect 37960 38640 37976 38704
rect 38040 38640 38056 38704
rect 38120 38640 38136 38704
rect 38200 38640 38216 38704
rect 38280 38640 38296 38704
rect 38360 38640 38376 38704
rect 38440 38640 38456 38704
rect 38520 38640 38536 38704
rect 38600 38640 38616 38704
rect 38680 38640 38696 38704
rect 38760 38640 38776 38704
rect 38840 38640 38856 38704
rect 38920 38640 38936 38704
rect 39000 38640 39016 38704
rect 39080 38640 39096 38704
rect 39160 38640 39176 38704
rect 39240 38640 39256 38704
rect 39320 38640 39336 38704
rect 39400 38640 39416 38704
rect 39480 38640 39496 38704
rect 39560 38640 39576 38704
rect 39640 38640 39656 38704
rect 39720 38640 39736 38704
rect 39800 38640 39816 38704
rect 39880 38640 39896 38704
rect 39960 38640 39976 38704
rect 40040 38640 40056 38704
rect 40120 38640 40136 38704
rect 40200 38640 40216 38704
rect 40280 38640 40296 38704
rect 40360 38640 40368 38704
rect 5000 38624 40368 38640
rect 5000 38560 5008 38624
rect 5072 38560 5088 38624
rect 5152 38560 5168 38624
rect 5232 38560 5248 38624
rect 5312 38560 5328 38624
rect 5392 38560 5408 38624
rect 5472 38560 5488 38624
rect 5552 38560 5568 38624
rect 5632 38560 5648 38624
rect 5712 38560 5728 38624
rect 5792 38560 5808 38624
rect 5872 38560 5888 38624
rect 5952 38560 5968 38624
rect 6032 38560 6048 38624
rect 6112 38560 6128 38624
rect 6192 38560 6208 38624
rect 6272 38560 6288 38624
rect 6352 38560 6368 38624
rect 6432 38560 6448 38624
rect 6512 38560 6528 38624
rect 6592 38560 6608 38624
rect 6672 38560 6688 38624
rect 6752 38560 6768 38624
rect 6832 38560 6848 38624
rect 6912 38560 6928 38624
rect 6992 38560 7008 38624
rect 7072 38560 7088 38624
rect 7152 38560 7168 38624
rect 7232 38560 7248 38624
rect 7312 38560 7328 38624
rect 7392 38560 7408 38624
rect 7472 38560 7488 38624
rect 7552 38560 7568 38624
rect 7632 38560 7648 38624
rect 7712 38560 7728 38624
rect 7792 38560 7808 38624
rect 7872 38560 7888 38624
rect 7952 38560 7968 38624
rect 8032 38560 8048 38624
rect 8112 38560 8128 38624
rect 8192 38560 8208 38624
rect 8272 38560 8288 38624
rect 8352 38560 8368 38624
rect 8432 38560 8448 38624
rect 8512 38560 8528 38624
rect 8592 38560 8608 38624
rect 8672 38560 8688 38624
rect 8752 38560 8768 38624
rect 8832 38560 8848 38624
rect 8912 38560 8928 38624
rect 8992 38560 14112 38624
rect 14176 38560 14192 38624
rect 14256 38560 14272 38624
rect 14336 38560 14352 38624
rect 14416 38560 24112 38624
rect 24176 38560 24192 38624
rect 24256 38560 24272 38624
rect 24336 38560 24352 38624
rect 24416 38560 36376 38624
rect 36440 38560 36456 38624
rect 36520 38560 36536 38624
rect 36600 38560 36616 38624
rect 36680 38560 36696 38624
rect 36760 38560 36776 38624
rect 36840 38560 36856 38624
rect 36920 38560 36936 38624
rect 37000 38560 37016 38624
rect 37080 38560 37096 38624
rect 37160 38560 37176 38624
rect 37240 38560 37256 38624
rect 37320 38560 37336 38624
rect 37400 38560 37416 38624
rect 37480 38560 37496 38624
rect 37560 38560 37576 38624
rect 37640 38560 37656 38624
rect 37720 38560 37736 38624
rect 37800 38560 37816 38624
rect 37880 38560 37896 38624
rect 37960 38560 37976 38624
rect 38040 38560 38056 38624
rect 38120 38560 38136 38624
rect 38200 38560 38216 38624
rect 38280 38560 38296 38624
rect 38360 38560 38376 38624
rect 38440 38560 38456 38624
rect 38520 38560 38536 38624
rect 38600 38560 38616 38624
rect 38680 38560 38696 38624
rect 38760 38560 38776 38624
rect 38840 38560 38856 38624
rect 38920 38560 38936 38624
rect 39000 38560 39016 38624
rect 39080 38560 39096 38624
rect 39160 38560 39176 38624
rect 39240 38560 39256 38624
rect 39320 38560 39336 38624
rect 39400 38560 39416 38624
rect 39480 38560 39496 38624
rect 39560 38560 39576 38624
rect 39640 38560 39656 38624
rect 39720 38560 39736 38624
rect 39800 38560 39816 38624
rect 39880 38560 39896 38624
rect 39960 38560 39976 38624
rect 40040 38560 40056 38624
rect 40120 38560 40136 38624
rect 40200 38560 40216 38624
rect 40280 38560 40296 38624
rect 40360 38560 40368 38624
rect 5000 38544 40368 38560
rect 5000 38480 5008 38544
rect 5072 38480 5088 38544
rect 5152 38480 5168 38544
rect 5232 38480 5248 38544
rect 5312 38480 5328 38544
rect 5392 38480 5408 38544
rect 5472 38480 5488 38544
rect 5552 38480 5568 38544
rect 5632 38480 5648 38544
rect 5712 38480 5728 38544
rect 5792 38480 5808 38544
rect 5872 38480 5888 38544
rect 5952 38480 5968 38544
rect 6032 38480 6048 38544
rect 6112 38480 6128 38544
rect 6192 38480 6208 38544
rect 6272 38480 6288 38544
rect 6352 38480 6368 38544
rect 6432 38480 6448 38544
rect 6512 38480 6528 38544
rect 6592 38480 6608 38544
rect 6672 38480 6688 38544
rect 6752 38480 6768 38544
rect 6832 38480 6848 38544
rect 6912 38480 6928 38544
rect 6992 38480 7008 38544
rect 7072 38480 7088 38544
rect 7152 38480 7168 38544
rect 7232 38480 7248 38544
rect 7312 38480 7328 38544
rect 7392 38480 7408 38544
rect 7472 38480 7488 38544
rect 7552 38480 7568 38544
rect 7632 38480 7648 38544
rect 7712 38480 7728 38544
rect 7792 38480 7808 38544
rect 7872 38480 7888 38544
rect 7952 38480 7968 38544
rect 8032 38480 8048 38544
rect 8112 38480 8128 38544
rect 8192 38480 8208 38544
rect 8272 38480 8288 38544
rect 8352 38480 8368 38544
rect 8432 38480 8448 38544
rect 8512 38480 8528 38544
rect 8592 38480 8608 38544
rect 8672 38480 8688 38544
rect 8752 38480 8768 38544
rect 8832 38480 8848 38544
rect 8912 38480 8928 38544
rect 8992 38480 14112 38544
rect 14176 38480 14192 38544
rect 14256 38480 14272 38544
rect 14336 38480 14352 38544
rect 14416 38480 24112 38544
rect 24176 38480 24192 38544
rect 24256 38480 24272 38544
rect 24336 38480 24352 38544
rect 24416 38480 36376 38544
rect 36440 38480 36456 38544
rect 36520 38480 36536 38544
rect 36600 38480 36616 38544
rect 36680 38480 36696 38544
rect 36760 38480 36776 38544
rect 36840 38480 36856 38544
rect 36920 38480 36936 38544
rect 37000 38480 37016 38544
rect 37080 38480 37096 38544
rect 37160 38480 37176 38544
rect 37240 38480 37256 38544
rect 37320 38480 37336 38544
rect 37400 38480 37416 38544
rect 37480 38480 37496 38544
rect 37560 38480 37576 38544
rect 37640 38480 37656 38544
rect 37720 38480 37736 38544
rect 37800 38480 37816 38544
rect 37880 38480 37896 38544
rect 37960 38480 37976 38544
rect 38040 38480 38056 38544
rect 38120 38480 38136 38544
rect 38200 38480 38216 38544
rect 38280 38480 38296 38544
rect 38360 38480 38376 38544
rect 38440 38480 38456 38544
rect 38520 38480 38536 38544
rect 38600 38480 38616 38544
rect 38680 38480 38696 38544
rect 38760 38480 38776 38544
rect 38840 38480 38856 38544
rect 38920 38480 38936 38544
rect 39000 38480 39016 38544
rect 39080 38480 39096 38544
rect 39160 38480 39176 38544
rect 39240 38480 39256 38544
rect 39320 38480 39336 38544
rect 39400 38480 39416 38544
rect 39480 38480 39496 38544
rect 39560 38480 39576 38544
rect 39640 38480 39656 38544
rect 39720 38480 39736 38544
rect 39800 38480 39816 38544
rect 39880 38480 39896 38544
rect 39960 38480 39976 38544
rect 40040 38480 40056 38544
rect 40120 38480 40136 38544
rect 40200 38480 40216 38544
rect 40280 38480 40296 38544
rect 40360 38480 40368 38544
rect 5000 38464 40368 38480
rect 5000 38400 5008 38464
rect 5072 38400 5088 38464
rect 5152 38400 5168 38464
rect 5232 38400 5248 38464
rect 5312 38400 5328 38464
rect 5392 38400 5408 38464
rect 5472 38400 5488 38464
rect 5552 38400 5568 38464
rect 5632 38400 5648 38464
rect 5712 38400 5728 38464
rect 5792 38400 5808 38464
rect 5872 38400 5888 38464
rect 5952 38400 5968 38464
rect 6032 38400 6048 38464
rect 6112 38400 6128 38464
rect 6192 38400 6208 38464
rect 6272 38400 6288 38464
rect 6352 38400 6368 38464
rect 6432 38400 6448 38464
rect 6512 38400 6528 38464
rect 6592 38400 6608 38464
rect 6672 38400 6688 38464
rect 6752 38400 6768 38464
rect 6832 38400 6848 38464
rect 6912 38400 6928 38464
rect 6992 38400 7008 38464
rect 7072 38400 7088 38464
rect 7152 38400 7168 38464
rect 7232 38400 7248 38464
rect 7312 38400 7328 38464
rect 7392 38400 7408 38464
rect 7472 38400 7488 38464
rect 7552 38400 7568 38464
rect 7632 38400 7648 38464
rect 7712 38400 7728 38464
rect 7792 38400 7808 38464
rect 7872 38400 7888 38464
rect 7952 38400 7968 38464
rect 8032 38400 8048 38464
rect 8112 38400 8128 38464
rect 8192 38400 8208 38464
rect 8272 38400 8288 38464
rect 8352 38400 8368 38464
rect 8432 38400 8448 38464
rect 8512 38400 8528 38464
rect 8592 38400 8608 38464
rect 8672 38400 8688 38464
rect 8752 38400 8768 38464
rect 8832 38400 8848 38464
rect 8912 38400 8928 38464
rect 8992 38400 14112 38464
rect 14176 38400 14192 38464
rect 14256 38400 14272 38464
rect 14336 38400 14352 38464
rect 14416 38400 24112 38464
rect 24176 38400 24192 38464
rect 24256 38400 24272 38464
rect 24336 38400 24352 38464
rect 24416 38400 36376 38464
rect 36440 38400 36456 38464
rect 36520 38400 36536 38464
rect 36600 38400 36616 38464
rect 36680 38400 36696 38464
rect 36760 38400 36776 38464
rect 36840 38400 36856 38464
rect 36920 38400 36936 38464
rect 37000 38400 37016 38464
rect 37080 38400 37096 38464
rect 37160 38400 37176 38464
rect 37240 38400 37256 38464
rect 37320 38400 37336 38464
rect 37400 38400 37416 38464
rect 37480 38400 37496 38464
rect 37560 38400 37576 38464
rect 37640 38400 37656 38464
rect 37720 38400 37736 38464
rect 37800 38400 37816 38464
rect 37880 38400 37896 38464
rect 37960 38400 37976 38464
rect 38040 38400 38056 38464
rect 38120 38400 38136 38464
rect 38200 38400 38216 38464
rect 38280 38400 38296 38464
rect 38360 38400 38376 38464
rect 38440 38400 38456 38464
rect 38520 38400 38536 38464
rect 38600 38400 38616 38464
rect 38680 38400 38696 38464
rect 38760 38400 38776 38464
rect 38840 38400 38856 38464
rect 38920 38400 38936 38464
rect 39000 38400 39016 38464
rect 39080 38400 39096 38464
rect 39160 38400 39176 38464
rect 39240 38400 39256 38464
rect 39320 38400 39336 38464
rect 39400 38400 39416 38464
rect 39480 38400 39496 38464
rect 39560 38400 39576 38464
rect 39640 38400 39656 38464
rect 39720 38400 39736 38464
rect 39800 38400 39816 38464
rect 39880 38400 39896 38464
rect 39960 38400 39976 38464
rect 40040 38400 40056 38464
rect 40120 38400 40136 38464
rect 40200 38400 40216 38464
rect 40280 38400 40296 38464
rect 40360 38400 40368 38464
rect 5000 38384 40368 38400
rect 5000 38320 5008 38384
rect 5072 38320 5088 38384
rect 5152 38320 5168 38384
rect 5232 38320 5248 38384
rect 5312 38320 5328 38384
rect 5392 38320 5408 38384
rect 5472 38320 5488 38384
rect 5552 38320 5568 38384
rect 5632 38320 5648 38384
rect 5712 38320 5728 38384
rect 5792 38320 5808 38384
rect 5872 38320 5888 38384
rect 5952 38320 5968 38384
rect 6032 38320 6048 38384
rect 6112 38320 6128 38384
rect 6192 38320 6208 38384
rect 6272 38320 6288 38384
rect 6352 38320 6368 38384
rect 6432 38320 6448 38384
rect 6512 38320 6528 38384
rect 6592 38320 6608 38384
rect 6672 38320 6688 38384
rect 6752 38320 6768 38384
rect 6832 38320 6848 38384
rect 6912 38320 6928 38384
rect 6992 38320 7008 38384
rect 7072 38320 7088 38384
rect 7152 38320 7168 38384
rect 7232 38320 7248 38384
rect 7312 38320 7328 38384
rect 7392 38320 7408 38384
rect 7472 38320 7488 38384
rect 7552 38320 7568 38384
rect 7632 38320 7648 38384
rect 7712 38320 7728 38384
rect 7792 38320 7808 38384
rect 7872 38320 7888 38384
rect 7952 38320 7968 38384
rect 8032 38320 8048 38384
rect 8112 38320 8128 38384
rect 8192 38320 8208 38384
rect 8272 38320 8288 38384
rect 8352 38320 8368 38384
rect 8432 38320 8448 38384
rect 8512 38320 8528 38384
rect 8592 38320 8608 38384
rect 8672 38320 8688 38384
rect 8752 38320 8768 38384
rect 8832 38320 8848 38384
rect 8912 38320 8928 38384
rect 8992 38320 14112 38384
rect 14176 38320 14192 38384
rect 14256 38320 14272 38384
rect 14336 38320 14352 38384
rect 14416 38320 24112 38384
rect 24176 38320 24192 38384
rect 24256 38320 24272 38384
rect 24336 38320 24352 38384
rect 24416 38320 36376 38384
rect 36440 38320 36456 38384
rect 36520 38320 36536 38384
rect 36600 38320 36616 38384
rect 36680 38320 36696 38384
rect 36760 38320 36776 38384
rect 36840 38320 36856 38384
rect 36920 38320 36936 38384
rect 37000 38320 37016 38384
rect 37080 38320 37096 38384
rect 37160 38320 37176 38384
rect 37240 38320 37256 38384
rect 37320 38320 37336 38384
rect 37400 38320 37416 38384
rect 37480 38320 37496 38384
rect 37560 38320 37576 38384
rect 37640 38320 37656 38384
rect 37720 38320 37736 38384
rect 37800 38320 37816 38384
rect 37880 38320 37896 38384
rect 37960 38320 37976 38384
rect 38040 38320 38056 38384
rect 38120 38320 38136 38384
rect 38200 38320 38216 38384
rect 38280 38320 38296 38384
rect 38360 38320 38376 38384
rect 38440 38320 38456 38384
rect 38520 38320 38536 38384
rect 38600 38320 38616 38384
rect 38680 38320 38696 38384
rect 38760 38320 38776 38384
rect 38840 38320 38856 38384
rect 38920 38320 38936 38384
rect 39000 38320 39016 38384
rect 39080 38320 39096 38384
rect 39160 38320 39176 38384
rect 39240 38320 39256 38384
rect 39320 38320 39336 38384
rect 39400 38320 39416 38384
rect 39480 38320 39496 38384
rect 39560 38320 39576 38384
rect 39640 38320 39656 38384
rect 39720 38320 39736 38384
rect 39800 38320 39816 38384
rect 39880 38320 39896 38384
rect 39960 38320 39976 38384
rect 40040 38320 40056 38384
rect 40120 38320 40136 38384
rect 40200 38320 40216 38384
rect 40280 38320 40296 38384
rect 40360 38320 40368 38384
rect 5000 38304 40368 38320
rect 5000 38240 5008 38304
rect 5072 38240 5088 38304
rect 5152 38240 5168 38304
rect 5232 38240 5248 38304
rect 5312 38240 5328 38304
rect 5392 38240 5408 38304
rect 5472 38240 5488 38304
rect 5552 38240 5568 38304
rect 5632 38240 5648 38304
rect 5712 38240 5728 38304
rect 5792 38240 5808 38304
rect 5872 38240 5888 38304
rect 5952 38240 5968 38304
rect 6032 38240 6048 38304
rect 6112 38240 6128 38304
rect 6192 38240 6208 38304
rect 6272 38240 6288 38304
rect 6352 38240 6368 38304
rect 6432 38240 6448 38304
rect 6512 38240 6528 38304
rect 6592 38240 6608 38304
rect 6672 38240 6688 38304
rect 6752 38240 6768 38304
rect 6832 38240 6848 38304
rect 6912 38240 6928 38304
rect 6992 38240 7008 38304
rect 7072 38240 7088 38304
rect 7152 38240 7168 38304
rect 7232 38240 7248 38304
rect 7312 38240 7328 38304
rect 7392 38240 7408 38304
rect 7472 38240 7488 38304
rect 7552 38240 7568 38304
rect 7632 38240 7648 38304
rect 7712 38240 7728 38304
rect 7792 38240 7808 38304
rect 7872 38240 7888 38304
rect 7952 38240 7968 38304
rect 8032 38240 8048 38304
rect 8112 38240 8128 38304
rect 8192 38240 8208 38304
rect 8272 38240 8288 38304
rect 8352 38240 8368 38304
rect 8432 38240 8448 38304
rect 8512 38240 8528 38304
rect 8592 38240 8608 38304
rect 8672 38240 8688 38304
rect 8752 38240 8768 38304
rect 8832 38240 8848 38304
rect 8912 38240 8928 38304
rect 8992 38240 14112 38304
rect 14176 38240 14192 38304
rect 14256 38240 14272 38304
rect 14336 38240 14352 38304
rect 14416 38240 24112 38304
rect 24176 38240 24192 38304
rect 24256 38240 24272 38304
rect 24336 38240 24352 38304
rect 24416 38240 36376 38304
rect 36440 38240 36456 38304
rect 36520 38240 36536 38304
rect 36600 38240 36616 38304
rect 36680 38240 36696 38304
rect 36760 38240 36776 38304
rect 36840 38240 36856 38304
rect 36920 38240 36936 38304
rect 37000 38240 37016 38304
rect 37080 38240 37096 38304
rect 37160 38240 37176 38304
rect 37240 38240 37256 38304
rect 37320 38240 37336 38304
rect 37400 38240 37416 38304
rect 37480 38240 37496 38304
rect 37560 38240 37576 38304
rect 37640 38240 37656 38304
rect 37720 38240 37736 38304
rect 37800 38240 37816 38304
rect 37880 38240 37896 38304
rect 37960 38240 37976 38304
rect 38040 38240 38056 38304
rect 38120 38240 38136 38304
rect 38200 38240 38216 38304
rect 38280 38240 38296 38304
rect 38360 38240 38376 38304
rect 38440 38240 38456 38304
rect 38520 38240 38536 38304
rect 38600 38240 38616 38304
rect 38680 38240 38696 38304
rect 38760 38240 38776 38304
rect 38840 38240 38856 38304
rect 38920 38240 38936 38304
rect 39000 38240 39016 38304
rect 39080 38240 39096 38304
rect 39160 38240 39176 38304
rect 39240 38240 39256 38304
rect 39320 38240 39336 38304
rect 39400 38240 39416 38304
rect 39480 38240 39496 38304
rect 39560 38240 39576 38304
rect 39640 38240 39656 38304
rect 39720 38240 39736 38304
rect 39800 38240 39816 38304
rect 39880 38240 39896 38304
rect 39960 38240 39976 38304
rect 40040 38240 40056 38304
rect 40120 38240 40136 38304
rect 40200 38240 40216 38304
rect 40280 38240 40296 38304
rect 40360 38240 40368 38304
rect 5000 38224 40368 38240
rect 5000 38160 5008 38224
rect 5072 38160 5088 38224
rect 5152 38160 5168 38224
rect 5232 38160 5248 38224
rect 5312 38160 5328 38224
rect 5392 38160 5408 38224
rect 5472 38160 5488 38224
rect 5552 38160 5568 38224
rect 5632 38160 5648 38224
rect 5712 38160 5728 38224
rect 5792 38160 5808 38224
rect 5872 38160 5888 38224
rect 5952 38160 5968 38224
rect 6032 38160 6048 38224
rect 6112 38160 6128 38224
rect 6192 38160 6208 38224
rect 6272 38160 6288 38224
rect 6352 38160 6368 38224
rect 6432 38160 6448 38224
rect 6512 38160 6528 38224
rect 6592 38160 6608 38224
rect 6672 38160 6688 38224
rect 6752 38160 6768 38224
rect 6832 38160 6848 38224
rect 6912 38160 6928 38224
rect 6992 38160 7008 38224
rect 7072 38160 7088 38224
rect 7152 38160 7168 38224
rect 7232 38160 7248 38224
rect 7312 38160 7328 38224
rect 7392 38160 7408 38224
rect 7472 38160 7488 38224
rect 7552 38160 7568 38224
rect 7632 38160 7648 38224
rect 7712 38160 7728 38224
rect 7792 38160 7808 38224
rect 7872 38160 7888 38224
rect 7952 38160 7968 38224
rect 8032 38160 8048 38224
rect 8112 38160 8128 38224
rect 8192 38160 8208 38224
rect 8272 38160 8288 38224
rect 8352 38160 8368 38224
rect 8432 38160 8448 38224
rect 8512 38160 8528 38224
rect 8592 38160 8608 38224
rect 8672 38160 8688 38224
rect 8752 38160 8768 38224
rect 8832 38160 8848 38224
rect 8912 38160 8928 38224
rect 8992 38160 14112 38224
rect 14176 38160 14192 38224
rect 14256 38160 14272 38224
rect 14336 38160 14352 38224
rect 14416 38160 24112 38224
rect 24176 38160 24192 38224
rect 24256 38160 24272 38224
rect 24336 38160 24352 38224
rect 24416 38160 36376 38224
rect 36440 38160 36456 38224
rect 36520 38160 36536 38224
rect 36600 38160 36616 38224
rect 36680 38160 36696 38224
rect 36760 38160 36776 38224
rect 36840 38160 36856 38224
rect 36920 38160 36936 38224
rect 37000 38160 37016 38224
rect 37080 38160 37096 38224
rect 37160 38160 37176 38224
rect 37240 38160 37256 38224
rect 37320 38160 37336 38224
rect 37400 38160 37416 38224
rect 37480 38160 37496 38224
rect 37560 38160 37576 38224
rect 37640 38160 37656 38224
rect 37720 38160 37736 38224
rect 37800 38160 37816 38224
rect 37880 38160 37896 38224
rect 37960 38160 37976 38224
rect 38040 38160 38056 38224
rect 38120 38160 38136 38224
rect 38200 38160 38216 38224
rect 38280 38160 38296 38224
rect 38360 38160 38376 38224
rect 38440 38160 38456 38224
rect 38520 38160 38536 38224
rect 38600 38160 38616 38224
rect 38680 38160 38696 38224
rect 38760 38160 38776 38224
rect 38840 38160 38856 38224
rect 38920 38160 38936 38224
rect 39000 38160 39016 38224
rect 39080 38160 39096 38224
rect 39160 38160 39176 38224
rect 39240 38160 39256 38224
rect 39320 38160 39336 38224
rect 39400 38160 39416 38224
rect 39480 38160 39496 38224
rect 39560 38160 39576 38224
rect 39640 38160 39656 38224
rect 39720 38160 39736 38224
rect 39800 38160 39816 38224
rect 39880 38160 39896 38224
rect 39960 38160 39976 38224
rect 40040 38160 40056 38224
rect 40120 38160 40136 38224
rect 40200 38160 40216 38224
rect 40280 38160 40296 38224
rect 40360 38160 40368 38224
rect 5000 38144 40368 38160
rect 5000 38080 5008 38144
rect 5072 38080 5088 38144
rect 5152 38080 5168 38144
rect 5232 38080 5248 38144
rect 5312 38080 5328 38144
rect 5392 38080 5408 38144
rect 5472 38080 5488 38144
rect 5552 38080 5568 38144
rect 5632 38080 5648 38144
rect 5712 38080 5728 38144
rect 5792 38080 5808 38144
rect 5872 38080 5888 38144
rect 5952 38080 5968 38144
rect 6032 38080 6048 38144
rect 6112 38080 6128 38144
rect 6192 38080 6208 38144
rect 6272 38080 6288 38144
rect 6352 38080 6368 38144
rect 6432 38080 6448 38144
rect 6512 38080 6528 38144
rect 6592 38080 6608 38144
rect 6672 38080 6688 38144
rect 6752 38080 6768 38144
rect 6832 38080 6848 38144
rect 6912 38080 6928 38144
rect 6992 38080 7008 38144
rect 7072 38080 7088 38144
rect 7152 38080 7168 38144
rect 7232 38080 7248 38144
rect 7312 38080 7328 38144
rect 7392 38080 7408 38144
rect 7472 38080 7488 38144
rect 7552 38080 7568 38144
rect 7632 38080 7648 38144
rect 7712 38080 7728 38144
rect 7792 38080 7808 38144
rect 7872 38080 7888 38144
rect 7952 38080 7968 38144
rect 8032 38080 8048 38144
rect 8112 38080 8128 38144
rect 8192 38080 8208 38144
rect 8272 38080 8288 38144
rect 8352 38080 8368 38144
rect 8432 38080 8448 38144
rect 8512 38080 8528 38144
rect 8592 38080 8608 38144
rect 8672 38080 8688 38144
rect 8752 38080 8768 38144
rect 8832 38080 8848 38144
rect 8912 38080 8928 38144
rect 8992 38080 14112 38144
rect 14176 38080 14192 38144
rect 14256 38080 14272 38144
rect 14336 38080 14352 38144
rect 14416 38080 24112 38144
rect 24176 38080 24192 38144
rect 24256 38080 24272 38144
rect 24336 38080 24352 38144
rect 24416 38080 36376 38144
rect 36440 38080 36456 38144
rect 36520 38080 36536 38144
rect 36600 38080 36616 38144
rect 36680 38080 36696 38144
rect 36760 38080 36776 38144
rect 36840 38080 36856 38144
rect 36920 38080 36936 38144
rect 37000 38080 37016 38144
rect 37080 38080 37096 38144
rect 37160 38080 37176 38144
rect 37240 38080 37256 38144
rect 37320 38080 37336 38144
rect 37400 38080 37416 38144
rect 37480 38080 37496 38144
rect 37560 38080 37576 38144
rect 37640 38080 37656 38144
rect 37720 38080 37736 38144
rect 37800 38080 37816 38144
rect 37880 38080 37896 38144
rect 37960 38080 37976 38144
rect 38040 38080 38056 38144
rect 38120 38080 38136 38144
rect 38200 38080 38216 38144
rect 38280 38080 38296 38144
rect 38360 38080 38376 38144
rect 38440 38080 38456 38144
rect 38520 38080 38536 38144
rect 38600 38080 38616 38144
rect 38680 38080 38696 38144
rect 38760 38080 38776 38144
rect 38840 38080 38856 38144
rect 38920 38080 38936 38144
rect 39000 38080 39016 38144
rect 39080 38080 39096 38144
rect 39160 38080 39176 38144
rect 39240 38080 39256 38144
rect 39320 38080 39336 38144
rect 39400 38080 39416 38144
rect 39480 38080 39496 38144
rect 39560 38080 39576 38144
rect 39640 38080 39656 38144
rect 39720 38080 39736 38144
rect 39800 38080 39816 38144
rect 39880 38080 39896 38144
rect 39960 38080 39976 38144
rect 40040 38080 40056 38144
rect 40120 38080 40136 38144
rect 40200 38080 40216 38144
rect 40280 38080 40296 38144
rect 40360 38080 40368 38144
rect 5000 38064 40368 38080
rect 5000 38000 5008 38064
rect 5072 38000 5088 38064
rect 5152 38000 5168 38064
rect 5232 38000 5248 38064
rect 5312 38000 5328 38064
rect 5392 38000 5408 38064
rect 5472 38000 5488 38064
rect 5552 38000 5568 38064
rect 5632 38000 5648 38064
rect 5712 38000 5728 38064
rect 5792 38000 5808 38064
rect 5872 38000 5888 38064
rect 5952 38000 5968 38064
rect 6032 38000 6048 38064
rect 6112 38000 6128 38064
rect 6192 38000 6208 38064
rect 6272 38000 6288 38064
rect 6352 38000 6368 38064
rect 6432 38000 6448 38064
rect 6512 38000 6528 38064
rect 6592 38000 6608 38064
rect 6672 38000 6688 38064
rect 6752 38000 6768 38064
rect 6832 38000 6848 38064
rect 6912 38000 6928 38064
rect 6992 38000 7008 38064
rect 7072 38000 7088 38064
rect 7152 38000 7168 38064
rect 7232 38000 7248 38064
rect 7312 38000 7328 38064
rect 7392 38000 7408 38064
rect 7472 38000 7488 38064
rect 7552 38000 7568 38064
rect 7632 38000 7648 38064
rect 7712 38000 7728 38064
rect 7792 38000 7808 38064
rect 7872 38000 7888 38064
rect 7952 38000 7968 38064
rect 8032 38000 8048 38064
rect 8112 38000 8128 38064
rect 8192 38000 8208 38064
rect 8272 38000 8288 38064
rect 8352 38000 8368 38064
rect 8432 38000 8448 38064
rect 8512 38000 8528 38064
rect 8592 38000 8608 38064
rect 8672 38000 8688 38064
rect 8752 38000 8768 38064
rect 8832 38000 8848 38064
rect 8912 38000 8928 38064
rect 8992 38000 14112 38064
rect 14176 38000 14192 38064
rect 14256 38000 14272 38064
rect 14336 38000 14352 38064
rect 14416 38000 24112 38064
rect 24176 38000 24192 38064
rect 24256 38000 24272 38064
rect 24336 38000 24352 38064
rect 24416 38000 36376 38064
rect 36440 38000 36456 38064
rect 36520 38000 36536 38064
rect 36600 38000 36616 38064
rect 36680 38000 36696 38064
rect 36760 38000 36776 38064
rect 36840 38000 36856 38064
rect 36920 38000 36936 38064
rect 37000 38000 37016 38064
rect 37080 38000 37096 38064
rect 37160 38000 37176 38064
rect 37240 38000 37256 38064
rect 37320 38000 37336 38064
rect 37400 38000 37416 38064
rect 37480 38000 37496 38064
rect 37560 38000 37576 38064
rect 37640 38000 37656 38064
rect 37720 38000 37736 38064
rect 37800 38000 37816 38064
rect 37880 38000 37896 38064
rect 37960 38000 37976 38064
rect 38040 38000 38056 38064
rect 38120 38000 38136 38064
rect 38200 38000 38216 38064
rect 38280 38000 38296 38064
rect 38360 38000 38376 38064
rect 38440 38000 38456 38064
rect 38520 38000 38536 38064
rect 38600 38000 38616 38064
rect 38680 38000 38696 38064
rect 38760 38000 38776 38064
rect 38840 38000 38856 38064
rect 38920 38000 38936 38064
rect 39000 38000 39016 38064
rect 39080 38000 39096 38064
rect 39160 38000 39176 38064
rect 39240 38000 39256 38064
rect 39320 38000 39336 38064
rect 39400 38000 39416 38064
rect 39480 38000 39496 38064
rect 39560 38000 39576 38064
rect 39640 38000 39656 38064
rect 39720 38000 39736 38064
rect 39800 38000 39816 38064
rect 39880 38000 39896 38064
rect 39960 38000 39976 38064
rect 40040 38000 40056 38064
rect 40120 38000 40136 38064
rect 40200 38000 40216 38064
rect 40280 38000 40296 38064
rect 40360 38000 40368 38064
rect 5000 37984 40368 38000
rect 5000 37920 5008 37984
rect 5072 37920 5088 37984
rect 5152 37920 5168 37984
rect 5232 37920 5248 37984
rect 5312 37920 5328 37984
rect 5392 37920 5408 37984
rect 5472 37920 5488 37984
rect 5552 37920 5568 37984
rect 5632 37920 5648 37984
rect 5712 37920 5728 37984
rect 5792 37920 5808 37984
rect 5872 37920 5888 37984
rect 5952 37920 5968 37984
rect 6032 37920 6048 37984
rect 6112 37920 6128 37984
rect 6192 37920 6208 37984
rect 6272 37920 6288 37984
rect 6352 37920 6368 37984
rect 6432 37920 6448 37984
rect 6512 37920 6528 37984
rect 6592 37920 6608 37984
rect 6672 37920 6688 37984
rect 6752 37920 6768 37984
rect 6832 37920 6848 37984
rect 6912 37920 6928 37984
rect 6992 37920 7008 37984
rect 7072 37920 7088 37984
rect 7152 37920 7168 37984
rect 7232 37920 7248 37984
rect 7312 37920 7328 37984
rect 7392 37920 7408 37984
rect 7472 37920 7488 37984
rect 7552 37920 7568 37984
rect 7632 37920 7648 37984
rect 7712 37920 7728 37984
rect 7792 37920 7808 37984
rect 7872 37920 7888 37984
rect 7952 37920 7968 37984
rect 8032 37920 8048 37984
rect 8112 37920 8128 37984
rect 8192 37920 8208 37984
rect 8272 37920 8288 37984
rect 8352 37920 8368 37984
rect 8432 37920 8448 37984
rect 8512 37920 8528 37984
rect 8592 37920 8608 37984
rect 8672 37920 8688 37984
rect 8752 37920 8768 37984
rect 8832 37920 8848 37984
rect 8912 37920 8928 37984
rect 8992 37920 14112 37984
rect 14176 37920 14192 37984
rect 14256 37920 14272 37984
rect 14336 37920 14352 37984
rect 14416 37920 24112 37984
rect 24176 37920 24192 37984
rect 24256 37920 24272 37984
rect 24336 37920 24352 37984
rect 24416 37920 36376 37984
rect 36440 37920 36456 37984
rect 36520 37920 36536 37984
rect 36600 37920 36616 37984
rect 36680 37920 36696 37984
rect 36760 37920 36776 37984
rect 36840 37920 36856 37984
rect 36920 37920 36936 37984
rect 37000 37920 37016 37984
rect 37080 37920 37096 37984
rect 37160 37920 37176 37984
rect 37240 37920 37256 37984
rect 37320 37920 37336 37984
rect 37400 37920 37416 37984
rect 37480 37920 37496 37984
rect 37560 37920 37576 37984
rect 37640 37920 37656 37984
rect 37720 37920 37736 37984
rect 37800 37920 37816 37984
rect 37880 37920 37896 37984
rect 37960 37920 37976 37984
rect 38040 37920 38056 37984
rect 38120 37920 38136 37984
rect 38200 37920 38216 37984
rect 38280 37920 38296 37984
rect 38360 37920 38376 37984
rect 38440 37920 38456 37984
rect 38520 37920 38536 37984
rect 38600 37920 38616 37984
rect 38680 37920 38696 37984
rect 38760 37920 38776 37984
rect 38840 37920 38856 37984
rect 38920 37920 38936 37984
rect 39000 37920 39016 37984
rect 39080 37920 39096 37984
rect 39160 37920 39176 37984
rect 39240 37920 39256 37984
rect 39320 37920 39336 37984
rect 39400 37920 39416 37984
rect 39480 37920 39496 37984
rect 39560 37920 39576 37984
rect 39640 37920 39656 37984
rect 39720 37920 39736 37984
rect 39800 37920 39816 37984
rect 39880 37920 39896 37984
rect 39960 37920 39976 37984
rect 40040 37920 40056 37984
rect 40120 37920 40136 37984
rect 40200 37920 40216 37984
rect 40280 37920 40296 37984
rect 40360 37920 40368 37984
rect 5000 37904 40368 37920
rect 5000 37840 5008 37904
rect 5072 37840 5088 37904
rect 5152 37840 5168 37904
rect 5232 37840 5248 37904
rect 5312 37840 5328 37904
rect 5392 37840 5408 37904
rect 5472 37840 5488 37904
rect 5552 37840 5568 37904
rect 5632 37840 5648 37904
rect 5712 37840 5728 37904
rect 5792 37840 5808 37904
rect 5872 37840 5888 37904
rect 5952 37840 5968 37904
rect 6032 37840 6048 37904
rect 6112 37840 6128 37904
rect 6192 37840 6208 37904
rect 6272 37840 6288 37904
rect 6352 37840 6368 37904
rect 6432 37840 6448 37904
rect 6512 37840 6528 37904
rect 6592 37840 6608 37904
rect 6672 37840 6688 37904
rect 6752 37840 6768 37904
rect 6832 37840 6848 37904
rect 6912 37840 6928 37904
rect 6992 37840 7008 37904
rect 7072 37840 7088 37904
rect 7152 37840 7168 37904
rect 7232 37840 7248 37904
rect 7312 37840 7328 37904
rect 7392 37840 7408 37904
rect 7472 37840 7488 37904
rect 7552 37840 7568 37904
rect 7632 37840 7648 37904
rect 7712 37840 7728 37904
rect 7792 37840 7808 37904
rect 7872 37840 7888 37904
rect 7952 37840 7968 37904
rect 8032 37840 8048 37904
rect 8112 37840 8128 37904
rect 8192 37840 8208 37904
rect 8272 37840 8288 37904
rect 8352 37840 8368 37904
rect 8432 37840 8448 37904
rect 8512 37840 8528 37904
rect 8592 37840 8608 37904
rect 8672 37840 8688 37904
rect 8752 37840 8768 37904
rect 8832 37840 8848 37904
rect 8912 37840 8928 37904
rect 8992 37840 14112 37904
rect 14176 37840 14192 37904
rect 14256 37840 14272 37904
rect 14336 37840 14352 37904
rect 14416 37840 24112 37904
rect 24176 37840 24192 37904
rect 24256 37840 24272 37904
rect 24336 37840 24352 37904
rect 24416 37840 36376 37904
rect 36440 37840 36456 37904
rect 36520 37840 36536 37904
rect 36600 37840 36616 37904
rect 36680 37840 36696 37904
rect 36760 37840 36776 37904
rect 36840 37840 36856 37904
rect 36920 37840 36936 37904
rect 37000 37840 37016 37904
rect 37080 37840 37096 37904
rect 37160 37840 37176 37904
rect 37240 37840 37256 37904
rect 37320 37840 37336 37904
rect 37400 37840 37416 37904
rect 37480 37840 37496 37904
rect 37560 37840 37576 37904
rect 37640 37840 37656 37904
rect 37720 37840 37736 37904
rect 37800 37840 37816 37904
rect 37880 37840 37896 37904
rect 37960 37840 37976 37904
rect 38040 37840 38056 37904
rect 38120 37840 38136 37904
rect 38200 37840 38216 37904
rect 38280 37840 38296 37904
rect 38360 37840 38376 37904
rect 38440 37840 38456 37904
rect 38520 37840 38536 37904
rect 38600 37840 38616 37904
rect 38680 37840 38696 37904
rect 38760 37840 38776 37904
rect 38840 37840 38856 37904
rect 38920 37840 38936 37904
rect 39000 37840 39016 37904
rect 39080 37840 39096 37904
rect 39160 37840 39176 37904
rect 39240 37840 39256 37904
rect 39320 37840 39336 37904
rect 39400 37840 39416 37904
rect 39480 37840 39496 37904
rect 39560 37840 39576 37904
rect 39640 37840 39656 37904
rect 39720 37840 39736 37904
rect 39800 37840 39816 37904
rect 39880 37840 39896 37904
rect 39960 37840 39976 37904
rect 40040 37840 40056 37904
rect 40120 37840 40136 37904
rect 40200 37840 40216 37904
rect 40280 37840 40296 37904
rect 40360 37840 40368 37904
rect 5000 37824 40368 37840
rect 5000 37760 5008 37824
rect 5072 37760 5088 37824
rect 5152 37760 5168 37824
rect 5232 37760 5248 37824
rect 5312 37760 5328 37824
rect 5392 37760 5408 37824
rect 5472 37760 5488 37824
rect 5552 37760 5568 37824
rect 5632 37760 5648 37824
rect 5712 37760 5728 37824
rect 5792 37760 5808 37824
rect 5872 37760 5888 37824
rect 5952 37760 5968 37824
rect 6032 37760 6048 37824
rect 6112 37760 6128 37824
rect 6192 37760 6208 37824
rect 6272 37760 6288 37824
rect 6352 37760 6368 37824
rect 6432 37760 6448 37824
rect 6512 37760 6528 37824
rect 6592 37760 6608 37824
rect 6672 37760 6688 37824
rect 6752 37760 6768 37824
rect 6832 37760 6848 37824
rect 6912 37760 6928 37824
rect 6992 37760 7008 37824
rect 7072 37760 7088 37824
rect 7152 37760 7168 37824
rect 7232 37760 7248 37824
rect 7312 37760 7328 37824
rect 7392 37760 7408 37824
rect 7472 37760 7488 37824
rect 7552 37760 7568 37824
rect 7632 37760 7648 37824
rect 7712 37760 7728 37824
rect 7792 37760 7808 37824
rect 7872 37760 7888 37824
rect 7952 37760 7968 37824
rect 8032 37760 8048 37824
rect 8112 37760 8128 37824
rect 8192 37760 8208 37824
rect 8272 37760 8288 37824
rect 8352 37760 8368 37824
rect 8432 37760 8448 37824
rect 8512 37760 8528 37824
rect 8592 37760 8608 37824
rect 8672 37760 8688 37824
rect 8752 37760 8768 37824
rect 8832 37760 8848 37824
rect 8912 37760 8928 37824
rect 8992 37760 14112 37824
rect 14176 37760 14192 37824
rect 14256 37760 14272 37824
rect 14336 37760 14352 37824
rect 14416 37760 24112 37824
rect 24176 37760 24192 37824
rect 24256 37760 24272 37824
rect 24336 37760 24352 37824
rect 24416 37760 36376 37824
rect 36440 37760 36456 37824
rect 36520 37760 36536 37824
rect 36600 37760 36616 37824
rect 36680 37760 36696 37824
rect 36760 37760 36776 37824
rect 36840 37760 36856 37824
rect 36920 37760 36936 37824
rect 37000 37760 37016 37824
rect 37080 37760 37096 37824
rect 37160 37760 37176 37824
rect 37240 37760 37256 37824
rect 37320 37760 37336 37824
rect 37400 37760 37416 37824
rect 37480 37760 37496 37824
rect 37560 37760 37576 37824
rect 37640 37760 37656 37824
rect 37720 37760 37736 37824
rect 37800 37760 37816 37824
rect 37880 37760 37896 37824
rect 37960 37760 37976 37824
rect 38040 37760 38056 37824
rect 38120 37760 38136 37824
rect 38200 37760 38216 37824
rect 38280 37760 38296 37824
rect 38360 37760 38376 37824
rect 38440 37760 38456 37824
rect 38520 37760 38536 37824
rect 38600 37760 38616 37824
rect 38680 37760 38696 37824
rect 38760 37760 38776 37824
rect 38840 37760 38856 37824
rect 38920 37760 38936 37824
rect 39000 37760 39016 37824
rect 39080 37760 39096 37824
rect 39160 37760 39176 37824
rect 39240 37760 39256 37824
rect 39320 37760 39336 37824
rect 39400 37760 39416 37824
rect 39480 37760 39496 37824
rect 39560 37760 39576 37824
rect 39640 37760 39656 37824
rect 39720 37760 39736 37824
rect 39800 37760 39816 37824
rect 39880 37760 39896 37824
rect 39960 37760 39976 37824
rect 40040 37760 40056 37824
rect 40120 37760 40136 37824
rect 40200 37760 40216 37824
rect 40280 37760 40296 37824
rect 40360 37760 40368 37824
rect 5000 37744 40368 37760
rect 5000 37680 5008 37744
rect 5072 37680 5088 37744
rect 5152 37680 5168 37744
rect 5232 37680 5248 37744
rect 5312 37680 5328 37744
rect 5392 37680 5408 37744
rect 5472 37680 5488 37744
rect 5552 37680 5568 37744
rect 5632 37680 5648 37744
rect 5712 37680 5728 37744
rect 5792 37680 5808 37744
rect 5872 37680 5888 37744
rect 5952 37680 5968 37744
rect 6032 37680 6048 37744
rect 6112 37680 6128 37744
rect 6192 37680 6208 37744
rect 6272 37680 6288 37744
rect 6352 37680 6368 37744
rect 6432 37680 6448 37744
rect 6512 37680 6528 37744
rect 6592 37680 6608 37744
rect 6672 37680 6688 37744
rect 6752 37680 6768 37744
rect 6832 37680 6848 37744
rect 6912 37680 6928 37744
rect 6992 37680 7008 37744
rect 7072 37680 7088 37744
rect 7152 37680 7168 37744
rect 7232 37680 7248 37744
rect 7312 37680 7328 37744
rect 7392 37680 7408 37744
rect 7472 37680 7488 37744
rect 7552 37680 7568 37744
rect 7632 37680 7648 37744
rect 7712 37680 7728 37744
rect 7792 37680 7808 37744
rect 7872 37680 7888 37744
rect 7952 37680 7968 37744
rect 8032 37680 8048 37744
rect 8112 37680 8128 37744
rect 8192 37680 8208 37744
rect 8272 37680 8288 37744
rect 8352 37680 8368 37744
rect 8432 37680 8448 37744
rect 8512 37680 8528 37744
rect 8592 37680 8608 37744
rect 8672 37680 8688 37744
rect 8752 37680 8768 37744
rect 8832 37680 8848 37744
rect 8912 37680 8928 37744
rect 8992 37680 14112 37744
rect 14176 37680 14192 37744
rect 14256 37680 14272 37744
rect 14336 37680 14352 37744
rect 14416 37680 24112 37744
rect 24176 37680 24192 37744
rect 24256 37680 24272 37744
rect 24336 37680 24352 37744
rect 24416 37680 36376 37744
rect 36440 37680 36456 37744
rect 36520 37680 36536 37744
rect 36600 37680 36616 37744
rect 36680 37680 36696 37744
rect 36760 37680 36776 37744
rect 36840 37680 36856 37744
rect 36920 37680 36936 37744
rect 37000 37680 37016 37744
rect 37080 37680 37096 37744
rect 37160 37680 37176 37744
rect 37240 37680 37256 37744
rect 37320 37680 37336 37744
rect 37400 37680 37416 37744
rect 37480 37680 37496 37744
rect 37560 37680 37576 37744
rect 37640 37680 37656 37744
rect 37720 37680 37736 37744
rect 37800 37680 37816 37744
rect 37880 37680 37896 37744
rect 37960 37680 37976 37744
rect 38040 37680 38056 37744
rect 38120 37680 38136 37744
rect 38200 37680 38216 37744
rect 38280 37680 38296 37744
rect 38360 37680 38376 37744
rect 38440 37680 38456 37744
rect 38520 37680 38536 37744
rect 38600 37680 38616 37744
rect 38680 37680 38696 37744
rect 38760 37680 38776 37744
rect 38840 37680 38856 37744
rect 38920 37680 38936 37744
rect 39000 37680 39016 37744
rect 39080 37680 39096 37744
rect 39160 37680 39176 37744
rect 39240 37680 39256 37744
rect 39320 37680 39336 37744
rect 39400 37680 39416 37744
rect 39480 37680 39496 37744
rect 39560 37680 39576 37744
rect 39640 37680 39656 37744
rect 39720 37680 39736 37744
rect 39800 37680 39816 37744
rect 39880 37680 39896 37744
rect 39960 37680 39976 37744
rect 40040 37680 40056 37744
rect 40120 37680 40136 37744
rect 40200 37680 40216 37744
rect 40280 37680 40296 37744
rect 40360 37680 40368 37744
rect 5000 37664 40368 37680
rect 5000 37600 5008 37664
rect 5072 37600 5088 37664
rect 5152 37600 5168 37664
rect 5232 37600 5248 37664
rect 5312 37600 5328 37664
rect 5392 37600 5408 37664
rect 5472 37600 5488 37664
rect 5552 37600 5568 37664
rect 5632 37600 5648 37664
rect 5712 37600 5728 37664
rect 5792 37600 5808 37664
rect 5872 37600 5888 37664
rect 5952 37600 5968 37664
rect 6032 37600 6048 37664
rect 6112 37600 6128 37664
rect 6192 37600 6208 37664
rect 6272 37600 6288 37664
rect 6352 37600 6368 37664
rect 6432 37600 6448 37664
rect 6512 37600 6528 37664
rect 6592 37600 6608 37664
rect 6672 37600 6688 37664
rect 6752 37600 6768 37664
rect 6832 37600 6848 37664
rect 6912 37600 6928 37664
rect 6992 37600 7008 37664
rect 7072 37600 7088 37664
rect 7152 37600 7168 37664
rect 7232 37600 7248 37664
rect 7312 37600 7328 37664
rect 7392 37600 7408 37664
rect 7472 37600 7488 37664
rect 7552 37600 7568 37664
rect 7632 37600 7648 37664
rect 7712 37600 7728 37664
rect 7792 37600 7808 37664
rect 7872 37600 7888 37664
rect 7952 37600 7968 37664
rect 8032 37600 8048 37664
rect 8112 37600 8128 37664
rect 8192 37600 8208 37664
rect 8272 37600 8288 37664
rect 8352 37600 8368 37664
rect 8432 37600 8448 37664
rect 8512 37600 8528 37664
rect 8592 37600 8608 37664
rect 8672 37600 8688 37664
rect 8752 37600 8768 37664
rect 8832 37600 8848 37664
rect 8912 37600 8928 37664
rect 8992 37600 14112 37664
rect 14176 37600 14192 37664
rect 14256 37600 14272 37664
rect 14336 37600 14352 37664
rect 14416 37600 24112 37664
rect 24176 37600 24192 37664
rect 24256 37600 24272 37664
rect 24336 37600 24352 37664
rect 24416 37600 36376 37664
rect 36440 37600 36456 37664
rect 36520 37600 36536 37664
rect 36600 37600 36616 37664
rect 36680 37600 36696 37664
rect 36760 37600 36776 37664
rect 36840 37600 36856 37664
rect 36920 37600 36936 37664
rect 37000 37600 37016 37664
rect 37080 37600 37096 37664
rect 37160 37600 37176 37664
rect 37240 37600 37256 37664
rect 37320 37600 37336 37664
rect 37400 37600 37416 37664
rect 37480 37600 37496 37664
rect 37560 37600 37576 37664
rect 37640 37600 37656 37664
rect 37720 37600 37736 37664
rect 37800 37600 37816 37664
rect 37880 37600 37896 37664
rect 37960 37600 37976 37664
rect 38040 37600 38056 37664
rect 38120 37600 38136 37664
rect 38200 37600 38216 37664
rect 38280 37600 38296 37664
rect 38360 37600 38376 37664
rect 38440 37600 38456 37664
rect 38520 37600 38536 37664
rect 38600 37600 38616 37664
rect 38680 37600 38696 37664
rect 38760 37600 38776 37664
rect 38840 37600 38856 37664
rect 38920 37600 38936 37664
rect 39000 37600 39016 37664
rect 39080 37600 39096 37664
rect 39160 37600 39176 37664
rect 39240 37600 39256 37664
rect 39320 37600 39336 37664
rect 39400 37600 39416 37664
rect 39480 37600 39496 37664
rect 39560 37600 39576 37664
rect 39640 37600 39656 37664
rect 39720 37600 39736 37664
rect 39800 37600 39816 37664
rect 39880 37600 39896 37664
rect 39960 37600 39976 37664
rect 40040 37600 40056 37664
rect 40120 37600 40136 37664
rect 40200 37600 40216 37664
rect 40280 37600 40296 37664
rect 40360 37600 40368 37664
rect 5000 37584 40368 37600
rect 5000 37520 5008 37584
rect 5072 37520 5088 37584
rect 5152 37520 5168 37584
rect 5232 37520 5248 37584
rect 5312 37520 5328 37584
rect 5392 37520 5408 37584
rect 5472 37520 5488 37584
rect 5552 37520 5568 37584
rect 5632 37520 5648 37584
rect 5712 37520 5728 37584
rect 5792 37520 5808 37584
rect 5872 37520 5888 37584
rect 5952 37520 5968 37584
rect 6032 37520 6048 37584
rect 6112 37520 6128 37584
rect 6192 37520 6208 37584
rect 6272 37520 6288 37584
rect 6352 37520 6368 37584
rect 6432 37520 6448 37584
rect 6512 37520 6528 37584
rect 6592 37520 6608 37584
rect 6672 37520 6688 37584
rect 6752 37520 6768 37584
rect 6832 37520 6848 37584
rect 6912 37520 6928 37584
rect 6992 37520 7008 37584
rect 7072 37520 7088 37584
rect 7152 37520 7168 37584
rect 7232 37520 7248 37584
rect 7312 37520 7328 37584
rect 7392 37520 7408 37584
rect 7472 37520 7488 37584
rect 7552 37520 7568 37584
rect 7632 37520 7648 37584
rect 7712 37520 7728 37584
rect 7792 37520 7808 37584
rect 7872 37520 7888 37584
rect 7952 37520 7968 37584
rect 8032 37520 8048 37584
rect 8112 37520 8128 37584
rect 8192 37520 8208 37584
rect 8272 37520 8288 37584
rect 8352 37520 8368 37584
rect 8432 37520 8448 37584
rect 8512 37520 8528 37584
rect 8592 37520 8608 37584
rect 8672 37520 8688 37584
rect 8752 37520 8768 37584
rect 8832 37520 8848 37584
rect 8912 37520 8928 37584
rect 8992 37520 14112 37584
rect 14176 37520 14192 37584
rect 14256 37520 14272 37584
rect 14336 37520 14352 37584
rect 14416 37520 24112 37584
rect 24176 37520 24192 37584
rect 24256 37520 24272 37584
rect 24336 37520 24352 37584
rect 24416 37520 36376 37584
rect 36440 37520 36456 37584
rect 36520 37520 36536 37584
rect 36600 37520 36616 37584
rect 36680 37520 36696 37584
rect 36760 37520 36776 37584
rect 36840 37520 36856 37584
rect 36920 37520 36936 37584
rect 37000 37520 37016 37584
rect 37080 37520 37096 37584
rect 37160 37520 37176 37584
rect 37240 37520 37256 37584
rect 37320 37520 37336 37584
rect 37400 37520 37416 37584
rect 37480 37520 37496 37584
rect 37560 37520 37576 37584
rect 37640 37520 37656 37584
rect 37720 37520 37736 37584
rect 37800 37520 37816 37584
rect 37880 37520 37896 37584
rect 37960 37520 37976 37584
rect 38040 37520 38056 37584
rect 38120 37520 38136 37584
rect 38200 37520 38216 37584
rect 38280 37520 38296 37584
rect 38360 37520 38376 37584
rect 38440 37520 38456 37584
rect 38520 37520 38536 37584
rect 38600 37520 38616 37584
rect 38680 37520 38696 37584
rect 38760 37520 38776 37584
rect 38840 37520 38856 37584
rect 38920 37520 38936 37584
rect 39000 37520 39016 37584
rect 39080 37520 39096 37584
rect 39160 37520 39176 37584
rect 39240 37520 39256 37584
rect 39320 37520 39336 37584
rect 39400 37520 39416 37584
rect 39480 37520 39496 37584
rect 39560 37520 39576 37584
rect 39640 37520 39656 37584
rect 39720 37520 39736 37584
rect 39800 37520 39816 37584
rect 39880 37520 39896 37584
rect 39960 37520 39976 37584
rect 40040 37520 40056 37584
rect 40120 37520 40136 37584
rect 40200 37520 40216 37584
rect 40280 37520 40296 37584
rect 40360 37520 40368 37584
rect 5000 37504 40368 37520
rect 5000 37440 5008 37504
rect 5072 37440 5088 37504
rect 5152 37440 5168 37504
rect 5232 37440 5248 37504
rect 5312 37440 5328 37504
rect 5392 37440 5408 37504
rect 5472 37440 5488 37504
rect 5552 37440 5568 37504
rect 5632 37440 5648 37504
rect 5712 37440 5728 37504
rect 5792 37440 5808 37504
rect 5872 37440 5888 37504
rect 5952 37440 5968 37504
rect 6032 37440 6048 37504
rect 6112 37440 6128 37504
rect 6192 37440 6208 37504
rect 6272 37440 6288 37504
rect 6352 37440 6368 37504
rect 6432 37440 6448 37504
rect 6512 37440 6528 37504
rect 6592 37440 6608 37504
rect 6672 37440 6688 37504
rect 6752 37440 6768 37504
rect 6832 37440 6848 37504
rect 6912 37440 6928 37504
rect 6992 37440 7008 37504
rect 7072 37440 7088 37504
rect 7152 37440 7168 37504
rect 7232 37440 7248 37504
rect 7312 37440 7328 37504
rect 7392 37440 7408 37504
rect 7472 37440 7488 37504
rect 7552 37440 7568 37504
rect 7632 37440 7648 37504
rect 7712 37440 7728 37504
rect 7792 37440 7808 37504
rect 7872 37440 7888 37504
rect 7952 37440 7968 37504
rect 8032 37440 8048 37504
rect 8112 37440 8128 37504
rect 8192 37440 8208 37504
rect 8272 37440 8288 37504
rect 8352 37440 8368 37504
rect 8432 37440 8448 37504
rect 8512 37440 8528 37504
rect 8592 37440 8608 37504
rect 8672 37440 8688 37504
rect 8752 37440 8768 37504
rect 8832 37440 8848 37504
rect 8912 37440 8928 37504
rect 8992 37440 14112 37504
rect 14176 37440 14192 37504
rect 14256 37440 14272 37504
rect 14336 37440 14352 37504
rect 14416 37440 24112 37504
rect 24176 37440 24192 37504
rect 24256 37440 24272 37504
rect 24336 37440 24352 37504
rect 24416 37440 36376 37504
rect 36440 37440 36456 37504
rect 36520 37440 36536 37504
rect 36600 37440 36616 37504
rect 36680 37440 36696 37504
rect 36760 37440 36776 37504
rect 36840 37440 36856 37504
rect 36920 37440 36936 37504
rect 37000 37440 37016 37504
rect 37080 37440 37096 37504
rect 37160 37440 37176 37504
rect 37240 37440 37256 37504
rect 37320 37440 37336 37504
rect 37400 37440 37416 37504
rect 37480 37440 37496 37504
rect 37560 37440 37576 37504
rect 37640 37440 37656 37504
rect 37720 37440 37736 37504
rect 37800 37440 37816 37504
rect 37880 37440 37896 37504
rect 37960 37440 37976 37504
rect 38040 37440 38056 37504
rect 38120 37440 38136 37504
rect 38200 37440 38216 37504
rect 38280 37440 38296 37504
rect 38360 37440 38376 37504
rect 38440 37440 38456 37504
rect 38520 37440 38536 37504
rect 38600 37440 38616 37504
rect 38680 37440 38696 37504
rect 38760 37440 38776 37504
rect 38840 37440 38856 37504
rect 38920 37440 38936 37504
rect 39000 37440 39016 37504
rect 39080 37440 39096 37504
rect 39160 37440 39176 37504
rect 39240 37440 39256 37504
rect 39320 37440 39336 37504
rect 39400 37440 39416 37504
rect 39480 37440 39496 37504
rect 39560 37440 39576 37504
rect 39640 37440 39656 37504
rect 39720 37440 39736 37504
rect 39800 37440 39816 37504
rect 39880 37440 39896 37504
rect 39960 37440 39976 37504
rect 40040 37440 40056 37504
rect 40120 37440 40136 37504
rect 40200 37440 40216 37504
rect 40280 37440 40296 37504
rect 40360 37440 40368 37504
rect 5000 37424 40368 37440
rect 5000 37360 5008 37424
rect 5072 37360 5088 37424
rect 5152 37360 5168 37424
rect 5232 37360 5248 37424
rect 5312 37360 5328 37424
rect 5392 37360 5408 37424
rect 5472 37360 5488 37424
rect 5552 37360 5568 37424
rect 5632 37360 5648 37424
rect 5712 37360 5728 37424
rect 5792 37360 5808 37424
rect 5872 37360 5888 37424
rect 5952 37360 5968 37424
rect 6032 37360 6048 37424
rect 6112 37360 6128 37424
rect 6192 37360 6208 37424
rect 6272 37360 6288 37424
rect 6352 37360 6368 37424
rect 6432 37360 6448 37424
rect 6512 37360 6528 37424
rect 6592 37360 6608 37424
rect 6672 37360 6688 37424
rect 6752 37360 6768 37424
rect 6832 37360 6848 37424
rect 6912 37360 6928 37424
rect 6992 37360 7008 37424
rect 7072 37360 7088 37424
rect 7152 37360 7168 37424
rect 7232 37360 7248 37424
rect 7312 37360 7328 37424
rect 7392 37360 7408 37424
rect 7472 37360 7488 37424
rect 7552 37360 7568 37424
rect 7632 37360 7648 37424
rect 7712 37360 7728 37424
rect 7792 37360 7808 37424
rect 7872 37360 7888 37424
rect 7952 37360 7968 37424
rect 8032 37360 8048 37424
rect 8112 37360 8128 37424
rect 8192 37360 8208 37424
rect 8272 37360 8288 37424
rect 8352 37360 8368 37424
rect 8432 37360 8448 37424
rect 8512 37360 8528 37424
rect 8592 37360 8608 37424
rect 8672 37360 8688 37424
rect 8752 37360 8768 37424
rect 8832 37360 8848 37424
rect 8912 37360 8928 37424
rect 8992 37360 14112 37424
rect 14176 37360 14192 37424
rect 14256 37360 14272 37424
rect 14336 37360 14352 37424
rect 14416 37360 24112 37424
rect 24176 37360 24192 37424
rect 24256 37360 24272 37424
rect 24336 37360 24352 37424
rect 24416 37360 36376 37424
rect 36440 37360 36456 37424
rect 36520 37360 36536 37424
rect 36600 37360 36616 37424
rect 36680 37360 36696 37424
rect 36760 37360 36776 37424
rect 36840 37360 36856 37424
rect 36920 37360 36936 37424
rect 37000 37360 37016 37424
rect 37080 37360 37096 37424
rect 37160 37360 37176 37424
rect 37240 37360 37256 37424
rect 37320 37360 37336 37424
rect 37400 37360 37416 37424
rect 37480 37360 37496 37424
rect 37560 37360 37576 37424
rect 37640 37360 37656 37424
rect 37720 37360 37736 37424
rect 37800 37360 37816 37424
rect 37880 37360 37896 37424
rect 37960 37360 37976 37424
rect 38040 37360 38056 37424
rect 38120 37360 38136 37424
rect 38200 37360 38216 37424
rect 38280 37360 38296 37424
rect 38360 37360 38376 37424
rect 38440 37360 38456 37424
rect 38520 37360 38536 37424
rect 38600 37360 38616 37424
rect 38680 37360 38696 37424
rect 38760 37360 38776 37424
rect 38840 37360 38856 37424
rect 38920 37360 38936 37424
rect 39000 37360 39016 37424
rect 39080 37360 39096 37424
rect 39160 37360 39176 37424
rect 39240 37360 39256 37424
rect 39320 37360 39336 37424
rect 39400 37360 39416 37424
rect 39480 37360 39496 37424
rect 39560 37360 39576 37424
rect 39640 37360 39656 37424
rect 39720 37360 39736 37424
rect 39800 37360 39816 37424
rect 39880 37360 39896 37424
rect 39960 37360 39976 37424
rect 40040 37360 40056 37424
rect 40120 37360 40136 37424
rect 40200 37360 40216 37424
rect 40280 37360 40296 37424
rect 40360 37360 40368 37424
rect 5000 37344 40368 37360
rect 5000 37280 5008 37344
rect 5072 37280 5088 37344
rect 5152 37280 5168 37344
rect 5232 37280 5248 37344
rect 5312 37280 5328 37344
rect 5392 37280 5408 37344
rect 5472 37280 5488 37344
rect 5552 37280 5568 37344
rect 5632 37280 5648 37344
rect 5712 37280 5728 37344
rect 5792 37280 5808 37344
rect 5872 37280 5888 37344
rect 5952 37280 5968 37344
rect 6032 37280 6048 37344
rect 6112 37280 6128 37344
rect 6192 37280 6208 37344
rect 6272 37280 6288 37344
rect 6352 37280 6368 37344
rect 6432 37280 6448 37344
rect 6512 37280 6528 37344
rect 6592 37280 6608 37344
rect 6672 37280 6688 37344
rect 6752 37280 6768 37344
rect 6832 37280 6848 37344
rect 6912 37280 6928 37344
rect 6992 37280 7008 37344
rect 7072 37280 7088 37344
rect 7152 37280 7168 37344
rect 7232 37280 7248 37344
rect 7312 37280 7328 37344
rect 7392 37280 7408 37344
rect 7472 37280 7488 37344
rect 7552 37280 7568 37344
rect 7632 37280 7648 37344
rect 7712 37280 7728 37344
rect 7792 37280 7808 37344
rect 7872 37280 7888 37344
rect 7952 37280 7968 37344
rect 8032 37280 8048 37344
rect 8112 37280 8128 37344
rect 8192 37280 8208 37344
rect 8272 37280 8288 37344
rect 8352 37280 8368 37344
rect 8432 37280 8448 37344
rect 8512 37280 8528 37344
rect 8592 37280 8608 37344
rect 8672 37280 8688 37344
rect 8752 37280 8768 37344
rect 8832 37280 8848 37344
rect 8912 37280 8928 37344
rect 8992 37280 14112 37344
rect 14176 37280 14192 37344
rect 14256 37280 14272 37344
rect 14336 37280 14352 37344
rect 14416 37280 24112 37344
rect 24176 37280 24192 37344
rect 24256 37280 24272 37344
rect 24336 37280 24352 37344
rect 24416 37280 36376 37344
rect 36440 37280 36456 37344
rect 36520 37280 36536 37344
rect 36600 37280 36616 37344
rect 36680 37280 36696 37344
rect 36760 37280 36776 37344
rect 36840 37280 36856 37344
rect 36920 37280 36936 37344
rect 37000 37280 37016 37344
rect 37080 37280 37096 37344
rect 37160 37280 37176 37344
rect 37240 37280 37256 37344
rect 37320 37280 37336 37344
rect 37400 37280 37416 37344
rect 37480 37280 37496 37344
rect 37560 37280 37576 37344
rect 37640 37280 37656 37344
rect 37720 37280 37736 37344
rect 37800 37280 37816 37344
rect 37880 37280 37896 37344
rect 37960 37280 37976 37344
rect 38040 37280 38056 37344
rect 38120 37280 38136 37344
rect 38200 37280 38216 37344
rect 38280 37280 38296 37344
rect 38360 37280 38376 37344
rect 38440 37280 38456 37344
rect 38520 37280 38536 37344
rect 38600 37280 38616 37344
rect 38680 37280 38696 37344
rect 38760 37280 38776 37344
rect 38840 37280 38856 37344
rect 38920 37280 38936 37344
rect 39000 37280 39016 37344
rect 39080 37280 39096 37344
rect 39160 37280 39176 37344
rect 39240 37280 39256 37344
rect 39320 37280 39336 37344
rect 39400 37280 39416 37344
rect 39480 37280 39496 37344
rect 39560 37280 39576 37344
rect 39640 37280 39656 37344
rect 39720 37280 39736 37344
rect 39800 37280 39816 37344
rect 39880 37280 39896 37344
rect 39960 37280 39976 37344
rect 40040 37280 40056 37344
rect 40120 37280 40136 37344
rect 40200 37280 40216 37344
rect 40280 37280 40296 37344
rect 40360 37280 40368 37344
rect 5000 37264 40368 37280
rect 5000 37200 5008 37264
rect 5072 37200 5088 37264
rect 5152 37200 5168 37264
rect 5232 37200 5248 37264
rect 5312 37200 5328 37264
rect 5392 37200 5408 37264
rect 5472 37200 5488 37264
rect 5552 37200 5568 37264
rect 5632 37200 5648 37264
rect 5712 37200 5728 37264
rect 5792 37200 5808 37264
rect 5872 37200 5888 37264
rect 5952 37200 5968 37264
rect 6032 37200 6048 37264
rect 6112 37200 6128 37264
rect 6192 37200 6208 37264
rect 6272 37200 6288 37264
rect 6352 37200 6368 37264
rect 6432 37200 6448 37264
rect 6512 37200 6528 37264
rect 6592 37200 6608 37264
rect 6672 37200 6688 37264
rect 6752 37200 6768 37264
rect 6832 37200 6848 37264
rect 6912 37200 6928 37264
rect 6992 37200 7008 37264
rect 7072 37200 7088 37264
rect 7152 37200 7168 37264
rect 7232 37200 7248 37264
rect 7312 37200 7328 37264
rect 7392 37200 7408 37264
rect 7472 37200 7488 37264
rect 7552 37200 7568 37264
rect 7632 37200 7648 37264
rect 7712 37200 7728 37264
rect 7792 37200 7808 37264
rect 7872 37200 7888 37264
rect 7952 37200 7968 37264
rect 8032 37200 8048 37264
rect 8112 37200 8128 37264
rect 8192 37200 8208 37264
rect 8272 37200 8288 37264
rect 8352 37200 8368 37264
rect 8432 37200 8448 37264
rect 8512 37200 8528 37264
rect 8592 37200 8608 37264
rect 8672 37200 8688 37264
rect 8752 37200 8768 37264
rect 8832 37200 8848 37264
rect 8912 37200 8928 37264
rect 8992 37200 14112 37264
rect 14176 37200 14192 37264
rect 14256 37200 14272 37264
rect 14336 37200 14352 37264
rect 14416 37200 24112 37264
rect 24176 37200 24192 37264
rect 24256 37200 24272 37264
rect 24336 37200 24352 37264
rect 24416 37200 36376 37264
rect 36440 37200 36456 37264
rect 36520 37200 36536 37264
rect 36600 37200 36616 37264
rect 36680 37200 36696 37264
rect 36760 37200 36776 37264
rect 36840 37200 36856 37264
rect 36920 37200 36936 37264
rect 37000 37200 37016 37264
rect 37080 37200 37096 37264
rect 37160 37200 37176 37264
rect 37240 37200 37256 37264
rect 37320 37200 37336 37264
rect 37400 37200 37416 37264
rect 37480 37200 37496 37264
rect 37560 37200 37576 37264
rect 37640 37200 37656 37264
rect 37720 37200 37736 37264
rect 37800 37200 37816 37264
rect 37880 37200 37896 37264
rect 37960 37200 37976 37264
rect 38040 37200 38056 37264
rect 38120 37200 38136 37264
rect 38200 37200 38216 37264
rect 38280 37200 38296 37264
rect 38360 37200 38376 37264
rect 38440 37200 38456 37264
rect 38520 37200 38536 37264
rect 38600 37200 38616 37264
rect 38680 37200 38696 37264
rect 38760 37200 38776 37264
rect 38840 37200 38856 37264
rect 38920 37200 38936 37264
rect 39000 37200 39016 37264
rect 39080 37200 39096 37264
rect 39160 37200 39176 37264
rect 39240 37200 39256 37264
rect 39320 37200 39336 37264
rect 39400 37200 39416 37264
rect 39480 37200 39496 37264
rect 39560 37200 39576 37264
rect 39640 37200 39656 37264
rect 39720 37200 39736 37264
rect 39800 37200 39816 37264
rect 39880 37200 39896 37264
rect 39960 37200 39976 37264
rect 40040 37200 40056 37264
rect 40120 37200 40136 37264
rect 40200 37200 40216 37264
rect 40280 37200 40296 37264
rect 40360 37200 40368 37264
rect 5000 37184 40368 37200
rect 5000 37120 5008 37184
rect 5072 37120 5088 37184
rect 5152 37120 5168 37184
rect 5232 37120 5248 37184
rect 5312 37120 5328 37184
rect 5392 37120 5408 37184
rect 5472 37120 5488 37184
rect 5552 37120 5568 37184
rect 5632 37120 5648 37184
rect 5712 37120 5728 37184
rect 5792 37120 5808 37184
rect 5872 37120 5888 37184
rect 5952 37120 5968 37184
rect 6032 37120 6048 37184
rect 6112 37120 6128 37184
rect 6192 37120 6208 37184
rect 6272 37120 6288 37184
rect 6352 37120 6368 37184
rect 6432 37120 6448 37184
rect 6512 37120 6528 37184
rect 6592 37120 6608 37184
rect 6672 37120 6688 37184
rect 6752 37120 6768 37184
rect 6832 37120 6848 37184
rect 6912 37120 6928 37184
rect 6992 37120 7008 37184
rect 7072 37120 7088 37184
rect 7152 37120 7168 37184
rect 7232 37120 7248 37184
rect 7312 37120 7328 37184
rect 7392 37120 7408 37184
rect 7472 37120 7488 37184
rect 7552 37120 7568 37184
rect 7632 37120 7648 37184
rect 7712 37120 7728 37184
rect 7792 37120 7808 37184
rect 7872 37120 7888 37184
rect 7952 37120 7968 37184
rect 8032 37120 8048 37184
rect 8112 37120 8128 37184
rect 8192 37120 8208 37184
rect 8272 37120 8288 37184
rect 8352 37120 8368 37184
rect 8432 37120 8448 37184
rect 8512 37120 8528 37184
rect 8592 37120 8608 37184
rect 8672 37120 8688 37184
rect 8752 37120 8768 37184
rect 8832 37120 8848 37184
rect 8912 37120 8928 37184
rect 8992 37120 14112 37184
rect 14176 37120 14192 37184
rect 14256 37120 14272 37184
rect 14336 37120 14352 37184
rect 14416 37120 24112 37184
rect 24176 37120 24192 37184
rect 24256 37120 24272 37184
rect 24336 37120 24352 37184
rect 24416 37120 36376 37184
rect 36440 37120 36456 37184
rect 36520 37120 36536 37184
rect 36600 37120 36616 37184
rect 36680 37120 36696 37184
rect 36760 37120 36776 37184
rect 36840 37120 36856 37184
rect 36920 37120 36936 37184
rect 37000 37120 37016 37184
rect 37080 37120 37096 37184
rect 37160 37120 37176 37184
rect 37240 37120 37256 37184
rect 37320 37120 37336 37184
rect 37400 37120 37416 37184
rect 37480 37120 37496 37184
rect 37560 37120 37576 37184
rect 37640 37120 37656 37184
rect 37720 37120 37736 37184
rect 37800 37120 37816 37184
rect 37880 37120 37896 37184
rect 37960 37120 37976 37184
rect 38040 37120 38056 37184
rect 38120 37120 38136 37184
rect 38200 37120 38216 37184
rect 38280 37120 38296 37184
rect 38360 37120 38376 37184
rect 38440 37120 38456 37184
rect 38520 37120 38536 37184
rect 38600 37120 38616 37184
rect 38680 37120 38696 37184
rect 38760 37120 38776 37184
rect 38840 37120 38856 37184
rect 38920 37120 38936 37184
rect 39000 37120 39016 37184
rect 39080 37120 39096 37184
rect 39160 37120 39176 37184
rect 39240 37120 39256 37184
rect 39320 37120 39336 37184
rect 39400 37120 39416 37184
rect 39480 37120 39496 37184
rect 39560 37120 39576 37184
rect 39640 37120 39656 37184
rect 39720 37120 39736 37184
rect 39800 37120 39816 37184
rect 39880 37120 39896 37184
rect 39960 37120 39976 37184
rect 40040 37120 40056 37184
rect 40120 37120 40136 37184
rect 40200 37120 40216 37184
rect 40280 37120 40296 37184
rect 40360 37120 40368 37184
rect 5000 37104 40368 37120
rect 5000 37040 5008 37104
rect 5072 37040 5088 37104
rect 5152 37040 5168 37104
rect 5232 37040 5248 37104
rect 5312 37040 5328 37104
rect 5392 37040 5408 37104
rect 5472 37040 5488 37104
rect 5552 37040 5568 37104
rect 5632 37040 5648 37104
rect 5712 37040 5728 37104
rect 5792 37040 5808 37104
rect 5872 37040 5888 37104
rect 5952 37040 5968 37104
rect 6032 37040 6048 37104
rect 6112 37040 6128 37104
rect 6192 37040 6208 37104
rect 6272 37040 6288 37104
rect 6352 37040 6368 37104
rect 6432 37040 6448 37104
rect 6512 37040 6528 37104
rect 6592 37040 6608 37104
rect 6672 37040 6688 37104
rect 6752 37040 6768 37104
rect 6832 37040 6848 37104
rect 6912 37040 6928 37104
rect 6992 37040 7008 37104
rect 7072 37040 7088 37104
rect 7152 37040 7168 37104
rect 7232 37040 7248 37104
rect 7312 37040 7328 37104
rect 7392 37040 7408 37104
rect 7472 37040 7488 37104
rect 7552 37040 7568 37104
rect 7632 37040 7648 37104
rect 7712 37040 7728 37104
rect 7792 37040 7808 37104
rect 7872 37040 7888 37104
rect 7952 37040 7968 37104
rect 8032 37040 8048 37104
rect 8112 37040 8128 37104
rect 8192 37040 8208 37104
rect 8272 37040 8288 37104
rect 8352 37040 8368 37104
rect 8432 37040 8448 37104
rect 8512 37040 8528 37104
rect 8592 37040 8608 37104
rect 8672 37040 8688 37104
rect 8752 37040 8768 37104
rect 8832 37040 8848 37104
rect 8912 37040 8928 37104
rect 8992 37040 14112 37104
rect 14176 37040 14192 37104
rect 14256 37040 14272 37104
rect 14336 37040 14352 37104
rect 14416 37040 24112 37104
rect 24176 37040 24192 37104
rect 24256 37040 24272 37104
rect 24336 37040 24352 37104
rect 24416 37040 36376 37104
rect 36440 37040 36456 37104
rect 36520 37040 36536 37104
rect 36600 37040 36616 37104
rect 36680 37040 36696 37104
rect 36760 37040 36776 37104
rect 36840 37040 36856 37104
rect 36920 37040 36936 37104
rect 37000 37040 37016 37104
rect 37080 37040 37096 37104
rect 37160 37040 37176 37104
rect 37240 37040 37256 37104
rect 37320 37040 37336 37104
rect 37400 37040 37416 37104
rect 37480 37040 37496 37104
rect 37560 37040 37576 37104
rect 37640 37040 37656 37104
rect 37720 37040 37736 37104
rect 37800 37040 37816 37104
rect 37880 37040 37896 37104
rect 37960 37040 37976 37104
rect 38040 37040 38056 37104
rect 38120 37040 38136 37104
rect 38200 37040 38216 37104
rect 38280 37040 38296 37104
rect 38360 37040 38376 37104
rect 38440 37040 38456 37104
rect 38520 37040 38536 37104
rect 38600 37040 38616 37104
rect 38680 37040 38696 37104
rect 38760 37040 38776 37104
rect 38840 37040 38856 37104
rect 38920 37040 38936 37104
rect 39000 37040 39016 37104
rect 39080 37040 39096 37104
rect 39160 37040 39176 37104
rect 39240 37040 39256 37104
rect 39320 37040 39336 37104
rect 39400 37040 39416 37104
rect 39480 37040 39496 37104
rect 39560 37040 39576 37104
rect 39640 37040 39656 37104
rect 39720 37040 39736 37104
rect 39800 37040 39816 37104
rect 39880 37040 39896 37104
rect 39960 37040 39976 37104
rect 40040 37040 40056 37104
rect 40120 37040 40136 37104
rect 40200 37040 40216 37104
rect 40280 37040 40296 37104
rect 40360 37040 40368 37104
rect 5000 37024 40368 37040
rect 5000 36960 5008 37024
rect 5072 36960 5088 37024
rect 5152 36960 5168 37024
rect 5232 36960 5248 37024
rect 5312 36960 5328 37024
rect 5392 36960 5408 37024
rect 5472 36960 5488 37024
rect 5552 36960 5568 37024
rect 5632 36960 5648 37024
rect 5712 36960 5728 37024
rect 5792 36960 5808 37024
rect 5872 36960 5888 37024
rect 5952 36960 5968 37024
rect 6032 36960 6048 37024
rect 6112 36960 6128 37024
rect 6192 36960 6208 37024
rect 6272 36960 6288 37024
rect 6352 36960 6368 37024
rect 6432 36960 6448 37024
rect 6512 36960 6528 37024
rect 6592 36960 6608 37024
rect 6672 36960 6688 37024
rect 6752 36960 6768 37024
rect 6832 36960 6848 37024
rect 6912 36960 6928 37024
rect 6992 36960 7008 37024
rect 7072 36960 7088 37024
rect 7152 36960 7168 37024
rect 7232 36960 7248 37024
rect 7312 36960 7328 37024
rect 7392 36960 7408 37024
rect 7472 36960 7488 37024
rect 7552 36960 7568 37024
rect 7632 36960 7648 37024
rect 7712 36960 7728 37024
rect 7792 36960 7808 37024
rect 7872 36960 7888 37024
rect 7952 36960 7968 37024
rect 8032 36960 8048 37024
rect 8112 36960 8128 37024
rect 8192 36960 8208 37024
rect 8272 36960 8288 37024
rect 8352 36960 8368 37024
rect 8432 36960 8448 37024
rect 8512 36960 8528 37024
rect 8592 36960 8608 37024
rect 8672 36960 8688 37024
rect 8752 36960 8768 37024
rect 8832 36960 8848 37024
rect 8912 36960 8928 37024
rect 8992 36960 14112 37024
rect 14176 36960 14192 37024
rect 14256 36960 14272 37024
rect 14336 36960 14352 37024
rect 14416 36960 24112 37024
rect 24176 36960 24192 37024
rect 24256 36960 24272 37024
rect 24336 36960 24352 37024
rect 24416 36960 36376 37024
rect 36440 36960 36456 37024
rect 36520 36960 36536 37024
rect 36600 36960 36616 37024
rect 36680 36960 36696 37024
rect 36760 36960 36776 37024
rect 36840 36960 36856 37024
rect 36920 36960 36936 37024
rect 37000 36960 37016 37024
rect 37080 36960 37096 37024
rect 37160 36960 37176 37024
rect 37240 36960 37256 37024
rect 37320 36960 37336 37024
rect 37400 36960 37416 37024
rect 37480 36960 37496 37024
rect 37560 36960 37576 37024
rect 37640 36960 37656 37024
rect 37720 36960 37736 37024
rect 37800 36960 37816 37024
rect 37880 36960 37896 37024
rect 37960 36960 37976 37024
rect 38040 36960 38056 37024
rect 38120 36960 38136 37024
rect 38200 36960 38216 37024
rect 38280 36960 38296 37024
rect 38360 36960 38376 37024
rect 38440 36960 38456 37024
rect 38520 36960 38536 37024
rect 38600 36960 38616 37024
rect 38680 36960 38696 37024
rect 38760 36960 38776 37024
rect 38840 36960 38856 37024
rect 38920 36960 38936 37024
rect 39000 36960 39016 37024
rect 39080 36960 39096 37024
rect 39160 36960 39176 37024
rect 39240 36960 39256 37024
rect 39320 36960 39336 37024
rect 39400 36960 39416 37024
rect 39480 36960 39496 37024
rect 39560 36960 39576 37024
rect 39640 36960 39656 37024
rect 39720 36960 39736 37024
rect 39800 36960 39816 37024
rect 39880 36960 39896 37024
rect 39960 36960 39976 37024
rect 40040 36960 40056 37024
rect 40120 36960 40136 37024
rect 40200 36960 40216 37024
rect 40280 36960 40296 37024
rect 40360 36960 40368 37024
rect 5000 36944 40368 36960
rect 5000 36880 5008 36944
rect 5072 36880 5088 36944
rect 5152 36880 5168 36944
rect 5232 36880 5248 36944
rect 5312 36880 5328 36944
rect 5392 36880 5408 36944
rect 5472 36880 5488 36944
rect 5552 36880 5568 36944
rect 5632 36880 5648 36944
rect 5712 36880 5728 36944
rect 5792 36880 5808 36944
rect 5872 36880 5888 36944
rect 5952 36880 5968 36944
rect 6032 36880 6048 36944
rect 6112 36880 6128 36944
rect 6192 36880 6208 36944
rect 6272 36880 6288 36944
rect 6352 36880 6368 36944
rect 6432 36880 6448 36944
rect 6512 36880 6528 36944
rect 6592 36880 6608 36944
rect 6672 36880 6688 36944
rect 6752 36880 6768 36944
rect 6832 36880 6848 36944
rect 6912 36880 6928 36944
rect 6992 36880 7008 36944
rect 7072 36880 7088 36944
rect 7152 36880 7168 36944
rect 7232 36880 7248 36944
rect 7312 36880 7328 36944
rect 7392 36880 7408 36944
rect 7472 36880 7488 36944
rect 7552 36880 7568 36944
rect 7632 36880 7648 36944
rect 7712 36880 7728 36944
rect 7792 36880 7808 36944
rect 7872 36880 7888 36944
rect 7952 36880 7968 36944
rect 8032 36880 8048 36944
rect 8112 36880 8128 36944
rect 8192 36880 8208 36944
rect 8272 36880 8288 36944
rect 8352 36880 8368 36944
rect 8432 36880 8448 36944
rect 8512 36880 8528 36944
rect 8592 36880 8608 36944
rect 8672 36880 8688 36944
rect 8752 36880 8768 36944
rect 8832 36880 8848 36944
rect 8912 36880 8928 36944
rect 8992 36880 14112 36944
rect 14176 36880 14192 36944
rect 14256 36880 14272 36944
rect 14336 36880 14352 36944
rect 14416 36880 24112 36944
rect 24176 36880 24192 36944
rect 24256 36880 24272 36944
rect 24336 36880 24352 36944
rect 24416 36880 36376 36944
rect 36440 36880 36456 36944
rect 36520 36880 36536 36944
rect 36600 36880 36616 36944
rect 36680 36880 36696 36944
rect 36760 36880 36776 36944
rect 36840 36880 36856 36944
rect 36920 36880 36936 36944
rect 37000 36880 37016 36944
rect 37080 36880 37096 36944
rect 37160 36880 37176 36944
rect 37240 36880 37256 36944
rect 37320 36880 37336 36944
rect 37400 36880 37416 36944
rect 37480 36880 37496 36944
rect 37560 36880 37576 36944
rect 37640 36880 37656 36944
rect 37720 36880 37736 36944
rect 37800 36880 37816 36944
rect 37880 36880 37896 36944
rect 37960 36880 37976 36944
rect 38040 36880 38056 36944
rect 38120 36880 38136 36944
rect 38200 36880 38216 36944
rect 38280 36880 38296 36944
rect 38360 36880 38376 36944
rect 38440 36880 38456 36944
rect 38520 36880 38536 36944
rect 38600 36880 38616 36944
rect 38680 36880 38696 36944
rect 38760 36880 38776 36944
rect 38840 36880 38856 36944
rect 38920 36880 38936 36944
rect 39000 36880 39016 36944
rect 39080 36880 39096 36944
rect 39160 36880 39176 36944
rect 39240 36880 39256 36944
rect 39320 36880 39336 36944
rect 39400 36880 39416 36944
rect 39480 36880 39496 36944
rect 39560 36880 39576 36944
rect 39640 36880 39656 36944
rect 39720 36880 39736 36944
rect 39800 36880 39816 36944
rect 39880 36880 39896 36944
rect 39960 36880 39976 36944
rect 40040 36880 40056 36944
rect 40120 36880 40136 36944
rect 40200 36880 40216 36944
rect 40280 36880 40296 36944
rect 40360 36880 40368 36944
rect 5000 36864 40368 36880
rect 5000 36800 5008 36864
rect 5072 36800 5088 36864
rect 5152 36800 5168 36864
rect 5232 36800 5248 36864
rect 5312 36800 5328 36864
rect 5392 36800 5408 36864
rect 5472 36800 5488 36864
rect 5552 36800 5568 36864
rect 5632 36800 5648 36864
rect 5712 36800 5728 36864
rect 5792 36800 5808 36864
rect 5872 36800 5888 36864
rect 5952 36800 5968 36864
rect 6032 36800 6048 36864
rect 6112 36800 6128 36864
rect 6192 36800 6208 36864
rect 6272 36800 6288 36864
rect 6352 36800 6368 36864
rect 6432 36800 6448 36864
rect 6512 36800 6528 36864
rect 6592 36800 6608 36864
rect 6672 36800 6688 36864
rect 6752 36800 6768 36864
rect 6832 36800 6848 36864
rect 6912 36800 6928 36864
rect 6992 36800 7008 36864
rect 7072 36800 7088 36864
rect 7152 36800 7168 36864
rect 7232 36800 7248 36864
rect 7312 36800 7328 36864
rect 7392 36800 7408 36864
rect 7472 36800 7488 36864
rect 7552 36800 7568 36864
rect 7632 36800 7648 36864
rect 7712 36800 7728 36864
rect 7792 36800 7808 36864
rect 7872 36800 7888 36864
rect 7952 36800 7968 36864
rect 8032 36800 8048 36864
rect 8112 36800 8128 36864
rect 8192 36800 8208 36864
rect 8272 36800 8288 36864
rect 8352 36800 8368 36864
rect 8432 36800 8448 36864
rect 8512 36800 8528 36864
rect 8592 36800 8608 36864
rect 8672 36800 8688 36864
rect 8752 36800 8768 36864
rect 8832 36800 8848 36864
rect 8912 36800 8928 36864
rect 8992 36800 14112 36864
rect 14176 36800 14192 36864
rect 14256 36800 14272 36864
rect 14336 36800 14352 36864
rect 14416 36800 24112 36864
rect 24176 36800 24192 36864
rect 24256 36800 24272 36864
rect 24336 36800 24352 36864
rect 24416 36800 36376 36864
rect 36440 36800 36456 36864
rect 36520 36800 36536 36864
rect 36600 36800 36616 36864
rect 36680 36800 36696 36864
rect 36760 36800 36776 36864
rect 36840 36800 36856 36864
rect 36920 36800 36936 36864
rect 37000 36800 37016 36864
rect 37080 36800 37096 36864
rect 37160 36800 37176 36864
rect 37240 36800 37256 36864
rect 37320 36800 37336 36864
rect 37400 36800 37416 36864
rect 37480 36800 37496 36864
rect 37560 36800 37576 36864
rect 37640 36800 37656 36864
rect 37720 36800 37736 36864
rect 37800 36800 37816 36864
rect 37880 36800 37896 36864
rect 37960 36800 37976 36864
rect 38040 36800 38056 36864
rect 38120 36800 38136 36864
rect 38200 36800 38216 36864
rect 38280 36800 38296 36864
rect 38360 36800 38376 36864
rect 38440 36800 38456 36864
rect 38520 36800 38536 36864
rect 38600 36800 38616 36864
rect 38680 36800 38696 36864
rect 38760 36800 38776 36864
rect 38840 36800 38856 36864
rect 38920 36800 38936 36864
rect 39000 36800 39016 36864
rect 39080 36800 39096 36864
rect 39160 36800 39176 36864
rect 39240 36800 39256 36864
rect 39320 36800 39336 36864
rect 39400 36800 39416 36864
rect 39480 36800 39496 36864
rect 39560 36800 39576 36864
rect 39640 36800 39656 36864
rect 39720 36800 39736 36864
rect 39800 36800 39816 36864
rect 39880 36800 39896 36864
rect 39960 36800 39976 36864
rect 40040 36800 40056 36864
rect 40120 36800 40136 36864
rect 40200 36800 40216 36864
rect 40280 36800 40296 36864
rect 40360 36800 40368 36864
rect 5000 36784 40368 36800
rect 5000 36720 5008 36784
rect 5072 36720 5088 36784
rect 5152 36720 5168 36784
rect 5232 36720 5248 36784
rect 5312 36720 5328 36784
rect 5392 36720 5408 36784
rect 5472 36720 5488 36784
rect 5552 36720 5568 36784
rect 5632 36720 5648 36784
rect 5712 36720 5728 36784
rect 5792 36720 5808 36784
rect 5872 36720 5888 36784
rect 5952 36720 5968 36784
rect 6032 36720 6048 36784
rect 6112 36720 6128 36784
rect 6192 36720 6208 36784
rect 6272 36720 6288 36784
rect 6352 36720 6368 36784
rect 6432 36720 6448 36784
rect 6512 36720 6528 36784
rect 6592 36720 6608 36784
rect 6672 36720 6688 36784
rect 6752 36720 6768 36784
rect 6832 36720 6848 36784
rect 6912 36720 6928 36784
rect 6992 36720 7008 36784
rect 7072 36720 7088 36784
rect 7152 36720 7168 36784
rect 7232 36720 7248 36784
rect 7312 36720 7328 36784
rect 7392 36720 7408 36784
rect 7472 36720 7488 36784
rect 7552 36720 7568 36784
rect 7632 36720 7648 36784
rect 7712 36720 7728 36784
rect 7792 36720 7808 36784
rect 7872 36720 7888 36784
rect 7952 36720 7968 36784
rect 8032 36720 8048 36784
rect 8112 36720 8128 36784
rect 8192 36720 8208 36784
rect 8272 36720 8288 36784
rect 8352 36720 8368 36784
rect 8432 36720 8448 36784
rect 8512 36720 8528 36784
rect 8592 36720 8608 36784
rect 8672 36720 8688 36784
rect 8752 36720 8768 36784
rect 8832 36720 8848 36784
rect 8912 36720 8928 36784
rect 8992 36720 14112 36784
rect 14176 36720 14192 36784
rect 14256 36720 14272 36784
rect 14336 36720 14352 36784
rect 14416 36720 24112 36784
rect 24176 36720 24192 36784
rect 24256 36720 24272 36784
rect 24336 36720 24352 36784
rect 24416 36720 36376 36784
rect 36440 36720 36456 36784
rect 36520 36720 36536 36784
rect 36600 36720 36616 36784
rect 36680 36720 36696 36784
rect 36760 36720 36776 36784
rect 36840 36720 36856 36784
rect 36920 36720 36936 36784
rect 37000 36720 37016 36784
rect 37080 36720 37096 36784
rect 37160 36720 37176 36784
rect 37240 36720 37256 36784
rect 37320 36720 37336 36784
rect 37400 36720 37416 36784
rect 37480 36720 37496 36784
rect 37560 36720 37576 36784
rect 37640 36720 37656 36784
rect 37720 36720 37736 36784
rect 37800 36720 37816 36784
rect 37880 36720 37896 36784
rect 37960 36720 37976 36784
rect 38040 36720 38056 36784
rect 38120 36720 38136 36784
rect 38200 36720 38216 36784
rect 38280 36720 38296 36784
rect 38360 36720 38376 36784
rect 38440 36720 38456 36784
rect 38520 36720 38536 36784
rect 38600 36720 38616 36784
rect 38680 36720 38696 36784
rect 38760 36720 38776 36784
rect 38840 36720 38856 36784
rect 38920 36720 38936 36784
rect 39000 36720 39016 36784
rect 39080 36720 39096 36784
rect 39160 36720 39176 36784
rect 39240 36720 39256 36784
rect 39320 36720 39336 36784
rect 39400 36720 39416 36784
rect 39480 36720 39496 36784
rect 39560 36720 39576 36784
rect 39640 36720 39656 36784
rect 39720 36720 39736 36784
rect 39800 36720 39816 36784
rect 39880 36720 39896 36784
rect 39960 36720 39976 36784
rect 40040 36720 40056 36784
rect 40120 36720 40136 36784
rect 40200 36720 40216 36784
rect 40280 36720 40296 36784
rect 40360 36720 40368 36784
rect 5000 36704 40368 36720
rect 5000 36640 5008 36704
rect 5072 36640 5088 36704
rect 5152 36640 5168 36704
rect 5232 36640 5248 36704
rect 5312 36640 5328 36704
rect 5392 36640 5408 36704
rect 5472 36640 5488 36704
rect 5552 36640 5568 36704
rect 5632 36640 5648 36704
rect 5712 36640 5728 36704
rect 5792 36640 5808 36704
rect 5872 36640 5888 36704
rect 5952 36640 5968 36704
rect 6032 36640 6048 36704
rect 6112 36640 6128 36704
rect 6192 36640 6208 36704
rect 6272 36640 6288 36704
rect 6352 36640 6368 36704
rect 6432 36640 6448 36704
rect 6512 36640 6528 36704
rect 6592 36640 6608 36704
rect 6672 36640 6688 36704
rect 6752 36640 6768 36704
rect 6832 36640 6848 36704
rect 6912 36640 6928 36704
rect 6992 36640 7008 36704
rect 7072 36640 7088 36704
rect 7152 36640 7168 36704
rect 7232 36640 7248 36704
rect 7312 36640 7328 36704
rect 7392 36640 7408 36704
rect 7472 36640 7488 36704
rect 7552 36640 7568 36704
rect 7632 36640 7648 36704
rect 7712 36640 7728 36704
rect 7792 36640 7808 36704
rect 7872 36640 7888 36704
rect 7952 36640 7968 36704
rect 8032 36640 8048 36704
rect 8112 36640 8128 36704
rect 8192 36640 8208 36704
rect 8272 36640 8288 36704
rect 8352 36640 8368 36704
rect 8432 36640 8448 36704
rect 8512 36640 8528 36704
rect 8592 36640 8608 36704
rect 8672 36640 8688 36704
rect 8752 36640 8768 36704
rect 8832 36640 8848 36704
rect 8912 36640 8928 36704
rect 8992 36640 14112 36704
rect 14176 36640 14192 36704
rect 14256 36640 14272 36704
rect 14336 36640 14352 36704
rect 14416 36640 24112 36704
rect 24176 36640 24192 36704
rect 24256 36640 24272 36704
rect 24336 36640 24352 36704
rect 24416 36640 36376 36704
rect 36440 36640 36456 36704
rect 36520 36640 36536 36704
rect 36600 36640 36616 36704
rect 36680 36640 36696 36704
rect 36760 36640 36776 36704
rect 36840 36640 36856 36704
rect 36920 36640 36936 36704
rect 37000 36640 37016 36704
rect 37080 36640 37096 36704
rect 37160 36640 37176 36704
rect 37240 36640 37256 36704
rect 37320 36640 37336 36704
rect 37400 36640 37416 36704
rect 37480 36640 37496 36704
rect 37560 36640 37576 36704
rect 37640 36640 37656 36704
rect 37720 36640 37736 36704
rect 37800 36640 37816 36704
rect 37880 36640 37896 36704
rect 37960 36640 37976 36704
rect 38040 36640 38056 36704
rect 38120 36640 38136 36704
rect 38200 36640 38216 36704
rect 38280 36640 38296 36704
rect 38360 36640 38376 36704
rect 38440 36640 38456 36704
rect 38520 36640 38536 36704
rect 38600 36640 38616 36704
rect 38680 36640 38696 36704
rect 38760 36640 38776 36704
rect 38840 36640 38856 36704
rect 38920 36640 38936 36704
rect 39000 36640 39016 36704
rect 39080 36640 39096 36704
rect 39160 36640 39176 36704
rect 39240 36640 39256 36704
rect 39320 36640 39336 36704
rect 39400 36640 39416 36704
rect 39480 36640 39496 36704
rect 39560 36640 39576 36704
rect 39640 36640 39656 36704
rect 39720 36640 39736 36704
rect 39800 36640 39816 36704
rect 39880 36640 39896 36704
rect 39960 36640 39976 36704
rect 40040 36640 40056 36704
rect 40120 36640 40136 36704
rect 40200 36640 40216 36704
rect 40280 36640 40296 36704
rect 40360 36640 40368 36704
rect 5000 36624 40368 36640
rect 5000 36560 5008 36624
rect 5072 36560 5088 36624
rect 5152 36560 5168 36624
rect 5232 36560 5248 36624
rect 5312 36560 5328 36624
rect 5392 36560 5408 36624
rect 5472 36560 5488 36624
rect 5552 36560 5568 36624
rect 5632 36560 5648 36624
rect 5712 36560 5728 36624
rect 5792 36560 5808 36624
rect 5872 36560 5888 36624
rect 5952 36560 5968 36624
rect 6032 36560 6048 36624
rect 6112 36560 6128 36624
rect 6192 36560 6208 36624
rect 6272 36560 6288 36624
rect 6352 36560 6368 36624
rect 6432 36560 6448 36624
rect 6512 36560 6528 36624
rect 6592 36560 6608 36624
rect 6672 36560 6688 36624
rect 6752 36560 6768 36624
rect 6832 36560 6848 36624
rect 6912 36560 6928 36624
rect 6992 36560 7008 36624
rect 7072 36560 7088 36624
rect 7152 36560 7168 36624
rect 7232 36560 7248 36624
rect 7312 36560 7328 36624
rect 7392 36560 7408 36624
rect 7472 36560 7488 36624
rect 7552 36560 7568 36624
rect 7632 36560 7648 36624
rect 7712 36560 7728 36624
rect 7792 36560 7808 36624
rect 7872 36560 7888 36624
rect 7952 36560 7968 36624
rect 8032 36560 8048 36624
rect 8112 36560 8128 36624
rect 8192 36560 8208 36624
rect 8272 36560 8288 36624
rect 8352 36560 8368 36624
rect 8432 36560 8448 36624
rect 8512 36560 8528 36624
rect 8592 36560 8608 36624
rect 8672 36560 8688 36624
rect 8752 36560 8768 36624
rect 8832 36560 8848 36624
rect 8912 36560 8928 36624
rect 8992 36560 14112 36624
rect 14176 36560 14192 36624
rect 14256 36560 14272 36624
rect 14336 36560 14352 36624
rect 14416 36560 24112 36624
rect 24176 36560 24192 36624
rect 24256 36560 24272 36624
rect 24336 36560 24352 36624
rect 24416 36560 36376 36624
rect 36440 36560 36456 36624
rect 36520 36560 36536 36624
rect 36600 36560 36616 36624
rect 36680 36560 36696 36624
rect 36760 36560 36776 36624
rect 36840 36560 36856 36624
rect 36920 36560 36936 36624
rect 37000 36560 37016 36624
rect 37080 36560 37096 36624
rect 37160 36560 37176 36624
rect 37240 36560 37256 36624
rect 37320 36560 37336 36624
rect 37400 36560 37416 36624
rect 37480 36560 37496 36624
rect 37560 36560 37576 36624
rect 37640 36560 37656 36624
rect 37720 36560 37736 36624
rect 37800 36560 37816 36624
rect 37880 36560 37896 36624
rect 37960 36560 37976 36624
rect 38040 36560 38056 36624
rect 38120 36560 38136 36624
rect 38200 36560 38216 36624
rect 38280 36560 38296 36624
rect 38360 36560 38376 36624
rect 38440 36560 38456 36624
rect 38520 36560 38536 36624
rect 38600 36560 38616 36624
rect 38680 36560 38696 36624
rect 38760 36560 38776 36624
rect 38840 36560 38856 36624
rect 38920 36560 38936 36624
rect 39000 36560 39016 36624
rect 39080 36560 39096 36624
rect 39160 36560 39176 36624
rect 39240 36560 39256 36624
rect 39320 36560 39336 36624
rect 39400 36560 39416 36624
rect 39480 36560 39496 36624
rect 39560 36560 39576 36624
rect 39640 36560 39656 36624
rect 39720 36560 39736 36624
rect 39800 36560 39816 36624
rect 39880 36560 39896 36624
rect 39960 36560 39976 36624
rect 40040 36560 40056 36624
rect 40120 36560 40136 36624
rect 40200 36560 40216 36624
rect 40280 36560 40296 36624
rect 40360 36560 40368 36624
rect 5000 36544 40368 36560
rect 5000 36480 5008 36544
rect 5072 36480 5088 36544
rect 5152 36480 5168 36544
rect 5232 36480 5248 36544
rect 5312 36480 5328 36544
rect 5392 36480 5408 36544
rect 5472 36480 5488 36544
rect 5552 36480 5568 36544
rect 5632 36480 5648 36544
rect 5712 36480 5728 36544
rect 5792 36480 5808 36544
rect 5872 36480 5888 36544
rect 5952 36480 5968 36544
rect 6032 36480 6048 36544
rect 6112 36480 6128 36544
rect 6192 36480 6208 36544
rect 6272 36480 6288 36544
rect 6352 36480 6368 36544
rect 6432 36480 6448 36544
rect 6512 36480 6528 36544
rect 6592 36480 6608 36544
rect 6672 36480 6688 36544
rect 6752 36480 6768 36544
rect 6832 36480 6848 36544
rect 6912 36480 6928 36544
rect 6992 36480 7008 36544
rect 7072 36480 7088 36544
rect 7152 36480 7168 36544
rect 7232 36480 7248 36544
rect 7312 36480 7328 36544
rect 7392 36480 7408 36544
rect 7472 36480 7488 36544
rect 7552 36480 7568 36544
rect 7632 36480 7648 36544
rect 7712 36480 7728 36544
rect 7792 36480 7808 36544
rect 7872 36480 7888 36544
rect 7952 36480 7968 36544
rect 8032 36480 8048 36544
rect 8112 36480 8128 36544
rect 8192 36480 8208 36544
rect 8272 36480 8288 36544
rect 8352 36480 8368 36544
rect 8432 36480 8448 36544
rect 8512 36480 8528 36544
rect 8592 36480 8608 36544
rect 8672 36480 8688 36544
rect 8752 36480 8768 36544
rect 8832 36480 8848 36544
rect 8912 36480 8928 36544
rect 8992 36480 14112 36544
rect 14176 36480 14192 36544
rect 14256 36480 14272 36544
rect 14336 36480 14352 36544
rect 14416 36480 24112 36544
rect 24176 36480 24192 36544
rect 24256 36480 24272 36544
rect 24336 36480 24352 36544
rect 24416 36480 36376 36544
rect 36440 36480 36456 36544
rect 36520 36480 36536 36544
rect 36600 36480 36616 36544
rect 36680 36480 36696 36544
rect 36760 36480 36776 36544
rect 36840 36480 36856 36544
rect 36920 36480 36936 36544
rect 37000 36480 37016 36544
rect 37080 36480 37096 36544
rect 37160 36480 37176 36544
rect 37240 36480 37256 36544
rect 37320 36480 37336 36544
rect 37400 36480 37416 36544
rect 37480 36480 37496 36544
rect 37560 36480 37576 36544
rect 37640 36480 37656 36544
rect 37720 36480 37736 36544
rect 37800 36480 37816 36544
rect 37880 36480 37896 36544
rect 37960 36480 37976 36544
rect 38040 36480 38056 36544
rect 38120 36480 38136 36544
rect 38200 36480 38216 36544
rect 38280 36480 38296 36544
rect 38360 36480 38376 36544
rect 38440 36480 38456 36544
rect 38520 36480 38536 36544
rect 38600 36480 38616 36544
rect 38680 36480 38696 36544
rect 38760 36480 38776 36544
rect 38840 36480 38856 36544
rect 38920 36480 38936 36544
rect 39000 36480 39016 36544
rect 39080 36480 39096 36544
rect 39160 36480 39176 36544
rect 39240 36480 39256 36544
rect 39320 36480 39336 36544
rect 39400 36480 39416 36544
rect 39480 36480 39496 36544
rect 39560 36480 39576 36544
rect 39640 36480 39656 36544
rect 39720 36480 39736 36544
rect 39800 36480 39816 36544
rect 39880 36480 39896 36544
rect 39960 36480 39976 36544
rect 40040 36480 40056 36544
rect 40120 36480 40136 36544
rect 40200 36480 40216 36544
rect 40280 36480 40296 36544
rect 40360 36480 40368 36544
rect 5000 36464 40368 36480
rect 5000 36400 5008 36464
rect 5072 36400 5088 36464
rect 5152 36400 5168 36464
rect 5232 36400 5248 36464
rect 5312 36400 5328 36464
rect 5392 36400 5408 36464
rect 5472 36400 5488 36464
rect 5552 36400 5568 36464
rect 5632 36400 5648 36464
rect 5712 36400 5728 36464
rect 5792 36400 5808 36464
rect 5872 36400 5888 36464
rect 5952 36400 5968 36464
rect 6032 36400 6048 36464
rect 6112 36400 6128 36464
rect 6192 36400 6208 36464
rect 6272 36400 6288 36464
rect 6352 36400 6368 36464
rect 6432 36400 6448 36464
rect 6512 36400 6528 36464
rect 6592 36400 6608 36464
rect 6672 36400 6688 36464
rect 6752 36400 6768 36464
rect 6832 36400 6848 36464
rect 6912 36400 6928 36464
rect 6992 36400 7008 36464
rect 7072 36400 7088 36464
rect 7152 36400 7168 36464
rect 7232 36400 7248 36464
rect 7312 36400 7328 36464
rect 7392 36400 7408 36464
rect 7472 36400 7488 36464
rect 7552 36400 7568 36464
rect 7632 36400 7648 36464
rect 7712 36400 7728 36464
rect 7792 36400 7808 36464
rect 7872 36400 7888 36464
rect 7952 36400 7968 36464
rect 8032 36400 8048 36464
rect 8112 36400 8128 36464
rect 8192 36400 8208 36464
rect 8272 36400 8288 36464
rect 8352 36400 8368 36464
rect 8432 36400 8448 36464
rect 8512 36400 8528 36464
rect 8592 36400 8608 36464
rect 8672 36400 8688 36464
rect 8752 36400 8768 36464
rect 8832 36400 8848 36464
rect 8912 36400 8928 36464
rect 8992 36400 14112 36464
rect 14176 36400 14192 36464
rect 14256 36400 14272 36464
rect 14336 36400 14352 36464
rect 14416 36400 24112 36464
rect 24176 36400 24192 36464
rect 24256 36400 24272 36464
rect 24336 36400 24352 36464
rect 24416 36400 36376 36464
rect 36440 36400 36456 36464
rect 36520 36400 36536 36464
rect 36600 36400 36616 36464
rect 36680 36400 36696 36464
rect 36760 36400 36776 36464
rect 36840 36400 36856 36464
rect 36920 36400 36936 36464
rect 37000 36400 37016 36464
rect 37080 36400 37096 36464
rect 37160 36400 37176 36464
rect 37240 36400 37256 36464
rect 37320 36400 37336 36464
rect 37400 36400 37416 36464
rect 37480 36400 37496 36464
rect 37560 36400 37576 36464
rect 37640 36400 37656 36464
rect 37720 36400 37736 36464
rect 37800 36400 37816 36464
rect 37880 36400 37896 36464
rect 37960 36400 37976 36464
rect 38040 36400 38056 36464
rect 38120 36400 38136 36464
rect 38200 36400 38216 36464
rect 38280 36400 38296 36464
rect 38360 36400 38376 36464
rect 38440 36400 38456 36464
rect 38520 36400 38536 36464
rect 38600 36400 38616 36464
rect 38680 36400 38696 36464
rect 38760 36400 38776 36464
rect 38840 36400 38856 36464
rect 38920 36400 38936 36464
rect 39000 36400 39016 36464
rect 39080 36400 39096 36464
rect 39160 36400 39176 36464
rect 39240 36400 39256 36464
rect 39320 36400 39336 36464
rect 39400 36400 39416 36464
rect 39480 36400 39496 36464
rect 39560 36400 39576 36464
rect 39640 36400 39656 36464
rect 39720 36400 39736 36464
rect 39800 36400 39816 36464
rect 39880 36400 39896 36464
rect 39960 36400 39976 36464
rect 40040 36400 40056 36464
rect 40120 36400 40136 36464
rect 40200 36400 40216 36464
rect 40280 36400 40296 36464
rect 40360 36400 40368 36464
rect 5000 36392 40368 36400
rect 19104 34424 19424 34425
rect 19104 34360 19112 34424
rect 19176 34360 19192 34424
rect 19256 34360 19272 34424
rect 19336 34360 19352 34424
rect 19416 34360 19424 34424
rect 19104 34359 19424 34360
rect 29104 34424 29424 34425
rect 29104 34360 29112 34424
rect 29176 34360 29192 34424
rect 29256 34360 29272 34424
rect 29336 34360 29352 34424
rect 29416 34360 29424 34424
rect 29104 34359 29424 34360
rect 31069 33946 31135 33949
rect 34737 33946 35537 33976
rect 31069 33944 35537 33946
rect 31069 33888 31074 33944
rect 31130 33888 35537 33944
rect 31069 33886 35537 33888
rect 31069 33883 31135 33886
rect 14104 33880 14424 33881
rect 14104 33816 14112 33880
rect 14176 33816 14192 33880
rect 14256 33816 14272 33880
rect 14336 33816 14352 33880
rect 14416 33816 14424 33880
rect 14104 33815 14424 33816
rect 24104 33880 24424 33881
rect 24104 33816 24112 33880
rect 24176 33816 24192 33880
rect 24256 33816 24272 33880
rect 24336 33816 24352 33880
rect 24416 33816 24424 33880
rect 34737 33856 35537 33886
rect 24104 33815 24424 33816
rect 19104 33336 19424 33337
rect 19104 33272 19112 33336
rect 19176 33272 19192 33336
rect 19256 33272 19272 33336
rect 19336 33272 19352 33336
rect 19416 33272 19424 33336
rect 19104 33271 19424 33272
rect 29104 33336 29424 33337
rect 29104 33272 29112 33336
rect 29176 33272 29192 33336
rect 29256 33272 29272 33336
rect 29336 33272 29352 33336
rect 29416 33272 29424 33336
rect 29104 33271 29424 33272
rect 9896 33130 10696 33160
rect 13957 33130 14023 33133
rect 9896 33128 14023 33130
rect 9896 33072 13962 33128
rect 14018 33072 14023 33128
rect 9896 33070 14023 33072
rect 9896 33040 10696 33070
rect 13957 33067 14023 33070
rect 14104 32792 14424 32793
rect 14104 32728 14112 32792
rect 14176 32728 14192 32792
rect 14256 32728 14272 32792
rect 14336 32728 14352 32792
rect 14416 32728 14424 32792
rect 14104 32727 14424 32728
rect 24104 32792 24424 32793
rect 24104 32728 24112 32792
rect 24176 32728 24192 32792
rect 24256 32728 24272 32792
rect 24336 32728 24352 32792
rect 24416 32728 24424 32792
rect 24104 32727 24424 32728
rect 19104 32248 19424 32249
rect 19104 32184 19112 32248
rect 19176 32184 19192 32248
rect 19256 32184 19272 32248
rect 19336 32184 19352 32248
rect 19416 32184 19424 32248
rect 19104 32183 19424 32184
rect 29104 32248 29424 32249
rect 29104 32184 29112 32248
rect 29176 32184 29192 32248
rect 29256 32184 29272 32248
rect 29336 32184 29352 32248
rect 29416 32184 29424 32248
rect 29104 32183 29424 32184
rect 14104 31704 14424 31705
rect 14104 31640 14112 31704
rect 14176 31640 14192 31704
rect 14256 31640 14272 31704
rect 14336 31640 14352 31704
rect 14416 31640 14424 31704
rect 14104 31639 14424 31640
rect 24104 31704 24424 31705
rect 24104 31640 24112 31704
rect 24176 31640 24192 31704
rect 24256 31640 24272 31704
rect 24336 31640 24352 31704
rect 24416 31640 24424 31704
rect 24104 31639 24424 31640
rect 19104 31160 19424 31161
rect 19104 31096 19112 31160
rect 19176 31096 19192 31160
rect 19256 31096 19272 31160
rect 19336 31096 19352 31160
rect 19416 31096 19424 31160
rect 19104 31095 19424 31096
rect 29104 31160 29424 31161
rect 29104 31096 29112 31160
rect 29176 31096 29192 31160
rect 29256 31096 29272 31160
rect 29336 31096 29352 31160
rect 29416 31096 29424 31160
rect 29104 31095 29424 31096
rect 31805 30682 31871 30685
rect 34737 30682 35537 30712
rect 31805 30680 35537 30682
rect 31805 30624 31810 30680
rect 31866 30624 35537 30680
rect 31805 30622 35537 30624
rect 31805 30619 31871 30622
rect 14104 30616 14424 30617
rect 14104 30552 14112 30616
rect 14176 30552 14192 30616
rect 14256 30552 14272 30616
rect 14336 30552 14352 30616
rect 14416 30552 14424 30616
rect 14104 30551 14424 30552
rect 24104 30616 24424 30617
rect 24104 30552 24112 30616
rect 24176 30552 24192 30616
rect 24256 30552 24272 30616
rect 24336 30552 24352 30616
rect 24416 30552 24424 30616
rect 34737 30592 35537 30622
rect 24104 30551 24424 30552
rect 19104 30072 19424 30073
rect 19104 30008 19112 30072
rect 19176 30008 19192 30072
rect 19256 30008 19272 30072
rect 19336 30008 19352 30072
rect 19416 30008 19424 30072
rect 19104 30007 19424 30008
rect 29104 30072 29424 30073
rect 29104 30008 29112 30072
rect 29176 30008 29192 30072
rect 29256 30008 29272 30072
rect 29336 30008 29352 30072
rect 29416 30008 29424 30072
rect 29104 30007 29424 30008
rect 9896 29866 10696 29896
rect 13957 29866 14023 29869
rect 9896 29864 14023 29866
rect 9896 29808 13962 29864
rect 14018 29808 14023 29864
rect 9896 29806 14023 29808
rect 9896 29776 10696 29806
rect 13957 29803 14023 29806
rect 14104 29528 14424 29529
rect 14104 29464 14112 29528
rect 14176 29464 14192 29528
rect 14256 29464 14272 29528
rect 14336 29464 14352 29528
rect 14416 29464 14424 29528
rect 14104 29463 14424 29464
rect 24104 29528 24424 29529
rect 24104 29464 24112 29528
rect 24176 29464 24192 29528
rect 24256 29464 24272 29528
rect 24336 29464 24352 29528
rect 24416 29464 24424 29528
rect 24104 29463 24424 29464
rect 19104 28984 19424 28985
rect 19104 28920 19112 28984
rect 19176 28920 19192 28984
rect 19256 28920 19272 28984
rect 19336 28920 19352 28984
rect 19416 28920 19424 28984
rect 19104 28919 19424 28920
rect 29104 28984 29424 28985
rect 29104 28920 29112 28984
rect 29176 28920 29192 28984
rect 29256 28920 29272 28984
rect 29336 28920 29352 28984
rect 29416 28920 29424 28984
rect 29104 28919 29424 28920
rect 14104 28440 14424 28441
rect 14104 28376 14112 28440
rect 14176 28376 14192 28440
rect 14256 28376 14272 28440
rect 14336 28376 14352 28440
rect 14416 28376 14424 28440
rect 14104 28375 14424 28376
rect 24104 28440 24424 28441
rect 24104 28376 24112 28440
rect 24176 28376 24192 28440
rect 24256 28376 24272 28440
rect 24336 28376 24352 28440
rect 24416 28376 24424 28440
rect 24104 28375 24424 28376
rect 19104 27896 19424 27897
rect 19104 27832 19112 27896
rect 19176 27832 19192 27896
rect 19256 27832 19272 27896
rect 19336 27832 19352 27896
rect 19416 27832 19424 27896
rect 19104 27831 19424 27832
rect 29104 27896 29424 27897
rect 29104 27832 29112 27896
rect 29176 27832 29192 27896
rect 29256 27832 29272 27896
rect 29336 27832 29352 27896
rect 29416 27832 29424 27896
rect 29104 27831 29424 27832
rect 31253 27418 31319 27421
rect 34737 27418 35537 27448
rect 31253 27416 35537 27418
rect 31253 27360 31258 27416
rect 31314 27360 35537 27416
rect 31253 27358 35537 27360
rect 31253 27355 31319 27358
rect 14104 27352 14424 27353
rect 14104 27288 14112 27352
rect 14176 27288 14192 27352
rect 14256 27288 14272 27352
rect 14336 27288 14352 27352
rect 14416 27288 14424 27352
rect 14104 27287 14424 27288
rect 24104 27352 24424 27353
rect 24104 27288 24112 27352
rect 24176 27288 24192 27352
rect 24256 27288 24272 27352
rect 24336 27288 24352 27352
rect 24416 27288 24424 27352
rect 34737 27328 35537 27358
rect 24104 27287 24424 27288
rect 19104 26808 19424 26809
rect 19104 26744 19112 26808
rect 19176 26744 19192 26808
rect 19256 26744 19272 26808
rect 19336 26744 19352 26808
rect 19416 26744 19424 26808
rect 19104 26743 19424 26744
rect 29104 26808 29424 26809
rect 29104 26744 29112 26808
rect 29176 26744 29192 26808
rect 29256 26744 29272 26808
rect 29336 26744 29352 26808
rect 29416 26744 29424 26808
rect 29104 26743 29424 26744
rect 9896 26330 10696 26360
rect 11933 26330 11999 26333
rect 9896 26328 11999 26330
rect 9896 26272 11938 26328
rect 11994 26272 11999 26328
rect 9896 26270 11999 26272
rect 9896 26240 10696 26270
rect 11933 26267 11999 26270
rect 14104 26264 14424 26265
rect 14104 26200 14112 26264
rect 14176 26200 14192 26264
rect 14256 26200 14272 26264
rect 14336 26200 14352 26264
rect 14416 26200 14424 26264
rect 14104 26199 14424 26200
rect 24104 26264 24424 26265
rect 24104 26200 24112 26264
rect 24176 26200 24192 26264
rect 24256 26200 24272 26264
rect 24336 26200 24352 26264
rect 24416 26200 24424 26264
rect 24104 26199 24424 26200
rect 19104 25720 19424 25721
rect 19104 25656 19112 25720
rect 19176 25656 19192 25720
rect 19256 25656 19272 25720
rect 19336 25656 19352 25720
rect 19416 25656 19424 25720
rect 19104 25655 19424 25656
rect 29104 25720 29424 25721
rect 29104 25656 29112 25720
rect 29176 25656 29192 25720
rect 29256 25656 29272 25720
rect 29336 25656 29352 25720
rect 29416 25656 29424 25720
rect 29104 25655 29424 25656
rect 14104 25176 14424 25177
rect 14104 25112 14112 25176
rect 14176 25112 14192 25176
rect 14256 25112 14272 25176
rect 14336 25112 14352 25176
rect 14416 25112 14424 25176
rect 14104 25111 14424 25112
rect 24104 25176 24424 25177
rect 24104 25112 24112 25176
rect 24176 25112 24192 25176
rect 24256 25112 24272 25176
rect 24336 25112 24352 25176
rect 24416 25112 24424 25176
rect 24104 25111 24424 25112
rect 22513 24834 22579 24837
rect 26469 24834 26535 24837
rect 27941 24834 28007 24837
rect 22513 24832 28007 24834
rect 22513 24776 22518 24832
rect 22574 24776 26474 24832
rect 26530 24776 27946 24832
rect 28002 24776 28007 24832
rect 22513 24774 28007 24776
rect 22513 24771 22579 24774
rect 26469 24771 26535 24774
rect 27941 24771 28007 24774
rect 19104 24632 19424 24633
rect 19104 24568 19112 24632
rect 19176 24568 19192 24632
rect 19256 24568 19272 24632
rect 19336 24568 19352 24632
rect 19416 24568 19424 24632
rect 19104 24567 19424 24568
rect 29104 24632 29424 24633
rect 29104 24568 29112 24632
rect 29176 24568 29192 24632
rect 29256 24568 29272 24632
rect 29336 24568 29352 24632
rect 29416 24568 29424 24632
rect 29104 24567 29424 24568
rect 14104 24088 14424 24089
rect 14104 24024 14112 24088
rect 14176 24024 14192 24088
rect 14256 24024 14272 24088
rect 14336 24024 14352 24088
rect 14416 24024 14424 24088
rect 14104 24023 14424 24024
rect 24104 24088 24424 24089
rect 24104 24024 24112 24088
rect 24176 24024 24192 24088
rect 24256 24024 24272 24088
rect 24336 24024 24352 24088
rect 24416 24024 24424 24088
rect 24104 24023 24424 24024
rect 30609 23882 30675 23885
rect 34737 23882 35537 23912
rect 30609 23880 35537 23882
rect 30609 23824 30614 23880
rect 30670 23824 35537 23880
rect 30609 23822 35537 23824
rect 30609 23819 30675 23822
rect 34737 23792 35537 23822
rect 19104 23544 19424 23545
rect 19104 23480 19112 23544
rect 19176 23480 19192 23544
rect 19256 23480 19272 23544
rect 19336 23480 19352 23544
rect 19416 23480 19424 23544
rect 19104 23479 19424 23480
rect 29104 23544 29424 23545
rect 29104 23480 29112 23544
rect 29176 23480 29192 23544
rect 29256 23480 29272 23544
rect 29336 23480 29352 23544
rect 29416 23480 29424 23544
rect 29104 23479 29424 23480
rect 18465 23202 18531 23205
rect 19477 23202 19543 23205
rect 18465 23200 19543 23202
rect 18465 23144 18470 23200
rect 18526 23144 19482 23200
rect 19538 23144 19543 23200
rect 18465 23142 19543 23144
rect 18465 23139 18531 23142
rect 19477 23139 19543 23142
rect 9896 23066 10696 23096
rect 13129 23066 13195 23069
rect 9896 23064 13195 23066
rect 9896 23008 13134 23064
rect 13190 23008 13195 23064
rect 9896 23006 13195 23008
rect 9896 22976 10696 23006
rect 13129 23003 13195 23006
rect 14104 23000 14424 23001
rect 14104 22936 14112 23000
rect 14176 22936 14192 23000
rect 14256 22936 14272 23000
rect 14336 22936 14352 23000
rect 14416 22936 14424 23000
rect 14104 22935 14424 22936
rect 24104 23000 24424 23001
rect 24104 22936 24112 23000
rect 24176 22936 24192 23000
rect 24256 22936 24272 23000
rect 24336 22936 24352 23000
rect 24416 22936 24424 23000
rect 24104 22935 24424 22936
rect 19569 22794 19635 22797
rect 25917 22794 25983 22797
rect 19569 22792 25983 22794
rect 19569 22736 19574 22792
rect 19630 22736 25922 22792
rect 25978 22736 25983 22792
rect 19569 22734 25983 22736
rect 19569 22731 19635 22734
rect 25917 22731 25983 22734
rect 19104 22456 19424 22457
rect 19104 22392 19112 22456
rect 19176 22392 19192 22456
rect 19256 22392 19272 22456
rect 19336 22392 19352 22456
rect 19416 22392 19424 22456
rect 19104 22391 19424 22392
rect 29104 22456 29424 22457
rect 29104 22392 29112 22456
rect 29176 22392 29192 22456
rect 29256 22392 29272 22456
rect 29336 22392 29352 22456
rect 29416 22392 29424 22456
rect 29104 22391 29424 22392
rect 14104 21912 14424 21913
rect 14104 21848 14112 21912
rect 14176 21848 14192 21912
rect 14256 21848 14272 21912
rect 14336 21848 14352 21912
rect 14416 21848 14424 21912
rect 14104 21847 14424 21848
rect 24104 21912 24424 21913
rect 24104 21848 24112 21912
rect 24176 21848 24192 21912
rect 24256 21848 24272 21912
rect 24336 21848 24352 21912
rect 24416 21848 24424 21912
rect 24104 21847 24424 21848
rect 19104 21368 19424 21369
rect 19104 21304 19112 21368
rect 19176 21304 19192 21368
rect 19256 21304 19272 21368
rect 19336 21304 19352 21368
rect 19416 21304 19424 21368
rect 19104 21303 19424 21304
rect 29104 21368 29424 21369
rect 29104 21304 29112 21368
rect 29176 21304 29192 21368
rect 29256 21304 29272 21368
rect 29336 21304 29352 21368
rect 29416 21304 29424 21368
rect 29104 21303 29424 21304
rect 14104 20824 14424 20825
rect 14104 20760 14112 20824
rect 14176 20760 14192 20824
rect 14256 20760 14272 20824
rect 14336 20760 14352 20824
rect 14416 20760 14424 20824
rect 14104 20759 14424 20760
rect 24104 20824 24424 20825
rect 24104 20760 24112 20824
rect 24176 20760 24192 20824
rect 24256 20760 24272 20824
rect 24336 20760 24352 20824
rect 24416 20760 24424 20824
rect 24104 20759 24424 20760
rect 32081 20618 32147 20621
rect 34737 20618 35537 20648
rect 32081 20616 35537 20618
rect 32081 20560 32086 20616
rect 32142 20560 35537 20616
rect 32081 20558 35537 20560
rect 32081 20555 32147 20558
rect 34737 20528 35537 20558
rect 19104 20280 19424 20281
rect 19104 20216 19112 20280
rect 19176 20216 19192 20280
rect 19256 20216 19272 20280
rect 19336 20216 19352 20280
rect 19416 20216 19424 20280
rect 19104 20215 19424 20216
rect 29104 20280 29424 20281
rect 29104 20216 29112 20280
rect 29176 20216 29192 20280
rect 29256 20216 29272 20280
rect 29336 20216 29352 20280
rect 29416 20216 29424 20280
rect 29104 20215 29424 20216
rect 9896 19802 10696 19832
rect 12669 19802 12735 19805
rect 9896 19800 12735 19802
rect 9896 19744 12674 19800
rect 12730 19744 12735 19800
rect 9896 19742 12735 19744
rect 9896 19712 10696 19742
rect 12669 19739 12735 19742
rect 14104 19736 14424 19737
rect 14104 19672 14112 19736
rect 14176 19672 14192 19736
rect 14256 19672 14272 19736
rect 14336 19672 14352 19736
rect 14416 19672 14424 19736
rect 14104 19671 14424 19672
rect 24104 19736 24424 19737
rect 24104 19672 24112 19736
rect 24176 19672 24192 19736
rect 24256 19672 24272 19736
rect 24336 19672 24352 19736
rect 24416 19672 24424 19736
rect 24104 19671 24424 19672
rect 19104 19192 19424 19193
rect 19104 19128 19112 19192
rect 19176 19128 19192 19192
rect 19256 19128 19272 19192
rect 19336 19128 19352 19192
rect 19416 19128 19424 19192
rect 19104 19127 19424 19128
rect 29104 19192 29424 19193
rect 29104 19128 29112 19192
rect 29176 19128 29192 19192
rect 29256 19128 29272 19192
rect 29336 19128 29352 19192
rect 29416 19128 29424 19192
rect 29104 19127 29424 19128
rect 14104 18648 14424 18649
rect 14104 18584 14112 18648
rect 14176 18584 14192 18648
rect 14256 18584 14272 18648
rect 14336 18584 14352 18648
rect 14416 18584 14424 18648
rect 14104 18583 14424 18584
rect 24104 18648 24424 18649
rect 24104 18584 24112 18648
rect 24176 18584 24192 18648
rect 24256 18584 24272 18648
rect 24336 18584 24352 18648
rect 24416 18584 24424 18648
rect 24104 18583 24424 18584
rect 19104 18104 19424 18105
rect 19104 18040 19112 18104
rect 19176 18040 19192 18104
rect 19256 18040 19272 18104
rect 19336 18040 19352 18104
rect 19416 18040 19424 18104
rect 19104 18039 19424 18040
rect 29104 18104 29424 18105
rect 29104 18040 29112 18104
rect 29176 18040 29192 18104
rect 29256 18040 29272 18104
rect 29336 18040 29352 18104
rect 29416 18040 29424 18104
rect 29104 18039 29424 18040
rect 14104 17560 14424 17561
rect 14104 17496 14112 17560
rect 14176 17496 14192 17560
rect 14256 17496 14272 17560
rect 14336 17496 14352 17560
rect 14416 17496 14424 17560
rect 14104 17495 14424 17496
rect 24104 17560 24424 17561
rect 24104 17496 24112 17560
rect 24176 17496 24192 17560
rect 24256 17496 24272 17560
rect 24336 17496 24352 17560
rect 24416 17496 24424 17560
rect 24104 17495 24424 17496
rect 30609 17082 30675 17085
rect 34737 17082 35537 17112
rect 30609 17080 35537 17082
rect 30609 17024 30614 17080
rect 30670 17024 35537 17080
rect 30609 17022 35537 17024
rect 30609 17019 30675 17022
rect 19104 17016 19424 17017
rect 19104 16952 19112 17016
rect 19176 16952 19192 17016
rect 19256 16952 19272 17016
rect 19336 16952 19352 17016
rect 19416 16952 19424 17016
rect 19104 16951 19424 16952
rect 29104 17016 29424 17017
rect 29104 16952 29112 17016
rect 29176 16952 29192 17016
rect 29256 16952 29272 17016
rect 29336 16952 29352 17016
rect 29416 16952 29424 17016
rect 34737 16992 35537 17022
rect 29104 16951 29424 16952
rect 14104 16472 14424 16473
rect 14104 16408 14112 16472
rect 14176 16408 14192 16472
rect 14256 16408 14272 16472
rect 14336 16408 14352 16472
rect 14416 16408 14424 16472
rect 14104 16407 14424 16408
rect 24104 16472 24424 16473
rect 24104 16408 24112 16472
rect 24176 16408 24192 16472
rect 24256 16408 24272 16472
rect 24336 16408 24352 16472
rect 24416 16408 24424 16472
rect 24104 16407 24424 16408
rect 9896 16266 10696 16296
rect 13957 16266 14023 16269
rect 9896 16264 14023 16266
rect 9896 16208 13962 16264
rect 14018 16208 14023 16264
rect 9896 16206 14023 16208
rect 9896 16176 10696 16206
rect 13957 16203 14023 16206
rect 19104 15928 19424 15929
rect 19104 15864 19112 15928
rect 19176 15864 19192 15928
rect 19256 15864 19272 15928
rect 19336 15864 19352 15928
rect 19416 15864 19424 15928
rect 19104 15863 19424 15864
rect 29104 15928 29424 15929
rect 29104 15864 29112 15928
rect 29176 15864 29192 15928
rect 29256 15864 29272 15928
rect 29336 15864 29352 15928
rect 29416 15864 29424 15928
rect 29104 15863 29424 15864
rect 14104 15384 14424 15385
rect 14104 15320 14112 15384
rect 14176 15320 14192 15384
rect 14256 15320 14272 15384
rect 14336 15320 14352 15384
rect 14416 15320 14424 15384
rect 14104 15319 14424 15320
rect 24104 15384 24424 15385
rect 24104 15320 24112 15384
rect 24176 15320 24192 15384
rect 24256 15320 24272 15384
rect 24336 15320 24352 15384
rect 24416 15320 24424 15384
rect 24104 15319 24424 15320
rect 19104 14840 19424 14841
rect 19104 14776 19112 14840
rect 19176 14776 19192 14840
rect 19256 14776 19272 14840
rect 19336 14776 19352 14840
rect 19416 14776 19424 14840
rect 19104 14775 19424 14776
rect 29104 14840 29424 14841
rect 29104 14776 29112 14840
rect 29176 14776 29192 14840
rect 29256 14776 29272 14840
rect 29336 14776 29352 14840
rect 29416 14776 29424 14840
rect 29104 14775 29424 14776
rect 14104 14296 14424 14297
rect 14104 14232 14112 14296
rect 14176 14232 14192 14296
rect 14256 14232 14272 14296
rect 14336 14232 14352 14296
rect 14416 14232 14424 14296
rect 14104 14231 14424 14232
rect 24104 14296 24424 14297
rect 24104 14232 24112 14296
rect 24176 14232 24192 14296
rect 24256 14232 24272 14296
rect 24336 14232 24352 14296
rect 24416 14232 24424 14296
rect 24104 14231 24424 14232
rect 30701 13818 30767 13821
rect 34737 13818 35537 13848
rect 30701 13816 35537 13818
rect 30701 13760 30706 13816
rect 30762 13760 35537 13816
rect 30701 13758 35537 13760
rect 30701 13755 30767 13758
rect 19104 13752 19424 13753
rect 19104 13688 19112 13752
rect 19176 13688 19192 13752
rect 19256 13688 19272 13752
rect 19336 13688 19352 13752
rect 19416 13688 19424 13752
rect 19104 13687 19424 13688
rect 29104 13752 29424 13753
rect 29104 13688 29112 13752
rect 29176 13688 29192 13752
rect 29256 13688 29272 13752
rect 29336 13688 29352 13752
rect 29416 13688 29424 13752
rect 34737 13728 35537 13758
rect 29104 13687 29424 13688
rect 14104 13208 14424 13209
rect 14104 13144 14112 13208
rect 14176 13144 14192 13208
rect 14256 13144 14272 13208
rect 14336 13144 14352 13208
rect 14416 13144 14424 13208
rect 14104 13143 14424 13144
rect 24104 13208 24424 13209
rect 24104 13144 24112 13208
rect 24176 13144 24192 13208
rect 24256 13144 24272 13208
rect 24336 13144 24352 13208
rect 24416 13144 24424 13208
rect 24104 13143 24424 13144
rect 9896 13002 10696 13032
rect 12669 13002 12735 13005
rect 9896 13000 12735 13002
rect 9896 12944 12674 13000
rect 12730 12944 12735 13000
rect 9896 12942 12735 12944
rect 9896 12912 10696 12942
rect 12669 12939 12735 12942
rect 19104 12664 19424 12665
rect 19104 12600 19112 12664
rect 19176 12600 19192 12664
rect 19256 12600 19272 12664
rect 19336 12600 19352 12664
rect 19416 12600 19424 12664
rect 19104 12599 19424 12600
rect 29104 12664 29424 12665
rect 29104 12600 29112 12664
rect 29176 12600 29192 12664
rect 29256 12600 29272 12664
rect 29336 12600 29352 12664
rect 29416 12600 29424 12664
rect 29104 12599 29424 12600
rect 14104 12120 14424 12121
rect 14104 12056 14112 12120
rect 14176 12056 14192 12120
rect 14256 12056 14272 12120
rect 14336 12056 14352 12120
rect 14416 12056 14424 12120
rect 14104 12055 14424 12056
rect 24104 12120 24424 12121
rect 24104 12056 24112 12120
rect 24176 12056 24192 12120
rect 24256 12056 24272 12120
rect 24336 12056 24352 12120
rect 24416 12056 24424 12120
rect 24104 12055 24424 12056
rect 19104 11576 19424 11577
rect 19104 11512 19112 11576
rect 19176 11512 19192 11576
rect 19256 11512 19272 11576
rect 19336 11512 19352 11576
rect 19416 11512 19424 11576
rect 19104 11511 19424 11512
rect 29104 11576 29424 11577
rect 29104 11512 29112 11576
rect 29176 11512 29192 11576
rect 29256 11512 29272 11576
rect 29336 11512 29352 11576
rect 29416 11512 29424 11576
rect 29104 11511 29424 11512
rect 14104 11032 14424 11033
rect 14104 10968 14112 11032
rect 14176 10968 14192 11032
rect 14256 10968 14272 11032
rect 14336 10968 14352 11032
rect 14416 10968 14424 11032
rect 14104 10967 14424 10968
rect 24104 11032 24424 11033
rect 24104 10968 24112 11032
rect 24176 10968 24192 11032
rect 24256 10968 24272 11032
rect 24336 10968 24352 11032
rect 24416 10968 24424 11032
rect 24104 10967 24424 10968
rect 30609 10554 30675 10557
rect 34737 10554 35537 10584
rect 30609 10552 35537 10554
rect 30609 10496 30614 10552
rect 30670 10496 35537 10552
rect 30609 10494 35537 10496
rect 30609 10491 30675 10494
rect 34737 10464 35537 10494
rect 5000 8992 40368 9000
rect 5000 8928 5008 8992
rect 5072 8928 5088 8992
rect 5152 8928 5168 8992
rect 5232 8928 5248 8992
rect 5312 8928 5328 8992
rect 5392 8928 5408 8992
rect 5472 8928 5488 8992
rect 5552 8928 5568 8992
rect 5632 8928 5648 8992
rect 5712 8928 5728 8992
rect 5792 8928 5808 8992
rect 5872 8928 5888 8992
rect 5952 8928 5968 8992
rect 6032 8928 6048 8992
rect 6112 8928 6128 8992
rect 6192 8928 6208 8992
rect 6272 8928 6288 8992
rect 6352 8928 6368 8992
rect 6432 8928 6448 8992
rect 6512 8928 6528 8992
rect 6592 8928 6608 8992
rect 6672 8928 6688 8992
rect 6752 8928 6768 8992
rect 6832 8928 6848 8992
rect 6912 8928 6928 8992
rect 6992 8928 7008 8992
rect 7072 8928 7088 8992
rect 7152 8928 7168 8992
rect 7232 8928 7248 8992
rect 7312 8928 7328 8992
rect 7392 8928 7408 8992
rect 7472 8928 7488 8992
rect 7552 8928 7568 8992
rect 7632 8928 7648 8992
rect 7712 8928 7728 8992
rect 7792 8928 7808 8992
rect 7872 8928 7888 8992
rect 7952 8928 7968 8992
rect 8032 8928 8048 8992
rect 8112 8928 8128 8992
rect 8192 8928 8208 8992
rect 8272 8928 8288 8992
rect 8352 8928 8368 8992
rect 8432 8928 8448 8992
rect 8512 8928 8528 8992
rect 8592 8928 8608 8992
rect 8672 8928 8688 8992
rect 8752 8928 8768 8992
rect 8832 8928 8848 8992
rect 8912 8928 8928 8992
rect 8992 8928 14112 8992
rect 14176 8928 14192 8992
rect 14256 8928 14272 8992
rect 14336 8928 14352 8992
rect 14416 8928 24112 8992
rect 24176 8928 24192 8992
rect 24256 8928 24272 8992
rect 24336 8928 24352 8992
rect 24416 8928 36376 8992
rect 36440 8928 36456 8992
rect 36520 8928 36536 8992
rect 36600 8928 36616 8992
rect 36680 8928 36696 8992
rect 36760 8928 36776 8992
rect 36840 8928 36856 8992
rect 36920 8928 36936 8992
rect 37000 8928 37016 8992
rect 37080 8928 37096 8992
rect 37160 8928 37176 8992
rect 37240 8928 37256 8992
rect 37320 8928 37336 8992
rect 37400 8928 37416 8992
rect 37480 8928 37496 8992
rect 37560 8928 37576 8992
rect 37640 8928 37656 8992
rect 37720 8928 37736 8992
rect 37800 8928 37816 8992
rect 37880 8928 37896 8992
rect 37960 8928 37976 8992
rect 38040 8928 38056 8992
rect 38120 8928 38136 8992
rect 38200 8928 38216 8992
rect 38280 8928 38296 8992
rect 38360 8928 38376 8992
rect 38440 8928 38456 8992
rect 38520 8928 38536 8992
rect 38600 8928 38616 8992
rect 38680 8928 38696 8992
rect 38760 8928 38776 8992
rect 38840 8928 38856 8992
rect 38920 8928 38936 8992
rect 39000 8928 39016 8992
rect 39080 8928 39096 8992
rect 39160 8928 39176 8992
rect 39240 8928 39256 8992
rect 39320 8928 39336 8992
rect 39400 8928 39416 8992
rect 39480 8928 39496 8992
rect 39560 8928 39576 8992
rect 39640 8928 39656 8992
rect 39720 8928 39736 8992
rect 39800 8928 39816 8992
rect 39880 8928 39896 8992
rect 39960 8928 39976 8992
rect 40040 8928 40056 8992
rect 40120 8928 40136 8992
rect 40200 8928 40216 8992
rect 40280 8928 40296 8992
rect 40360 8928 40368 8992
rect 5000 8912 40368 8928
rect 5000 8848 5008 8912
rect 5072 8848 5088 8912
rect 5152 8848 5168 8912
rect 5232 8848 5248 8912
rect 5312 8848 5328 8912
rect 5392 8848 5408 8912
rect 5472 8848 5488 8912
rect 5552 8848 5568 8912
rect 5632 8848 5648 8912
rect 5712 8848 5728 8912
rect 5792 8848 5808 8912
rect 5872 8848 5888 8912
rect 5952 8848 5968 8912
rect 6032 8848 6048 8912
rect 6112 8848 6128 8912
rect 6192 8848 6208 8912
rect 6272 8848 6288 8912
rect 6352 8848 6368 8912
rect 6432 8848 6448 8912
rect 6512 8848 6528 8912
rect 6592 8848 6608 8912
rect 6672 8848 6688 8912
rect 6752 8848 6768 8912
rect 6832 8848 6848 8912
rect 6912 8848 6928 8912
rect 6992 8848 7008 8912
rect 7072 8848 7088 8912
rect 7152 8848 7168 8912
rect 7232 8848 7248 8912
rect 7312 8848 7328 8912
rect 7392 8848 7408 8912
rect 7472 8848 7488 8912
rect 7552 8848 7568 8912
rect 7632 8848 7648 8912
rect 7712 8848 7728 8912
rect 7792 8848 7808 8912
rect 7872 8848 7888 8912
rect 7952 8848 7968 8912
rect 8032 8848 8048 8912
rect 8112 8848 8128 8912
rect 8192 8848 8208 8912
rect 8272 8848 8288 8912
rect 8352 8848 8368 8912
rect 8432 8848 8448 8912
rect 8512 8848 8528 8912
rect 8592 8848 8608 8912
rect 8672 8848 8688 8912
rect 8752 8848 8768 8912
rect 8832 8848 8848 8912
rect 8912 8848 8928 8912
rect 8992 8848 14112 8912
rect 14176 8848 14192 8912
rect 14256 8848 14272 8912
rect 14336 8848 14352 8912
rect 14416 8848 24112 8912
rect 24176 8848 24192 8912
rect 24256 8848 24272 8912
rect 24336 8848 24352 8912
rect 24416 8848 36376 8912
rect 36440 8848 36456 8912
rect 36520 8848 36536 8912
rect 36600 8848 36616 8912
rect 36680 8848 36696 8912
rect 36760 8848 36776 8912
rect 36840 8848 36856 8912
rect 36920 8848 36936 8912
rect 37000 8848 37016 8912
rect 37080 8848 37096 8912
rect 37160 8848 37176 8912
rect 37240 8848 37256 8912
rect 37320 8848 37336 8912
rect 37400 8848 37416 8912
rect 37480 8848 37496 8912
rect 37560 8848 37576 8912
rect 37640 8848 37656 8912
rect 37720 8848 37736 8912
rect 37800 8848 37816 8912
rect 37880 8848 37896 8912
rect 37960 8848 37976 8912
rect 38040 8848 38056 8912
rect 38120 8848 38136 8912
rect 38200 8848 38216 8912
rect 38280 8848 38296 8912
rect 38360 8848 38376 8912
rect 38440 8848 38456 8912
rect 38520 8848 38536 8912
rect 38600 8848 38616 8912
rect 38680 8848 38696 8912
rect 38760 8848 38776 8912
rect 38840 8848 38856 8912
rect 38920 8848 38936 8912
rect 39000 8848 39016 8912
rect 39080 8848 39096 8912
rect 39160 8848 39176 8912
rect 39240 8848 39256 8912
rect 39320 8848 39336 8912
rect 39400 8848 39416 8912
rect 39480 8848 39496 8912
rect 39560 8848 39576 8912
rect 39640 8848 39656 8912
rect 39720 8848 39736 8912
rect 39800 8848 39816 8912
rect 39880 8848 39896 8912
rect 39960 8848 39976 8912
rect 40040 8848 40056 8912
rect 40120 8848 40136 8912
rect 40200 8848 40216 8912
rect 40280 8848 40296 8912
rect 40360 8848 40368 8912
rect 5000 8832 40368 8848
rect 5000 8768 5008 8832
rect 5072 8768 5088 8832
rect 5152 8768 5168 8832
rect 5232 8768 5248 8832
rect 5312 8768 5328 8832
rect 5392 8768 5408 8832
rect 5472 8768 5488 8832
rect 5552 8768 5568 8832
rect 5632 8768 5648 8832
rect 5712 8768 5728 8832
rect 5792 8768 5808 8832
rect 5872 8768 5888 8832
rect 5952 8768 5968 8832
rect 6032 8768 6048 8832
rect 6112 8768 6128 8832
rect 6192 8768 6208 8832
rect 6272 8768 6288 8832
rect 6352 8768 6368 8832
rect 6432 8768 6448 8832
rect 6512 8768 6528 8832
rect 6592 8768 6608 8832
rect 6672 8768 6688 8832
rect 6752 8768 6768 8832
rect 6832 8768 6848 8832
rect 6912 8768 6928 8832
rect 6992 8768 7008 8832
rect 7072 8768 7088 8832
rect 7152 8768 7168 8832
rect 7232 8768 7248 8832
rect 7312 8768 7328 8832
rect 7392 8768 7408 8832
rect 7472 8768 7488 8832
rect 7552 8768 7568 8832
rect 7632 8768 7648 8832
rect 7712 8768 7728 8832
rect 7792 8768 7808 8832
rect 7872 8768 7888 8832
rect 7952 8768 7968 8832
rect 8032 8768 8048 8832
rect 8112 8768 8128 8832
rect 8192 8768 8208 8832
rect 8272 8768 8288 8832
rect 8352 8768 8368 8832
rect 8432 8768 8448 8832
rect 8512 8768 8528 8832
rect 8592 8768 8608 8832
rect 8672 8768 8688 8832
rect 8752 8768 8768 8832
rect 8832 8768 8848 8832
rect 8912 8768 8928 8832
rect 8992 8768 14112 8832
rect 14176 8768 14192 8832
rect 14256 8768 14272 8832
rect 14336 8768 14352 8832
rect 14416 8768 24112 8832
rect 24176 8768 24192 8832
rect 24256 8768 24272 8832
rect 24336 8768 24352 8832
rect 24416 8768 36376 8832
rect 36440 8768 36456 8832
rect 36520 8768 36536 8832
rect 36600 8768 36616 8832
rect 36680 8768 36696 8832
rect 36760 8768 36776 8832
rect 36840 8768 36856 8832
rect 36920 8768 36936 8832
rect 37000 8768 37016 8832
rect 37080 8768 37096 8832
rect 37160 8768 37176 8832
rect 37240 8768 37256 8832
rect 37320 8768 37336 8832
rect 37400 8768 37416 8832
rect 37480 8768 37496 8832
rect 37560 8768 37576 8832
rect 37640 8768 37656 8832
rect 37720 8768 37736 8832
rect 37800 8768 37816 8832
rect 37880 8768 37896 8832
rect 37960 8768 37976 8832
rect 38040 8768 38056 8832
rect 38120 8768 38136 8832
rect 38200 8768 38216 8832
rect 38280 8768 38296 8832
rect 38360 8768 38376 8832
rect 38440 8768 38456 8832
rect 38520 8768 38536 8832
rect 38600 8768 38616 8832
rect 38680 8768 38696 8832
rect 38760 8768 38776 8832
rect 38840 8768 38856 8832
rect 38920 8768 38936 8832
rect 39000 8768 39016 8832
rect 39080 8768 39096 8832
rect 39160 8768 39176 8832
rect 39240 8768 39256 8832
rect 39320 8768 39336 8832
rect 39400 8768 39416 8832
rect 39480 8768 39496 8832
rect 39560 8768 39576 8832
rect 39640 8768 39656 8832
rect 39720 8768 39736 8832
rect 39800 8768 39816 8832
rect 39880 8768 39896 8832
rect 39960 8768 39976 8832
rect 40040 8768 40056 8832
rect 40120 8768 40136 8832
rect 40200 8768 40216 8832
rect 40280 8768 40296 8832
rect 40360 8768 40368 8832
rect 5000 8752 40368 8768
rect 5000 8688 5008 8752
rect 5072 8688 5088 8752
rect 5152 8688 5168 8752
rect 5232 8688 5248 8752
rect 5312 8688 5328 8752
rect 5392 8688 5408 8752
rect 5472 8688 5488 8752
rect 5552 8688 5568 8752
rect 5632 8688 5648 8752
rect 5712 8688 5728 8752
rect 5792 8688 5808 8752
rect 5872 8688 5888 8752
rect 5952 8688 5968 8752
rect 6032 8688 6048 8752
rect 6112 8688 6128 8752
rect 6192 8688 6208 8752
rect 6272 8688 6288 8752
rect 6352 8688 6368 8752
rect 6432 8688 6448 8752
rect 6512 8688 6528 8752
rect 6592 8688 6608 8752
rect 6672 8688 6688 8752
rect 6752 8688 6768 8752
rect 6832 8688 6848 8752
rect 6912 8688 6928 8752
rect 6992 8688 7008 8752
rect 7072 8688 7088 8752
rect 7152 8688 7168 8752
rect 7232 8688 7248 8752
rect 7312 8688 7328 8752
rect 7392 8688 7408 8752
rect 7472 8688 7488 8752
rect 7552 8688 7568 8752
rect 7632 8688 7648 8752
rect 7712 8688 7728 8752
rect 7792 8688 7808 8752
rect 7872 8688 7888 8752
rect 7952 8688 7968 8752
rect 8032 8688 8048 8752
rect 8112 8688 8128 8752
rect 8192 8688 8208 8752
rect 8272 8688 8288 8752
rect 8352 8688 8368 8752
rect 8432 8688 8448 8752
rect 8512 8688 8528 8752
rect 8592 8688 8608 8752
rect 8672 8688 8688 8752
rect 8752 8688 8768 8752
rect 8832 8688 8848 8752
rect 8912 8688 8928 8752
rect 8992 8688 14112 8752
rect 14176 8688 14192 8752
rect 14256 8688 14272 8752
rect 14336 8688 14352 8752
rect 14416 8688 24112 8752
rect 24176 8688 24192 8752
rect 24256 8688 24272 8752
rect 24336 8688 24352 8752
rect 24416 8688 36376 8752
rect 36440 8688 36456 8752
rect 36520 8688 36536 8752
rect 36600 8688 36616 8752
rect 36680 8688 36696 8752
rect 36760 8688 36776 8752
rect 36840 8688 36856 8752
rect 36920 8688 36936 8752
rect 37000 8688 37016 8752
rect 37080 8688 37096 8752
rect 37160 8688 37176 8752
rect 37240 8688 37256 8752
rect 37320 8688 37336 8752
rect 37400 8688 37416 8752
rect 37480 8688 37496 8752
rect 37560 8688 37576 8752
rect 37640 8688 37656 8752
rect 37720 8688 37736 8752
rect 37800 8688 37816 8752
rect 37880 8688 37896 8752
rect 37960 8688 37976 8752
rect 38040 8688 38056 8752
rect 38120 8688 38136 8752
rect 38200 8688 38216 8752
rect 38280 8688 38296 8752
rect 38360 8688 38376 8752
rect 38440 8688 38456 8752
rect 38520 8688 38536 8752
rect 38600 8688 38616 8752
rect 38680 8688 38696 8752
rect 38760 8688 38776 8752
rect 38840 8688 38856 8752
rect 38920 8688 38936 8752
rect 39000 8688 39016 8752
rect 39080 8688 39096 8752
rect 39160 8688 39176 8752
rect 39240 8688 39256 8752
rect 39320 8688 39336 8752
rect 39400 8688 39416 8752
rect 39480 8688 39496 8752
rect 39560 8688 39576 8752
rect 39640 8688 39656 8752
rect 39720 8688 39736 8752
rect 39800 8688 39816 8752
rect 39880 8688 39896 8752
rect 39960 8688 39976 8752
rect 40040 8688 40056 8752
rect 40120 8688 40136 8752
rect 40200 8688 40216 8752
rect 40280 8688 40296 8752
rect 40360 8688 40368 8752
rect 5000 8672 40368 8688
rect 5000 8608 5008 8672
rect 5072 8608 5088 8672
rect 5152 8608 5168 8672
rect 5232 8608 5248 8672
rect 5312 8608 5328 8672
rect 5392 8608 5408 8672
rect 5472 8608 5488 8672
rect 5552 8608 5568 8672
rect 5632 8608 5648 8672
rect 5712 8608 5728 8672
rect 5792 8608 5808 8672
rect 5872 8608 5888 8672
rect 5952 8608 5968 8672
rect 6032 8608 6048 8672
rect 6112 8608 6128 8672
rect 6192 8608 6208 8672
rect 6272 8608 6288 8672
rect 6352 8608 6368 8672
rect 6432 8608 6448 8672
rect 6512 8608 6528 8672
rect 6592 8608 6608 8672
rect 6672 8608 6688 8672
rect 6752 8608 6768 8672
rect 6832 8608 6848 8672
rect 6912 8608 6928 8672
rect 6992 8608 7008 8672
rect 7072 8608 7088 8672
rect 7152 8608 7168 8672
rect 7232 8608 7248 8672
rect 7312 8608 7328 8672
rect 7392 8608 7408 8672
rect 7472 8608 7488 8672
rect 7552 8608 7568 8672
rect 7632 8608 7648 8672
rect 7712 8608 7728 8672
rect 7792 8608 7808 8672
rect 7872 8608 7888 8672
rect 7952 8608 7968 8672
rect 8032 8608 8048 8672
rect 8112 8608 8128 8672
rect 8192 8608 8208 8672
rect 8272 8608 8288 8672
rect 8352 8608 8368 8672
rect 8432 8608 8448 8672
rect 8512 8608 8528 8672
rect 8592 8608 8608 8672
rect 8672 8608 8688 8672
rect 8752 8608 8768 8672
rect 8832 8608 8848 8672
rect 8912 8608 8928 8672
rect 8992 8608 14112 8672
rect 14176 8608 14192 8672
rect 14256 8608 14272 8672
rect 14336 8608 14352 8672
rect 14416 8608 24112 8672
rect 24176 8608 24192 8672
rect 24256 8608 24272 8672
rect 24336 8608 24352 8672
rect 24416 8608 36376 8672
rect 36440 8608 36456 8672
rect 36520 8608 36536 8672
rect 36600 8608 36616 8672
rect 36680 8608 36696 8672
rect 36760 8608 36776 8672
rect 36840 8608 36856 8672
rect 36920 8608 36936 8672
rect 37000 8608 37016 8672
rect 37080 8608 37096 8672
rect 37160 8608 37176 8672
rect 37240 8608 37256 8672
rect 37320 8608 37336 8672
rect 37400 8608 37416 8672
rect 37480 8608 37496 8672
rect 37560 8608 37576 8672
rect 37640 8608 37656 8672
rect 37720 8608 37736 8672
rect 37800 8608 37816 8672
rect 37880 8608 37896 8672
rect 37960 8608 37976 8672
rect 38040 8608 38056 8672
rect 38120 8608 38136 8672
rect 38200 8608 38216 8672
rect 38280 8608 38296 8672
rect 38360 8608 38376 8672
rect 38440 8608 38456 8672
rect 38520 8608 38536 8672
rect 38600 8608 38616 8672
rect 38680 8608 38696 8672
rect 38760 8608 38776 8672
rect 38840 8608 38856 8672
rect 38920 8608 38936 8672
rect 39000 8608 39016 8672
rect 39080 8608 39096 8672
rect 39160 8608 39176 8672
rect 39240 8608 39256 8672
rect 39320 8608 39336 8672
rect 39400 8608 39416 8672
rect 39480 8608 39496 8672
rect 39560 8608 39576 8672
rect 39640 8608 39656 8672
rect 39720 8608 39736 8672
rect 39800 8608 39816 8672
rect 39880 8608 39896 8672
rect 39960 8608 39976 8672
rect 40040 8608 40056 8672
rect 40120 8608 40136 8672
rect 40200 8608 40216 8672
rect 40280 8608 40296 8672
rect 40360 8608 40368 8672
rect 5000 8592 40368 8608
rect 5000 8528 5008 8592
rect 5072 8528 5088 8592
rect 5152 8528 5168 8592
rect 5232 8528 5248 8592
rect 5312 8528 5328 8592
rect 5392 8528 5408 8592
rect 5472 8528 5488 8592
rect 5552 8528 5568 8592
rect 5632 8528 5648 8592
rect 5712 8528 5728 8592
rect 5792 8528 5808 8592
rect 5872 8528 5888 8592
rect 5952 8528 5968 8592
rect 6032 8528 6048 8592
rect 6112 8528 6128 8592
rect 6192 8528 6208 8592
rect 6272 8528 6288 8592
rect 6352 8528 6368 8592
rect 6432 8528 6448 8592
rect 6512 8528 6528 8592
rect 6592 8528 6608 8592
rect 6672 8528 6688 8592
rect 6752 8528 6768 8592
rect 6832 8528 6848 8592
rect 6912 8528 6928 8592
rect 6992 8528 7008 8592
rect 7072 8528 7088 8592
rect 7152 8528 7168 8592
rect 7232 8528 7248 8592
rect 7312 8528 7328 8592
rect 7392 8528 7408 8592
rect 7472 8528 7488 8592
rect 7552 8528 7568 8592
rect 7632 8528 7648 8592
rect 7712 8528 7728 8592
rect 7792 8528 7808 8592
rect 7872 8528 7888 8592
rect 7952 8528 7968 8592
rect 8032 8528 8048 8592
rect 8112 8528 8128 8592
rect 8192 8528 8208 8592
rect 8272 8528 8288 8592
rect 8352 8528 8368 8592
rect 8432 8528 8448 8592
rect 8512 8528 8528 8592
rect 8592 8528 8608 8592
rect 8672 8528 8688 8592
rect 8752 8528 8768 8592
rect 8832 8528 8848 8592
rect 8912 8528 8928 8592
rect 8992 8528 14112 8592
rect 14176 8528 14192 8592
rect 14256 8528 14272 8592
rect 14336 8528 14352 8592
rect 14416 8528 24112 8592
rect 24176 8528 24192 8592
rect 24256 8528 24272 8592
rect 24336 8528 24352 8592
rect 24416 8528 36376 8592
rect 36440 8528 36456 8592
rect 36520 8528 36536 8592
rect 36600 8528 36616 8592
rect 36680 8528 36696 8592
rect 36760 8528 36776 8592
rect 36840 8528 36856 8592
rect 36920 8528 36936 8592
rect 37000 8528 37016 8592
rect 37080 8528 37096 8592
rect 37160 8528 37176 8592
rect 37240 8528 37256 8592
rect 37320 8528 37336 8592
rect 37400 8528 37416 8592
rect 37480 8528 37496 8592
rect 37560 8528 37576 8592
rect 37640 8528 37656 8592
rect 37720 8528 37736 8592
rect 37800 8528 37816 8592
rect 37880 8528 37896 8592
rect 37960 8528 37976 8592
rect 38040 8528 38056 8592
rect 38120 8528 38136 8592
rect 38200 8528 38216 8592
rect 38280 8528 38296 8592
rect 38360 8528 38376 8592
rect 38440 8528 38456 8592
rect 38520 8528 38536 8592
rect 38600 8528 38616 8592
rect 38680 8528 38696 8592
rect 38760 8528 38776 8592
rect 38840 8528 38856 8592
rect 38920 8528 38936 8592
rect 39000 8528 39016 8592
rect 39080 8528 39096 8592
rect 39160 8528 39176 8592
rect 39240 8528 39256 8592
rect 39320 8528 39336 8592
rect 39400 8528 39416 8592
rect 39480 8528 39496 8592
rect 39560 8528 39576 8592
rect 39640 8528 39656 8592
rect 39720 8528 39736 8592
rect 39800 8528 39816 8592
rect 39880 8528 39896 8592
rect 39960 8528 39976 8592
rect 40040 8528 40056 8592
rect 40120 8528 40136 8592
rect 40200 8528 40216 8592
rect 40280 8528 40296 8592
rect 40360 8528 40368 8592
rect 5000 8512 40368 8528
rect 5000 8448 5008 8512
rect 5072 8448 5088 8512
rect 5152 8448 5168 8512
rect 5232 8448 5248 8512
rect 5312 8448 5328 8512
rect 5392 8448 5408 8512
rect 5472 8448 5488 8512
rect 5552 8448 5568 8512
rect 5632 8448 5648 8512
rect 5712 8448 5728 8512
rect 5792 8448 5808 8512
rect 5872 8448 5888 8512
rect 5952 8448 5968 8512
rect 6032 8448 6048 8512
rect 6112 8448 6128 8512
rect 6192 8448 6208 8512
rect 6272 8448 6288 8512
rect 6352 8448 6368 8512
rect 6432 8448 6448 8512
rect 6512 8448 6528 8512
rect 6592 8448 6608 8512
rect 6672 8448 6688 8512
rect 6752 8448 6768 8512
rect 6832 8448 6848 8512
rect 6912 8448 6928 8512
rect 6992 8448 7008 8512
rect 7072 8448 7088 8512
rect 7152 8448 7168 8512
rect 7232 8448 7248 8512
rect 7312 8448 7328 8512
rect 7392 8448 7408 8512
rect 7472 8448 7488 8512
rect 7552 8448 7568 8512
rect 7632 8448 7648 8512
rect 7712 8448 7728 8512
rect 7792 8448 7808 8512
rect 7872 8448 7888 8512
rect 7952 8448 7968 8512
rect 8032 8448 8048 8512
rect 8112 8448 8128 8512
rect 8192 8448 8208 8512
rect 8272 8448 8288 8512
rect 8352 8448 8368 8512
rect 8432 8448 8448 8512
rect 8512 8448 8528 8512
rect 8592 8448 8608 8512
rect 8672 8448 8688 8512
rect 8752 8448 8768 8512
rect 8832 8448 8848 8512
rect 8912 8448 8928 8512
rect 8992 8448 14112 8512
rect 14176 8448 14192 8512
rect 14256 8448 14272 8512
rect 14336 8448 14352 8512
rect 14416 8448 24112 8512
rect 24176 8448 24192 8512
rect 24256 8448 24272 8512
rect 24336 8448 24352 8512
rect 24416 8448 36376 8512
rect 36440 8448 36456 8512
rect 36520 8448 36536 8512
rect 36600 8448 36616 8512
rect 36680 8448 36696 8512
rect 36760 8448 36776 8512
rect 36840 8448 36856 8512
rect 36920 8448 36936 8512
rect 37000 8448 37016 8512
rect 37080 8448 37096 8512
rect 37160 8448 37176 8512
rect 37240 8448 37256 8512
rect 37320 8448 37336 8512
rect 37400 8448 37416 8512
rect 37480 8448 37496 8512
rect 37560 8448 37576 8512
rect 37640 8448 37656 8512
rect 37720 8448 37736 8512
rect 37800 8448 37816 8512
rect 37880 8448 37896 8512
rect 37960 8448 37976 8512
rect 38040 8448 38056 8512
rect 38120 8448 38136 8512
rect 38200 8448 38216 8512
rect 38280 8448 38296 8512
rect 38360 8448 38376 8512
rect 38440 8448 38456 8512
rect 38520 8448 38536 8512
rect 38600 8448 38616 8512
rect 38680 8448 38696 8512
rect 38760 8448 38776 8512
rect 38840 8448 38856 8512
rect 38920 8448 38936 8512
rect 39000 8448 39016 8512
rect 39080 8448 39096 8512
rect 39160 8448 39176 8512
rect 39240 8448 39256 8512
rect 39320 8448 39336 8512
rect 39400 8448 39416 8512
rect 39480 8448 39496 8512
rect 39560 8448 39576 8512
rect 39640 8448 39656 8512
rect 39720 8448 39736 8512
rect 39800 8448 39816 8512
rect 39880 8448 39896 8512
rect 39960 8448 39976 8512
rect 40040 8448 40056 8512
rect 40120 8448 40136 8512
rect 40200 8448 40216 8512
rect 40280 8448 40296 8512
rect 40360 8448 40368 8512
rect 5000 8432 40368 8448
rect 5000 8368 5008 8432
rect 5072 8368 5088 8432
rect 5152 8368 5168 8432
rect 5232 8368 5248 8432
rect 5312 8368 5328 8432
rect 5392 8368 5408 8432
rect 5472 8368 5488 8432
rect 5552 8368 5568 8432
rect 5632 8368 5648 8432
rect 5712 8368 5728 8432
rect 5792 8368 5808 8432
rect 5872 8368 5888 8432
rect 5952 8368 5968 8432
rect 6032 8368 6048 8432
rect 6112 8368 6128 8432
rect 6192 8368 6208 8432
rect 6272 8368 6288 8432
rect 6352 8368 6368 8432
rect 6432 8368 6448 8432
rect 6512 8368 6528 8432
rect 6592 8368 6608 8432
rect 6672 8368 6688 8432
rect 6752 8368 6768 8432
rect 6832 8368 6848 8432
rect 6912 8368 6928 8432
rect 6992 8368 7008 8432
rect 7072 8368 7088 8432
rect 7152 8368 7168 8432
rect 7232 8368 7248 8432
rect 7312 8368 7328 8432
rect 7392 8368 7408 8432
rect 7472 8368 7488 8432
rect 7552 8368 7568 8432
rect 7632 8368 7648 8432
rect 7712 8368 7728 8432
rect 7792 8368 7808 8432
rect 7872 8368 7888 8432
rect 7952 8368 7968 8432
rect 8032 8368 8048 8432
rect 8112 8368 8128 8432
rect 8192 8368 8208 8432
rect 8272 8368 8288 8432
rect 8352 8368 8368 8432
rect 8432 8368 8448 8432
rect 8512 8368 8528 8432
rect 8592 8368 8608 8432
rect 8672 8368 8688 8432
rect 8752 8368 8768 8432
rect 8832 8368 8848 8432
rect 8912 8368 8928 8432
rect 8992 8368 14112 8432
rect 14176 8368 14192 8432
rect 14256 8368 14272 8432
rect 14336 8368 14352 8432
rect 14416 8368 24112 8432
rect 24176 8368 24192 8432
rect 24256 8368 24272 8432
rect 24336 8368 24352 8432
rect 24416 8368 36376 8432
rect 36440 8368 36456 8432
rect 36520 8368 36536 8432
rect 36600 8368 36616 8432
rect 36680 8368 36696 8432
rect 36760 8368 36776 8432
rect 36840 8368 36856 8432
rect 36920 8368 36936 8432
rect 37000 8368 37016 8432
rect 37080 8368 37096 8432
rect 37160 8368 37176 8432
rect 37240 8368 37256 8432
rect 37320 8368 37336 8432
rect 37400 8368 37416 8432
rect 37480 8368 37496 8432
rect 37560 8368 37576 8432
rect 37640 8368 37656 8432
rect 37720 8368 37736 8432
rect 37800 8368 37816 8432
rect 37880 8368 37896 8432
rect 37960 8368 37976 8432
rect 38040 8368 38056 8432
rect 38120 8368 38136 8432
rect 38200 8368 38216 8432
rect 38280 8368 38296 8432
rect 38360 8368 38376 8432
rect 38440 8368 38456 8432
rect 38520 8368 38536 8432
rect 38600 8368 38616 8432
rect 38680 8368 38696 8432
rect 38760 8368 38776 8432
rect 38840 8368 38856 8432
rect 38920 8368 38936 8432
rect 39000 8368 39016 8432
rect 39080 8368 39096 8432
rect 39160 8368 39176 8432
rect 39240 8368 39256 8432
rect 39320 8368 39336 8432
rect 39400 8368 39416 8432
rect 39480 8368 39496 8432
rect 39560 8368 39576 8432
rect 39640 8368 39656 8432
rect 39720 8368 39736 8432
rect 39800 8368 39816 8432
rect 39880 8368 39896 8432
rect 39960 8368 39976 8432
rect 40040 8368 40056 8432
rect 40120 8368 40136 8432
rect 40200 8368 40216 8432
rect 40280 8368 40296 8432
rect 40360 8368 40368 8432
rect 5000 8352 40368 8368
rect 5000 8288 5008 8352
rect 5072 8288 5088 8352
rect 5152 8288 5168 8352
rect 5232 8288 5248 8352
rect 5312 8288 5328 8352
rect 5392 8288 5408 8352
rect 5472 8288 5488 8352
rect 5552 8288 5568 8352
rect 5632 8288 5648 8352
rect 5712 8288 5728 8352
rect 5792 8288 5808 8352
rect 5872 8288 5888 8352
rect 5952 8288 5968 8352
rect 6032 8288 6048 8352
rect 6112 8288 6128 8352
rect 6192 8288 6208 8352
rect 6272 8288 6288 8352
rect 6352 8288 6368 8352
rect 6432 8288 6448 8352
rect 6512 8288 6528 8352
rect 6592 8288 6608 8352
rect 6672 8288 6688 8352
rect 6752 8288 6768 8352
rect 6832 8288 6848 8352
rect 6912 8288 6928 8352
rect 6992 8288 7008 8352
rect 7072 8288 7088 8352
rect 7152 8288 7168 8352
rect 7232 8288 7248 8352
rect 7312 8288 7328 8352
rect 7392 8288 7408 8352
rect 7472 8288 7488 8352
rect 7552 8288 7568 8352
rect 7632 8288 7648 8352
rect 7712 8288 7728 8352
rect 7792 8288 7808 8352
rect 7872 8288 7888 8352
rect 7952 8288 7968 8352
rect 8032 8288 8048 8352
rect 8112 8288 8128 8352
rect 8192 8288 8208 8352
rect 8272 8288 8288 8352
rect 8352 8288 8368 8352
rect 8432 8288 8448 8352
rect 8512 8288 8528 8352
rect 8592 8288 8608 8352
rect 8672 8288 8688 8352
rect 8752 8288 8768 8352
rect 8832 8288 8848 8352
rect 8912 8288 8928 8352
rect 8992 8288 14112 8352
rect 14176 8288 14192 8352
rect 14256 8288 14272 8352
rect 14336 8288 14352 8352
rect 14416 8288 24112 8352
rect 24176 8288 24192 8352
rect 24256 8288 24272 8352
rect 24336 8288 24352 8352
rect 24416 8288 36376 8352
rect 36440 8288 36456 8352
rect 36520 8288 36536 8352
rect 36600 8288 36616 8352
rect 36680 8288 36696 8352
rect 36760 8288 36776 8352
rect 36840 8288 36856 8352
rect 36920 8288 36936 8352
rect 37000 8288 37016 8352
rect 37080 8288 37096 8352
rect 37160 8288 37176 8352
rect 37240 8288 37256 8352
rect 37320 8288 37336 8352
rect 37400 8288 37416 8352
rect 37480 8288 37496 8352
rect 37560 8288 37576 8352
rect 37640 8288 37656 8352
rect 37720 8288 37736 8352
rect 37800 8288 37816 8352
rect 37880 8288 37896 8352
rect 37960 8288 37976 8352
rect 38040 8288 38056 8352
rect 38120 8288 38136 8352
rect 38200 8288 38216 8352
rect 38280 8288 38296 8352
rect 38360 8288 38376 8352
rect 38440 8288 38456 8352
rect 38520 8288 38536 8352
rect 38600 8288 38616 8352
rect 38680 8288 38696 8352
rect 38760 8288 38776 8352
rect 38840 8288 38856 8352
rect 38920 8288 38936 8352
rect 39000 8288 39016 8352
rect 39080 8288 39096 8352
rect 39160 8288 39176 8352
rect 39240 8288 39256 8352
rect 39320 8288 39336 8352
rect 39400 8288 39416 8352
rect 39480 8288 39496 8352
rect 39560 8288 39576 8352
rect 39640 8288 39656 8352
rect 39720 8288 39736 8352
rect 39800 8288 39816 8352
rect 39880 8288 39896 8352
rect 39960 8288 39976 8352
rect 40040 8288 40056 8352
rect 40120 8288 40136 8352
rect 40200 8288 40216 8352
rect 40280 8288 40296 8352
rect 40360 8288 40368 8352
rect 5000 8272 40368 8288
rect 5000 8208 5008 8272
rect 5072 8208 5088 8272
rect 5152 8208 5168 8272
rect 5232 8208 5248 8272
rect 5312 8208 5328 8272
rect 5392 8208 5408 8272
rect 5472 8208 5488 8272
rect 5552 8208 5568 8272
rect 5632 8208 5648 8272
rect 5712 8208 5728 8272
rect 5792 8208 5808 8272
rect 5872 8208 5888 8272
rect 5952 8208 5968 8272
rect 6032 8208 6048 8272
rect 6112 8208 6128 8272
rect 6192 8208 6208 8272
rect 6272 8208 6288 8272
rect 6352 8208 6368 8272
rect 6432 8208 6448 8272
rect 6512 8208 6528 8272
rect 6592 8208 6608 8272
rect 6672 8208 6688 8272
rect 6752 8208 6768 8272
rect 6832 8208 6848 8272
rect 6912 8208 6928 8272
rect 6992 8208 7008 8272
rect 7072 8208 7088 8272
rect 7152 8208 7168 8272
rect 7232 8208 7248 8272
rect 7312 8208 7328 8272
rect 7392 8208 7408 8272
rect 7472 8208 7488 8272
rect 7552 8208 7568 8272
rect 7632 8208 7648 8272
rect 7712 8208 7728 8272
rect 7792 8208 7808 8272
rect 7872 8208 7888 8272
rect 7952 8208 7968 8272
rect 8032 8208 8048 8272
rect 8112 8208 8128 8272
rect 8192 8208 8208 8272
rect 8272 8208 8288 8272
rect 8352 8208 8368 8272
rect 8432 8208 8448 8272
rect 8512 8208 8528 8272
rect 8592 8208 8608 8272
rect 8672 8208 8688 8272
rect 8752 8208 8768 8272
rect 8832 8208 8848 8272
rect 8912 8208 8928 8272
rect 8992 8208 14112 8272
rect 14176 8208 14192 8272
rect 14256 8208 14272 8272
rect 14336 8208 14352 8272
rect 14416 8208 24112 8272
rect 24176 8208 24192 8272
rect 24256 8208 24272 8272
rect 24336 8208 24352 8272
rect 24416 8208 36376 8272
rect 36440 8208 36456 8272
rect 36520 8208 36536 8272
rect 36600 8208 36616 8272
rect 36680 8208 36696 8272
rect 36760 8208 36776 8272
rect 36840 8208 36856 8272
rect 36920 8208 36936 8272
rect 37000 8208 37016 8272
rect 37080 8208 37096 8272
rect 37160 8208 37176 8272
rect 37240 8208 37256 8272
rect 37320 8208 37336 8272
rect 37400 8208 37416 8272
rect 37480 8208 37496 8272
rect 37560 8208 37576 8272
rect 37640 8208 37656 8272
rect 37720 8208 37736 8272
rect 37800 8208 37816 8272
rect 37880 8208 37896 8272
rect 37960 8208 37976 8272
rect 38040 8208 38056 8272
rect 38120 8208 38136 8272
rect 38200 8208 38216 8272
rect 38280 8208 38296 8272
rect 38360 8208 38376 8272
rect 38440 8208 38456 8272
rect 38520 8208 38536 8272
rect 38600 8208 38616 8272
rect 38680 8208 38696 8272
rect 38760 8208 38776 8272
rect 38840 8208 38856 8272
rect 38920 8208 38936 8272
rect 39000 8208 39016 8272
rect 39080 8208 39096 8272
rect 39160 8208 39176 8272
rect 39240 8208 39256 8272
rect 39320 8208 39336 8272
rect 39400 8208 39416 8272
rect 39480 8208 39496 8272
rect 39560 8208 39576 8272
rect 39640 8208 39656 8272
rect 39720 8208 39736 8272
rect 39800 8208 39816 8272
rect 39880 8208 39896 8272
rect 39960 8208 39976 8272
rect 40040 8208 40056 8272
rect 40120 8208 40136 8272
rect 40200 8208 40216 8272
rect 40280 8208 40296 8272
rect 40360 8208 40368 8272
rect 5000 8192 40368 8208
rect 5000 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5168 8192
rect 5232 8128 5248 8192
rect 5312 8128 5328 8192
rect 5392 8128 5408 8192
rect 5472 8128 5488 8192
rect 5552 8128 5568 8192
rect 5632 8128 5648 8192
rect 5712 8128 5728 8192
rect 5792 8128 5808 8192
rect 5872 8128 5888 8192
rect 5952 8128 5968 8192
rect 6032 8128 6048 8192
rect 6112 8128 6128 8192
rect 6192 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6528 8192
rect 6592 8128 6608 8192
rect 6672 8128 6688 8192
rect 6752 8128 6768 8192
rect 6832 8128 6848 8192
rect 6912 8128 6928 8192
rect 6992 8128 7008 8192
rect 7072 8128 7088 8192
rect 7152 8128 7168 8192
rect 7232 8128 7248 8192
rect 7312 8128 7328 8192
rect 7392 8128 7408 8192
rect 7472 8128 7488 8192
rect 7552 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7888 8192
rect 7952 8128 7968 8192
rect 8032 8128 8048 8192
rect 8112 8128 8128 8192
rect 8192 8128 8208 8192
rect 8272 8128 8288 8192
rect 8352 8128 8368 8192
rect 8432 8128 8448 8192
rect 8512 8128 8528 8192
rect 8592 8128 8608 8192
rect 8672 8128 8688 8192
rect 8752 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14272 8192
rect 14336 8128 14352 8192
rect 14416 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 36376 8192
rect 36440 8128 36456 8192
rect 36520 8128 36536 8192
rect 36600 8128 36616 8192
rect 36680 8128 36696 8192
rect 36760 8128 36776 8192
rect 36840 8128 36856 8192
rect 36920 8128 36936 8192
rect 37000 8128 37016 8192
rect 37080 8128 37096 8192
rect 37160 8128 37176 8192
rect 37240 8128 37256 8192
rect 37320 8128 37336 8192
rect 37400 8128 37416 8192
rect 37480 8128 37496 8192
rect 37560 8128 37576 8192
rect 37640 8128 37656 8192
rect 37720 8128 37736 8192
rect 37800 8128 37816 8192
rect 37880 8128 37896 8192
rect 37960 8128 37976 8192
rect 38040 8128 38056 8192
rect 38120 8128 38136 8192
rect 38200 8128 38216 8192
rect 38280 8128 38296 8192
rect 38360 8128 38376 8192
rect 38440 8128 38456 8192
rect 38520 8128 38536 8192
rect 38600 8128 38616 8192
rect 38680 8128 38696 8192
rect 38760 8128 38776 8192
rect 38840 8128 38856 8192
rect 38920 8128 38936 8192
rect 39000 8128 39016 8192
rect 39080 8128 39096 8192
rect 39160 8128 39176 8192
rect 39240 8128 39256 8192
rect 39320 8128 39336 8192
rect 39400 8128 39416 8192
rect 39480 8128 39496 8192
rect 39560 8128 39576 8192
rect 39640 8128 39656 8192
rect 39720 8128 39736 8192
rect 39800 8128 39816 8192
rect 39880 8128 39896 8192
rect 39960 8128 39976 8192
rect 40040 8128 40056 8192
rect 40120 8128 40136 8192
rect 40200 8128 40216 8192
rect 40280 8128 40296 8192
rect 40360 8128 40368 8192
rect 5000 8112 40368 8128
rect 5000 8048 5008 8112
rect 5072 8048 5088 8112
rect 5152 8048 5168 8112
rect 5232 8048 5248 8112
rect 5312 8048 5328 8112
rect 5392 8048 5408 8112
rect 5472 8048 5488 8112
rect 5552 8048 5568 8112
rect 5632 8048 5648 8112
rect 5712 8048 5728 8112
rect 5792 8048 5808 8112
rect 5872 8048 5888 8112
rect 5952 8048 5968 8112
rect 6032 8048 6048 8112
rect 6112 8048 6128 8112
rect 6192 8048 6208 8112
rect 6272 8048 6288 8112
rect 6352 8048 6368 8112
rect 6432 8048 6448 8112
rect 6512 8048 6528 8112
rect 6592 8048 6608 8112
rect 6672 8048 6688 8112
rect 6752 8048 6768 8112
rect 6832 8048 6848 8112
rect 6912 8048 6928 8112
rect 6992 8048 7008 8112
rect 7072 8048 7088 8112
rect 7152 8048 7168 8112
rect 7232 8048 7248 8112
rect 7312 8048 7328 8112
rect 7392 8048 7408 8112
rect 7472 8048 7488 8112
rect 7552 8048 7568 8112
rect 7632 8048 7648 8112
rect 7712 8048 7728 8112
rect 7792 8048 7808 8112
rect 7872 8048 7888 8112
rect 7952 8048 7968 8112
rect 8032 8048 8048 8112
rect 8112 8048 8128 8112
rect 8192 8048 8208 8112
rect 8272 8048 8288 8112
rect 8352 8048 8368 8112
rect 8432 8048 8448 8112
rect 8512 8048 8528 8112
rect 8592 8048 8608 8112
rect 8672 8048 8688 8112
rect 8752 8048 8768 8112
rect 8832 8048 8848 8112
rect 8912 8048 8928 8112
rect 8992 8048 14112 8112
rect 14176 8048 14192 8112
rect 14256 8048 14272 8112
rect 14336 8048 14352 8112
rect 14416 8048 24112 8112
rect 24176 8048 24192 8112
rect 24256 8048 24272 8112
rect 24336 8048 24352 8112
rect 24416 8048 36376 8112
rect 36440 8048 36456 8112
rect 36520 8048 36536 8112
rect 36600 8048 36616 8112
rect 36680 8048 36696 8112
rect 36760 8048 36776 8112
rect 36840 8048 36856 8112
rect 36920 8048 36936 8112
rect 37000 8048 37016 8112
rect 37080 8048 37096 8112
rect 37160 8048 37176 8112
rect 37240 8048 37256 8112
rect 37320 8048 37336 8112
rect 37400 8048 37416 8112
rect 37480 8048 37496 8112
rect 37560 8048 37576 8112
rect 37640 8048 37656 8112
rect 37720 8048 37736 8112
rect 37800 8048 37816 8112
rect 37880 8048 37896 8112
rect 37960 8048 37976 8112
rect 38040 8048 38056 8112
rect 38120 8048 38136 8112
rect 38200 8048 38216 8112
rect 38280 8048 38296 8112
rect 38360 8048 38376 8112
rect 38440 8048 38456 8112
rect 38520 8048 38536 8112
rect 38600 8048 38616 8112
rect 38680 8048 38696 8112
rect 38760 8048 38776 8112
rect 38840 8048 38856 8112
rect 38920 8048 38936 8112
rect 39000 8048 39016 8112
rect 39080 8048 39096 8112
rect 39160 8048 39176 8112
rect 39240 8048 39256 8112
rect 39320 8048 39336 8112
rect 39400 8048 39416 8112
rect 39480 8048 39496 8112
rect 39560 8048 39576 8112
rect 39640 8048 39656 8112
rect 39720 8048 39736 8112
rect 39800 8048 39816 8112
rect 39880 8048 39896 8112
rect 39960 8048 39976 8112
rect 40040 8048 40056 8112
rect 40120 8048 40136 8112
rect 40200 8048 40216 8112
rect 40280 8048 40296 8112
rect 40360 8048 40368 8112
rect 5000 8032 40368 8048
rect 5000 7968 5008 8032
rect 5072 7968 5088 8032
rect 5152 7968 5168 8032
rect 5232 7968 5248 8032
rect 5312 7968 5328 8032
rect 5392 7968 5408 8032
rect 5472 7968 5488 8032
rect 5552 7968 5568 8032
rect 5632 7968 5648 8032
rect 5712 7968 5728 8032
rect 5792 7968 5808 8032
rect 5872 7968 5888 8032
rect 5952 7968 5968 8032
rect 6032 7968 6048 8032
rect 6112 7968 6128 8032
rect 6192 7968 6208 8032
rect 6272 7968 6288 8032
rect 6352 7968 6368 8032
rect 6432 7968 6448 8032
rect 6512 7968 6528 8032
rect 6592 7968 6608 8032
rect 6672 7968 6688 8032
rect 6752 7968 6768 8032
rect 6832 7968 6848 8032
rect 6912 7968 6928 8032
rect 6992 7968 7008 8032
rect 7072 7968 7088 8032
rect 7152 7968 7168 8032
rect 7232 7968 7248 8032
rect 7312 7968 7328 8032
rect 7392 7968 7408 8032
rect 7472 7968 7488 8032
rect 7552 7968 7568 8032
rect 7632 7968 7648 8032
rect 7712 7968 7728 8032
rect 7792 7968 7808 8032
rect 7872 7968 7888 8032
rect 7952 7968 7968 8032
rect 8032 7968 8048 8032
rect 8112 7968 8128 8032
rect 8192 7968 8208 8032
rect 8272 7968 8288 8032
rect 8352 7968 8368 8032
rect 8432 7968 8448 8032
rect 8512 7968 8528 8032
rect 8592 7968 8608 8032
rect 8672 7968 8688 8032
rect 8752 7968 8768 8032
rect 8832 7968 8848 8032
rect 8912 7968 8928 8032
rect 8992 7968 14112 8032
rect 14176 7968 14192 8032
rect 14256 7968 14272 8032
rect 14336 7968 14352 8032
rect 14416 7968 24112 8032
rect 24176 7968 24192 8032
rect 24256 7968 24272 8032
rect 24336 7968 24352 8032
rect 24416 7968 36376 8032
rect 36440 7968 36456 8032
rect 36520 7968 36536 8032
rect 36600 7968 36616 8032
rect 36680 7968 36696 8032
rect 36760 7968 36776 8032
rect 36840 7968 36856 8032
rect 36920 7968 36936 8032
rect 37000 7968 37016 8032
rect 37080 7968 37096 8032
rect 37160 7968 37176 8032
rect 37240 7968 37256 8032
rect 37320 7968 37336 8032
rect 37400 7968 37416 8032
rect 37480 7968 37496 8032
rect 37560 7968 37576 8032
rect 37640 7968 37656 8032
rect 37720 7968 37736 8032
rect 37800 7968 37816 8032
rect 37880 7968 37896 8032
rect 37960 7968 37976 8032
rect 38040 7968 38056 8032
rect 38120 7968 38136 8032
rect 38200 7968 38216 8032
rect 38280 7968 38296 8032
rect 38360 7968 38376 8032
rect 38440 7968 38456 8032
rect 38520 7968 38536 8032
rect 38600 7968 38616 8032
rect 38680 7968 38696 8032
rect 38760 7968 38776 8032
rect 38840 7968 38856 8032
rect 38920 7968 38936 8032
rect 39000 7968 39016 8032
rect 39080 7968 39096 8032
rect 39160 7968 39176 8032
rect 39240 7968 39256 8032
rect 39320 7968 39336 8032
rect 39400 7968 39416 8032
rect 39480 7968 39496 8032
rect 39560 7968 39576 8032
rect 39640 7968 39656 8032
rect 39720 7968 39736 8032
rect 39800 7968 39816 8032
rect 39880 7968 39896 8032
rect 39960 7968 39976 8032
rect 40040 7968 40056 8032
rect 40120 7968 40136 8032
rect 40200 7968 40216 8032
rect 40280 7968 40296 8032
rect 40360 7968 40368 8032
rect 5000 7952 40368 7968
rect 5000 7888 5008 7952
rect 5072 7888 5088 7952
rect 5152 7888 5168 7952
rect 5232 7888 5248 7952
rect 5312 7888 5328 7952
rect 5392 7888 5408 7952
rect 5472 7888 5488 7952
rect 5552 7888 5568 7952
rect 5632 7888 5648 7952
rect 5712 7888 5728 7952
rect 5792 7888 5808 7952
rect 5872 7888 5888 7952
rect 5952 7888 5968 7952
rect 6032 7888 6048 7952
rect 6112 7888 6128 7952
rect 6192 7888 6208 7952
rect 6272 7888 6288 7952
rect 6352 7888 6368 7952
rect 6432 7888 6448 7952
rect 6512 7888 6528 7952
rect 6592 7888 6608 7952
rect 6672 7888 6688 7952
rect 6752 7888 6768 7952
rect 6832 7888 6848 7952
rect 6912 7888 6928 7952
rect 6992 7888 7008 7952
rect 7072 7888 7088 7952
rect 7152 7888 7168 7952
rect 7232 7888 7248 7952
rect 7312 7888 7328 7952
rect 7392 7888 7408 7952
rect 7472 7888 7488 7952
rect 7552 7888 7568 7952
rect 7632 7888 7648 7952
rect 7712 7888 7728 7952
rect 7792 7888 7808 7952
rect 7872 7888 7888 7952
rect 7952 7888 7968 7952
rect 8032 7888 8048 7952
rect 8112 7888 8128 7952
rect 8192 7888 8208 7952
rect 8272 7888 8288 7952
rect 8352 7888 8368 7952
rect 8432 7888 8448 7952
rect 8512 7888 8528 7952
rect 8592 7888 8608 7952
rect 8672 7888 8688 7952
rect 8752 7888 8768 7952
rect 8832 7888 8848 7952
rect 8912 7888 8928 7952
rect 8992 7888 14112 7952
rect 14176 7888 14192 7952
rect 14256 7888 14272 7952
rect 14336 7888 14352 7952
rect 14416 7888 24112 7952
rect 24176 7888 24192 7952
rect 24256 7888 24272 7952
rect 24336 7888 24352 7952
rect 24416 7888 36376 7952
rect 36440 7888 36456 7952
rect 36520 7888 36536 7952
rect 36600 7888 36616 7952
rect 36680 7888 36696 7952
rect 36760 7888 36776 7952
rect 36840 7888 36856 7952
rect 36920 7888 36936 7952
rect 37000 7888 37016 7952
rect 37080 7888 37096 7952
rect 37160 7888 37176 7952
rect 37240 7888 37256 7952
rect 37320 7888 37336 7952
rect 37400 7888 37416 7952
rect 37480 7888 37496 7952
rect 37560 7888 37576 7952
rect 37640 7888 37656 7952
rect 37720 7888 37736 7952
rect 37800 7888 37816 7952
rect 37880 7888 37896 7952
rect 37960 7888 37976 7952
rect 38040 7888 38056 7952
rect 38120 7888 38136 7952
rect 38200 7888 38216 7952
rect 38280 7888 38296 7952
rect 38360 7888 38376 7952
rect 38440 7888 38456 7952
rect 38520 7888 38536 7952
rect 38600 7888 38616 7952
rect 38680 7888 38696 7952
rect 38760 7888 38776 7952
rect 38840 7888 38856 7952
rect 38920 7888 38936 7952
rect 39000 7888 39016 7952
rect 39080 7888 39096 7952
rect 39160 7888 39176 7952
rect 39240 7888 39256 7952
rect 39320 7888 39336 7952
rect 39400 7888 39416 7952
rect 39480 7888 39496 7952
rect 39560 7888 39576 7952
rect 39640 7888 39656 7952
rect 39720 7888 39736 7952
rect 39800 7888 39816 7952
rect 39880 7888 39896 7952
rect 39960 7888 39976 7952
rect 40040 7888 40056 7952
rect 40120 7888 40136 7952
rect 40200 7888 40216 7952
rect 40280 7888 40296 7952
rect 40360 7888 40368 7952
rect 5000 7872 40368 7888
rect 5000 7808 5008 7872
rect 5072 7808 5088 7872
rect 5152 7808 5168 7872
rect 5232 7808 5248 7872
rect 5312 7808 5328 7872
rect 5392 7808 5408 7872
rect 5472 7808 5488 7872
rect 5552 7808 5568 7872
rect 5632 7808 5648 7872
rect 5712 7808 5728 7872
rect 5792 7808 5808 7872
rect 5872 7808 5888 7872
rect 5952 7808 5968 7872
rect 6032 7808 6048 7872
rect 6112 7808 6128 7872
rect 6192 7808 6208 7872
rect 6272 7808 6288 7872
rect 6352 7808 6368 7872
rect 6432 7808 6448 7872
rect 6512 7808 6528 7872
rect 6592 7808 6608 7872
rect 6672 7808 6688 7872
rect 6752 7808 6768 7872
rect 6832 7808 6848 7872
rect 6912 7808 6928 7872
rect 6992 7808 7008 7872
rect 7072 7808 7088 7872
rect 7152 7808 7168 7872
rect 7232 7808 7248 7872
rect 7312 7808 7328 7872
rect 7392 7808 7408 7872
rect 7472 7808 7488 7872
rect 7552 7808 7568 7872
rect 7632 7808 7648 7872
rect 7712 7808 7728 7872
rect 7792 7808 7808 7872
rect 7872 7808 7888 7872
rect 7952 7808 7968 7872
rect 8032 7808 8048 7872
rect 8112 7808 8128 7872
rect 8192 7808 8208 7872
rect 8272 7808 8288 7872
rect 8352 7808 8368 7872
rect 8432 7808 8448 7872
rect 8512 7808 8528 7872
rect 8592 7808 8608 7872
rect 8672 7808 8688 7872
rect 8752 7808 8768 7872
rect 8832 7808 8848 7872
rect 8912 7808 8928 7872
rect 8992 7808 14112 7872
rect 14176 7808 14192 7872
rect 14256 7808 14272 7872
rect 14336 7808 14352 7872
rect 14416 7808 24112 7872
rect 24176 7808 24192 7872
rect 24256 7808 24272 7872
rect 24336 7808 24352 7872
rect 24416 7808 36376 7872
rect 36440 7808 36456 7872
rect 36520 7808 36536 7872
rect 36600 7808 36616 7872
rect 36680 7808 36696 7872
rect 36760 7808 36776 7872
rect 36840 7808 36856 7872
rect 36920 7808 36936 7872
rect 37000 7808 37016 7872
rect 37080 7808 37096 7872
rect 37160 7808 37176 7872
rect 37240 7808 37256 7872
rect 37320 7808 37336 7872
rect 37400 7808 37416 7872
rect 37480 7808 37496 7872
rect 37560 7808 37576 7872
rect 37640 7808 37656 7872
rect 37720 7808 37736 7872
rect 37800 7808 37816 7872
rect 37880 7808 37896 7872
rect 37960 7808 37976 7872
rect 38040 7808 38056 7872
rect 38120 7808 38136 7872
rect 38200 7808 38216 7872
rect 38280 7808 38296 7872
rect 38360 7808 38376 7872
rect 38440 7808 38456 7872
rect 38520 7808 38536 7872
rect 38600 7808 38616 7872
rect 38680 7808 38696 7872
rect 38760 7808 38776 7872
rect 38840 7808 38856 7872
rect 38920 7808 38936 7872
rect 39000 7808 39016 7872
rect 39080 7808 39096 7872
rect 39160 7808 39176 7872
rect 39240 7808 39256 7872
rect 39320 7808 39336 7872
rect 39400 7808 39416 7872
rect 39480 7808 39496 7872
rect 39560 7808 39576 7872
rect 39640 7808 39656 7872
rect 39720 7808 39736 7872
rect 39800 7808 39816 7872
rect 39880 7808 39896 7872
rect 39960 7808 39976 7872
rect 40040 7808 40056 7872
rect 40120 7808 40136 7872
rect 40200 7808 40216 7872
rect 40280 7808 40296 7872
rect 40360 7808 40368 7872
rect 5000 7792 40368 7808
rect 5000 7728 5008 7792
rect 5072 7728 5088 7792
rect 5152 7728 5168 7792
rect 5232 7728 5248 7792
rect 5312 7728 5328 7792
rect 5392 7728 5408 7792
rect 5472 7728 5488 7792
rect 5552 7728 5568 7792
rect 5632 7728 5648 7792
rect 5712 7728 5728 7792
rect 5792 7728 5808 7792
rect 5872 7728 5888 7792
rect 5952 7728 5968 7792
rect 6032 7728 6048 7792
rect 6112 7728 6128 7792
rect 6192 7728 6208 7792
rect 6272 7728 6288 7792
rect 6352 7728 6368 7792
rect 6432 7728 6448 7792
rect 6512 7728 6528 7792
rect 6592 7728 6608 7792
rect 6672 7728 6688 7792
rect 6752 7728 6768 7792
rect 6832 7728 6848 7792
rect 6912 7728 6928 7792
rect 6992 7728 7008 7792
rect 7072 7728 7088 7792
rect 7152 7728 7168 7792
rect 7232 7728 7248 7792
rect 7312 7728 7328 7792
rect 7392 7728 7408 7792
rect 7472 7728 7488 7792
rect 7552 7728 7568 7792
rect 7632 7728 7648 7792
rect 7712 7728 7728 7792
rect 7792 7728 7808 7792
rect 7872 7728 7888 7792
rect 7952 7728 7968 7792
rect 8032 7728 8048 7792
rect 8112 7728 8128 7792
rect 8192 7728 8208 7792
rect 8272 7728 8288 7792
rect 8352 7728 8368 7792
rect 8432 7728 8448 7792
rect 8512 7728 8528 7792
rect 8592 7728 8608 7792
rect 8672 7728 8688 7792
rect 8752 7728 8768 7792
rect 8832 7728 8848 7792
rect 8912 7728 8928 7792
rect 8992 7728 14112 7792
rect 14176 7728 14192 7792
rect 14256 7728 14272 7792
rect 14336 7728 14352 7792
rect 14416 7728 24112 7792
rect 24176 7728 24192 7792
rect 24256 7728 24272 7792
rect 24336 7728 24352 7792
rect 24416 7728 36376 7792
rect 36440 7728 36456 7792
rect 36520 7728 36536 7792
rect 36600 7728 36616 7792
rect 36680 7728 36696 7792
rect 36760 7728 36776 7792
rect 36840 7728 36856 7792
rect 36920 7728 36936 7792
rect 37000 7728 37016 7792
rect 37080 7728 37096 7792
rect 37160 7728 37176 7792
rect 37240 7728 37256 7792
rect 37320 7728 37336 7792
rect 37400 7728 37416 7792
rect 37480 7728 37496 7792
rect 37560 7728 37576 7792
rect 37640 7728 37656 7792
rect 37720 7728 37736 7792
rect 37800 7728 37816 7792
rect 37880 7728 37896 7792
rect 37960 7728 37976 7792
rect 38040 7728 38056 7792
rect 38120 7728 38136 7792
rect 38200 7728 38216 7792
rect 38280 7728 38296 7792
rect 38360 7728 38376 7792
rect 38440 7728 38456 7792
rect 38520 7728 38536 7792
rect 38600 7728 38616 7792
rect 38680 7728 38696 7792
rect 38760 7728 38776 7792
rect 38840 7728 38856 7792
rect 38920 7728 38936 7792
rect 39000 7728 39016 7792
rect 39080 7728 39096 7792
rect 39160 7728 39176 7792
rect 39240 7728 39256 7792
rect 39320 7728 39336 7792
rect 39400 7728 39416 7792
rect 39480 7728 39496 7792
rect 39560 7728 39576 7792
rect 39640 7728 39656 7792
rect 39720 7728 39736 7792
rect 39800 7728 39816 7792
rect 39880 7728 39896 7792
rect 39960 7728 39976 7792
rect 40040 7728 40056 7792
rect 40120 7728 40136 7792
rect 40200 7728 40216 7792
rect 40280 7728 40296 7792
rect 40360 7728 40368 7792
rect 5000 7712 40368 7728
rect 5000 7648 5008 7712
rect 5072 7648 5088 7712
rect 5152 7648 5168 7712
rect 5232 7648 5248 7712
rect 5312 7648 5328 7712
rect 5392 7648 5408 7712
rect 5472 7648 5488 7712
rect 5552 7648 5568 7712
rect 5632 7648 5648 7712
rect 5712 7648 5728 7712
rect 5792 7648 5808 7712
rect 5872 7648 5888 7712
rect 5952 7648 5968 7712
rect 6032 7648 6048 7712
rect 6112 7648 6128 7712
rect 6192 7648 6208 7712
rect 6272 7648 6288 7712
rect 6352 7648 6368 7712
rect 6432 7648 6448 7712
rect 6512 7648 6528 7712
rect 6592 7648 6608 7712
rect 6672 7648 6688 7712
rect 6752 7648 6768 7712
rect 6832 7648 6848 7712
rect 6912 7648 6928 7712
rect 6992 7648 7008 7712
rect 7072 7648 7088 7712
rect 7152 7648 7168 7712
rect 7232 7648 7248 7712
rect 7312 7648 7328 7712
rect 7392 7648 7408 7712
rect 7472 7648 7488 7712
rect 7552 7648 7568 7712
rect 7632 7648 7648 7712
rect 7712 7648 7728 7712
rect 7792 7648 7808 7712
rect 7872 7648 7888 7712
rect 7952 7648 7968 7712
rect 8032 7648 8048 7712
rect 8112 7648 8128 7712
rect 8192 7648 8208 7712
rect 8272 7648 8288 7712
rect 8352 7648 8368 7712
rect 8432 7648 8448 7712
rect 8512 7648 8528 7712
rect 8592 7648 8608 7712
rect 8672 7648 8688 7712
rect 8752 7648 8768 7712
rect 8832 7648 8848 7712
rect 8912 7648 8928 7712
rect 8992 7648 14112 7712
rect 14176 7648 14192 7712
rect 14256 7648 14272 7712
rect 14336 7648 14352 7712
rect 14416 7648 24112 7712
rect 24176 7648 24192 7712
rect 24256 7648 24272 7712
rect 24336 7648 24352 7712
rect 24416 7648 36376 7712
rect 36440 7648 36456 7712
rect 36520 7648 36536 7712
rect 36600 7648 36616 7712
rect 36680 7648 36696 7712
rect 36760 7648 36776 7712
rect 36840 7648 36856 7712
rect 36920 7648 36936 7712
rect 37000 7648 37016 7712
rect 37080 7648 37096 7712
rect 37160 7648 37176 7712
rect 37240 7648 37256 7712
rect 37320 7648 37336 7712
rect 37400 7648 37416 7712
rect 37480 7648 37496 7712
rect 37560 7648 37576 7712
rect 37640 7648 37656 7712
rect 37720 7648 37736 7712
rect 37800 7648 37816 7712
rect 37880 7648 37896 7712
rect 37960 7648 37976 7712
rect 38040 7648 38056 7712
rect 38120 7648 38136 7712
rect 38200 7648 38216 7712
rect 38280 7648 38296 7712
rect 38360 7648 38376 7712
rect 38440 7648 38456 7712
rect 38520 7648 38536 7712
rect 38600 7648 38616 7712
rect 38680 7648 38696 7712
rect 38760 7648 38776 7712
rect 38840 7648 38856 7712
rect 38920 7648 38936 7712
rect 39000 7648 39016 7712
rect 39080 7648 39096 7712
rect 39160 7648 39176 7712
rect 39240 7648 39256 7712
rect 39320 7648 39336 7712
rect 39400 7648 39416 7712
rect 39480 7648 39496 7712
rect 39560 7648 39576 7712
rect 39640 7648 39656 7712
rect 39720 7648 39736 7712
rect 39800 7648 39816 7712
rect 39880 7648 39896 7712
rect 39960 7648 39976 7712
rect 40040 7648 40056 7712
rect 40120 7648 40136 7712
rect 40200 7648 40216 7712
rect 40280 7648 40296 7712
rect 40360 7648 40368 7712
rect 5000 7632 40368 7648
rect 5000 7568 5008 7632
rect 5072 7568 5088 7632
rect 5152 7568 5168 7632
rect 5232 7568 5248 7632
rect 5312 7568 5328 7632
rect 5392 7568 5408 7632
rect 5472 7568 5488 7632
rect 5552 7568 5568 7632
rect 5632 7568 5648 7632
rect 5712 7568 5728 7632
rect 5792 7568 5808 7632
rect 5872 7568 5888 7632
rect 5952 7568 5968 7632
rect 6032 7568 6048 7632
rect 6112 7568 6128 7632
rect 6192 7568 6208 7632
rect 6272 7568 6288 7632
rect 6352 7568 6368 7632
rect 6432 7568 6448 7632
rect 6512 7568 6528 7632
rect 6592 7568 6608 7632
rect 6672 7568 6688 7632
rect 6752 7568 6768 7632
rect 6832 7568 6848 7632
rect 6912 7568 6928 7632
rect 6992 7568 7008 7632
rect 7072 7568 7088 7632
rect 7152 7568 7168 7632
rect 7232 7568 7248 7632
rect 7312 7568 7328 7632
rect 7392 7568 7408 7632
rect 7472 7568 7488 7632
rect 7552 7568 7568 7632
rect 7632 7568 7648 7632
rect 7712 7568 7728 7632
rect 7792 7568 7808 7632
rect 7872 7568 7888 7632
rect 7952 7568 7968 7632
rect 8032 7568 8048 7632
rect 8112 7568 8128 7632
rect 8192 7568 8208 7632
rect 8272 7568 8288 7632
rect 8352 7568 8368 7632
rect 8432 7568 8448 7632
rect 8512 7568 8528 7632
rect 8592 7568 8608 7632
rect 8672 7568 8688 7632
rect 8752 7568 8768 7632
rect 8832 7568 8848 7632
rect 8912 7568 8928 7632
rect 8992 7568 14112 7632
rect 14176 7568 14192 7632
rect 14256 7568 14272 7632
rect 14336 7568 14352 7632
rect 14416 7568 24112 7632
rect 24176 7568 24192 7632
rect 24256 7568 24272 7632
rect 24336 7568 24352 7632
rect 24416 7568 36376 7632
rect 36440 7568 36456 7632
rect 36520 7568 36536 7632
rect 36600 7568 36616 7632
rect 36680 7568 36696 7632
rect 36760 7568 36776 7632
rect 36840 7568 36856 7632
rect 36920 7568 36936 7632
rect 37000 7568 37016 7632
rect 37080 7568 37096 7632
rect 37160 7568 37176 7632
rect 37240 7568 37256 7632
rect 37320 7568 37336 7632
rect 37400 7568 37416 7632
rect 37480 7568 37496 7632
rect 37560 7568 37576 7632
rect 37640 7568 37656 7632
rect 37720 7568 37736 7632
rect 37800 7568 37816 7632
rect 37880 7568 37896 7632
rect 37960 7568 37976 7632
rect 38040 7568 38056 7632
rect 38120 7568 38136 7632
rect 38200 7568 38216 7632
rect 38280 7568 38296 7632
rect 38360 7568 38376 7632
rect 38440 7568 38456 7632
rect 38520 7568 38536 7632
rect 38600 7568 38616 7632
rect 38680 7568 38696 7632
rect 38760 7568 38776 7632
rect 38840 7568 38856 7632
rect 38920 7568 38936 7632
rect 39000 7568 39016 7632
rect 39080 7568 39096 7632
rect 39160 7568 39176 7632
rect 39240 7568 39256 7632
rect 39320 7568 39336 7632
rect 39400 7568 39416 7632
rect 39480 7568 39496 7632
rect 39560 7568 39576 7632
rect 39640 7568 39656 7632
rect 39720 7568 39736 7632
rect 39800 7568 39816 7632
rect 39880 7568 39896 7632
rect 39960 7568 39976 7632
rect 40040 7568 40056 7632
rect 40120 7568 40136 7632
rect 40200 7568 40216 7632
rect 40280 7568 40296 7632
rect 40360 7568 40368 7632
rect 5000 7552 40368 7568
rect 5000 7488 5008 7552
rect 5072 7488 5088 7552
rect 5152 7488 5168 7552
rect 5232 7488 5248 7552
rect 5312 7488 5328 7552
rect 5392 7488 5408 7552
rect 5472 7488 5488 7552
rect 5552 7488 5568 7552
rect 5632 7488 5648 7552
rect 5712 7488 5728 7552
rect 5792 7488 5808 7552
rect 5872 7488 5888 7552
rect 5952 7488 5968 7552
rect 6032 7488 6048 7552
rect 6112 7488 6128 7552
rect 6192 7488 6208 7552
rect 6272 7488 6288 7552
rect 6352 7488 6368 7552
rect 6432 7488 6448 7552
rect 6512 7488 6528 7552
rect 6592 7488 6608 7552
rect 6672 7488 6688 7552
rect 6752 7488 6768 7552
rect 6832 7488 6848 7552
rect 6912 7488 6928 7552
rect 6992 7488 7008 7552
rect 7072 7488 7088 7552
rect 7152 7488 7168 7552
rect 7232 7488 7248 7552
rect 7312 7488 7328 7552
rect 7392 7488 7408 7552
rect 7472 7488 7488 7552
rect 7552 7488 7568 7552
rect 7632 7488 7648 7552
rect 7712 7488 7728 7552
rect 7792 7488 7808 7552
rect 7872 7488 7888 7552
rect 7952 7488 7968 7552
rect 8032 7488 8048 7552
rect 8112 7488 8128 7552
rect 8192 7488 8208 7552
rect 8272 7488 8288 7552
rect 8352 7488 8368 7552
rect 8432 7488 8448 7552
rect 8512 7488 8528 7552
rect 8592 7488 8608 7552
rect 8672 7488 8688 7552
rect 8752 7488 8768 7552
rect 8832 7488 8848 7552
rect 8912 7488 8928 7552
rect 8992 7488 14112 7552
rect 14176 7488 14192 7552
rect 14256 7488 14272 7552
rect 14336 7488 14352 7552
rect 14416 7488 24112 7552
rect 24176 7488 24192 7552
rect 24256 7488 24272 7552
rect 24336 7488 24352 7552
rect 24416 7488 36376 7552
rect 36440 7488 36456 7552
rect 36520 7488 36536 7552
rect 36600 7488 36616 7552
rect 36680 7488 36696 7552
rect 36760 7488 36776 7552
rect 36840 7488 36856 7552
rect 36920 7488 36936 7552
rect 37000 7488 37016 7552
rect 37080 7488 37096 7552
rect 37160 7488 37176 7552
rect 37240 7488 37256 7552
rect 37320 7488 37336 7552
rect 37400 7488 37416 7552
rect 37480 7488 37496 7552
rect 37560 7488 37576 7552
rect 37640 7488 37656 7552
rect 37720 7488 37736 7552
rect 37800 7488 37816 7552
rect 37880 7488 37896 7552
rect 37960 7488 37976 7552
rect 38040 7488 38056 7552
rect 38120 7488 38136 7552
rect 38200 7488 38216 7552
rect 38280 7488 38296 7552
rect 38360 7488 38376 7552
rect 38440 7488 38456 7552
rect 38520 7488 38536 7552
rect 38600 7488 38616 7552
rect 38680 7488 38696 7552
rect 38760 7488 38776 7552
rect 38840 7488 38856 7552
rect 38920 7488 38936 7552
rect 39000 7488 39016 7552
rect 39080 7488 39096 7552
rect 39160 7488 39176 7552
rect 39240 7488 39256 7552
rect 39320 7488 39336 7552
rect 39400 7488 39416 7552
rect 39480 7488 39496 7552
rect 39560 7488 39576 7552
rect 39640 7488 39656 7552
rect 39720 7488 39736 7552
rect 39800 7488 39816 7552
rect 39880 7488 39896 7552
rect 39960 7488 39976 7552
rect 40040 7488 40056 7552
rect 40120 7488 40136 7552
rect 40200 7488 40216 7552
rect 40280 7488 40296 7552
rect 40360 7488 40368 7552
rect 5000 7472 40368 7488
rect 5000 7408 5008 7472
rect 5072 7408 5088 7472
rect 5152 7408 5168 7472
rect 5232 7408 5248 7472
rect 5312 7408 5328 7472
rect 5392 7408 5408 7472
rect 5472 7408 5488 7472
rect 5552 7408 5568 7472
rect 5632 7408 5648 7472
rect 5712 7408 5728 7472
rect 5792 7408 5808 7472
rect 5872 7408 5888 7472
rect 5952 7408 5968 7472
rect 6032 7408 6048 7472
rect 6112 7408 6128 7472
rect 6192 7408 6208 7472
rect 6272 7408 6288 7472
rect 6352 7408 6368 7472
rect 6432 7408 6448 7472
rect 6512 7408 6528 7472
rect 6592 7408 6608 7472
rect 6672 7408 6688 7472
rect 6752 7408 6768 7472
rect 6832 7408 6848 7472
rect 6912 7408 6928 7472
rect 6992 7408 7008 7472
rect 7072 7408 7088 7472
rect 7152 7408 7168 7472
rect 7232 7408 7248 7472
rect 7312 7408 7328 7472
rect 7392 7408 7408 7472
rect 7472 7408 7488 7472
rect 7552 7408 7568 7472
rect 7632 7408 7648 7472
rect 7712 7408 7728 7472
rect 7792 7408 7808 7472
rect 7872 7408 7888 7472
rect 7952 7408 7968 7472
rect 8032 7408 8048 7472
rect 8112 7408 8128 7472
rect 8192 7408 8208 7472
rect 8272 7408 8288 7472
rect 8352 7408 8368 7472
rect 8432 7408 8448 7472
rect 8512 7408 8528 7472
rect 8592 7408 8608 7472
rect 8672 7408 8688 7472
rect 8752 7408 8768 7472
rect 8832 7408 8848 7472
rect 8912 7408 8928 7472
rect 8992 7408 14112 7472
rect 14176 7408 14192 7472
rect 14256 7408 14272 7472
rect 14336 7408 14352 7472
rect 14416 7408 24112 7472
rect 24176 7408 24192 7472
rect 24256 7408 24272 7472
rect 24336 7408 24352 7472
rect 24416 7408 36376 7472
rect 36440 7408 36456 7472
rect 36520 7408 36536 7472
rect 36600 7408 36616 7472
rect 36680 7408 36696 7472
rect 36760 7408 36776 7472
rect 36840 7408 36856 7472
rect 36920 7408 36936 7472
rect 37000 7408 37016 7472
rect 37080 7408 37096 7472
rect 37160 7408 37176 7472
rect 37240 7408 37256 7472
rect 37320 7408 37336 7472
rect 37400 7408 37416 7472
rect 37480 7408 37496 7472
rect 37560 7408 37576 7472
rect 37640 7408 37656 7472
rect 37720 7408 37736 7472
rect 37800 7408 37816 7472
rect 37880 7408 37896 7472
rect 37960 7408 37976 7472
rect 38040 7408 38056 7472
rect 38120 7408 38136 7472
rect 38200 7408 38216 7472
rect 38280 7408 38296 7472
rect 38360 7408 38376 7472
rect 38440 7408 38456 7472
rect 38520 7408 38536 7472
rect 38600 7408 38616 7472
rect 38680 7408 38696 7472
rect 38760 7408 38776 7472
rect 38840 7408 38856 7472
rect 38920 7408 38936 7472
rect 39000 7408 39016 7472
rect 39080 7408 39096 7472
rect 39160 7408 39176 7472
rect 39240 7408 39256 7472
rect 39320 7408 39336 7472
rect 39400 7408 39416 7472
rect 39480 7408 39496 7472
rect 39560 7408 39576 7472
rect 39640 7408 39656 7472
rect 39720 7408 39736 7472
rect 39800 7408 39816 7472
rect 39880 7408 39896 7472
rect 39960 7408 39976 7472
rect 40040 7408 40056 7472
rect 40120 7408 40136 7472
rect 40200 7408 40216 7472
rect 40280 7408 40296 7472
rect 40360 7408 40368 7472
rect 5000 7392 40368 7408
rect 5000 7328 5008 7392
rect 5072 7328 5088 7392
rect 5152 7328 5168 7392
rect 5232 7328 5248 7392
rect 5312 7328 5328 7392
rect 5392 7328 5408 7392
rect 5472 7328 5488 7392
rect 5552 7328 5568 7392
rect 5632 7328 5648 7392
rect 5712 7328 5728 7392
rect 5792 7328 5808 7392
rect 5872 7328 5888 7392
rect 5952 7328 5968 7392
rect 6032 7328 6048 7392
rect 6112 7328 6128 7392
rect 6192 7328 6208 7392
rect 6272 7328 6288 7392
rect 6352 7328 6368 7392
rect 6432 7328 6448 7392
rect 6512 7328 6528 7392
rect 6592 7328 6608 7392
rect 6672 7328 6688 7392
rect 6752 7328 6768 7392
rect 6832 7328 6848 7392
rect 6912 7328 6928 7392
rect 6992 7328 7008 7392
rect 7072 7328 7088 7392
rect 7152 7328 7168 7392
rect 7232 7328 7248 7392
rect 7312 7328 7328 7392
rect 7392 7328 7408 7392
rect 7472 7328 7488 7392
rect 7552 7328 7568 7392
rect 7632 7328 7648 7392
rect 7712 7328 7728 7392
rect 7792 7328 7808 7392
rect 7872 7328 7888 7392
rect 7952 7328 7968 7392
rect 8032 7328 8048 7392
rect 8112 7328 8128 7392
rect 8192 7328 8208 7392
rect 8272 7328 8288 7392
rect 8352 7328 8368 7392
rect 8432 7328 8448 7392
rect 8512 7328 8528 7392
rect 8592 7328 8608 7392
rect 8672 7328 8688 7392
rect 8752 7328 8768 7392
rect 8832 7328 8848 7392
rect 8912 7328 8928 7392
rect 8992 7328 14112 7392
rect 14176 7328 14192 7392
rect 14256 7328 14272 7392
rect 14336 7328 14352 7392
rect 14416 7328 24112 7392
rect 24176 7328 24192 7392
rect 24256 7328 24272 7392
rect 24336 7328 24352 7392
rect 24416 7328 36376 7392
rect 36440 7328 36456 7392
rect 36520 7328 36536 7392
rect 36600 7328 36616 7392
rect 36680 7328 36696 7392
rect 36760 7328 36776 7392
rect 36840 7328 36856 7392
rect 36920 7328 36936 7392
rect 37000 7328 37016 7392
rect 37080 7328 37096 7392
rect 37160 7328 37176 7392
rect 37240 7328 37256 7392
rect 37320 7328 37336 7392
rect 37400 7328 37416 7392
rect 37480 7328 37496 7392
rect 37560 7328 37576 7392
rect 37640 7328 37656 7392
rect 37720 7328 37736 7392
rect 37800 7328 37816 7392
rect 37880 7328 37896 7392
rect 37960 7328 37976 7392
rect 38040 7328 38056 7392
rect 38120 7328 38136 7392
rect 38200 7328 38216 7392
rect 38280 7328 38296 7392
rect 38360 7328 38376 7392
rect 38440 7328 38456 7392
rect 38520 7328 38536 7392
rect 38600 7328 38616 7392
rect 38680 7328 38696 7392
rect 38760 7328 38776 7392
rect 38840 7328 38856 7392
rect 38920 7328 38936 7392
rect 39000 7328 39016 7392
rect 39080 7328 39096 7392
rect 39160 7328 39176 7392
rect 39240 7328 39256 7392
rect 39320 7328 39336 7392
rect 39400 7328 39416 7392
rect 39480 7328 39496 7392
rect 39560 7328 39576 7392
rect 39640 7328 39656 7392
rect 39720 7328 39736 7392
rect 39800 7328 39816 7392
rect 39880 7328 39896 7392
rect 39960 7328 39976 7392
rect 40040 7328 40056 7392
rect 40120 7328 40136 7392
rect 40200 7328 40216 7392
rect 40280 7328 40296 7392
rect 40360 7328 40368 7392
rect 5000 7312 40368 7328
rect 5000 7248 5008 7312
rect 5072 7248 5088 7312
rect 5152 7248 5168 7312
rect 5232 7248 5248 7312
rect 5312 7248 5328 7312
rect 5392 7248 5408 7312
rect 5472 7248 5488 7312
rect 5552 7248 5568 7312
rect 5632 7248 5648 7312
rect 5712 7248 5728 7312
rect 5792 7248 5808 7312
rect 5872 7248 5888 7312
rect 5952 7248 5968 7312
rect 6032 7248 6048 7312
rect 6112 7248 6128 7312
rect 6192 7248 6208 7312
rect 6272 7248 6288 7312
rect 6352 7248 6368 7312
rect 6432 7248 6448 7312
rect 6512 7248 6528 7312
rect 6592 7248 6608 7312
rect 6672 7248 6688 7312
rect 6752 7248 6768 7312
rect 6832 7248 6848 7312
rect 6912 7248 6928 7312
rect 6992 7248 7008 7312
rect 7072 7248 7088 7312
rect 7152 7248 7168 7312
rect 7232 7248 7248 7312
rect 7312 7248 7328 7312
rect 7392 7248 7408 7312
rect 7472 7248 7488 7312
rect 7552 7248 7568 7312
rect 7632 7248 7648 7312
rect 7712 7248 7728 7312
rect 7792 7248 7808 7312
rect 7872 7248 7888 7312
rect 7952 7248 7968 7312
rect 8032 7248 8048 7312
rect 8112 7248 8128 7312
rect 8192 7248 8208 7312
rect 8272 7248 8288 7312
rect 8352 7248 8368 7312
rect 8432 7248 8448 7312
rect 8512 7248 8528 7312
rect 8592 7248 8608 7312
rect 8672 7248 8688 7312
rect 8752 7248 8768 7312
rect 8832 7248 8848 7312
rect 8912 7248 8928 7312
rect 8992 7248 14112 7312
rect 14176 7248 14192 7312
rect 14256 7248 14272 7312
rect 14336 7248 14352 7312
rect 14416 7248 24112 7312
rect 24176 7248 24192 7312
rect 24256 7248 24272 7312
rect 24336 7248 24352 7312
rect 24416 7248 36376 7312
rect 36440 7248 36456 7312
rect 36520 7248 36536 7312
rect 36600 7248 36616 7312
rect 36680 7248 36696 7312
rect 36760 7248 36776 7312
rect 36840 7248 36856 7312
rect 36920 7248 36936 7312
rect 37000 7248 37016 7312
rect 37080 7248 37096 7312
rect 37160 7248 37176 7312
rect 37240 7248 37256 7312
rect 37320 7248 37336 7312
rect 37400 7248 37416 7312
rect 37480 7248 37496 7312
rect 37560 7248 37576 7312
rect 37640 7248 37656 7312
rect 37720 7248 37736 7312
rect 37800 7248 37816 7312
rect 37880 7248 37896 7312
rect 37960 7248 37976 7312
rect 38040 7248 38056 7312
rect 38120 7248 38136 7312
rect 38200 7248 38216 7312
rect 38280 7248 38296 7312
rect 38360 7248 38376 7312
rect 38440 7248 38456 7312
rect 38520 7248 38536 7312
rect 38600 7248 38616 7312
rect 38680 7248 38696 7312
rect 38760 7248 38776 7312
rect 38840 7248 38856 7312
rect 38920 7248 38936 7312
rect 39000 7248 39016 7312
rect 39080 7248 39096 7312
rect 39160 7248 39176 7312
rect 39240 7248 39256 7312
rect 39320 7248 39336 7312
rect 39400 7248 39416 7312
rect 39480 7248 39496 7312
rect 39560 7248 39576 7312
rect 39640 7248 39656 7312
rect 39720 7248 39736 7312
rect 39800 7248 39816 7312
rect 39880 7248 39896 7312
rect 39960 7248 39976 7312
rect 40040 7248 40056 7312
rect 40120 7248 40136 7312
rect 40200 7248 40216 7312
rect 40280 7248 40296 7312
rect 40360 7248 40368 7312
rect 5000 7232 40368 7248
rect 5000 7168 5008 7232
rect 5072 7168 5088 7232
rect 5152 7168 5168 7232
rect 5232 7168 5248 7232
rect 5312 7168 5328 7232
rect 5392 7168 5408 7232
rect 5472 7168 5488 7232
rect 5552 7168 5568 7232
rect 5632 7168 5648 7232
rect 5712 7168 5728 7232
rect 5792 7168 5808 7232
rect 5872 7168 5888 7232
rect 5952 7168 5968 7232
rect 6032 7168 6048 7232
rect 6112 7168 6128 7232
rect 6192 7168 6208 7232
rect 6272 7168 6288 7232
rect 6352 7168 6368 7232
rect 6432 7168 6448 7232
rect 6512 7168 6528 7232
rect 6592 7168 6608 7232
rect 6672 7168 6688 7232
rect 6752 7168 6768 7232
rect 6832 7168 6848 7232
rect 6912 7168 6928 7232
rect 6992 7168 7008 7232
rect 7072 7168 7088 7232
rect 7152 7168 7168 7232
rect 7232 7168 7248 7232
rect 7312 7168 7328 7232
rect 7392 7168 7408 7232
rect 7472 7168 7488 7232
rect 7552 7168 7568 7232
rect 7632 7168 7648 7232
rect 7712 7168 7728 7232
rect 7792 7168 7808 7232
rect 7872 7168 7888 7232
rect 7952 7168 7968 7232
rect 8032 7168 8048 7232
rect 8112 7168 8128 7232
rect 8192 7168 8208 7232
rect 8272 7168 8288 7232
rect 8352 7168 8368 7232
rect 8432 7168 8448 7232
rect 8512 7168 8528 7232
rect 8592 7168 8608 7232
rect 8672 7168 8688 7232
rect 8752 7168 8768 7232
rect 8832 7168 8848 7232
rect 8912 7168 8928 7232
rect 8992 7168 14112 7232
rect 14176 7168 14192 7232
rect 14256 7168 14272 7232
rect 14336 7168 14352 7232
rect 14416 7168 24112 7232
rect 24176 7168 24192 7232
rect 24256 7168 24272 7232
rect 24336 7168 24352 7232
rect 24416 7168 36376 7232
rect 36440 7168 36456 7232
rect 36520 7168 36536 7232
rect 36600 7168 36616 7232
rect 36680 7168 36696 7232
rect 36760 7168 36776 7232
rect 36840 7168 36856 7232
rect 36920 7168 36936 7232
rect 37000 7168 37016 7232
rect 37080 7168 37096 7232
rect 37160 7168 37176 7232
rect 37240 7168 37256 7232
rect 37320 7168 37336 7232
rect 37400 7168 37416 7232
rect 37480 7168 37496 7232
rect 37560 7168 37576 7232
rect 37640 7168 37656 7232
rect 37720 7168 37736 7232
rect 37800 7168 37816 7232
rect 37880 7168 37896 7232
rect 37960 7168 37976 7232
rect 38040 7168 38056 7232
rect 38120 7168 38136 7232
rect 38200 7168 38216 7232
rect 38280 7168 38296 7232
rect 38360 7168 38376 7232
rect 38440 7168 38456 7232
rect 38520 7168 38536 7232
rect 38600 7168 38616 7232
rect 38680 7168 38696 7232
rect 38760 7168 38776 7232
rect 38840 7168 38856 7232
rect 38920 7168 38936 7232
rect 39000 7168 39016 7232
rect 39080 7168 39096 7232
rect 39160 7168 39176 7232
rect 39240 7168 39256 7232
rect 39320 7168 39336 7232
rect 39400 7168 39416 7232
rect 39480 7168 39496 7232
rect 39560 7168 39576 7232
rect 39640 7168 39656 7232
rect 39720 7168 39736 7232
rect 39800 7168 39816 7232
rect 39880 7168 39896 7232
rect 39960 7168 39976 7232
rect 40040 7168 40056 7232
rect 40120 7168 40136 7232
rect 40200 7168 40216 7232
rect 40280 7168 40296 7232
rect 40360 7168 40368 7232
rect 5000 7152 40368 7168
rect 5000 7088 5008 7152
rect 5072 7088 5088 7152
rect 5152 7088 5168 7152
rect 5232 7088 5248 7152
rect 5312 7088 5328 7152
rect 5392 7088 5408 7152
rect 5472 7088 5488 7152
rect 5552 7088 5568 7152
rect 5632 7088 5648 7152
rect 5712 7088 5728 7152
rect 5792 7088 5808 7152
rect 5872 7088 5888 7152
rect 5952 7088 5968 7152
rect 6032 7088 6048 7152
rect 6112 7088 6128 7152
rect 6192 7088 6208 7152
rect 6272 7088 6288 7152
rect 6352 7088 6368 7152
rect 6432 7088 6448 7152
rect 6512 7088 6528 7152
rect 6592 7088 6608 7152
rect 6672 7088 6688 7152
rect 6752 7088 6768 7152
rect 6832 7088 6848 7152
rect 6912 7088 6928 7152
rect 6992 7088 7008 7152
rect 7072 7088 7088 7152
rect 7152 7088 7168 7152
rect 7232 7088 7248 7152
rect 7312 7088 7328 7152
rect 7392 7088 7408 7152
rect 7472 7088 7488 7152
rect 7552 7088 7568 7152
rect 7632 7088 7648 7152
rect 7712 7088 7728 7152
rect 7792 7088 7808 7152
rect 7872 7088 7888 7152
rect 7952 7088 7968 7152
rect 8032 7088 8048 7152
rect 8112 7088 8128 7152
rect 8192 7088 8208 7152
rect 8272 7088 8288 7152
rect 8352 7088 8368 7152
rect 8432 7088 8448 7152
rect 8512 7088 8528 7152
rect 8592 7088 8608 7152
rect 8672 7088 8688 7152
rect 8752 7088 8768 7152
rect 8832 7088 8848 7152
rect 8912 7088 8928 7152
rect 8992 7088 14112 7152
rect 14176 7088 14192 7152
rect 14256 7088 14272 7152
rect 14336 7088 14352 7152
rect 14416 7088 24112 7152
rect 24176 7088 24192 7152
rect 24256 7088 24272 7152
rect 24336 7088 24352 7152
rect 24416 7088 36376 7152
rect 36440 7088 36456 7152
rect 36520 7088 36536 7152
rect 36600 7088 36616 7152
rect 36680 7088 36696 7152
rect 36760 7088 36776 7152
rect 36840 7088 36856 7152
rect 36920 7088 36936 7152
rect 37000 7088 37016 7152
rect 37080 7088 37096 7152
rect 37160 7088 37176 7152
rect 37240 7088 37256 7152
rect 37320 7088 37336 7152
rect 37400 7088 37416 7152
rect 37480 7088 37496 7152
rect 37560 7088 37576 7152
rect 37640 7088 37656 7152
rect 37720 7088 37736 7152
rect 37800 7088 37816 7152
rect 37880 7088 37896 7152
rect 37960 7088 37976 7152
rect 38040 7088 38056 7152
rect 38120 7088 38136 7152
rect 38200 7088 38216 7152
rect 38280 7088 38296 7152
rect 38360 7088 38376 7152
rect 38440 7088 38456 7152
rect 38520 7088 38536 7152
rect 38600 7088 38616 7152
rect 38680 7088 38696 7152
rect 38760 7088 38776 7152
rect 38840 7088 38856 7152
rect 38920 7088 38936 7152
rect 39000 7088 39016 7152
rect 39080 7088 39096 7152
rect 39160 7088 39176 7152
rect 39240 7088 39256 7152
rect 39320 7088 39336 7152
rect 39400 7088 39416 7152
rect 39480 7088 39496 7152
rect 39560 7088 39576 7152
rect 39640 7088 39656 7152
rect 39720 7088 39736 7152
rect 39800 7088 39816 7152
rect 39880 7088 39896 7152
rect 39960 7088 39976 7152
rect 40040 7088 40056 7152
rect 40120 7088 40136 7152
rect 40200 7088 40216 7152
rect 40280 7088 40296 7152
rect 40360 7088 40368 7152
rect 5000 7072 40368 7088
rect 5000 7008 5008 7072
rect 5072 7008 5088 7072
rect 5152 7008 5168 7072
rect 5232 7008 5248 7072
rect 5312 7008 5328 7072
rect 5392 7008 5408 7072
rect 5472 7008 5488 7072
rect 5552 7008 5568 7072
rect 5632 7008 5648 7072
rect 5712 7008 5728 7072
rect 5792 7008 5808 7072
rect 5872 7008 5888 7072
rect 5952 7008 5968 7072
rect 6032 7008 6048 7072
rect 6112 7008 6128 7072
rect 6192 7008 6208 7072
rect 6272 7008 6288 7072
rect 6352 7008 6368 7072
rect 6432 7008 6448 7072
rect 6512 7008 6528 7072
rect 6592 7008 6608 7072
rect 6672 7008 6688 7072
rect 6752 7008 6768 7072
rect 6832 7008 6848 7072
rect 6912 7008 6928 7072
rect 6992 7008 7008 7072
rect 7072 7008 7088 7072
rect 7152 7008 7168 7072
rect 7232 7008 7248 7072
rect 7312 7008 7328 7072
rect 7392 7008 7408 7072
rect 7472 7008 7488 7072
rect 7552 7008 7568 7072
rect 7632 7008 7648 7072
rect 7712 7008 7728 7072
rect 7792 7008 7808 7072
rect 7872 7008 7888 7072
rect 7952 7008 7968 7072
rect 8032 7008 8048 7072
rect 8112 7008 8128 7072
rect 8192 7008 8208 7072
rect 8272 7008 8288 7072
rect 8352 7008 8368 7072
rect 8432 7008 8448 7072
rect 8512 7008 8528 7072
rect 8592 7008 8608 7072
rect 8672 7008 8688 7072
rect 8752 7008 8768 7072
rect 8832 7008 8848 7072
rect 8912 7008 8928 7072
rect 8992 7008 14112 7072
rect 14176 7008 14192 7072
rect 14256 7008 14272 7072
rect 14336 7008 14352 7072
rect 14416 7008 24112 7072
rect 24176 7008 24192 7072
rect 24256 7008 24272 7072
rect 24336 7008 24352 7072
rect 24416 7008 36376 7072
rect 36440 7008 36456 7072
rect 36520 7008 36536 7072
rect 36600 7008 36616 7072
rect 36680 7008 36696 7072
rect 36760 7008 36776 7072
rect 36840 7008 36856 7072
rect 36920 7008 36936 7072
rect 37000 7008 37016 7072
rect 37080 7008 37096 7072
rect 37160 7008 37176 7072
rect 37240 7008 37256 7072
rect 37320 7008 37336 7072
rect 37400 7008 37416 7072
rect 37480 7008 37496 7072
rect 37560 7008 37576 7072
rect 37640 7008 37656 7072
rect 37720 7008 37736 7072
rect 37800 7008 37816 7072
rect 37880 7008 37896 7072
rect 37960 7008 37976 7072
rect 38040 7008 38056 7072
rect 38120 7008 38136 7072
rect 38200 7008 38216 7072
rect 38280 7008 38296 7072
rect 38360 7008 38376 7072
rect 38440 7008 38456 7072
rect 38520 7008 38536 7072
rect 38600 7008 38616 7072
rect 38680 7008 38696 7072
rect 38760 7008 38776 7072
rect 38840 7008 38856 7072
rect 38920 7008 38936 7072
rect 39000 7008 39016 7072
rect 39080 7008 39096 7072
rect 39160 7008 39176 7072
rect 39240 7008 39256 7072
rect 39320 7008 39336 7072
rect 39400 7008 39416 7072
rect 39480 7008 39496 7072
rect 39560 7008 39576 7072
rect 39640 7008 39656 7072
rect 39720 7008 39736 7072
rect 39800 7008 39816 7072
rect 39880 7008 39896 7072
rect 39960 7008 39976 7072
rect 40040 7008 40056 7072
rect 40120 7008 40136 7072
rect 40200 7008 40216 7072
rect 40280 7008 40296 7072
rect 40360 7008 40368 7072
rect 5000 6992 40368 7008
rect 5000 6928 5008 6992
rect 5072 6928 5088 6992
rect 5152 6928 5168 6992
rect 5232 6928 5248 6992
rect 5312 6928 5328 6992
rect 5392 6928 5408 6992
rect 5472 6928 5488 6992
rect 5552 6928 5568 6992
rect 5632 6928 5648 6992
rect 5712 6928 5728 6992
rect 5792 6928 5808 6992
rect 5872 6928 5888 6992
rect 5952 6928 5968 6992
rect 6032 6928 6048 6992
rect 6112 6928 6128 6992
rect 6192 6928 6208 6992
rect 6272 6928 6288 6992
rect 6352 6928 6368 6992
rect 6432 6928 6448 6992
rect 6512 6928 6528 6992
rect 6592 6928 6608 6992
rect 6672 6928 6688 6992
rect 6752 6928 6768 6992
rect 6832 6928 6848 6992
rect 6912 6928 6928 6992
rect 6992 6928 7008 6992
rect 7072 6928 7088 6992
rect 7152 6928 7168 6992
rect 7232 6928 7248 6992
rect 7312 6928 7328 6992
rect 7392 6928 7408 6992
rect 7472 6928 7488 6992
rect 7552 6928 7568 6992
rect 7632 6928 7648 6992
rect 7712 6928 7728 6992
rect 7792 6928 7808 6992
rect 7872 6928 7888 6992
rect 7952 6928 7968 6992
rect 8032 6928 8048 6992
rect 8112 6928 8128 6992
rect 8192 6928 8208 6992
rect 8272 6928 8288 6992
rect 8352 6928 8368 6992
rect 8432 6928 8448 6992
rect 8512 6928 8528 6992
rect 8592 6928 8608 6992
rect 8672 6928 8688 6992
rect 8752 6928 8768 6992
rect 8832 6928 8848 6992
rect 8912 6928 8928 6992
rect 8992 6928 14112 6992
rect 14176 6928 14192 6992
rect 14256 6928 14272 6992
rect 14336 6928 14352 6992
rect 14416 6928 24112 6992
rect 24176 6928 24192 6992
rect 24256 6928 24272 6992
rect 24336 6928 24352 6992
rect 24416 6928 36376 6992
rect 36440 6928 36456 6992
rect 36520 6928 36536 6992
rect 36600 6928 36616 6992
rect 36680 6928 36696 6992
rect 36760 6928 36776 6992
rect 36840 6928 36856 6992
rect 36920 6928 36936 6992
rect 37000 6928 37016 6992
rect 37080 6928 37096 6992
rect 37160 6928 37176 6992
rect 37240 6928 37256 6992
rect 37320 6928 37336 6992
rect 37400 6928 37416 6992
rect 37480 6928 37496 6992
rect 37560 6928 37576 6992
rect 37640 6928 37656 6992
rect 37720 6928 37736 6992
rect 37800 6928 37816 6992
rect 37880 6928 37896 6992
rect 37960 6928 37976 6992
rect 38040 6928 38056 6992
rect 38120 6928 38136 6992
rect 38200 6928 38216 6992
rect 38280 6928 38296 6992
rect 38360 6928 38376 6992
rect 38440 6928 38456 6992
rect 38520 6928 38536 6992
rect 38600 6928 38616 6992
rect 38680 6928 38696 6992
rect 38760 6928 38776 6992
rect 38840 6928 38856 6992
rect 38920 6928 38936 6992
rect 39000 6928 39016 6992
rect 39080 6928 39096 6992
rect 39160 6928 39176 6992
rect 39240 6928 39256 6992
rect 39320 6928 39336 6992
rect 39400 6928 39416 6992
rect 39480 6928 39496 6992
rect 39560 6928 39576 6992
rect 39640 6928 39656 6992
rect 39720 6928 39736 6992
rect 39800 6928 39816 6992
rect 39880 6928 39896 6992
rect 39960 6928 39976 6992
rect 40040 6928 40056 6992
rect 40120 6928 40136 6992
rect 40200 6928 40216 6992
rect 40280 6928 40296 6992
rect 40360 6928 40368 6992
rect 5000 6912 40368 6928
rect 5000 6848 5008 6912
rect 5072 6848 5088 6912
rect 5152 6848 5168 6912
rect 5232 6848 5248 6912
rect 5312 6848 5328 6912
rect 5392 6848 5408 6912
rect 5472 6848 5488 6912
rect 5552 6848 5568 6912
rect 5632 6848 5648 6912
rect 5712 6848 5728 6912
rect 5792 6848 5808 6912
rect 5872 6848 5888 6912
rect 5952 6848 5968 6912
rect 6032 6848 6048 6912
rect 6112 6848 6128 6912
rect 6192 6848 6208 6912
rect 6272 6848 6288 6912
rect 6352 6848 6368 6912
rect 6432 6848 6448 6912
rect 6512 6848 6528 6912
rect 6592 6848 6608 6912
rect 6672 6848 6688 6912
rect 6752 6848 6768 6912
rect 6832 6848 6848 6912
rect 6912 6848 6928 6912
rect 6992 6848 7008 6912
rect 7072 6848 7088 6912
rect 7152 6848 7168 6912
rect 7232 6848 7248 6912
rect 7312 6848 7328 6912
rect 7392 6848 7408 6912
rect 7472 6848 7488 6912
rect 7552 6848 7568 6912
rect 7632 6848 7648 6912
rect 7712 6848 7728 6912
rect 7792 6848 7808 6912
rect 7872 6848 7888 6912
rect 7952 6848 7968 6912
rect 8032 6848 8048 6912
rect 8112 6848 8128 6912
rect 8192 6848 8208 6912
rect 8272 6848 8288 6912
rect 8352 6848 8368 6912
rect 8432 6848 8448 6912
rect 8512 6848 8528 6912
rect 8592 6848 8608 6912
rect 8672 6848 8688 6912
rect 8752 6848 8768 6912
rect 8832 6848 8848 6912
rect 8912 6848 8928 6912
rect 8992 6848 14112 6912
rect 14176 6848 14192 6912
rect 14256 6848 14272 6912
rect 14336 6848 14352 6912
rect 14416 6848 24112 6912
rect 24176 6848 24192 6912
rect 24256 6848 24272 6912
rect 24336 6848 24352 6912
rect 24416 6848 36376 6912
rect 36440 6848 36456 6912
rect 36520 6848 36536 6912
rect 36600 6848 36616 6912
rect 36680 6848 36696 6912
rect 36760 6848 36776 6912
rect 36840 6848 36856 6912
rect 36920 6848 36936 6912
rect 37000 6848 37016 6912
rect 37080 6848 37096 6912
rect 37160 6848 37176 6912
rect 37240 6848 37256 6912
rect 37320 6848 37336 6912
rect 37400 6848 37416 6912
rect 37480 6848 37496 6912
rect 37560 6848 37576 6912
rect 37640 6848 37656 6912
rect 37720 6848 37736 6912
rect 37800 6848 37816 6912
rect 37880 6848 37896 6912
rect 37960 6848 37976 6912
rect 38040 6848 38056 6912
rect 38120 6848 38136 6912
rect 38200 6848 38216 6912
rect 38280 6848 38296 6912
rect 38360 6848 38376 6912
rect 38440 6848 38456 6912
rect 38520 6848 38536 6912
rect 38600 6848 38616 6912
rect 38680 6848 38696 6912
rect 38760 6848 38776 6912
rect 38840 6848 38856 6912
rect 38920 6848 38936 6912
rect 39000 6848 39016 6912
rect 39080 6848 39096 6912
rect 39160 6848 39176 6912
rect 39240 6848 39256 6912
rect 39320 6848 39336 6912
rect 39400 6848 39416 6912
rect 39480 6848 39496 6912
rect 39560 6848 39576 6912
rect 39640 6848 39656 6912
rect 39720 6848 39736 6912
rect 39800 6848 39816 6912
rect 39880 6848 39896 6912
rect 39960 6848 39976 6912
rect 40040 6848 40056 6912
rect 40120 6848 40136 6912
rect 40200 6848 40216 6912
rect 40280 6848 40296 6912
rect 40360 6848 40368 6912
rect 5000 6832 40368 6848
rect 5000 6768 5008 6832
rect 5072 6768 5088 6832
rect 5152 6768 5168 6832
rect 5232 6768 5248 6832
rect 5312 6768 5328 6832
rect 5392 6768 5408 6832
rect 5472 6768 5488 6832
rect 5552 6768 5568 6832
rect 5632 6768 5648 6832
rect 5712 6768 5728 6832
rect 5792 6768 5808 6832
rect 5872 6768 5888 6832
rect 5952 6768 5968 6832
rect 6032 6768 6048 6832
rect 6112 6768 6128 6832
rect 6192 6768 6208 6832
rect 6272 6768 6288 6832
rect 6352 6768 6368 6832
rect 6432 6768 6448 6832
rect 6512 6768 6528 6832
rect 6592 6768 6608 6832
rect 6672 6768 6688 6832
rect 6752 6768 6768 6832
rect 6832 6768 6848 6832
rect 6912 6768 6928 6832
rect 6992 6768 7008 6832
rect 7072 6768 7088 6832
rect 7152 6768 7168 6832
rect 7232 6768 7248 6832
rect 7312 6768 7328 6832
rect 7392 6768 7408 6832
rect 7472 6768 7488 6832
rect 7552 6768 7568 6832
rect 7632 6768 7648 6832
rect 7712 6768 7728 6832
rect 7792 6768 7808 6832
rect 7872 6768 7888 6832
rect 7952 6768 7968 6832
rect 8032 6768 8048 6832
rect 8112 6768 8128 6832
rect 8192 6768 8208 6832
rect 8272 6768 8288 6832
rect 8352 6768 8368 6832
rect 8432 6768 8448 6832
rect 8512 6768 8528 6832
rect 8592 6768 8608 6832
rect 8672 6768 8688 6832
rect 8752 6768 8768 6832
rect 8832 6768 8848 6832
rect 8912 6768 8928 6832
rect 8992 6768 14112 6832
rect 14176 6768 14192 6832
rect 14256 6768 14272 6832
rect 14336 6768 14352 6832
rect 14416 6768 24112 6832
rect 24176 6768 24192 6832
rect 24256 6768 24272 6832
rect 24336 6768 24352 6832
rect 24416 6768 36376 6832
rect 36440 6768 36456 6832
rect 36520 6768 36536 6832
rect 36600 6768 36616 6832
rect 36680 6768 36696 6832
rect 36760 6768 36776 6832
rect 36840 6768 36856 6832
rect 36920 6768 36936 6832
rect 37000 6768 37016 6832
rect 37080 6768 37096 6832
rect 37160 6768 37176 6832
rect 37240 6768 37256 6832
rect 37320 6768 37336 6832
rect 37400 6768 37416 6832
rect 37480 6768 37496 6832
rect 37560 6768 37576 6832
rect 37640 6768 37656 6832
rect 37720 6768 37736 6832
rect 37800 6768 37816 6832
rect 37880 6768 37896 6832
rect 37960 6768 37976 6832
rect 38040 6768 38056 6832
rect 38120 6768 38136 6832
rect 38200 6768 38216 6832
rect 38280 6768 38296 6832
rect 38360 6768 38376 6832
rect 38440 6768 38456 6832
rect 38520 6768 38536 6832
rect 38600 6768 38616 6832
rect 38680 6768 38696 6832
rect 38760 6768 38776 6832
rect 38840 6768 38856 6832
rect 38920 6768 38936 6832
rect 39000 6768 39016 6832
rect 39080 6768 39096 6832
rect 39160 6768 39176 6832
rect 39240 6768 39256 6832
rect 39320 6768 39336 6832
rect 39400 6768 39416 6832
rect 39480 6768 39496 6832
rect 39560 6768 39576 6832
rect 39640 6768 39656 6832
rect 39720 6768 39736 6832
rect 39800 6768 39816 6832
rect 39880 6768 39896 6832
rect 39960 6768 39976 6832
rect 40040 6768 40056 6832
rect 40120 6768 40136 6832
rect 40200 6768 40216 6832
rect 40280 6768 40296 6832
rect 40360 6768 40368 6832
rect 5000 6752 40368 6768
rect 5000 6688 5008 6752
rect 5072 6688 5088 6752
rect 5152 6688 5168 6752
rect 5232 6688 5248 6752
rect 5312 6688 5328 6752
rect 5392 6688 5408 6752
rect 5472 6688 5488 6752
rect 5552 6688 5568 6752
rect 5632 6688 5648 6752
rect 5712 6688 5728 6752
rect 5792 6688 5808 6752
rect 5872 6688 5888 6752
rect 5952 6688 5968 6752
rect 6032 6688 6048 6752
rect 6112 6688 6128 6752
rect 6192 6688 6208 6752
rect 6272 6688 6288 6752
rect 6352 6688 6368 6752
rect 6432 6688 6448 6752
rect 6512 6688 6528 6752
rect 6592 6688 6608 6752
rect 6672 6688 6688 6752
rect 6752 6688 6768 6752
rect 6832 6688 6848 6752
rect 6912 6688 6928 6752
rect 6992 6688 7008 6752
rect 7072 6688 7088 6752
rect 7152 6688 7168 6752
rect 7232 6688 7248 6752
rect 7312 6688 7328 6752
rect 7392 6688 7408 6752
rect 7472 6688 7488 6752
rect 7552 6688 7568 6752
rect 7632 6688 7648 6752
rect 7712 6688 7728 6752
rect 7792 6688 7808 6752
rect 7872 6688 7888 6752
rect 7952 6688 7968 6752
rect 8032 6688 8048 6752
rect 8112 6688 8128 6752
rect 8192 6688 8208 6752
rect 8272 6688 8288 6752
rect 8352 6688 8368 6752
rect 8432 6688 8448 6752
rect 8512 6688 8528 6752
rect 8592 6688 8608 6752
rect 8672 6688 8688 6752
rect 8752 6688 8768 6752
rect 8832 6688 8848 6752
rect 8912 6688 8928 6752
rect 8992 6688 14112 6752
rect 14176 6688 14192 6752
rect 14256 6688 14272 6752
rect 14336 6688 14352 6752
rect 14416 6688 24112 6752
rect 24176 6688 24192 6752
rect 24256 6688 24272 6752
rect 24336 6688 24352 6752
rect 24416 6688 36376 6752
rect 36440 6688 36456 6752
rect 36520 6688 36536 6752
rect 36600 6688 36616 6752
rect 36680 6688 36696 6752
rect 36760 6688 36776 6752
rect 36840 6688 36856 6752
rect 36920 6688 36936 6752
rect 37000 6688 37016 6752
rect 37080 6688 37096 6752
rect 37160 6688 37176 6752
rect 37240 6688 37256 6752
rect 37320 6688 37336 6752
rect 37400 6688 37416 6752
rect 37480 6688 37496 6752
rect 37560 6688 37576 6752
rect 37640 6688 37656 6752
rect 37720 6688 37736 6752
rect 37800 6688 37816 6752
rect 37880 6688 37896 6752
rect 37960 6688 37976 6752
rect 38040 6688 38056 6752
rect 38120 6688 38136 6752
rect 38200 6688 38216 6752
rect 38280 6688 38296 6752
rect 38360 6688 38376 6752
rect 38440 6688 38456 6752
rect 38520 6688 38536 6752
rect 38600 6688 38616 6752
rect 38680 6688 38696 6752
rect 38760 6688 38776 6752
rect 38840 6688 38856 6752
rect 38920 6688 38936 6752
rect 39000 6688 39016 6752
rect 39080 6688 39096 6752
rect 39160 6688 39176 6752
rect 39240 6688 39256 6752
rect 39320 6688 39336 6752
rect 39400 6688 39416 6752
rect 39480 6688 39496 6752
rect 39560 6688 39576 6752
rect 39640 6688 39656 6752
rect 39720 6688 39736 6752
rect 39800 6688 39816 6752
rect 39880 6688 39896 6752
rect 39960 6688 39976 6752
rect 40040 6688 40056 6752
rect 40120 6688 40136 6752
rect 40200 6688 40216 6752
rect 40280 6688 40296 6752
rect 40360 6688 40368 6752
rect 5000 6672 40368 6688
rect 5000 6608 5008 6672
rect 5072 6608 5088 6672
rect 5152 6608 5168 6672
rect 5232 6608 5248 6672
rect 5312 6608 5328 6672
rect 5392 6608 5408 6672
rect 5472 6608 5488 6672
rect 5552 6608 5568 6672
rect 5632 6608 5648 6672
rect 5712 6608 5728 6672
rect 5792 6608 5808 6672
rect 5872 6608 5888 6672
rect 5952 6608 5968 6672
rect 6032 6608 6048 6672
rect 6112 6608 6128 6672
rect 6192 6608 6208 6672
rect 6272 6608 6288 6672
rect 6352 6608 6368 6672
rect 6432 6608 6448 6672
rect 6512 6608 6528 6672
rect 6592 6608 6608 6672
rect 6672 6608 6688 6672
rect 6752 6608 6768 6672
rect 6832 6608 6848 6672
rect 6912 6608 6928 6672
rect 6992 6608 7008 6672
rect 7072 6608 7088 6672
rect 7152 6608 7168 6672
rect 7232 6608 7248 6672
rect 7312 6608 7328 6672
rect 7392 6608 7408 6672
rect 7472 6608 7488 6672
rect 7552 6608 7568 6672
rect 7632 6608 7648 6672
rect 7712 6608 7728 6672
rect 7792 6608 7808 6672
rect 7872 6608 7888 6672
rect 7952 6608 7968 6672
rect 8032 6608 8048 6672
rect 8112 6608 8128 6672
rect 8192 6608 8208 6672
rect 8272 6608 8288 6672
rect 8352 6608 8368 6672
rect 8432 6608 8448 6672
rect 8512 6608 8528 6672
rect 8592 6608 8608 6672
rect 8672 6608 8688 6672
rect 8752 6608 8768 6672
rect 8832 6608 8848 6672
rect 8912 6608 8928 6672
rect 8992 6608 14112 6672
rect 14176 6608 14192 6672
rect 14256 6608 14272 6672
rect 14336 6608 14352 6672
rect 14416 6608 24112 6672
rect 24176 6608 24192 6672
rect 24256 6608 24272 6672
rect 24336 6608 24352 6672
rect 24416 6608 36376 6672
rect 36440 6608 36456 6672
rect 36520 6608 36536 6672
rect 36600 6608 36616 6672
rect 36680 6608 36696 6672
rect 36760 6608 36776 6672
rect 36840 6608 36856 6672
rect 36920 6608 36936 6672
rect 37000 6608 37016 6672
rect 37080 6608 37096 6672
rect 37160 6608 37176 6672
rect 37240 6608 37256 6672
rect 37320 6608 37336 6672
rect 37400 6608 37416 6672
rect 37480 6608 37496 6672
rect 37560 6608 37576 6672
rect 37640 6608 37656 6672
rect 37720 6608 37736 6672
rect 37800 6608 37816 6672
rect 37880 6608 37896 6672
rect 37960 6608 37976 6672
rect 38040 6608 38056 6672
rect 38120 6608 38136 6672
rect 38200 6608 38216 6672
rect 38280 6608 38296 6672
rect 38360 6608 38376 6672
rect 38440 6608 38456 6672
rect 38520 6608 38536 6672
rect 38600 6608 38616 6672
rect 38680 6608 38696 6672
rect 38760 6608 38776 6672
rect 38840 6608 38856 6672
rect 38920 6608 38936 6672
rect 39000 6608 39016 6672
rect 39080 6608 39096 6672
rect 39160 6608 39176 6672
rect 39240 6608 39256 6672
rect 39320 6608 39336 6672
rect 39400 6608 39416 6672
rect 39480 6608 39496 6672
rect 39560 6608 39576 6672
rect 39640 6608 39656 6672
rect 39720 6608 39736 6672
rect 39800 6608 39816 6672
rect 39880 6608 39896 6672
rect 39960 6608 39976 6672
rect 40040 6608 40056 6672
rect 40120 6608 40136 6672
rect 40200 6608 40216 6672
rect 40280 6608 40296 6672
rect 40360 6608 40368 6672
rect 5000 6592 40368 6608
rect 5000 6528 5008 6592
rect 5072 6528 5088 6592
rect 5152 6528 5168 6592
rect 5232 6528 5248 6592
rect 5312 6528 5328 6592
rect 5392 6528 5408 6592
rect 5472 6528 5488 6592
rect 5552 6528 5568 6592
rect 5632 6528 5648 6592
rect 5712 6528 5728 6592
rect 5792 6528 5808 6592
rect 5872 6528 5888 6592
rect 5952 6528 5968 6592
rect 6032 6528 6048 6592
rect 6112 6528 6128 6592
rect 6192 6528 6208 6592
rect 6272 6528 6288 6592
rect 6352 6528 6368 6592
rect 6432 6528 6448 6592
rect 6512 6528 6528 6592
rect 6592 6528 6608 6592
rect 6672 6528 6688 6592
rect 6752 6528 6768 6592
rect 6832 6528 6848 6592
rect 6912 6528 6928 6592
rect 6992 6528 7008 6592
rect 7072 6528 7088 6592
rect 7152 6528 7168 6592
rect 7232 6528 7248 6592
rect 7312 6528 7328 6592
rect 7392 6528 7408 6592
rect 7472 6528 7488 6592
rect 7552 6528 7568 6592
rect 7632 6528 7648 6592
rect 7712 6528 7728 6592
rect 7792 6528 7808 6592
rect 7872 6528 7888 6592
rect 7952 6528 7968 6592
rect 8032 6528 8048 6592
rect 8112 6528 8128 6592
rect 8192 6528 8208 6592
rect 8272 6528 8288 6592
rect 8352 6528 8368 6592
rect 8432 6528 8448 6592
rect 8512 6528 8528 6592
rect 8592 6528 8608 6592
rect 8672 6528 8688 6592
rect 8752 6528 8768 6592
rect 8832 6528 8848 6592
rect 8912 6528 8928 6592
rect 8992 6528 14112 6592
rect 14176 6528 14192 6592
rect 14256 6528 14272 6592
rect 14336 6528 14352 6592
rect 14416 6528 24112 6592
rect 24176 6528 24192 6592
rect 24256 6528 24272 6592
rect 24336 6528 24352 6592
rect 24416 6528 36376 6592
rect 36440 6528 36456 6592
rect 36520 6528 36536 6592
rect 36600 6528 36616 6592
rect 36680 6528 36696 6592
rect 36760 6528 36776 6592
rect 36840 6528 36856 6592
rect 36920 6528 36936 6592
rect 37000 6528 37016 6592
rect 37080 6528 37096 6592
rect 37160 6528 37176 6592
rect 37240 6528 37256 6592
rect 37320 6528 37336 6592
rect 37400 6528 37416 6592
rect 37480 6528 37496 6592
rect 37560 6528 37576 6592
rect 37640 6528 37656 6592
rect 37720 6528 37736 6592
rect 37800 6528 37816 6592
rect 37880 6528 37896 6592
rect 37960 6528 37976 6592
rect 38040 6528 38056 6592
rect 38120 6528 38136 6592
rect 38200 6528 38216 6592
rect 38280 6528 38296 6592
rect 38360 6528 38376 6592
rect 38440 6528 38456 6592
rect 38520 6528 38536 6592
rect 38600 6528 38616 6592
rect 38680 6528 38696 6592
rect 38760 6528 38776 6592
rect 38840 6528 38856 6592
rect 38920 6528 38936 6592
rect 39000 6528 39016 6592
rect 39080 6528 39096 6592
rect 39160 6528 39176 6592
rect 39240 6528 39256 6592
rect 39320 6528 39336 6592
rect 39400 6528 39416 6592
rect 39480 6528 39496 6592
rect 39560 6528 39576 6592
rect 39640 6528 39656 6592
rect 39720 6528 39736 6592
rect 39800 6528 39816 6592
rect 39880 6528 39896 6592
rect 39960 6528 39976 6592
rect 40040 6528 40056 6592
rect 40120 6528 40136 6592
rect 40200 6528 40216 6592
rect 40280 6528 40296 6592
rect 40360 6528 40368 6592
rect 5000 6512 40368 6528
rect 5000 6448 5008 6512
rect 5072 6448 5088 6512
rect 5152 6448 5168 6512
rect 5232 6448 5248 6512
rect 5312 6448 5328 6512
rect 5392 6448 5408 6512
rect 5472 6448 5488 6512
rect 5552 6448 5568 6512
rect 5632 6448 5648 6512
rect 5712 6448 5728 6512
rect 5792 6448 5808 6512
rect 5872 6448 5888 6512
rect 5952 6448 5968 6512
rect 6032 6448 6048 6512
rect 6112 6448 6128 6512
rect 6192 6448 6208 6512
rect 6272 6448 6288 6512
rect 6352 6448 6368 6512
rect 6432 6448 6448 6512
rect 6512 6448 6528 6512
rect 6592 6448 6608 6512
rect 6672 6448 6688 6512
rect 6752 6448 6768 6512
rect 6832 6448 6848 6512
rect 6912 6448 6928 6512
rect 6992 6448 7008 6512
rect 7072 6448 7088 6512
rect 7152 6448 7168 6512
rect 7232 6448 7248 6512
rect 7312 6448 7328 6512
rect 7392 6448 7408 6512
rect 7472 6448 7488 6512
rect 7552 6448 7568 6512
rect 7632 6448 7648 6512
rect 7712 6448 7728 6512
rect 7792 6448 7808 6512
rect 7872 6448 7888 6512
rect 7952 6448 7968 6512
rect 8032 6448 8048 6512
rect 8112 6448 8128 6512
rect 8192 6448 8208 6512
rect 8272 6448 8288 6512
rect 8352 6448 8368 6512
rect 8432 6448 8448 6512
rect 8512 6448 8528 6512
rect 8592 6448 8608 6512
rect 8672 6448 8688 6512
rect 8752 6448 8768 6512
rect 8832 6448 8848 6512
rect 8912 6448 8928 6512
rect 8992 6448 14112 6512
rect 14176 6448 14192 6512
rect 14256 6448 14272 6512
rect 14336 6448 14352 6512
rect 14416 6448 24112 6512
rect 24176 6448 24192 6512
rect 24256 6448 24272 6512
rect 24336 6448 24352 6512
rect 24416 6448 36376 6512
rect 36440 6448 36456 6512
rect 36520 6448 36536 6512
rect 36600 6448 36616 6512
rect 36680 6448 36696 6512
rect 36760 6448 36776 6512
rect 36840 6448 36856 6512
rect 36920 6448 36936 6512
rect 37000 6448 37016 6512
rect 37080 6448 37096 6512
rect 37160 6448 37176 6512
rect 37240 6448 37256 6512
rect 37320 6448 37336 6512
rect 37400 6448 37416 6512
rect 37480 6448 37496 6512
rect 37560 6448 37576 6512
rect 37640 6448 37656 6512
rect 37720 6448 37736 6512
rect 37800 6448 37816 6512
rect 37880 6448 37896 6512
rect 37960 6448 37976 6512
rect 38040 6448 38056 6512
rect 38120 6448 38136 6512
rect 38200 6448 38216 6512
rect 38280 6448 38296 6512
rect 38360 6448 38376 6512
rect 38440 6448 38456 6512
rect 38520 6448 38536 6512
rect 38600 6448 38616 6512
rect 38680 6448 38696 6512
rect 38760 6448 38776 6512
rect 38840 6448 38856 6512
rect 38920 6448 38936 6512
rect 39000 6448 39016 6512
rect 39080 6448 39096 6512
rect 39160 6448 39176 6512
rect 39240 6448 39256 6512
rect 39320 6448 39336 6512
rect 39400 6448 39416 6512
rect 39480 6448 39496 6512
rect 39560 6448 39576 6512
rect 39640 6448 39656 6512
rect 39720 6448 39736 6512
rect 39800 6448 39816 6512
rect 39880 6448 39896 6512
rect 39960 6448 39976 6512
rect 40040 6448 40056 6512
rect 40120 6448 40136 6512
rect 40200 6448 40216 6512
rect 40280 6448 40296 6512
rect 40360 6448 40368 6512
rect 5000 6432 40368 6448
rect 5000 6368 5008 6432
rect 5072 6368 5088 6432
rect 5152 6368 5168 6432
rect 5232 6368 5248 6432
rect 5312 6368 5328 6432
rect 5392 6368 5408 6432
rect 5472 6368 5488 6432
rect 5552 6368 5568 6432
rect 5632 6368 5648 6432
rect 5712 6368 5728 6432
rect 5792 6368 5808 6432
rect 5872 6368 5888 6432
rect 5952 6368 5968 6432
rect 6032 6368 6048 6432
rect 6112 6368 6128 6432
rect 6192 6368 6208 6432
rect 6272 6368 6288 6432
rect 6352 6368 6368 6432
rect 6432 6368 6448 6432
rect 6512 6368 6528 6432
rect 6592 6368 6608 6432
rect 6672 6368 6688 6432
rect 6752 6368 6768 6432
rect 6832 6368 6848 6432
rect 6912 6368 6928 6432
rect 6992 6368 7008 6432
rect 7072 6368 7088 6432
rect 7152 6368 7168 6432
rect 7232 6368 7248 6432
rect 7312 6368 7328 6432
rect 7392 6368 7408 6432
rect 7472 6368 7488 6432
rect 7552 6368 7568 6432
rect 7632 6368 7648 6432
rect 7712 6368 7728 6432
rect 7792 6368 7808 6432
rect 7872 6368 7888 6432
rect 7952 6368 7968 6432
rect 8032 6368 8048 6432
rect 8112 6368 8128 6432
rect 8192 6368 8208 6432
rect 8272 6368 8288 6432
rect 8352 6368 8368 6432
rect 8432 6368 8448 6432
rect 8512 6368 8528 6432
rect 8592 6368 8608 6432
rect 8672 6368 8688 6432
rect 8752 6368 8768 6432
rect 8832 6368 8848 6432
rect 8912 6368 8928 6432
rect 8992 6368 14112 6432
rect 14176 6368 14192 6432
rect 14256 6368 14272 6432
rect 14336 6368 14352 6432
rect 14416 6368 24112 6432
rect 24176 6368 24192 6432
rect 24256 6368 24272 6432
rect 24336 6368 24352 6432
rect 24416 6368 36376 6432
rect 36440 6368 36456 6432
rect 36520 6368 36536 6432
rect 36600 6368 36616 6432
rect 36680 6368 36696 6432
rect 36760 6368 36776 6432
rect 36840 6368 36856 6432
rect 36920 6368 36936 6432
rect 37000 6368 37016 6432
rect 37080 6368 37096 6432
rect 37160 6368 37176 6432
rect 37240 6368 37256 6432
rect 37320 6368 37336 6432
rect 37400 6368 37416 6432
rect 37480 6368 37496 6432
rect 37560 6368 37576 6432
rect 37640 6368 37656 6432
rect 37720 6368 37736 6432
rect 37800 6368 37816 6432
rect 37880 6368 37896 6432
rect 37960 6368 37976 6432
rect 38040 6368 38056 6432
rect 38120 6368 38136 6432
rect 38200 6368 38216 6432
rect 38280 6368 38296 6432
rect 38360 6368 38376 6432
rect 38440 6368 38456 6432
rect 38520 6368 38536 6432
rect 38600 6368 38616 6432
rect 38680 6368 38696 6432
rect 38760 6368 38776 6432
rect 38840 6368 38856 6432
rect 38920 6368 38936 6432
rect 39000 6368 39016 6432
rect 39080 6368 39096 6432
rect 39160 6368 39176 6432
rect 39240 6368 39256 6432
rect 39320 6368 39336 6432
rect 39400 6368 39416 6432
rect 39480 6368 39496 6432
rect 39560 6368 39576 6432
rect 39640 6368 39656 6432
rect 39720 6368 39736 6432
rect 39800 6368 39816 6432
rect 39880 6368 39896 6432
rect 39960 6368 39976 6432
rect 40040 6368 40056 6432
rect 40120 6368 40136 6432
rect 40200 6368 40216 6432
rect 40280 6368 40296 6432
rect 40360 6368 40368 6432
rect 5000 6352 40368 6368
rect 5000 6288 5008 6352
rect 5072 6288 5088 6352
rect 5152 6288 5168 6352
rect 5232 6288 5248 6352
rect 5312 6288 5328 6352
rect 5392 6288 5408 6352
rect 5472 6288 5488 6352
rect 5552 6288 5568 6352
rect 5632 6288 5648 6352
rect 5712 6288 5728 6352
rect 5792 6288 5808 6352
rect 5872 6288 5888 6352
rect 5952 6288 5968 6352
rect 6032 6288 6048 6352
rect 6112 6288 6128 6352
rect 6192 6288 6208 6352
rect 6272 6288 6288 6352
rect 6352 6288 6368 6352
rect 6432 6288 6448 6352
rect 6512 6288 6528 6352
rect 6592 6288 6608 6352
rect 6672 6288 6688 6352
rect 6752 6288 6768 6352
rect 6832 6288 6848 6352
rect 6912 6288 6928 6352
rect 6992 6288 7008 6352
rect 7072 6288 7088 6352
rect 7152 6288 7168 6352
rect 7232 6288 7248 6352
rect 7312 6288 7328 6352
rect 7392 6288 7408 6352
rect 7472 6288 7488 6352
rect 7552 6288 7568 6352
rect 7632 6288 7648 6352
rect 7712 6288 7728 6352
rect 7792 6288 7808 6352
rect 7872 6288 7888 6352
rect 7952 6288 7968 6352
rect 8032 6288 8048 6352
rect 8112 6288 8128 6352
rect 8192 6288 8208 6352
rect 8272 6288 8288 6352
rect 8352 6288 8368 6352
rect 8432 6288 8448 6352
rect 8512 6288 8528 6352
rect 8592 6288 8608 6352
rect 8672 6288 8688 6352
rect 8752 6288 8768 6352
rect 8832 6288 8848 6352
rect 8912 6288 8928 6352
rect 8992 6288 14112 6352
rect 14176 6288 14192 6352
rect 14256 6288 14272 6352
rect 14336 6288 14352 6352
rect 14416 6288 24112 6352
rect 24176 6288 24192 6352
rect 24256 6288 24272 6352
rect 24336 6288 24352 6352
rect 24416 6288 36376 6352
rect 36440 6288 36456 6352
rect 36520 6288 36536 6352
rect 36600 6288 36616 6352
rect 36680 6288 36696 6352
rect 36760 6288 36776 6352
rect 36840 6288 36856 6352
rect 36920 6288 36936 6352
rect 37000 6288 37016 6352
rect 37080 6288 37096 6352
rect 37160 6288 37176 6352
rect 37240 6288 37256 6352
rect 37320 6288 37336 6352
rect 37400 6288 37416 6352
rect 37480 6288 37496 6352
rect 37560 6288 37576 6352
rect 37640 6288 37656 6352
rect 37720 6288 37736 6352
rect 37800 6288 37816 6352
rect 37880 6288 37896 6352
rect 37960 6288 37976 6352
rect 38040 6288 38056 6352
rect 38120 6288 38136 6352
rect 38200 6288 38216 6352
rect 38280 6288 38296 6352
rect 38360 6288 38376 6352
rect 38440 6288 38456 6352
rect 38520 6288 38536 6352
rect 38600 6288 38616 6352
rect 38680 6288 38696 6352
rect 38760 6288 38776 6352
rect 38840 6288 38856 6352
rect 38920 6288 38936 6352
rect 39000 6288 39016 6352
rect 39080 6288 39096 6352
rect 39160 6288 39176 6352
rect 39240 6288 39256 6352
rect 39320 6288 39336 6352
rect 39400 6288 39416 6352
rect 39480 6288 39496 6352
rect 39560 6288 39576 6352
rect 39640 6288 39656 6352
rect 39720 6288 39736 6352
rect 39800 6288 39816 6352
rect 39880 6288 39896 6352
rect 39960 6288 39976 6352
rect 40040 6288 40056 6352
rect 40120 6288 40136 6352
rect 40200 6288 40216 6352
rect 40280 6288 40296 6352
rect 40360 6288 40368 6352
rect 5000 6272 40368 6288
rect 5000 6208 5008 6272
rect 5072 6208 5088 6272
rect 5152 6208 5168 6272
rect 5232 6208 5248 6272
rect 5312 6208 5328 6272
rect 5392 6208 5408 6272
rect 5472 6208 5488 6272
rect 5552 6208 5568 6272
rect 5632 6208 5648 6272
rect 5712 6208 5728 6272
rect 5792 6208 5808 6272
rect 5872 6208 5888 6272
rect 5952 6208 5968 6272
rect 6032 6208 6048 6272
rect 6112 6208 6128 6272
rect 6192 6208 6208 6272
rect 6272 6208 6288 6272
rect 6352 6208 6368 6272
rect 6432 6208 6448 6272
rect 6512 6208 6528 6272
rect 6592 6208 6608 6272
rect 6672 6208 6688 6272
rect 6752 6208 6768 6272
rect 6832 6208 6848 6272
rect 6912 6208 6928 6272
rect 6992 6208 7008 6272
rect 7072 6208 7088 6272
rect 7152 6208 7168 6272
rect 7232 6208 7248 6272
rect 7312 6208 7328 6272
rect 7392 6208 7408 6272
rect 7472 6208 7488 6272
rect 7552 6208 7568 6272
rect 7632 6208 7648 6272
rect 7712 6208 7728 6272
rect 7792 6208 7808 6272
rect 7872 6208 7888 6272
rect 7952 6208 7968 6272
rect 8032 6208 8048 6272
rect 8112 6208 8128 6272
rect 8192 6208 8208 6272
rect 8272 6208 8288 6272
rect 8352 6208 8368 6272
rect 8432 6208 8448 6272
rect 8512 6208 8528 6272
rect 8592 6208 8608 6272
rect 8672 6208 8688 6272
rect 8752 6208 8768 6272
rect 8832 6208 8848 6272
rect 8912 6208 8928 6272
rect 8992 6208 14112 6272
rect 14176 6208 14192 6272
rect 14256 6208 14272 6272
rect 14336 6208 14352 6272
rect 14416 6208 24112 6272
rect 24176 6208 24192 6272
rect 24256 6208 24272 6272
rect 24336 6208 24352 6272
rect 24416 6208 36376 6272
rect 36440 6208 36456 6272
rect 36520 6208 36536 6272
rect 36600 6208 36616 6272
rect 36680 6208 36696 6272
rect 36760 6208 36776 6272
rect 36840 6208 36856 6272
rect 36920 6208 36936 6272
rect 37000 6208 37016 6272
rect 37080 6208 37096 6272
rect 37160 6208 37176 6272
rect 37240 6208 37256 6272
rect 37320 6208 37336 6272
rect 37400 6208 37416 6272
rect 37480 6208 37496 6272
rect 37560 6208 37576 6272
rect 37640 6208 37656 6272
rect 37720 6208 37736 6272
rect 37800 6208 37816 6272
rect 37880 6208 37896 6272
rect 37960 6208 37976 6272
rect 38040 6208 38056 6272
rect 38120 6208 38136 6272
rect 38200 6208 38216 6272
rect 38280 6208 38296 6272
rect 38360 6208 38376 6272
rect 38440 6208 38456 6272
rect 38520 6208 38536 6272
rect 38600 6208 38616 6272
rect 38680 6208 38696 6272
rect 38760 6208 38776 6272
rect 38840 6208 38856 6272
rect 38920 6208 38936 6272
rect 39000 6208 39016 6272
rect 39080 6208 39096 6272
rect 39160 6208 39176 6272
rect 39240 6208 39256 6272
rect 39320 6208 39336 6272
rect 39400 6208 39416 6272
rect 39480 6208 39496 6272
rect 39560 6208 39576 6272
rect 39640 6208 39656 6272
rect 39720 6208 39736 6272
rect 39800 6208 39816 6272
rect 39880 6208 39896 6272
rect 39960 6208 39976 6272
rect 40040 6208 40056 6272
rect 40120 6208 40136 6272
rect 40200 6208 40216 6272
rect 40280 6208 40296 6272
rect 40360 6208 40368 6272
rect 5000 6192 40368 6208
rect 5000 6128 5008 6192
rect 5072 6128 5088 6192
rect 5152 6128 5168 6192
rect 5232 6128 5248 6192
rect 5312 6128 5328 6192
rect 5392 6128 5408 6192
rect 5472 6128 5488 6192
rect 5552 6128 5568 6192
rect 5632 6128 5648 6192
rect 5712 6128 5728 6192
rect 5792 6128 5808 6192
rect 5872 6128 5888 6192
rect 5952 6128 5968 6192
rect 6032 6128 6048 6192
rect 6112 6128 6128 6192
rect 6192 6128 6208 6192
rect 6272 6128 6288 6192
rect 6352 6128 6368 6192
rect 6432 6128 6448 6192
rect 6512 6128 6528 6192
rect 6592 6128 6608 6192
rect 6672 6128 6688 6192
rect 6752 6128 6768 6192
rect 6832 6128 6848 6192
rect 6912 6128 6928 6192
rect 6992 6128 7008 6192
rect 7072 6128 7088 6192
rect 7152 6128 7168 6192
rect 7232 6128 7248 6192
rect 7312 6128 7328 6192
rect 7392 6128 7408 6192
rect 7472 6128 7488 6192
rect 7552 6128 7568 6192
rect 7632 6128 7648 6192
rect 7712 6128 7728 6192
rect 7792 6128 7808 6192
rect 7872 6128 7888 6192
rect 7952 6128 7968 6192
rect 8032 6128 8048 6192
rect 8112 6128 8128 6192
rect 8192 6128 8208 6192
rect 8272 6128 8288 6192
rect 8352 6128 8368 6192
rect 8432 6128 8448 6192
rect 8512 6128 8528 6192
rect 8592 6128 8608 6192
rect 8672 6128 8688 6192
rect 8752 6128 8768 6192
rect 8832 6128 8848 6192
rect 8912 6128 8928 6192
rect 8992 6128 14112 6192
rect 14176 6128 14192 6192
rect 14256 6128 14272 6192
rect 14336 6128 14352 6192
rect 14416 6128 24112 6192
rect 24176 6128 24192 6192
rect 24256 6128 24272 6192
rect 24336 6128 24352 6192
rect 24416 6128 36376 6192
rect 36440 6128 36456 6192
rect 36520 6128 36536 6192
rect 36600 6128 36616 6192
rect 36680 6128 36696 6192
rect 36760 6128 36776 6192
rect 36840 6128 36856 6192
rect 36920 6128 36936 6192
rect 37000 6128 37016 6192
rect 37080 6128 37096 6192
rect 37160 6128 37176 6192
rect 37240 6128 37256 6192
rect 37320 6128 37336 6192
rect 37400 6128 37416 6192
rect 37480 6128 37496 6192
rect 37560 6128 37576 6192
rect 37640 6128 37656 6192
rect 37720 6128 37736 6192
rect 37800 6128 37816 6192
rect 37880 6128 37896 6192
rect 37960 6128 37976 6192
rect 38040 6128 38056 6192
rect 38120 6128 38136 6192
rect 38200 6128 38216 6192
rect 38280 6128 38296 6192
rect 38360 6128 38376 6192
rect 38440 6128 38456 6192
rect 38520 6128 38536 6192
rect 38600 6128 38616 6192
rect 38680 6128 38696 6192
rect 38760 6128 38776 6192
rect 38840 6128 38856 6192
rect 38920 6128 38936 6192
rect 39000 6128 39016 6192
rect 39080 6128 39096 6192
rect 39160 6128 39176 6192
rect 39240 6128 39256 6192
rect 39320 6128 39336 6192
rect 39400 6128 39416 6192
rect 39480 6128 39496 6192
rect 39560 6128 39576 6192
rect 39640 6128 39656 6192
rect 39720 6128 39736 6192
rect 39800 6128 39816 6192
rect 39880 6128 39896 6192
rect 39960 6128 39976 6192
rect 40040 6128 40056 6192
rect 40120 6128 40136 6192
rect 40200 6128 40216 6192
rect 40280 6128 40296 6192
rect 40360 6128 40368 6192
rect 5000 6112 40368 6128
rect 5000 6048 5008 6112
rect 5072 6048 5088 6112
rect 5152 6048 5168 6112
rect 5232 6048 5248 6112
rect 5312 6048 5328 6112
rect 5392 6048 5408 6112
rect 5472 6048 5488 6112
rect 5552 6048 5568 6112
rect 5632 6048 5648 6112
rect 5712 6048 5728 6112
rect 5792 6048 5808 6112
rect 5872 6048 5888 6112
rect 5952 6048 5968 6112
rect 6032 6048 6048 6112
rect 6112 6048 6128 6112
rect 6192 6048 6208 6112
rect 6272 6048 6288 6112
rect 6352 6048 6368 6112
rect 6432 6048 6448 6112
rect 6512 6048 6528 6112
rect 6592 6048 6608 6112
rect 6672 6048 6688 6112
rect 6752 6048 6768 6112
rect 6832 6048 6848 6112
rect 6912 6048 6928 6112
rect 6992 6048 7008 6112
rect 7072 6048 7088 6112
rect 7152 6048 7168 6112
rect 7232 6048 7248 6112
rect 7312 6048 7328 6112
rect 7392 6048 7408 6112
rect 7472 6048 7488 6112
rect 7552 6048 7568 6112
rect 7632 6048 7648 6112
rect 7712 6048 7728 6112
rect 7792 6048 7808 6112
rect 7872 6048 7888 6112
rect 7952 6048 7968 6112
rect 8032 6048 8048 6112
rect 8112 6048 8128 6112
rect 8192 6048 8208 6112
rect 8272 6048 8288 6112
rect 8352 6048 8368 6112
rect 8432 6048 8448 6112
rect 8512 6048 8528 6112
rect 8592 6048 8608 6112
rect 8672 6048 8688 6112
rect 8752 6048 8768 6112
rect 8832 6048 8848 6112
rect 8912 6048 8928 6112
rect 8992 6048 14112 6112
rect 14176 6048 14192 6112
rect 14256 6048 14272 6112
rect 14336 6048 14352 6112
rect 14416 6048 24112 6112
rect 24176 6048 24192 6112
rect 24256 6048 24272 6112
rect 24336 6048 24352 6112
rect 24416 6048 36376 6112
rect 36440 6048 36456 6112
rect 36520 6048 36536 6112
rect 36600 6048 36616 6112
rect 36680 6048 36696 6112
rect 36760 6048 36776 6112
rect 36840 6048 36856 6112
rect 36920 6048 36936 6112
rect 37000 6048 37016 6112
rect 37080 6048 37096 6112
rect 37160 6048 37176 6112
rect 37240 6048 37256 6112
rect 37320 6048 37336 6112
rect 37400 6048 37416 6112
rect 37480 6048 37496 6112
rect 37560 6048 37576 6112
rect 37640 6048 37656 6112
rect 37720 6048 37736 6112
rect 37800 6048 37816 6112
rect 37880 6048 37896 6112
rect 37960 6048 37976 6112
rect 38040 6048 38056 6112
rect 38120 6048 38136 6112
rect 38200 6048 38216 6112
rect 38280 6048 38296 6112
rect 38360 6048 38376 6112
rect 38440 6048 38456 6112
rect 38520 6048 38536 6112
rect 38600 6048 38616 6112
rect 38680 6048 38696 6112
rect 38760 6048 38776 6112
rect 38840 6048 38856 6112
rect 38920 6048 38936 6112
rect 39000 6048 39016 6112
rect 39080 6048 39096 6112
rect 39160 6048 39176 6112
rect 39240 6048 39256 6112
rect 39320 6048 39336 6112
rect 39400 6048 39416 6112
rect 39480 6048 39496 6112
rect 39560 6048 39576 6112
rect 39640 6048 39656 6112
rect 39720 6048 39736 6112
rect 39800 6048 39816 6112
rect 39880 6048 39896 6112
rect 39960 6048 39976 6112
rect 40040 6048 40056 6112
rect 40120 6048 40136 6112
rect 40200 6048 40216 6112
rect 40280 6048 40296 6112
rect 40360 6048 40368 6112
rect 5000 6032 40368 6048
rect 5000 5968 5008 6032
rect 5072 5968 5088 6032
rect 5152 5968 5168 6032
rect 5232 5968 5248 6032
rect 5312 5968 5328 6032
rect 5392 5968 5408 6032
rect 5472 5968 5488 6032
rect 5552 5968 5568 6032
rect 5632 5968 5648 6032
rect 5712 5968 5728 6032
rect 5792 5968 5808 6032
rect 5872 5968 5888 6032
rect 5952 5968 5968 6032
rect 6032 5968 6048 6032
rect 6112 5968 6128 6032
rect 6192 5968 6208 6032
rect 6272 5968 6288 6032
rect 6352 5968 6368 6032
rect 6432 5968 6448 6032
rect 6512 5968 6528 6032
rect 6592 5968 6608 6032
rect 6672 5968 6688 6032
rect 6752 5968 6768 6032
rect 6832 5968 6848 6032
rect 6912 5968 6928 6032
rect 6992 5968 7008 6032
rect 7072 5968 7088 6032
rect 7152 5968 7168 6032
rect 7232 5968 7248 6032
rect 7312 5968 7328 6032
rect 7392 5968 7408 6032
rect 7472 5968 7488 6032
rect 7552 5968 7568 6032
rect 7632 5968 7648 6032
rect 7712 5968 7728 6032
rect 7792 5968 7808 6032
rect 7872 5968 7888 6032
rect 7952 5968 7968 6032
rect 8032 5968 8048 6032
rect 8112 5968 8128 6032
rect 8192 5968 8208 6032
rect 8272 5968 8288 6032
rect 8352 5968 8368 6032
rect 8432 5968 8448 6032
rect 8512 5968 8528 6032
rect 8592 5968 8608 6032
rect 8672 5968 8688 6032
rect 8752 5968 8768 6032
rect 8832 5968 8848 6032
rect 8912 5968 8928 6032
rect 8992 5968 14112 6032
rect 14176 5968 14192 6032
rect 14256 5968 14272 6032
rect 14336 5968 14352 6032
rect 14416 5968 24112 6032
rect 24176 5968 24192 6032
rect 24256 5968 24272 6032
rect 24336 5968 24352 6032
rect 24416 5968 36376 6032
rect 36440 5968 36456 6032
rect 36520 5968 36536 6032
rect 36600 5968 36616 6032
rect 36680 5968 36696 6032
rect 36760 5968 36776 6032
rect 36840 5968 36856 6032
rect 36920 5968 36936 6032
rect 37000 5968 37016 6032
rect 37080 5968 37096 6032
rect 37160 5968 37176 6032
rect 37240 5968 37256 6032
rect 37320 5968 37336 6032
rect 37400 5968 37416 6032
rect 37480 5968 37496 6032
rect 37560 5968 37576 6032
rect 37640 5968 37656 6032
rect 37720 5968 37736 6032
rect 37800 5968 37816 6032
rect 37880 5968 37896 6032
rect 37960 5968 37976 6032
rect 38040 5968 38056 6032
rect 38120 5968 38136 6032
rect 38200 5968 38216 6032
rect 38280 5968 38296 6032
rect 38360 5968 38376 6032
rect 38440 5968 38456 6032
rect 38520 5968 38536 6032
rect 38600 5968 38616 6032
rect 38680 5968 38696 6032
rect 38760 5968 38776 6032
rect 38840 5968 38856 6032
rect 38920 5968 38936 6032
rect 39000 5968 39016 6032
rect 39080 5968 39096 6032
rect 39160 5968 39176 6032
rect 39240 5968 39256 6032
rect 39320 5968 39336 6032
rect 39400 5968 39416 6032
rect 39480 5968 39496 6032
rect 39560 5968 39576 6032
rect 39640 5968 39656 6032
rect 39720 5968 39736 6032
rect 39800 5968 39816 6032
rect 39880 5968 39896 6032
rect 39960 5968 39976 6032
rect 40040 5968 40056 6032
rect 40120 5968 40136 6032
rect 40200 5968 40216 6032
rect 40280 5968 40296 6032
rect 40360 5968 40368 6032
rect 5000 5952 40368 5968
rect 5000 5888 5008 5952
rect 5072 5888 5088 5952
rect 5152 5888 5168 5952
rect 5232 5888 5248 5952
rect 5312 5888 5328 5952
rect 5392 5888 5408 5952
rect 5472 5888 5488 5952
rect 5552 5888 5568 5952
rect 5632 5888 5648 5952
rect 5712 5888 5728 5952
rect 5792 5888 5808 5952
rect 5872 5888 5888 5952
rect 5952 5888 5968 5952
rect 6032 5888 6048 5952
rect 6112 5888 6128 5952
rect 6192 5888 6208 5952
rect 6272 5888 6288 5952
rect 6352 5888 6368 5952
rect 6432 5888 6448 5952
rect 6512 5888 6528 5952
rect 6592 5888 6608 5952
rect 6672 5888 6688 5952
rect 6752 5888 6768 5952
rect 6832 5888 6848 5952
rect 6912 5888 6928 5952
rect 6992 5888 7008 5952
rect 7072 5888 7088 5952
rect 7152 5888 7168 5952
rect 7232 5888 7248 5952
rect 7312 5888 7328 5952
rect 7392 5888 7408 5952
rect 7472 5888 7488 5952
rect 7552 5888 7568 5952
rect 7632 5888 7648 5952
rect 7712 5888 7728 5952
rect 7792 5888 7808 5952
rect 7872 5888 7888 5952
rect 7952 5888 7968 5952
rect 8032 5888 8048 5952
rect 8112 5888 8128 5952
rect 8192 5888 8208 5952
rect 8272 5888 8288 5952
rect 8352 5888 8368 5952
rect 8432 5888 8448 5952
rect 8512 5888 8528 5952
rect 8592 5888 8608 5952
rect 8672 5888 8688 5952
rect 8752 5888 8768 5952
rect 8832 5888 8848 5952
rect 8912 5888 8928 5952
rect 8992 5888 14112 5952
rect 14176 5888 14192 5952
rect 14256 5888 14272 5952
rect 14336 5888 14352 5952
rect 14416 5888 24112 5952
rect 24176 5888 24192 5952
rect 24256 5888 24272 5952
rect 24336 5888 24352 5952
rect 24416 5888 36376 5952
rect 36440 5888 36456 5952
rect 36520 5888 36536 5952
rect 36600 5888 36616 5952
rect 36680 5888 36696 5952
rect 36760 5888 36776 5952
rect 36840 5888 36856 5952
rect 36920 5888 36936 5952
rect 37000 5888 37016 5952
rect 37080 5888 37096 5952
rect 37160 5888 37176 5952
rect 37240 5888 37256 5952
rect 37320 5888 37336 5952
rect 37400 5888 37416 5952
rect 37480 5888 37496 5952
rect 37560 5888 37576 5952
rect 37640 5888 37656 5952
rect 37720 5888 37736 5952
rect 37800 5888 37816 5952
rect 37880 5888 37896 5952
rect 37960 5888 37976 5952
rect 38040 5888 38056 5952
rect 38120 5888 38136 5952
rect 38200 5888 38216 5952
rect 38280 5888 38296 5952
rect 38360 5888 38376 5952
rect 38440 5888 38456 5952
rect 38520 5888 38536 5952
rect 38600 5888 38616 5952
rect 38680 5888 38696 5952
rect 38760 5888 38776 5952
rect 38840 5888 38856 5952
rect 38920 5888 38936 5952
rect 39000 5888 39016 5952
rect 39080 5888 39096 5952
rect 39160 5888 39176 5952
rect 39240 5888 39256 5952
rect 39320 5888 39336 5952
rect 39400 5888 39416 5952
rect 39480 5888 39496 5952
rect 39560 5888 39576 5952
rect 39640 5888 39656 5952
rect 39720 5888 39736 5952
rect 39800 5888 39816 5952
rect 39880 5888 39896 5952
rect 39960 5888 39976 5952
rect 40040 5888 40056 5952
rect 40120 5888 40136 5952
rect 40200 5888 40216 5952
rect 40280 5888 40296 5952
rect 40360 5888 40368 5952
rect 5000 5872 40368 5888
rect 5000 5808 5008 5872
rect 5072 5808 5088 5872
rect 5152 5808 5168 5872
rect 5232 5808 5248 5872
rect 5312 5808 5328 5872
rect 5392 5808 5408 5872
rect 5472 5808 5488 5872
rect 5552 5808 5568 5872
rect 5632 5808 5648 5872
rect 5712 5808 5728 5872
rect 5792 5808 5808 5872
rect 5872 5808 5888 5872
rect 5952 5808 5968 5872
rect 6032 5808 6048 5872
rect 6112 5808 6128 5872
rect 6192 5808 6208 5872
rect 6272 5808 6288 5872
rect 6352 5808 6368 5872
rect 6432 5808 6448 5872
rect 6512 5808 6528 5872
rect 6592 5808 6608 5872
rect 6672 5808 6688 5872
rect 6752 5808 6768 5872
rect 6832 5808 6848 5872
rect 6912 5808 6928 5872
rect 6992 5808 7008 5872
rect 7072 5808 7088 5872
rect 7152 5808 7168 5872
rect 7232 5808 7248 5872
rect 7312 5808 7328 5872
rect 7392 5808 7408 5872
rect 7472 5808 7488 5872
rect 7552 5808 7568 5872
rect 7632 5808 7648 5872
rect 7712 5808 7728 5872
rect 7792 5808 7808 5872
rect 7872 5808 7888 5872
rect 7952 5808 7968 5872
rect 8032 5808 8048 5872
rect 8112 5808 8128 5872
rect 8192 5808 8208 5872
rect 8272 5808 8288 5872
rect 8352 5808 8368 5872
rect 8432 5808 8448 5872
rect 8512 5808 8528 5872
rect 8592 5808 8608 5872
rect 8672 5808 8688 5872
rect 8752 5808 8768 5872
rect 8832 5808 8848 5872
rect 8912 5808 8928 5872
rect 8992 5808 14112 5872
rect 14176 5808 14192 5872
rect 14256 5808 14272 5872
rect 14336 5808 14352 5872
rect 14416 5808 24112 5872
rect 24176 5808 24192 5872
rect 24256 5808 24272 5872
rect 24336 5808 24352 5872
rect 24416 5808 36376 5872
rect 36440 5808 36456 5872
rect 36520 5808 36536 5872
rect 36600 5808 36616 5872
rect 36680 5808 36696 5872
rect 36760 5808 36776 5872
rect 36840 5808 36856 5872
rect 36920 5808 36936 5872
rect 37000 5808 37016 5872
rect 37080 5808 37096 5872
rect 37160 5808 37176 5872
rect 37240 5808 37256 5872
rect 37320 5808 37336 5872
rect 37400 5808 37416 5872
rect 37480 5808 37496 5872
rect 37560 5808 37576 5872
rect 37640 5808 37656 5872
rect 37720 5808 37736 5872
rect 37800 5808 37816 5872
rect 37880 5808 37896 5872
rect 37960 5808 37976 5872
rect 38040 5808 38056 5872
rect 38120 5808 38136 5872
rect 38200 5808 38216 5872
rect 38280 5808 38296 5872
rect 38360 5808 38376 5872
rect 38440 5808 38456 5872
rect 38520 5808 38536 5872
rect 38600 5808 38616 5872
rect 38680 5808 38696 5872
rect 38760 5808 38776 5872
rect 38840 5808 38856 5872
rect 38920 5808 38936 5872
rect 39000 5808 39016 5872
rect 39080 5808 39096 5872
rect 39160 5808 39176 5872
rect 39240 5808 39256 5872
rect 39320 5808 39336 5872
rect 39400 5808 39416 5872
rect 39480 5808 39496 5872
rect 39560 5808 39576 5872
rect 39640 5808 39656 5872
rect 39720 5808 39736 5872
rect 39800 5808 39816 5872
rect 39880 5808 39896 5872
rect 39960 5808 39976 5872
rect 40040 5808 40056 5872
rect 40120 5808 40136 5872
rect 40200 5808 40216 5872
rect 40280 5808 40296 5872
rect 40360 5808 40368 5872
rect 5000 5792 40368 5808
rect 5000 5728 5008 5792
rect 5072 5728 5088 5792
rect 5152 5728 5168 5792
rect 5232 5728 5248 5792
rect 5312 5728 5328 5792
rect 5392 5728 5408 5792
rect 5472 5728 5488 5792
rect 5552 5728 5568 5792
rect 5632 5728 5648 5792
rect 5712 5728 5728 5792
rect 5792 5728 5808 5792
rect 5872 5728 5888 5792
rect 5952 5728 5968 5792
rect 6032 5728 6048 5792
rect 6112 5728 6128 5792
rect 6192 5728 6208 5792
rect 6272 5728 6288 5792
rect 6352 5728 6368 5792
rect 6432 5728 6448 5792
rect 6512 5728 6528 5792
rect 6592 5728 6608 5792
rect 6672 5728 6688 5792
rect 6752 5728 6768 5792
rect 6832 5728 6848 5792
rect 6912 5728 6928 5792
rect 6992 5728 7008 5792
rect 7072 5728 7088 5792
rect 7152 5728 7168 5792
rect 7232 5728 7248 5792
rect 7312 5728 7328 5792
rect 7392 5728 7408 5792
rect 7472 5728 7488 5792
rect 7552 5728 7568 5792
rect 7632 5728 7648 5792
rect 7712 5728 7728 5792
rect 7792 5728 7808 5792
rect 7872 5728 7888 5792
rect 7952 5728 7968 5792
rect 8032 5728 8048 5792
rect 8112 5728 8128 5792
rect 8192 5728 8208 5792
rect 8272 5728 8288 5792
rect 8352 5728 8368 5792
rect 8432 5728 8448 5792
rect 8512 5728 8528 5792
rect 8592 5728 8608 5792
rect 8672 5728 8688 5792
rect 8752 5728 8768 5792
rect 8832 5728 8848 5792
rect 8912 5728 8928 5792
rect 8992 5728 14112 5792
rect 14176 5728 14192 5792
rect 14256 5728 14272 5792
rect 14336 5728 14352 5792
rect 14416 5728 24112 5792
rect 24176 5728 24192 5792
rect 24256 5728 24272 5792
rect 24336 5728 24352 5792
rect 24416 5728 36376 5792
rect 36440 5728 36456 5792
rect 36520 5728 36536 5792
rect 36600 5728 36616 5792
rect 36680 5728 36696 5792
rect 36760 5728 36776 5792
rect 36840 5728 36856 5792
rect 36920 5728 36936 5792
rect 37000 5728 37016 5792
rect 37080 5728 37096 5792
rect 37160 5728 37176 5792
rect 37240 5728 37256 5792
rect 37320 5728 37336 5792
rect 37400 5728 37416 5792
rect 37480 5728 37496 5792
rect 37560 5728 37576 5792
rect 37640 5728 37656 5792
rect 37720 5728 37736 5792
rect 37800 5728 37816 5792
rect 37880 5728 37896 5792
rect 37960 5728 37976 5792
rect 38040 5728 38056 5792
rect 38120 5728 38136 5792
rect 38200 5728 38216 5792
rect 38280 5728 38296 5792
rect 38360 5728 38376 5792
rect 38440 5728 38456 5792
rect 38520 5728 38536 5792
rect 38600 5728 38616 5792
rect 38680 5728 38696 5792
rect 38760 5728 38776 5792
rect 38840 5728 38856 5792
rect 38920 5728 38936 5792
rect 39000 5728 39016 5792
rect 39080 5728 39096 5792
rect 39160 5728 39176 5792
rect 39240 5728 39256 5792
rect 39320 5728 39336 5792
rect 39400 5728 39416 5792
rect 39480 5728 39496 5792
rect 39560 5728 39576 5792
rect 39640 5728 39656 5792
rect 39720 5728 39736 5792
rect 39800 5728 39816 5792
rect 39880 5728 39896 5792
rect 39960 5728 39976 5792
rect 40040 5728 40056 5792
rect 40120 5728 40136 5792
rect 40200 5728 40216 5792
rect 40280 5728 40296 5792
rect 40360 5728 40368 5792
rect 5000 5712 40368 5728
rect 5000 5648 5008 5712
rect 5072 5648 5088 5712
rect 5152 5648 5168 5712
rect 5232 5648 5248 5712
rect 5312 5648 5328 5712
rect 5392 5648 5408 5712
rect 5472 5648 5488 5712
rect 5552 5648 5568 5712
rect 5632 5648 5648 5712
rect 5712 5648 5728 5712
rect 5792 5648 5808 5712
rect 5872 5648 5888 5712
rect 5952 5648 5968 5712
rect 6032 5648 6048 5712
rect 6112 5648 6128 5712
rect 6192 5648 6208 5712
rect 6272 5648 6288 5712
rect 6352 5648 6368 5712
rect 6432 5648 6448 5712
rect 6512 5648 6528 5712
rect 6592 5648 6608 5712
rect 6672 5648 6688 5712
rect 6752 5648 6768 5712
rect 6832 5648 6848 5712
rect 6912 5648 6928 5712
rect 6992 5648 7008 5712
rect 7072 5648 7088 5712
rect 7152 5648 7168 5712
rect 7232 5648 7248 5712
rect 7312 5648 7328 5712
rect 7392 5648 7408 5712
rect 7472 5648 7488 5712
rect 7552 5648 7568 5712
rect 7632 5648 7648 5712
rect 7712 5648 7728 5712
rect 7792 5648 7808 5712
rect 7872 5648 7888 5712
rect 7952 5648 7968 5712
rect 8032 5648 8048 5712
rect 8112 5648 8128 5712
rect 8192 5648 8208 5712
rect 8272 5648 8288 5712
rect 8352 5648 8368 5712
rect 8432 5648 8448 5712
rect 8512 5648 8528 5712
rect 8592 5648 8608 5712
rect 8672 5648 8688 5712
rect 8752 5648 8768 5712
rect 8832 5648 8848 5712
rect 8912 5648 8928 5712
rect 8992 5648 14112 5712
rect 14176 5648 14192 5712
rect 14256 5648 14272 5712
rect 14336 5648 14352 5712
rect 14416 5648 24112 5712
rect 24176 5648 24192 5712
rect 24256 5648 24272 5712
rect 24336 5648 24352 5712
rect 24416 5648 36376 5712
rect 36440 5648 36456 5712
rect 36520 5648 36536 5712
rect 36600 5648 36616 5712
rect 36680 5648 36696 5712
rect 36760 5648 36776 5712
rect 36840 5648 36856 5712
rect 36920 5648 36936 5712
rect 37000 5648 37016 5712
rect 37080 5648 37096 5712
rect 37160 5648 37176 5712
rect 37240 5648 37256 5712
rect 37320 5648 37336 5712
rect 37400 5648 37416 5712
rect 37480 5648 37496 5712
rect 37560 5648 37576 5712
rect 37640 5648 37656 5712
rect 37720 5648 37736 5712
rect 37800 5648 37816 5712
rect 37880 5648 37896 5712
rect 37960 5648 37976 5712
rect 38040 5648 38056 5712
rect 38120 5648 38136 5712
rect 38200 5648 38216 5712
rect 38280 5648 38296 5712
rect 38360 5648 38376 5712
rect 38440 5648 38456 5712
rect 38520 5648 38536 5712
rect 38600 5648 38616 5712
rect 38680 5648 38696 5712
rect 38760 5648 38776 5712
rect 38840 5648 38856 5712
rect 38920 5648 38936 5712
rect 39000 5648 39016 5712
rect 39080 5648 39096 5712
rect 39160 5648 39176 5712
rect 39240 5648 39256 5712
rect 39320 5648 39336 5712
rect 39400 5648 39416 5712
rect 39480 5648 39496 5712
rect 39560 5648 39576 5712
rect 39640 5648 39656 5712
rect 39720 5648 39736 5712
rect 39800 5648 39816 5712
rect 39880 5648 39896 5712
rect 39960 5648 39976 5712
rect 40040 5648 40056 5712
rect 40120 5648 40136 5712
rect 40200 5648 40216 5712
rect 40280 5648 40296 5712
rect 40360 5648 40368 5712
rect 5000 5632 40368 5648
rect 5000 5568 5008 5632
rect 5072 5568 5088 5632
rect 5152 5568 5168 5632
rect 5232 5568 5248 5632
rect 5312 5568 5328 5632
rect 5392 5568 5408 5632
rect 5472 5568 5488 5632
rect 5552 5568 5568 5632
rect 5632 5568 5648 5632
rect 5712 5568 5728 5632
rect 5792 5568 5808 5632
rect 5872 5568 5888 5632
rect 5952 5568 5968 5632
rect 6032 5568 6048 5632
rect 6112 5568 6128 5632
rect 6192 5568 6208 5632
rect 6272 5568 6288 5632
rect 6352 5568 6368 5632
rect 6432 5568 6448 5632
rect 6512 5568 6528 5632
rect 6592 5568 6608 5632
rect 6672 5568 6688 5632
rect 6752 5568 6768 5632
rect 6832 5568 6848 5632
rect 6912 5568 6928 5632
rect 6992 5568 7008 5632
rect 7072 5568 7088 5632
rect 7152 5568 7168 5632
rect 7232 5568 7248 5632
rect 7312 5568 7328 5632
rect 7392 5568 7408 5632
rect 7472 5568 7488 5632
rect 7552 5568 7568 5632
rect 7632 5568 7648 5632
rect 7712 5568 7728 5632
rect 7792 5568 7808 5632
rect 7872 5568 7888 5632
rect 7952 5568 7968 5632
rect 8032 5568 8048 5632
rect 8112 5568 8128 5632
rect 8192 5568 8208 5632
rect 8272 5568 8288 5632
rect 8352 5568 8368 5632
rect 8432 5568 8448 5632
rect 8512 5568 8528 5632
rect 8592 5568 8608 5632
rect 8672 5568 8688 5632
rect 8752 5568 8768 5632
rect 8832 5568 8848 5632
rect 8912 5568 8928 5632
rect 8992 5568 14112 5632
rect 14176 5568 14192 5632
rect 14256 5568 14272 5632
rect 14336 5568 14352 5632
rect 14416 5568 24112 5632
rect 24176 5568 24192 5632
rect 24256 5568 24272 5632
rect 24336 5568 24352 5632
rect 24416 5568 36376 5632
rect 36440 5568 36456 5632
rect 36520 5568 36536 5632
rect 36600 5568 36616 5632
rect 36680 5568 36696 5632
rect 36760 5568 36776 5632
rect 36840 5568 36856 5632
rect 36920 5568 36936 5632
rect 37000 5568 37016 5632
rect 37080 5568 37096 5632
rect 37160 5568 37176 5632
rect 37240 5568 37256 5632
rect 37320 5568 37336 5632
rect 37400 5568 37416 5632
rect 37480 5568 37496 5632
rect 37560 5568 37576 5632
rect 37640 5568 37656 5632
rect 37720 5568 37736 5632
rect 37800 5568 37816 5632
rect 37880 5568 37896 5632
rect 37960 5568 37976 5632
rect 38040 5568 38056 5632
rect 38120 5568 38136 5632
rect 38200 5568 38216 5632
rect 38280 5568 38296 5632
rect 38360 5568 38376 5632
rect 38440 5568 38456 5632
rect 38520 5568 38536 5632
rect 38600 5568 38616 5632
rect 38680 5568 38696 5632
rect 38760 5568 38776 5632
rect 38840 5568 38856 5632
rect 38920 5568 38936 5632
rect 39000 5568 39016 5632
rect 39080 5568 39096 5632
rect 39160 5568 39176 5632
rect 39240 5568 39256 5632
rect 39320 5568 39336 5632
rect 39400 5568 39416 5632
rect 39480 5568 39496 5632
rect 39560 5568 39576 5632
rect 39640 5568 39656 5632
rect 39720 5568 39736 5632
rect 39800 5568 39816 5632
rect 39880 5568 39896 5632
rect 39960 5568 39976 5632
rect 40040 5568 40056 5632
rect 40120 5568 40136 5632
rect 40200 5568 40216 5632
rect 40280 5568 40296 5632
rect 40360 5568 40368 5632
rect 5000 5552 40368 5568
rect 5000 5488 5008 5552
rect 5072 5488 5088 5552
rect 5152 5488 5168 5552
rect 5232 5488 5248 5552
rect 5312 5488 5328 5552
rect 5392 5488 5408 5552
rect 5472 5488 5488 5552
rect 5552 5488 5568 5552
rect 5632 5488 5648 5552
rect 5712 5488 5728 5552
rect 5792 5488 5808 5552
rect 5872 5488 5888 5552
rect 5952 5488 5968 5552
rect 6032 5488 6048 5552
rect 6112 5488 6128 5552
rect 6192 5488 6208 5552
rect 6272 5488 6288 5552
rect 6352 5488 6368 5552
rect 6432 5488 6448 5552
rect 6512 5488 6528 5552
rect 6592 5488 6608 5552
rect 6672 5488 6688 5552
rect 6752 5488 6768 5552
rect 6832 5488 6848 5552
rect 6912 5488 6928 5552
rect 6992 5488 7008 5552
rect 7072 5488 7088 5552
rect 7152 5488 7168 5552
rect 7232 5488 7248 5552
rect 7312 5488 7328 5552
rect 7392 5488 7408 5552
rect 7472 5488 7488 5552
rect 7552 5488 7568 5552
rect 7632 5488 7648 5552
rect 7712 5488 7728 5552
rect 7792 5488 7808 5552
rect 7872 5488 7888 5552
rect 7952 5488 7968 5552
rect 8032 5488 8048 5552
rect 8112 5488 8128 5552
rect 8192 5488 8208 5552
rect 8272 5488 8288 5552
rect 8352 5488 8368 5552
rect 8432 5488 8448 5552
rect 8512 5488 8528 5552
rect 8592 5488 8608 5552
rect 8672 5488 8688 5552
rect 8752 5488 8768 5552
rect 8832 5488 8848 5552
rect 8912 5488 8928 5552
rect 8992 5488 14112 5552
rect 14176 5488 14192 5552
rect 14256 5488 14272 5552
rect 14336 5488 14352 5552
rect 14416 5488 24112 5552
rect 24176 5488 24192 5552
rect 24256 5488 24272 5552
rect 24336 5488 24352 5552
rect 24416 5488 36376 5552
rect 36440 5488 36456 5552
rect 36520 5488 36536 5552
rect 36600 5488 36616 5552
rect 36680 5488 36696 5552
rect 36760 5488 36776 5552
rect 36840 5488 36856 5552
rect 36920 5488 36936 5552
rect 37000 5488 37016 5552
rect 37080 5488 37096 5552
rect 37160 5488 37176 5552
rect 37240 5488 37256 5552
rect 37320 5488 37336 5552
rect 37400 5488 37416 5552
rect 37480 5488 37496 5552
rect 37560 5488 37576 5552
rect 37640 5488 37656 5552
rect 37720 5488 37736 5552
rect 37800 5488 37816 5552
rect 37880 5488 37896 5552
rect 37960 5488 37976 5552
rect 38040 5488 38056 5552
rect 38120 5488 38136 5552
rect 38200 5488 38216 5552
rect 38280 5488 38296 5552
rect 38360 5488 38376 5552
rect 38440 5488 38456 5552
rect 38520 5488 38536 5552
rect 38600 5488 38616 5552
rect 38680 5488 38696 5552
rect 38760 5488 38776 5552
rect 38840 5488 38856 5552
rect 38920 5488 38936 5552
rect 39000 5488 39016 5552
rect 39080 5488 39096 5552
rect 39160 5488 39176 5552
rect 39240 5488 39256 5552
rect 39320 5488 39336 5552
rect 39400 5488 39416 5552
rect 39480 5488 39496 5552
rect 39560 5488 39576 5552
rect 39640 5488 39656 5552
rect 39720 5488 39736 5552
rect 39800 5488 39816 5552
rect 39880 5488 39896 5552
rect 39960 5488 39976 5552
rect 40040 5488 40056 5552
rect 40120 5488 40136 5552
rect 40200 5488 40216 5552
rect 40280 5488 40296 5552
rect 40360 5488 40368 5552
rect 5000 5472 40368 5488
rect 5000 5408 5008 5472
rect 5072 5408 5088 5472
rect 5152 5408 5168 5472
rect 5232 5408 5248 5472
rect 5312 5408 5328 5472
rect 5392 5408 5408 5472
rect 5472 5408 5488 5472
rect 5552 5408 5568 5472
rect 5632 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5968 5472
rect 6032 5408 6048 5472
rect 6112 5408 6128 5472
rect 6192 5408 6208 5472
rect 6272 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6608 5472
rect 6672 5408 6688 5472
rect 6752 5408 6768 5472
rect 6832 5408 6848 5472
rect 6912 5408 6928 5472
rect 6992 5408 7008 5472
rect 7072 5408 7088 5472
rect 7152 5408 7168 5472
rect 7232 5408 7248 5472
rect 7312 5408 7328 5472
rect 7392 5408 7408 5472
rect 7472 5408 7488 5472
rect 7552 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7888 5472
rect 7952 5408 7968 5472
rect 8032 5408 8048 5472
rect 8112 5408 8128 5472
rect 8192 5408 8208 5472
rect 8272 5408 8288 5472
rect 8352 5408 8368 5472
rect 8432 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8768 5472
rect 8832 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 24112 5472
rect 24176 5408 24192 5472
rect 24256 5408 24272 5472
rect 24336 5408 24352 5472
rect 24416 5408 36376 5472
rect 36440 5408 36456 5472
rect 36520 5408 36536 5472
rect 36600 5408 36616 5472
rect 36680 5408 36696 5472
rect 36760 5408 36776 5472
rect 36840 5408 36856 5472
rect 36920 5408 36936 5472
rect 37000 5408 37016 5472
rect 37080 5408 37096 5472
rect 37160 5408 37176 5472
rect 37240 5408 37256 5472
rect 37320 5408 37336 5472
rect 37400 5408 37416 5472
rect 37480 5408 37496 5472
rect 37560 5408 37576 5472
rect 37640 5408 37656 5472
rect 37720 5408 37736 5472
rect 37800 5408 37816 5472
rect 37880 5408 37896 5472
rect 37960 5408 37976 5472
rect 38040 5408 38056 5472
rect 38120 5408 38136 5472
rect 38200 5408 38216 5472
rect 38280 5408 38296 5472
rect 38360 5408 38376 5472
rect 38440 5408 38456 5472
rect 38520 5408 38536 5472
rect 38600 5408 38616 5472
rect 38680 5408 38696 5472
rect 38760 5408 38776 5472
rect 38840 5408 38856 5472
rect 38920 5408 38936 5472
rect 39000 5408 39016 5472
rect 39080 5408 39096 5472
rect 39160 5408 39176 5472
rect 39240 5408 39256 5472
rect 39320 5408 39336 5472
rect 39400 5408 39416 5472
rect 39480 5408 39496 5472
rect 39560 5408 39576 5472
rect 39640 5408 39656 5472
rect 39720 5408 39736 5472
rect 39800 5408 39816 5472
rect 39880 5408 39896 5472
rect 39960 5408 39976 5472
rect 40040 5408 40056 5472
rect 40120 5408 40136 5472
rect 40200 5408 40216 5472
rect 40280 5408 40296 5472
rect 40360 5408 40368 5472
rect 5000 5392 40368 5408
rect 5000 5328 5008 5392
rect 5072 5328 5088 5392
rect 5152 5328 5168 5392
rect 5232 5328 5248 5392
rect 5312 5328 5328 5392
rect 5392 5328 5408 5392
rect 5472 5328 5488 5392
rect 5552 5328 5568 5392
rect 5632 5328 5648 5392
rect 5712 5328 5728 5392
rect 5792 5328 5808 5392
rect 5872 5328 5888 5392
rect 5952 5328 5968 5392
rect 6032 5328 6048 5392
rect 6112 5328 6128 5392
rect 6192 5328 6208 5392
rect 6272 5328 6288 5392
rect 6352 5328 6368 5392
rect 6432 5328 6448 5392
rect 6512 5328 6528 5392
rect 6592 5328 6608 5392
rect 6672 5328 6688 5392
rect 6752 5328 6768 5392
rect 6832 5328 6848 5392
rect 6912 5328 6928 5392
rect 6992 5328 7008 5392
rect 7072 5328 7088 5392
rect 7152 5328 7168 5392
rect 7232 5328 7248 5392
rect 7312 5328 7328 5392
rect 7392 5328 7408 5392
rect 7472 5328 7488 5392
rect 7552 5328 7568 5392
rect 7632 5328 7648 5392
rect 7712 5328 7728 5392
rect 7792 5328 7808 5392
rect 7872 5328 7888 5392
rect 7952 5328 7968 5392
rect 8032 5328 8048 5392
rect 8112 5328 8128 5392
rect 8192 5328 8208 5392
rect 8272 5328 8288 5392
rect 8352 5328 8368 5392
rect 8432 5328 8448 5392
rect 8512 5328 8528 5392
rect 8592 5328 8608 5392
rect 8672 5328 8688 5392
rect 8752 5328 8768 5392
rect 8832 5328 8848 5392
rect 8912 5328 8928 5392
rect 8992 5328 14112 5392
rect 14176 5328 14192 5392
rect 14256 5328 14272 5392
rect 14336 5328 14352 5392
rect 14416 5328 24112 5392
rect 24176 5328 24192 5392
rect 24256 5328 24272 5392
rect 24336 5328 24352 5392
rect 24416 5328 36376 5392
rect 36440 5328 36456 5392
rect 36520 5328 36536 5392
rect 36600 5328 36616 5392
rect 36680 5328 36696 5392
rect 36760 5328 36776 5392
rect 36840 5328 36856 5392
rect 36920 5328 36936 5392
rect 37000 5328 37016 5392
rect 37080 5328 37096 5392
rect 37160 5328 37176 5392
rect 37240 5328 37256 5392
rect 37320 5328 37336 5392
rect 37400 5328 37416 5392
rect 37480 5328 37496 5392
rect 37560 5328 37576 5392
rect 37640 5328 37656 5392
rect 37720 5328 37736 5392
rect 37800 5328 37816 5392
rect 37880 5328 37896 5392
rect 37960 5328 37976 5392
rect 38040 5328 38056 5392
rect 38120 5328 38136 5392
rect 38200 5328 38216 5392
rect 38280 5328 38296 5392
rect 38360 5328 38376 5392
rect 38440 5328 38456 5392
rect 38520 5328 38536 5392
rect 38600 5328 38616 5392
rect 38680 5328 38696 5392
rect 38760 5328 38776 5392
rect 38840 5328 38856 5392
rect 38920 5328 38936 5392
rect 39000 5328 39016 5392
rect 39080 5328 39096 5392
rect 39160 5328 39176 5392
rect 39240 5328 39256 5392
rect 39320 5328 39336 5392
rect 39400 5328 39416 5392
rect 39480 5328 39496 5392
rect 39560 5328 39576 5392
rect 39640 5328 39656 5392
rect 39720 5328 39736 5392
rect 39800 5328 39816 5392
rect 39880 5328 39896 5392
rect 39960 5328 39976 5392
rect 40040 5328 40056 5392
rect 40120 5328 40136 5392
rect 40200 5328 40216 5392
rect 40280 5328 40296 5392
rect 40360 5328 40368 5392
rect 5000 5312 40368 5328
rect 5000 5248 5008 5312
rect 5072 5248 5088 5312
rect 5152 5248 5168 5312
rect 5232 5248 5248 5312
rect 5312 5248 5328 5312
rect 5392 5248 5408 5312
rect 5472 5248 5488 5312
rect 5552 5248 5568 5312
rect 5632 5248 5648 5312
rect 5712 5248 5728 5312
rect 5792 5248 5808 5312
rect 5872 5248 5888 5312
rect 5952 5248 5968 5312
rect 6032 5248 6048 5312
rect 6112 5248 6128 5312
rect 6192 5248 6208 5312
rect 6272 5248 6288 5312
rect 6352 5248 6368 5312
rect 6432 5248 6448 5312
rect 6512 5248 6528 5312
rect 6592 5248 6608 5312
rect 6672 5248 6688 5312
rect 6752 5248 6768 5312
rect 6832 5248 6848 5312
rect 6912 5248 6928 5312
rect 6992 5248 7008 5312
rect 7072 5248 7088 5312
rect 7152 5248 7168 5312
rect 7232 5248 7248 5312
rect 7312 5248 7328 5312
rect 7392 5248 7408 5312
rect 7472 5248 7488 5312
rect 7552 5248 7568 5312
rect 7632 5248 7648 5312
rect 7712 5248 7728 5312
rect 7792 5248 7808 5312
rect 7872 5248 7888 5312
rect 7952 5248 7968 5312
rect 8032 5248 8048 5312
rect 8112 5248 8128 5312
rect 8192 5248 8208 5312
rect 8272 5248 8288 5312
rect 8352 5248 8368 5312
rect 8432 5248 8448 5312
rect 8512 5248 8528 5312
rect 8592 5248 8608 5312
rect 8672 5248 8688 5312
rect 8752 5248 8768 5312
rect 8832 5248 8848 5312
rect 8912 5248 8928 5312
rect 8992 5248 14112 5312
rect 14176 5248 14192 5312
rect 14256 5248 14272 5312
rect 14336 5248 14352 5312
rect 14416 5248 24112 5312
rect 24176 5248 24192 5312
rect 24256 5248 24272 5312
rect 24336 5248 24352 5312
rect 24416 5248 36376 5312
rect 36440 5248 36456 5312
rect 36520 5248 36536 5312
rect 36600 5248 36616 5312
rect 36680 5248 36696 5312
rect 36760 5248 36776 5312
rect 36840 5248 36856 5312
rect 36920 5248 36936 5312
rect 37000 5248 37016 5312
rect 37080 5248 37096 5312
rect 37160 5248 37176 5312
rect 37240 5248 37256 5312
rect 37320 5248 37336 5312
rect 37400 5248 37416 5312
rect 37480 5248 37496 5312
rect 37560 5248 37576 5312
rect 37640 5248 37656 5312
rect 37720 5248 37736 5312
rect 37800 5248 37816 5312
rect 37880 5248 37896 5312
rect 37960 5248 37976 5312
rect 38040 5248 38056 5312
rect 38120 5248 38136 5312
rect 38200 5248 38216 5312
rect 38280 5248 38296 5312
rect 38360 5248 38376 5312
rect 38440 5248 38456 5312
rect 38520 5248 38536 5312
rect 38600 5248 38616 5312
rect 38680 5248 38696 5312
rect 38760 5248 38776 5312
rect 38840 5248 38856 5312
rect 38920 5248 38936 5312
rect 39000 5248 39016 5312
rect 39080 5248 39096 5312
rect 39160 5248 39176 5312
rect 39240 5248 39256 5312
rect 39320 5248 39336 5312
rect 39400 5248 39416 5312
rect 39480 5248 39496 5312
rect 39560 5248 39576 5312
rect 39640 5248 39656 5312
rect 39720 5248 39736 5312
rect 39800 5248 39816 5312
rect 39880 5248 39896 5312
rect 39960 5248 39976 5312
rect 40040 5248 40056 5312
rect 40120 5248 40136 5312
rect 40200 5248 40216 5312
rect 40280 5248 40296 5312
rect 40360 5248 40368 5312
rect 5000 5232 40368 5248
rect 5000 5168 5008 5232
rect 5072 5168 5088 5232
rect 5152 5168 5168 5232
rect 5232 5168 5248 5232
rect 5312 5168 5328 5232
rect 5392 5168 5408 5232
rect 5472 5168 5488 5232
rect 5552 5168 5568 5232
rect 5632 5168 5648 5232
rect 5712 5168 5728 5232
rect 5792 5168 5808 5232
rect 5872 5168 5888 5232
rect 5952 5168 5968 5232
rect 6032 5168 6048 5232
rect 6112 5168 6128 5232
rect 6192 5168 6208 5232
rect 6272 5168 6288 5232
rect 6352 5168 6368 5232
rect 6432 5168 6448 5232
rect 6512 5168 6528 5232
rect 6592 5168 6608 5232
rect 6672 5168 6688 5232
rect 6752 5168 6768 5232
rect 6832 5168 6848 5232
rect 6912 5168 6928 5232
rect 6992 5168 7008 5232
rect 7072 5168 7088 5232
rect 7152 5168 7168 5232
rect 7232 5168 7248 5232
rect 7312 5168 7328 5232
rect 7392 5168 7408 5232
rect 7472 5168 7488 5232
rect 7552 5168 7568 5232
rect 7632 5168 7648 5232
rect 7712 5168 7728 5232
rect 7792 5168 7808 5232
rect 7872 5168 7888 5232
rect 7952 5168 7968 5232
rect 8032 5168 8048 5232
rect 8112 5168 8128 5232
rect 8192 5168 8208 5232
rect 8272 5168 8288 5232
rect 8352 5168 8368 5232
rect 8432 5168 8448 5232
rect 8512 5168 8528 5232
rect 8592 5168 8608 5232
rect 8672 5168 8688 5232
rect 8752 5168 8768 5232
rect 8832 5168 8848 5232
rect 8912 5168 8928 5232
rect 8992 5168 14112 5232
rect 14176 5168 14192 5232
rect 14256 5168 14272 5232
rect 14336 5168 14352 5232
rect 14416 5168 24112 5232
rect 24176 5168 24192 5232
rect 24256 5168 24272 5232
rect 24336 5168 24352 5232
rect 24416 5168 36376 5232
rect 36440 5168 36456 5232
rect 36520 5168 36536 5232
rect 36600 5168 36616 5232
rect 36680 5168 36696 5232
rect 36760 5168 36776 5232
rect 36840 5168 36856 5232
rect 36920 5168 36936 5232
rect 37000 5168 37016 5232
rect 37080 5168 37096 5232
rect 37160 5168 37176 5232
rect 37240 5168 37256 5232
rect 37320 5168 37336 5232
rect 37400 5168 37416 5232
rect 37480 5168 37496 5232
rect 37560 5168 37576 5232
rect 37640 5168 37656 5232
rect 37720 5168 37736 5232
rect 37800 5168 37816 5232
rect 37880 5168 37896 5232
rect 37960 5168 37976 5232
rect 38040 5168 38056 5232
rect 38120 5168 38136 5232
rect 38200 5168 38216 5232
rect 38280 5168 38296 5232
rect 38360 5168 38376 5232
rect 38440 5168 38456 5232
rect 38520 5168 38536 5232
rect 38600 5168 38616 5232
rect 38680 5168 38696 5232
rect 38760 5168 38776 5232
rect 38840 5168 38856 5232
rect 38920 5168 38936 5232
rect 39000 5168 39016 5232
rect 39080 5168 39096 5232
rect 39160 5168 39176 5232
rect 39240 5168 39256 5232
rect 39320 5168 39336 5232
rect 39400 5168 39416 5232
rect 39480 5168 39496 5232
rect 39560 5168 39576 5232
rect 39640 5168 39656 5232
rect 39720 5168 39736 5232
rect 39800 5168 39816 5232
rect 39880 5168 39896 5232
rect 39960 5168 39976 5232
rect 40040 5168 40056 5232
rect 40120 5168 40136 5232
rect 40200 5168 40216 5232
rect 40280 5168 40296 5232
rect 40360 5168 40368 5232
rect 5000 5152 40368 5168
rect 5000 5088 5008 5152
rect 5072 5088 5088 5152
rect 5152 5088 5168 5152
rect 5232 5088 5248 5152
rect 5312 5088 5328 5152
rect 5392 5088 5408 5152
rect 5472 5088 5488 5152
rect 5552 5088 5568 5152
rect 5632 5088 5648 5152
rect 5712 5088 5728 5152
rect 5792 5088 5808 5152
rect 5872 5088 5888 5152
rect 5952 5088 5968 5152
rect 6032 5088 6048 5152
rect 6112 5088 6128 5152
rect 6192 5088 6208 5152
rect 6272 5088 6288 5152
rect 6352 5088 6368 5152
rect 6432 5088 6448 5152
rect 6512 5088 6528 5152
rect 6592 5088 6608 5152
rect 6672 5088 6688 5152
rect 6752 5088 6768 5152
rect 6832 5088 6848 5152
rect 6912 5088 6928 5152
rect 6992 5088 7008 5152
rect 7072 5088 7088 5152
rect 7152 5088 7168 5152
rect 7232 5088 7248 5152
rect 7312 5088 7328 5152
rect 7392 5088 7408 5152
rect 7472 5088 7488 5152
rect 7552 5088 7568 5152
rect 7632 5088 7648 5152
rect 7712 5088 7728 5152
rect 7792 5088 7808 5152
rect 7872 5088 7888 5152
rect 7952 5088 7968 5152
rect 8032 5088 8048 5152
rect 8112 5088 8128 5152
rect 8192 5088 8208 5152
rect 8272 5088 8288 5152
rect 8352 5088 8368 5152
rect 8432 5088 8448 5152
rect 8512 5088 8528 5152
rect 8592 5088 8608 5152
rect 8672 5088 8688 5152
rect 8752 5088 8768 5152
rect 8832 5088 8848 5152
rect 8912 5088 8928 5152
rect 8992 5088 14112 5152
rect 14176 5088 14192 5152
rect 14256 5088 14272 5152
rect 14336 5088 14352 5152
rect 14416 5088 24112 5152
rect 24176 5088 24192 5152
rect 24256 5088 24272 5152
rect 24336 5088 24352 5152
rect 24416 5088 36376 5152
rect 36440 5088 36456 5152
rect 36520 5088 36536 5152
rect 36600 5088 36616 5152
rect 36680 5088 36696 5152
rect 36760 5088 36776 5152
rect 36840 5088 36856 5152
rect 36920 5088 36936 5152
rect 37000 5088 37016 5152
rect 37080 5088 37096 5152
rect 37160 5088 37176 5152
rect 37240 5088 37256 5152
rect 37320 5088 37336 5152
rect 37400 5088 37416 5152
rect 37480 5088 37496 5152
rect 37560 5088 37576 5152
rect 37640 5088 37656 5152
rect 37720 5088 37736 5152
rect 37800 5088 37816 5152
rect 37880 5088 37896 5152
rect 37960 5088 37976 5152
rect 38040 5088 38056 5152
rect 38120 5088 38136 5152
rect 38200 5088 38216 5152
rect 38280 5088 38296 5152
rect 38360 5088 38376 5152
rect 38440 5088 38456 5152
rect 38520 5088 38536 5152
rect 38600 5088 38616 5152
rect 38680 5088 38696 5152
rect 38760 5088 38776 5152
rect 38840 5088 38856 5152
rect 38920 5088 38936 5152
rect 39000 5088 39016 5152
rect 39080 5088 39096 5152
rect 39160 5088 39176 5152
rect 39240 5088 39256 5152
rect 39320 5088 39336 5152
rect 39400 5088 39416 5152
rect 39480 5088 39496 5152
rect 39560 5088 39576 5152
rect 39640 5088 39656 5152
rect 39720 5088 39736 5152
rect 39800 5088 39816 5152
rect 39880 5088 39896 5152
rect 39960 5088 39976 5152
rect 40040 5088 40056 5152
rect 40120 5088 40136 5152
rect 40200 5088 40216 5152
rect 40280 5088 40296 5152
rect 40360 5088 40368 5152
rect 5000 5072 40368 5088
rect 5000 5008 5008 5072
rect 5072 5008 5088 5072
rect 5152 5008 5168 5072
rect 5232 5008 5248 5072
rect 5312 5008 5328 5072
rect 5392 5008 5408 5072
rect 5472 5008 5488 5072
rect 5552 5008 5568 5072
rect 5632 5008 5648 5072
rect 5712 5008 5728 5072
rect 5792 5008 5808 5072
rect 5872 5008 5888 5072
rect 5952 5008 5968 5072
rect 6032 5008 6048 5072
rect 6112 5008 6128 5072
rect 6192 5008 6208 5072
rect 6272 5008 6288 5072
rect 6352 5008 6368 5072
rect 6432 5008 6448 5072
rect 6512 5008 6528 5072
rect 6592 5008 6608 5072
rect 6672 5008 6688 5072
rect 6752 5008 6768 5072
rect 6832 5008 6848 5072
rect 6912 5008 6928 5072
rect 6992 5008 7008 5072
rect 7072 5008 7088 5072
rect 7152 5008 7168 5072
rect 7232 5008 7248 5072
rect 7312 5008 7328 5072
rect 7392 5008 7408 5072
rect 7472 5008 7488 5072
rect 7552 5008 7568 5072
rect 7632 5008 7648 5072
rect 7712 5008 7728 5072
rect 7792 5008 7808 5072
rect 7872 5008 7888 5072
rect 7952 5008 7968 5072
rect 8032 5008 8048 5072
rect 8112 5008 8128 5072
rect 8192 5008 8208 5072
rect 8272 5008 8288 5072
rect 8352 5008 8368 5072
rect 8432 5008 8448 5072
rect 8512 5008 8528 5072
rect 8592 5008 8608 5072
rect 8672 5008 8688 5072
rect 8752 5008 8768 5072
rect 8832 5008 8848 5072
rect 8912 5008 8928 5072
rect 8992 5008 14112 5072
rect 14176 5008 14192 5072
rect 14256 5008 14272 5072
rect 14336 5008 14352 5072
rect 14416 5008 24112 5072
rect 24176 5008 24192 5072
rect 24256 5008 24272 5072
rect 24336 5008 24352 5072
rect 24416 5008 36376 5072
rect 36440 5008 36456 5072
rect 36520 5008 36536 5072
rect 36600 5008 36616 5072
rect 36680 5008 36696 5072
rect 36760 5008 36776 5072
rect 36840 5008 36856 5072
rect 36920 5008 36936 5072
rect 37000 5008 37016 5072
rect 37080 5008 37096 5072
rect 37160 5008 37176 5072
rect 37240 5008 37256 5072
rect 37320 5008 37336 5072
rect 37400 5008 37416 5072
rect 37480 5008 37496 5072
rect 37560 5008 37576 5072
rect 37640 5008 37656 5072
rect 37720 5008 37736 5072
rect 37800 5008 37816 5072
rect 37880 5008 37896 5072
rect 37960 5008 37976 5072
rect 38040 5008 38056 5072
rect 38120 5008 38136 5072
rect 38200 5008 38216 5072
rect 38280 5008 38296 5072
rect 38360 5008 38376 5072
rect 38440 5008 38456 5072
rect 38520 5008 38536 5072
rect 38600 5008 38616 5072
rect 38680 5008 38696 5072
rect 38760 5008 38776 5072
rect 38840 5008 38856 5072
rect 38920 5008 38936 5072
rect 39000 5008 39016 5072
rect 39080 5008 39096 5072
rect 39160 5008 39176 5072
rect 39240 5008 39256 5072
rect 39320 5008 39336 5072
rect 39400 5008 39416 5072
rect 39480 5008 39496 5072
rect 39560 5008 39576 5072
rect 39640 5008 39656 5072
rect 39720 5008 39736 5072
rect 39800 5008 39816 5072
rect 39880 5008 39896 5072
rect 39960 5008 39976 5072
rect 40040 5008 40056 5072
rect 40120 5008 40136 5072
rect 40200 5008 40216 5072
rect 40280 5008 40296 5072
rect 40360 5008 40368 5072
rect 5000 5000 40368 5008
rect 0 3992 45368 4000
rect 0 3928 8 3992
rect 72 3928 88 3992
rect 152 3928 168 3992
rect 232 3928 248 3992
rect 312 3928 328 3992
rect 392 3928 408 3992
rect 472 3928 488 3992
rect 552 3928 568 3992
rect 632 3928 648 3992
rect 712 3928 728 3992
rect 792 3928 808 3992
rect 872 3928 888 3992
rect 952 3928 968 3992
rect 1032 3928 1048 3992
rect 1112 3928 1128 3992
rect 1192 3928 1208 3992
rect 1272 3928 1288 3992
rect 1352 3928 1368 3992
rect 1432 3928 1448 3992
rect 1512 3928 1528 3992
rect 1592 3928 1608 3992
rect 1672 3928 1688 3992
rect 1752 3928 1768 3992
rect 1832 3928 1848 3992
rect 1912 3928 1928 3992
rect 1992 3928 2008 3992
rect 2072 3928 2088 3992
rect 2152 3928 2168 3992
rect 2232 3928 2248 3992
rect 2312 3928 2328 3992
rect 2392 3928 2408 3992
rect 2472 3928 2488 3992
rect 2552 3928 2568 3992
rect 2632 3928 2648 3992
rect 2712 3928 2728 3992
rect 2792 3928 2808 3992
rect 2872 3928 2888 3992
rect 2952 3928 2968 3992
rect 3032 3928 3048 3992
rect 3112 3928 3128 3992
rect 3192 3928 3208 3992
rect 3272 3928 3288 3992
rect 3352 3928 3368 3992
rect 3432 3928 3448 3992
rect 3512 3928 3528 3992
rect 3592 3928 3608 3992
rect 3672 3928 3688 3992
rect 3752 3928 3768 3992
rect 3832 3928 3848 3992
rect 3912 3928 3928 3992
rect 3992 3928 19112 3992
rect 19176 3928 19192 3992
rect 19256 3928 19272 3992
rect 19336 3928 19352 3992
rect 19416 3928 29112 3992
rect 29176 3928 29192 3992
rect 29256 3928 29272 3992
rect 29336 3928 29352 3992
rect 29416 3928 41376 3992
rect 41440 3928 41456 3992
rect 41520 3928 41536 3992
rect 41600 3928 41616 3992
rect 41680 3928 41696 3992
rect 41760 3928 41776 3992
rect 41840 3928 41856 3992
rect 41920 3928 41936 3992
rect 42000 3928 42016 3992
rect 42080 3928 42096 3992
rect 42160 3928 42176 3992
rect 42240 3928 42256 3992
rect 42320 3928 42336 3992
rect 42400 3928 42416 3992
rect 42480 3928 42496 3992
rect 42560 3928 42576 3992
rect 42640 3928 42656 3992
rect 42720 3928 42736 3992
rect 42800 3928 42816 3992
rect 42880 3928 42896 3992
rect 42960 3928 42976 3992
rect 43040 3928 43056 3992
rect 43120 3928 43136 3992
rect 43200 3928 43216 3992
rect 43280 3928 43296 3992
rect 43360 3928 43376 3992
rect 43440 3928 43456 3992
rect 43520 3928 43536 3992
rect 43600 3928 43616 3992
rect 43680 3928 43696 3992
rect 43760 3928 43776 3992
rect 43840 3928 43856 3992
rect 43920 3928 43936 3992
rect 44000 3928 44016 3992
rect 44080 3928 44096 3992
rect 44160 3928 44176 3992
rect 44240 3928 44256 3992
rect 44320 3928 44336 3992
rect 44400 3928 44416 3992
rect 44480 3928 44496 3992
rect 44560 3928 44576 3992
rect 44640 3928 44656 3992
rect 44720 3928 44736 3992
rect 44800 3928 44816 3992
rect 44880 3928 44896 3992
rect 44960 3928 44976 3992
rect 45040 3928 45056 3992
rect 45120 3928 45136 3992
rect 45200 3928 45216 3992
rect 45280 3928 45296 3992
rect 45360 3928 45368 3992
rect 0 3912 45368 3928
rect 0 3848 8 3912
rect 72 3848 88 3912
rect 152 3848 168 3912
rect 232 3848 248 3912
rect 312 3848 328 3912
rect 392 3848 408 3912
rect 472 3848 488 3912
rect 552 3848 568 3912
rect 632 3848 648 3912
rect 712 3848 728 3912
rect 792 3848 808 3912
rect 872 3848 888 3912
rect 952 3848 968 3912
rect 1032 3848 1048 3912
rect 1112 3848 1128 3912
rect 1192 3848 1208 3912
rect 1272 3848 1288 3912
rect 1352 3848 1368 3912
rect 1432 3848 1448 3912
rect 1512 3848 1528 3912
rect 1592 3848 1608 3912
rect 1672 3848 1688 3912
rect 1752 3848 1768 3912
rect 1832 3848 1848 3912
rect 1912 3848 1928 3912
rect 1992 3848 2008 3912
rect 2072 3848 2088 3912
rect 2152 3848 2168 3912
rect 2232 3848 2248 3912
rect 2312 3848 2328 3912
rect 2392 3848 2408 3912
rect 2472 3848 2488 3912
rect 2552 3848 2568 3912
rect 2632 3848 2648 3912
rect 2712 3848 2728 3912
rect 2792 3848 2808 3912
rect 2872 3848 2888 3912
rect 2952 3848 2968 3912
rect 3032 3848 3048 3912
rect 3112 3848 3128 3912
rect 3192 3848 3208 3912
rect 3272 3848 3288 3912
rect 3352 3848 3368 3912
rect 3432 3848 3448 3912
rect 3512 3848 3528 3912
rect 3592 3848 3608 3912
rect 3672 3848 3688 3912
rect 3752 3848 3768 3912
rect 3832 3848 3848 3912
rect 3912 3848 3928 3912
rect 3992 3848 19112 3912
rect 19176 3848 19192 3912
rect 19256 3848 19272 3912
rect 19336 3848 19352 3912
rect 19416 3848 29112 3912
rect 29176 3848 29192 3912
rect 29256 3848 29272 3912
rect 29336 3848 29352 3912
rect 29416 3848 41376 3912
rect 41440 3848 41456 3912
rect 41520 3848 41536 3912
rect 41600 3848 41616 3912
rect 41680 3848 41696 3912
rect 41760 3848 41776 3912
rect 41840 3848 41856 3912
rect 41920 3848 41936 3912
rect 42000 3848 42016 3912
rect 42080 3848 42096 3912
rect 42160 3848 42176 3912
rect 42240 3848 42256 3912
rect 42320 3848 42336 3912
rect 42400 3848 42416 3912
rect 42480 3848 42496 3912
rect 42560 3848 42576 3912
rect 42640 3848 42656 3912
rect 42720 3848 42736 3912
rect 42800 3848 42816 3912
rect 42880 3848 42896 3912
rect 42960 3848 42976 3912
rect 43040 3848 43056 3912
rect 43120 3848 43136 3912
rect 43200 3848 43216 3912
rect 43280 3848 43296 3912
rect 43360 3848 43376 3912
rect 43440 3848 43456 3912
rect 43520 3848 43536 3912
rect 43600 3848 43616 3912
rect 43680 3848 43696 3912
rect 43760 3848 43776 3912
rect 43840 3848 43856 3912
rect 43920 3848 43936 3912
rect 44000 3848 44016 3912
rect 44080 3848 44096 3912
rect 44160 3848 44176 3912
rect 44240 3848 44256 3912
rect 44320 3848 44336 3912
rect 44400 3848 44416 3912
rect 44480 3848 44496 3912
rect 44560 3848 44576 3912
rect 44640 3848 44656 3912
rect 44720 3848 44736 3912
rect 44800 3848 44816 3912
rect 44880 3848 44896 3912
rect 44960 3848 44976 3912
rect 45040 3848 45056 3912
rect 45120 3848 45136 3912
rect 45200 3848 45216 3912
rect 45280 3848 45296 3912
rect 45360 3848 45368 3912
rect 0 3832 45368 3848
rect 0 3768 8 3832
rect 72 3768 88 3832
rect 152 3768 168 3832
rect 232 3768 248 3832
rect 312 3768 328 3832
rect 392 3768 408 3832
rect 472 3768 488 3832
rect 552 3768 568 3832
rect 632 3768 648 3832
rect 712 3768 728 3832
rect 792 3768 808 3832
rect 872 3768 888 3832
rect 952 3768 968 3832
rect 1032 3768 1048 3832
rect 1112 3768 1128 3832
rect 1192 3768 1208 3832
rect 1272 3768 1288 3832
rect 1352 3768 1368 3832
rect 1432 3768 1448 3832
rect 1512 3768 1528 3832
rect 1592 3768 1608 3832
rect 1672 3768 1688 3832
rect 1752 3768 1768 3832
rect 1832 3768 1848 3832
rect 1912 3768 1928 3832
rect 1992 3768 2008 3832
rect 2072 3768 2088 3832
rect 2152 3768 2168 3832
rect 2232 3768 2248 3832
rect 2312 3768 2328 3832
rect 2392 3768 2408 3832
rect 2472 3768 2488 3832
rect 2552 3768 2568 3832
rect 2632 3768 2648 3832
rect 2712 3768 2728 3832
rect 2792 3768 2808 3832
rect 2872 3768 2888 3832
rect 2952 3768 2968 3832
rect 3032 3768 3048 3832
rect 3112 3768 3128 3832
rect 3192 3768 3208 3832
rect 3272 3768 3288 3832
rect 3352 3768 3368 3832
rect 3432 3768 3448 3832
rect 3512 3768 3528 3832
rect 3592 3768 3608 3832
rect 3672 3768 3688 3832
rect 3752 3768 3768 3832
rect 3832 3768 3848 3832
rect 3912 3768 3928 3832
rect 3992 3768 19112 3832
rect 19176 3768 19192 3832
rect 19256 3768 19272 3832
rect 19336 3768 19352 3832
rect 19416 3768 29112 3832
rect 29176 3768 29192 3832
rect 29256 3768 29272 3832
rect 29336 3768 29352 3832
rect 29416 3768 41376 3832
rect 41440 3768 41456 3832
rect 41520 3768 41536 3832
rect 41600 3768 41616 3832
rect 41680 3768 41696 3832
rect 41760 3768 41776 3832
rect 41840 3768 41856 3832
rect 41920 3768 41936 3832
rect 42000 3768 42016 3832
rect 42080 3768 42096 3832
rect 42160 3768 42176 3832
rect 42240 3768 42256 3832
rect 42320 3768 42336 3832
rect 42400 3768 42416 3832
rect 42480 3768 42496 3832
rect 42560 3768 42576 3832
rect 42640 3768 42656 3832
rect 42720 3768 42736 3832
rect 42800 3768 42816 3832
rect 42880 3768 42896 3832
rect 42960 3768 42976 3832
rect 43040 3768 43056 3832
rect 43120 3768 43136 3832
rect 43200 3768 43216 3832
rect 43280 3768 43296 3832
rect 43360 3768 43376 3832
rect 43440 3768 43456 3832
rect 43520 3768 43536 3832
rect 43600 3768 43616 3832
rect 43680 3768 43696 3832
rect 43760 3768 43776 3832
rect 43840 3768 43856 3832
rect 43920 3768 43936 3832
rect 44000 3768 44016 3832
rect 44080 3768 44096 3832
rect 44160 3768 44176 3832
rect 44240 3768 44256 3832
rect 44320 3768 44336 3832
rect 44400 3768 44416 3832
rect 44480 3768 44496 3832
rect 44560 3768 44576 3832
rect 44640 3768 44656 3832
rect 44720 3768 44736 3832
rect 44800 3768 44816 3832
rect 44880 3768 44896 3832
rect 44960 3768 44976 3832
rect 45040 3768 45056 3832
rect 45120 3768 45136 3832
rect 45200 3768 45216 3832
rect 45280 3768 45296 3832
rect 45360 3768 45368 3832
rect 0 3752 45368 3768
rect 0 3688 8 3752
rect 72 3688 88 3752
rect 152 3688 168 3752
rect 232 3688 248 3752
rect 312 3688 328 3752
rect 392 3688 408 3752
rect 472 3688 488 3752
rect 552 3688 568 3752
rect 632 3688 648 3752
rect 712 3688 728 3752
rect 792 3688 808 3752
rect 872 3688 888 3752
rect 952 3688 968 3752
rect 1032 3688 1048 3752
rect 1112 3688 1128 3752
rect 1192 3688 1208 3752
rect 1272 3688 1288 3752
rect 1352 3688 1368 3752
rect 1432 3688 1448 3752
rect 1512 3688 1528 3752
rect 1592 3688 1608 3752
rect 1672 3688 1688 3752
rect 1752 3688 1768 3752
rect 1832 3688 1848 3752
rect 1912 3688 1928 3752
rect 1992 3688 2008 3752
rect 2072 3688 2088 3752
rect 2152 3688 2168 3752
rect 2232 3688 2248 3752
rect 2312 3688 2328 3752
rect 2392 3688 2408 3752
rect 2472 3688 2488 3752
rect 2552 3688 2568 3752
rect 2632 3688 2648 3752
rect 2712 3688 2728 3752
rect 2792 3688 2808 3752
rect 2872 3688 2888 3752
rect 2952 3688 2968 3752
rect 3032 3688 3048 3752
rect 3112 3688 3128 3752
rect 3192 3688 3208 3752
rect 3272 3688 3288 3752
rect 3352 3688 3368 3752
rect 3432 3688 3448 3752
rect 3512 3688 3528 3752
rect 3592 3688 3608 3752
rect 3672 3688 3688 3752
rect 3752 3688 3768 3752
rect 3832 3688 3848 3752
rect 3912 3688 3928 3752
rect 3992 3688 19112 3752
rect 19176 3688 19192 3752
rect 19256 3688 19272 3752
rect 19336 3688 19352 3752
rect 19416 3688 29112 3752
rect 29176 3688 29192 3752
rect 29256 3688 29272 3752
rect 29336 3688 29352 3752
rect 29416 3688 41376 3752
rect 41440 3688 41456 3752
rect 41520 3688 41536 3752
rect 41600 3688 41616 3752
rect 41680 3688 41696 3752
rect 41760 3688 41776 3752
rect 41840 3688 41856 3752
rect 41920 3688 41936 3752
rect 42000 3688 42016 3752
rect 42080 3688 42096 3752
rect 42160 3688 42176 3752
rect 42240 3688 42256 3752
rect 42320 3688 42336 3752
rect 42400 3688 42416 3752
rect 42480 3688 42496 3752
rect 42560 3688 42576 3752
rect 42640 3688 42656 3752
rect 42720 3688 42736 3752
rect 42800 3688 42816 3752
rect 42880 3688 42896 3752
rect 42960 3688 42976 3752
rect 43040 3688 43056 3752
rect 43120 3688 43136 3752
rect 43200 3688 43216 3752
rect 43280 3688 43296 3752
rect 43360 3688 43376 3752
rect 43440 3688 43456 3752
rect 43520 3688 43536 3752
rect 43600 3688 43616 3752
rect 43680 3688 43696 3752
rect 43760 3688 43776 3752
rect 43840 3688 43856 3752
rect 43920 3688 43936 3752
rect 44000 3688 44016 3752
rect 44080 3688 44096 3752
rect 44160 3688 44176 3752
rect 44240 3688 44256 3752
rect 44320 3688 44336 3752
rect 44400 3688 44416 3752
rect 44480 3688 44496 3752
rect 44560 3688 44576 3752
rect 44640 3688 44656 3752
rect 44720 3688 44736 3752
rect 44800 3688 44816 3752
rect 44880 3688 44896 3752
rect 44960 3688 44976 3752
rect 45040 3688 45056 3752
rect 45120 3688 45136 3752
rect 45200 3688 45216 3752
rect 45280 3688 45296 3752
rect 45360 3688 45368 3752
rect 0 3672 45368 3688
rect 0 3608 8 3672
rect 72 3608 88 3672
rect 152 3608 168 3672
rect 232 3608 248 3672
rect 312 3608 328 3672
rect 392 3608 408 3672
rect 472 3608 488 3672
rect 552 3608 568 3672
rect 632 3608 648 3672
rect 712 3608 728 3672
rect 792 3608 808 3672
rect 872 3608 888 3672
rect 952 3608 968 3672
rect 1032 3608 1048 3672
rect 1112 3608 1128 3672
rect 1192 3608 1208 3672
rect 1272 3608 1288 3672
rect 1352 3608 1368 3672
rect 1432 3608 1448 3672
rect 1512 3608 1528 3672
rect 1592 3608 1608 3672
rect 1672 3608 1688 3672
rect 1752 3608 1768 3672
rect 1832 3608 1848 3672
rect 1912 3608 1928 3672
rect 1992 3608 2008 3672
rect 2072 3608 2088 3672
rect 2152 3608 2168 3672
rect 2232 3608 2248 3672
rect 2312 3608 2328 3672
rect 2392 3608 2408 3672
rect 2472 3608 2488 3672
rect 2552 3608 2568 3672
rect 2632 3608 2648 3672
rect 2712 3608 2728 3672
rect 2792 3608 2808 3672
rect 2872 3608 2888 3672
rect 2952 3608 2968 3672
rect 3032 3608 3048 3672
rect 3112 3608 3128 3672
rect 3192 3608 3208 3672
rect 3272 3608 3288 3672
rect 3352 3608 3368 3672
rect 3432 3608 3448 3672
rect 3512 3608 3528 3672
rect 3592 3608 3608 3672
rect 3672 3608 3688 3672
rect 3752 3608 3768 3672
rect 3832 3608 3848 3672
rect 3912 3608 3928 3672
rect 3992 3608 19112 3672
rect 19176 3608 19192 3672
rect 19256 3608 19272 3672
rect 19336 3608 19352 3672
rect 19416 3608 29112 3672
rect 29176 3608 29192 3672
rect 29256 3608 29272 3672
rect 29336 3608 29352 3672
rect 29416 3608 41376 3672
rect 41440 3608 41456 3672
rect 41520 3608 41536 3672
rect 41600 3608 41616 3672
rect 41680 3608 41696 3672
rect 41760 3608 41776 3672
rect 41840 3608 41856 3672
rect 41920 3608 41936 3672
rect 42000 3608 42016 3672
rect 42080 3608 42096 3672
rect 42160 3608 42176 3672
rect 42240 3608 42256 3672
rect 42320 3608 42336 3672
rect 42400 3608 42416 3672
rect 42480 3608 42496 3672
rect 42560 3608 42576 3672
rect 42640 3608 42656 3672
rect 42720 3608 42736 3672
rect 42800 3608 42816 3672
rect 42880 3608 42896 3672
rect 42960 3608 42976 3672
rect 43040 3608 43056 3672
rect 43120 3608 43136 3672
rect 43200 3608 43216 3672
rect 43280 3608 43296 3672
rect 43360 3608 43376 3672
rect 43440 3608 43456 3672
rect 43520 3608 43536 3672
rect 43600 3608 43616 3672
rect 43680 3608 43696 3672
rect 43760 3608 43776 3672
rect 43840 3608 43856 3672
rect 43920 3608 43936 3672
rect 44000 3608 44016 3672
rect 44080 3608 44096 3672
rect 44160 3608 44176 3672
rect 44240 3608 44256 3672
rect 44320 3608 44336 3672
rect 44400 3608 44416 3672
rect 44480 3608 44496 3672
rect 44560 3608 44576 3672
rect 44640 3608 44656 3672
rect 44720 3608 44736 3672
rect 44800 3608 44816 3672
rect 44880 3608 44896 3672
rect 44960 3608 44976 3672
rect 45040 3608 45056 3672
rect 45120 3608 45136 3672
rect 45200 3608 45216 3672
rect 45280 3608 45296 3672
rect 45360 3608 45368 3672
rect 0 3592 45368 3608
rect 0 3528 8 3592
rect 72 3528 88 3592
rect 152 3528 168 3592
rect 232 3528 248 3592
rect 312 3528 328 3592
rect 392 3528 408 3592
rect 472 3528 488 3592
rect 552 3528 568 3592
rect 632 3528 648 3592
rect 712 3528 728 3592
rect 792 3528 808 3592
rect 872 3528 888 3592
rect 952 3528 968 3592
rect 1032 3528 1048 3592
rect 1112 3528 1128 3592
rect 1192 3528 1208 3592
rect 1272 3528 1288 3592
rect 1352 3528 1368 3592
rect 1432 3528 1448 3592
rect 1512 3528 1528 3592
rect 1592 3528 1608 3592
rect 1672 3528 1688 3592
rect 1752 3528 1768 3592
rect 1832 3528 1848 3592
rect 1912 3528 1928 3592
rect 1992 3528 2008 3592
rect 2072 3528 2088 3592
rect 2152 3528 2168 3592
rect 2232 3528 2248 3592
rect 2312 3528 2328 3592
rect 2392 3528 2408 3592
rect 2472 3528 2488 3592
rect 2552 3528 2568 3592
rect 2632 3528 2648 3592
rect 2712 3528 2728 3592
rect 2792 3528 2808 3592
rect 2872 3528 2888 3592
rect 2952 3528 2968 3592
rect 3032 3528 3048 3592
rect 3112 3528 3128 3592
rect 3192 3528 3208 3592
rect 3272 3528 3288 3592
rect 3352 3528 3368 3592
rect 3432 3528 3448 3592
rect 3512 3528 3528 3592
rect 3592 3528 3608 3592
rect 3672 3528 3688 3592
rect 3752 3528 3768 3592
rect 3832 3528 3848 3592
rect 3912 3528 3928 3592
rect 3992 3528 19112 3592
rect 19176 3528 19192 3592
rect 19256 3528 19272 3592
rect 19336 3528 19352 3592
rect 19416 3528 29112 3592
rect 29176 3528 29192 3592
rect 29256 3528 29272 3592
rect 29336 3528 29352 3592
rect 29416 3528 41376 3592
rect 41440 3528 41456 3592
rect 41520 3528 41536 3592
rect 41600 3528 41616 3592
rect 41680 3528 41696 3592
rect 41760 3528 41776 3592
rect 41840 3528 41856 3592
rect 41920 3528 41936 3592
rect 42000 3528 42016 3592
rect 42080 3528 42096 3592
rect 42160 3528 42176 3592
rect 42240 3528 42256 3592
rect 42320 3528 42336 3592
rect 42400 3528 42416 3592
rect 42480 3528 42496 3592
rect 42560 3528 42576 3592
rect 42640 3528 42656 3592
rect 42720 3528 42736 3592
rect 42800 3528 42816 3592
rect 42880 3528 42896 3592
rect 42960 3528 42976 3592
rect 43040 3528 43056 3592
rect 43120 3528 43136 3592
rect 43200 3528 43216 3592
rect 43280 3528 43296 3592
rect 43360 3528 43376 3592
rect 43440 3528 43456 3592
rect 43520 3528 43536 3592
rect 43600 3528 43616 3592
rect 43680 3528 43696 3592
rect 43760 3528 43776 3592
rect 43840 3528 43856 3592
rect 43920 3528 43936 3592
rect 44000 3528 44016 3592
rect 44080 3528 44096 3592
rect 44160 3528 44176 3592
rect 44240 3528 44256 3592
rect 44320 3528 44336 3592
rect 44400 3528 44416 3592
rect 44480 3528 44496 3592
rect 44560 3528 44576 3592
rect 44640 3528 44656 3592
rect 44720 3528 44736 3592
rect 44800 3528 44816 3592
rect 44880 3528 44896 3592
rect 44960 3528 44976 3592
rect 45040 3528 45056 3592
rect 45120 3528 45136 3592
rect 45200 3528 45216 3592
rect 45280 3528 45296 3592
rect 45360 3528 45368 3592
rect 0 3512 45368 3528
rect 0 3448 8 3512
rect 72 3448 88 3512
rect 152 3448 168 3512
rect 232 3448 248 3512
rect 312 3448 328 3512
rect 392 3448 408 3512
rect 472 3448 488 3512
rect 552 3448 568 3512
rect 632 3448 648 3512
rect 712 3448 728 3512
rect 792 3448 808 3512
rect 872 3448 888 3512
rect 952 3448 968 3512
rect 1032 3448 1048 3512
rect 1112 3448 1128 3512
rect 1192 3448 1208 3512
rect 1272 3448 1288 3512
rect 1352 3448 1368 3512
rect 1432 3448 1448 3512
rect 1512 3448 1528 3512
rect 1592 3448 1608 3512
rect 1672 3448 1688 3512
rect 1752 3448 1768 3512
rect 1832 3448 1848 3512
rect 1912 3448 1928 3512
rect 1992 3448 2008 3512
rect 2072 3448 2088 3512
rect 2152 3448 2168 3512
rect 2232 3448 2248 3512
rect 2312 3448 2328 3512
rect 2392 3448 2408 3512
rect 2472 3448 2488 3512
rect 2552 3448 2568 3512
rect 2632 3448 2648 3512
rect 2712 3448 2728 3512
rect 2792 3448 2808 3512
rect 2872 3448 2888 3512
rect 2952 3448 2968 3512
rect 3032 3448 3048 3512
rect 3112 3448 3128 3512
rect 3192 3448 3208 3512
rect 3272 3448 3288 3512
rect 3352 3448 3368 3512
rect 3432 3448 3448 3512
rect 3512 3448 3528 3512
rect 3592 3448 3608 3512
rect 3672 3448 3688 3512
rect 3752 3448 3768 3512
rect 3832 3448 3848 3512
rect 3912 3448 3928 3512
rect 3992 3448 19112 3512
rect 19176 3448 19192 3512
rect 19256 3448 19272 3512
rect 19336 3448 19352 3512
rect 19416 3448 29112 3512
rect 29176 3448 29192 3512
rect 29256 3448 29272 3512
rect 29336 3448 29352 3512
rect 29416 3448 41376 3512
rect 41440 3448 41456 3512
rect 41520 3448 41536 3512
rect 41600 3448 41616 3512
rect 41680 3448 41696 3512
rect 41760 3448 41776 3512
rect 41840 3448 41856 3512
rect 41920 3448 41936 3512
rect 42000 3448 42016 3512
rect 42080 3448 42096 3512
rect 42160 3448 42176 3512
rect 42240 3448 42256 3512
rect 42320 3448 42336 3512
rect 42400 3448 42416 3512
rect 42480 3448 42496 3512
rect 42560 3448 42576 3512
rect 42640 3448 42656 3512
rect 42720 3448 42736 3512
rect 42800 3448 42816 3512
rect 42880 3448 42896 3512
rect 42960 3448 42976 3512
rect 43040 3448 43056 3512
rect 43120 3448 43136 3512
rect 43200 3448 43216 3512
rect 43280 3448 43296 3512
rect 43360 3448 43376 3512
rect 43440 3448 43456 3512
rect 43520 3448 43536 3512
rect 43600 3448 43616 3512
rect 43680 3448 43696 3512
rect 43760 3448 43776 3512
rect 43840 3448 43856 3512
rect 43920 3448 43936 3512
rect 44000 3448 44016 3512
rect 44080 3448 44096 3512
rect 44160 3448 44176 3512
rect 44240 3448 44256 3512
rect 44320 3448 44336 3512
rect 44400 3448 44416 3512
rect 44480 3448 44496 3512
rect 44560 3448 44576 3512
rect 44640 3448 44656 3512
rect 44720 3448 44736 3512
rect 44800 3448 44816 3512
rect 44880 3448 44896 3512
rect 44960 3448 44976 3512
rect 45040 3448 45056 3512
rect 45120 3448 45136 3512
rect 45200 3448 45216 3512
rect 45280 3448 45296 3512
rect 45360 3448 45368 3512
rect 0 3432 45368 3448
rect 0 3368 8 3432
rect 72 3368 88 3432
rect 152 3368 168 3432
rect 232 3368 248 3432
rect 312 3368 328 3432
rect 392 3368 408 3432
rect 472 3368 488 3432
rect 552 3368 568 3432
rect 632 3368 648 3432
rect 712 3368 728 3432
rect 792 3368 808 3432
rect 872 3368 888 3432
rect 952 3368 968 3432
rect 1032 3368 1048 3432
rect 1112 3368 1128 3432
rect 1192 3368 1208 3432
rect 1272 3368 1288 3432
rect 1352 3368 1368 3432
rect 1432 3368 1448 3432
rect 1512 3368 1528 3432
rect 1592 3368 1608 3432
rect 1672 3368 1688 3432
rect 1752 3368 1768 3432
rect 1832 3368 1848 3432
rect 1912 3368 1928 3432
rect 1992 3368 2008 3432
rect 2072 3368 2088 3432
rect 2152 3368 2168 3432
rect 2232 3368 2248 3432
rect 2312 3368 2328 3432
rect 2392 3368 2408 3432
rect 2472 3368 2488 3432
rect 2552 3368 2568 3432
rect 2632 3368 2648 3432
rect 2712 3368 2728 3432
rect 2792 3368 2808 3432
rect 2872 3368 2888 3432
rect 2952 3368 2968 3432
rect 3032 3368 3048 3432
rect 3112 3368 3128 3432
rect 3192 3368 3208 3432
rect 3272 3368 3288 3432
rect 3352 3368 3368 3432
rect 3432 3368 3448 3432
rect 3512 3368 3528 3432
rect 3592 3368 3608 3432
rect 3672 3368 3688 3432
rect 3752 3368 3768 3432
rect 3832 3368 3848 3432
rect 3912 3368 3928 3432
rect 3992 3368 19112 3432
rect 19176 3368 19192 3432
rect 19256 3368 19272 3432
rect 19336 3368 19352 3432
rect 19416 3368 29112 3432
rect 29176 3368 29192 3432
rect 29256 3368 29272 3432
rect 29336 3368 29352 3432
rect 29416 3368 41376 3432
rect 41440 3368 41456 3432
rect 41520 3368 41536 3432
rect 41600 3368 41616 3432
rect 41680 3368 41696 3432
rect 41760 3368 41776 3432
rect 41840 3368 41856 3432
rect 41920 3368 41936 3432
rect 42000 3368 42016 3432
rect 42080 3368 42096 3432
rect 42160 3368 42176 3432
rect 42240 3368 42256 3432
rect 42320 3368 42336 3432
rect 42400 3368 42416 3432
rect 42480 3368 42496 3432
rect 42560 3368 42576 3432
rect 42640 3368 42656 3432
rect 42720 3368 42736 3432
rect 42800 3368 42816 3432
rect 42880 3368 42896 3432
rect 42960 3368 42976 3432
rect 43040 3368 43056 3432
rect 43120 3368 43136 3432
rect 43200 3368 43216 3432
rect 43280 3368 43296 3432
rect 43360 3368 43376 3432
rect 43440 3368 43456 3432
rect 43520 3368 43536 3432
rect 43600 3368 43616 3432
rect 43680 3368 43696 3432
rect 43760 3368 43776 3432
rect 43840 3368 43856 3432
rect 43920 3368 43936 3432
rect 44000 3368 44016 3432
rect 44080 3368 44096 3432
rect 44160 3368 44176 3432
rect 44240 3368 44256 3432
rect 44320 3368 44336 3432
rect 44400 3368 44416 3432
rect 44480 3368 44496 3432
rect 44560 3368 44576 3432
rect 44640 3368 44656 3432
rect 44720 3368 44736 3432
rect 44800 3368 44816 3432
rect 44880 3368 44896 3432
rect 44960 3368 44976 3432
rect 45040 3368 45056 3432
rect 45120 3368 45136 3432
rect 45200 3368 45216 3432
rect 45280 3368 45296 3432
rect 45360 3368 45368 3432
rect 0 3352 45368 3368
rect 0 3288 8 3352
rect 72 3288 88 3352
rect 152 3288 168 3352
rect 232 3288 248 3352
rect 312 3288 328 3352
rect 392 3288 408 3352
rect 472 3288 488 3352
rect 552 3288 568 3352
rect 632 3288 648 3352
rect 712 3288 728 3352
rect 792 3288 808 3352
rect 872 3288 888 3352
rect 952 3288 968 3352
rect 1032 3288 1048 3352
rect 1112 3288 1128 3352
rect 1192 3288 1208 3352
rect 1272 3288 1288 3352
rect 1352 3288 1368 3352
rect 1432 3288 1448 3352
rect 1512 3288 1528 3352
rect 1592 3288 1608 3352
rect 1672 3288 1688 3352
rect 1752 3288 1768 3352
rect 1832 3288 1848 3352
rect 1912 3288 1928 3352
rect 1992 3288 2008 3352
rect 2072 3288 2088 3352
rect 2152 3288 2168 3352
rect 2232 3288 2248 3352
rect 2312 3288 2328 3352
rect 2392 3288 2408 3352
rect 2472 3288 2488 3352
rect 2552 3288 2568 3352
rect 2632 3288 2648 3352
rect 2712 3288 2728 3352
rect 2792 3288 2808 3352
rect 2872 3288 2888 3352
rect 2952 3288 2968 3352
rect 3032 3288 3048 3352
rect 3112 3288 3128 3352
rect 3192 3288 3208 3352
rect 3272 3288 3288 3352
rect 3352 3288 3368 3352
rect 3432 3288 3448 3352
rect 3512 3288 3528 3352
rect 3592 3288 3608 3352
rect 3672 3288 3688 3352
rect 3752 3288 3768 3352
rect 3832 3288 3848 3352
rect 3912 3288 3928 3352
rect 3992 3288 19112 3352
rect 19176 3288 19192 3352
rect 19256 3288 19272 3352
rect 19336 3288 19352 3352
rect 19416 3288 29112 3352
rect 29176 3288 29192 3352
rect 29256 3288 29272 3352
rect 29336 3288 29352 3352
rect 29416 3288 41376 3352
rect 41440 3288 41456 3352
rect 41520 3288 41536 3352
rect 41600 3288 41616 3352
rect 41680 3288 41696 3352
rect 41760 3288 41776 3352
rect 41840 3288 41856 3352
rect 41920 3288 41936 3352
rect 42000 3288 42016 3352
rect 42080 3288 42096 3352
rect 42160 3288 42176 3352
rect 42240 3288 42256 3352
rect 42320 3288 42336 3352
rect 42400 3288 42416 3352
rect 42480 3288 42496 3352
rect 42560 3288 42576 3352
rect 42640 3288 42656 3352
rect 42720 3288 42736 3352
rect 42800 3288 42816 3352
rect 42880 3288 42896 3352
rect 42960 3288 42976 3352
rect 43040 3288 43056 3352
rect 43120 3288 43136 3352
rect 43200 3288 43216 3352
rect 43280 3288 43296 3352
rect 43360 3288 43376 3352
rect 43440 3288 43456 3352
rect 43520 3288 43536 3352
rect 43600 3288 43616 3352
rect 43680 3288 43696 3352
rect 43760 3288 43776 3352
rect 43840 3288 43856 3352
rect 43920 3288 43936 3352
rect 44000 3288 44016 3352
rect 44080 3288 44096 3352
rect 44160 3288 44176 3352
rect 44240 3288 44256 3352
rect 44320 3288 44336 3352
rect 44400 3288 44416 3352
rect 44480 3288 44496 3352
rect 44560 3288 44576 3352
rect 44640 3288 44656 3352
rect 44720 3288 44736 3352
rect 44800 3288 44816 3352
rect 44880 3288 44896 3352
rect 44960 3288 44976 3352
rect 45040 3288 45056 3352
rect 45120 3288 45136 3352
rect 45200 3288 45216 3352
rect 45280 3288 45296 3352
rect 45360 3288 45368 3352
rect 0 3272 45368 3288
rect 0 3208 8 3272
rect 72 3208 88 3272
rect 152 3208 168 3272
rect 232 3208 248 3272
rect 312 3208 328 3272
rect 392 3208 408 3272
rect 472 3208 488 3272
rect 552 3208 568 3272
rect 632 3208 648 3272
rect 712 3208 728 3272
rect 792 3208 808 3272
rect 872 3208 888 3272
rect 952 3208 968 3272
rect 1032 3208 1048 3272
rect 1112 3208 1128 3272
rect 1192 3208 1208 3272
rect 1272 3208 1288 3272
rect 1352 3208 1368 3272
rect 1432 3208 1448 3272
rect 1512 3208 1528 3272
rect 1592 3208 1608 3272
rect 1672 3208 1688 3272
rect 1752 3208 1768 3272
rect 1832 3208 1848 3272
rect 1912 3208 1928 3272
rect 1992 3208 2008 3272
rect 2072 3208 2088 3272
rect 2152 3208 2168 3272
rect 2232 3208 2248 3272
rect 2312 3208 2328 3272
rect 2392 3208 2408 3272
rect 2472 3208 2488 3272
rect 2552 3208 2568 3272
rect 2632 3208 2648 3272
rect 2712 3208 2728 3272
rect 2792 3208 2808 3272
rect 2872 3208 2888 3272
rect 2952 3208 2968 3272
rect 3032 3208 3048 3272
rect 3112 3208 3128 3272
rect 3192 3208 3208 3272
rect 3272 3208 3288 3272
rect 3352 3208 3368 3272
rect 3432 3208 3448 3272
rect 3512 3208 3528 3272
rect 3592 3208 3608 3272
rect 3672 3208 3688 3272
rect 3752 3208 3768 3272
rect 3832 3208 3848 3272
rect 3912 3208 3928 3272
rect 3992 3208 19112 3272
rect 19176 3208 19192 3272
rect 19256 3208 19272 3272
rect 19336 3208 19352 3272
rect 19416 3208 29112 3272
rect 29176 3208 29192 3272
rect 29256 3208 29272 3272
rect 29336 3208 29352 3272
rect 29416 3208 41376 3272
rect 41440 3208 41456 3272
rect 41520 3208 41536 3272
rect 41600 3208 41616 3272
rect 41680 3208 41696 3272
rect 41760 3208 41776 3272
rect 41840 3208 41856 3272
rect 41920 3208 41936 3272
rect 42000 3208 42016 3272
rect 42080 3208 42096 3272
rect 42160 3208 42176 3272
rect 42240 3208 42256 3272
rect 42320 3208 42336 3272
rect 42400 3208 42416 3272
rect 42480 3208 42496 3272
rect 42560 3208 42576 3272
rect 42640 3208 42656 3272
rect 42720 3208 42736 3272
rect 42800 3208 42816 3272
rect 42880 3208 42896 3272
rect 42960 3208 42976 3272
rect 43040 3208 43056 3272
rect 43120 3208 43136 3272
rect 43200 3208 43216 3272
rect 43280 3208 43296 3272
rect 43360 3208 43376 3272
rect 43440 3208 43456 3272
rect 43520 3208 43536 3272
rect 43600 3208 43616 3272
rect 43680 3208 43696 3272
rect 43760 3208 43776 3272
rect 43840 3208 43856 3272
rect 43920 3208 43936 3272
rect 44000 3208 44016 3272
rect 44080 3208 44096 3272
rect 44160 3208 44176 3272
rect 44240 3208 44256 3272
rect 44320 3208 44336 3272
rect 44400 3208 44416 3272
rect 44480 3208 44496 3272
rect 44560 3208 44576 3272
rect 44640 3208 44656 3272
rect 44720 3208 44736 3272
rect 44800 3208 44816 3272
rect 44880 3208 44896 3272
rect 44960 3208 44976 3272
rect 45040 3208 45056 3272
rect 45120 3208 45136 3272
rect 45200 3208 45216 3272
rect 45280 3208 45296 3272
rect 45360 3208 45368 3272
rect 0 3192 45368 3208
rect 0 3128 8 3192
rect 72 3128 88 3192
rect 152 3128 168 3192
rect 232 3128 248 3192
rect 312 3128 328 3192
rect 392 3128 408 3192
rect 472 3128 488 3192
rect 552 3128 568 3192
rect 632 3128 648 3192
rect 712 3128 728 3192
rect 792 3128 808 3192
rect 872 3128 888 3192
rect 952 3128 968 3192
rect 1032 3128 1048 3192
rect 1112 3128 1128 3192
rect 1192 3128 1208 3192
rect 1272 3128 1288 3192
rect 1352 3128 1368 3192
rect 1432 3128 1448 3192
rect 1512 3128 1528 3192
rect 1592 3128 1608 3192
rect 1672 3128 1688 3192
rect 1752 3128 1768 3192
rect 1832 3128 1848 3192
rect 1912 3128 1928 3192
rect 1992 3128 2008 3192
rect 2072 3128 2088 3192
rect 2152 3128 2168 3192
rect 2232 3128 2248 3192
rect 2312 3128 2328 3192
rect 2392 3128 2408 3192
rect 2472 3128 2488 3192
rect 2552 3128 2568 3192
rect 2632 3128 2648 3192
rect 2712 3128 2728 3192
rect 2792 3128 2808 3192
rect 2872 3128 2888 3192
rect 2952 3128 2968 3192
rect 3032 3128 3048 3192
rect 3112 3128 3128 3192
rect 3192 3128 3208 3192
rect 3272 3128 3288 3192
rect 3352 3128 3368 3192
rect 3432 3128 3448 3192
rect 3512 3128 3528 3192
rect 3592 3128 3608 3192
rect 3672 3128 3688 3192
rect 3752 3128 3768 3192
rect 3832 3128 3848 3192
rect 3912 3128 3928 3192
rect 3992 3128 19112 3192
rect 19176 3128 19192 3192
rect 19256 3128 19272 3192
rect 19336 3128 19352 3192
rect 19416 3128 29112 3192
rect 29176 3128 29192 3192
rect 29256 3128 29272 3192
rect 29336 3128 29352 3192
rect 29416 3128 41376 3192
rect 41440 3128 41456 3192
rect 41520 3128 41536 3192
rect 41600 3128 41616 3192
rect 41680 3128 41696 3192
rect 41760 3128 41776 3192
rect 41840 3128 41856 3192
rect 41920 3128 41936 3192
rect 42000 3128 42016 3192
rect 42080 3128 42096 3192
rect 42160 3128 42176 3192
rect 42240 3128 42256 3192
rect 42320 3128 42336 3192
rect 42400 3128 42416 3192
rect 42480 3128 42496 3192
rect 42560 3128 42576 3192
rect 42640 3128 42656 3192
rect 42720 3128 42736 3192
rect 42800 3128 42816 3192
rect 42880 3128 42896 3192
rect 42960 3128 42976 3192
rect 43040 3128 43056 3192
rect 43120 3128 43136 3192
rect 43200 3128 43216 3192
rect 43280 3128 43296 3192
rect 43360 3128 43376 3192
rect 43440 3128 43456 3192
rect 43520 3128 43536 3192
rect 43600 3128 43616 3192
rect 43680 3128 43696 3192
rect 43760 3128 43776 3192
rect 43840 3128 43856 3192
rect 43920 3128 43936 3192
rect 44000 3128 44016 3192
rect 44080 3128 44096 3192
rect 44160 3128 44176 3192
rect 44240 3128 44256 3192
rect 44320 3128 44336 3192
rect 44400 3128 44416 3192
rect 44480 3128 44496 3192
rect 44560 3128 44576 3192
rect 44640 3128 44656 3192
rect 44720 3128 44736 3192
rect 44800 3128 44816 3192
rect 44880 3128 44896 3192
rect 44960 3128 44976 3192
rect 45040 3128 45056 3192
rect 45120 3128 45136 3192
rect 45200 3128 45216 3192
rect 45280 3128 45296 3192
rect 45360 3128 45368 3192
rect 0 3112 45368 3128
rect 0 3048 8 3112
rect 72 3048 88 3112
rect 152 3048 168 3112
rect 232 3048 248 3112
rect 312 3048 328 3112
rect 392 3048 408 3112
rect 472 3048 488 3112
rect 552 3048 568 3112
rect 632 3048 648 3112
rect 712 3048 728 3112
rect 792 3048 808 3112
rect 872 3048 888 3112
rect 952 3048 968 3112
rect 1032 3048 1048 3112
rect 1112 3048 1128 3112
rect 1192 3048 1208 3112
rect 1272 3048 1288 3112
rect 1352 3048 1368 3112
rect 1432 3048 1448 3112
rect 1512 3048 1528 3112
rect 1592 3048 1608 3112
rect 1672 3048 1688 3112
rect 1752 3048 1768 3112
rect 1832 3048 1848 3112
rect 1912 3048 1928 3112
rect 1992 3048 2008 3112
rect 2072 3048 2088 3112
rect 2152 3048 2168 3112
rect 2232 3048 2248 3112
rect 2312 3048 2328 3112
rect 2392 3048 2408 3112
rect 2472 3048 2488 3112
rect 2552 3048 2568 3112
rect 2632 3048 2648 3112
rect 2712 3048 2728 3112
rect 2792 3048 2808 3112
rect 2872 3048 2888 3112
rect 2952 3048 2968 3112
rect 3032 3048 3048 3112
rect 3112 3048 3128 3112
rect 3192 3048 3208 3112
rect 3272 3048 3288 3112
rect 3352 3048 3368 3112
rect 3432 3048 3448 3112
rect 3512 3048 3528 3112
rect 3592 3048 3608 3112
rect 3672 3048 3688 3112
rect 3752 3048 3768 3112
rect 3832 3048 3848 3112
rect 3912 3048 3928 3112
rect 3992 3048 19112 3112
rect 19176 3048 19192 3112
rect 19256 3048 19272 3112
rect 19336 3048 19352 3112
rect 19416 3048 29112 3112
rect 29176 3048 29192 3112
rect 29256 3048 29272 3112
rect 29336 3048 29352 3112
rect 29416 3048 41376 3112
rect 41440 3048 41456 3112
rect 41520 3048 41536 3112
rect 41600 3048 41616 3112
rect 41680 3048 41696 3112
rect 41760 3048 41776 3112
rect 41840 3048 41856 3112
rect 41920 3048 41936 3112
rect 42000 3048 42016 3112
rect 42080 3048 42096 3112
rect 42160 3048 42176 3112
rect 42240 3048 42256 3112
rect 42320 3048 42336 3112
rect 42400 3048 42416 3112
rect 42480 3048 42496 3112
rect 42560 3048 42576 3112
rect 42640 3048 42656 3112
rect 42720 3048 42736 3112
rect 42800 3048 42816 3112
rect 42880 3048 42896 3112
rect 42960 3048 42976 3112
rect 43040 3048 43056 3112
rect 43120 3048 43136 3112
rect 43200 3048 43216 3112
rect 43280 3048 43296 3112
rect 43360 3048 43376 3112
rect 43440 3048 43456 3112
rect 43520 3048 43536 3112
rect 43600 3048 43616 3112
rect 43680 3048 43696 3112
rect 43760 3048 43776 3112
rect 43840 3048 43856 3112
rect 43920 3048 43936 3112
rect 44000 3048 44016 3112
rect 44080 3048 44096 3112
rect 44160 3048 44176 3112
rect 44240 3048 44256 3112
rect 44320 3048 44336 3112
rect 44400 3048 44416 3112
rect 44480 3048 44496 3112
rect 44560 3048 44576 3112
rect 44640 3048 44656 3112
rect 44720 3048 44736 3112
rect 44800 3048 44816 3112
rect 44880 3048 44896 3112
rect 44960 3048 44976 3112
rect 45040 3048 45056 3112
rect 45120 3048 45136 3112
rect 45200 3048 45216 3112
rect 45280 3048 45296 3112
rect 45360 3048 45368 3112
rect 0 3032 45368 3048
rect 0 2968 8 3032
rect 72 2968 88 3032
rect 152 2968 168 3032
rect 232 2968 248 3032
rect 312 2968 328 3032
rect 392 2968 408 3032
rect 472 2968 488 3032
rect 552 2968 568 3032
rect 632 2968 648 3032
rect 712 2968 728 3032
rect 792 2968 808 3032
rect 872 2968 888 3032
rect 952 2968 968 3032
rect 1032 2968 1048 3032
rect 1112 2968 1128 3032
rect 1192 2968 1208 3032
rect 1272 2968 1288 3032
rect 1352 2968 1368 3032
rect 1432 2968 1448 3032
rect 1512 2968 1528 3032
rect 1592 2968 1608 3032
rect 1672 2968 1688 3032
rect 1752 2968 1768 3032
rect 1832 2968 1848 3032
rect 1912 2968 1928 3032
rect 1992 2968 2008 3032
rect 2072 2968 2088 3032
rect 2152 2968 2168 3032
rect 2232 2968 2248 3032
rect 2312 2968 2328 3032
rect 2392 2968 2408 3032
rect 2472 2968 2488 3032
rect 2552 2968 2568 3032
rect 2632 2968 2648 3032
rect 2712 2968 2728 3032
rect 2792 2968 2808 3032
rect 2872 2968 2888 3032
rect 2952 2968 2968 3032
rect 3032 2968 3048 3032
rect 3112 2968 3128 3032
rect 3192 2968 3208 3032
rect 3272 2968 3288 3032
rect 3352 2968 3368 3032
rect 3432 2968 3448 3032
rect 3512 2968 3528 3032
rect 3592 2968 3608 3032
rect 3672 2968 3688 3032
rect 3752 2968 3768 3032
rect 3832 2968 3848 3032
rect 3912 2968 3928 3032
rect 3992 2968 19112 3032
rect 19176 2968 19192 3032
rect 19256 2968 19272 3032
rect 19336 2968 19352 3032
rect 19416 2968 29112 3032
rect 29176 2968 29192 3032
rect 29256 2968 29272 3032
rect 29336 2968 29352 3032
rect 29416 2968 41376 3032
rect 41440 2968 41456 3032
rect 41520 2968 41536 3032
rect 41600 2968 41616 3032
rect 41680 2968 41696 3032
rect 41760 2968 41776 3032
rect 41840 2968 41856 3032
rect 41920 2968 41936 3032
rect 42000 2968 42016 3032
rect 42080 2968 42096 3032
rect 42160 2968 42176 3032
rect 42240 2968 42256 3032
rect 42320 2968 42336 3032
rect 42400 2968 42416 3032
rect 42480 2968 42496 3032
rect 42560 2968 42576 3032
rect 42640 2968 42656 3032
rect 42720 2968 42736 3032
rect 42800 2968 42816 3032
rect 42880 2968 42896 3032
rect 42960 2968 42976 3032
rect 43040 2968 43056 3032
rect 43120 2968 43136 3032
rect 43200 2968 43216 3032
rect 43280 2968 43296 3032
rect 43360 2968 43376 3032
rect 43440 2968 43456 3032
rect 43520 2968 43536 3032
rect 43600 2968 43616 3032
rect 43680 2968 43696 3032
rect 43760 2968 43776 3032
rect 43840 2968 43856 3032
rect 43920 2968 43936 3032
rect 44000 2968 44016 3032
rect 44080 2968 44096 3032
rect 44160 2968 44176 3032
rect 44240 2968 44256 3032
rect 44320 2968 44336 3032
rect 44400 2968 44416 3032
rect 44480 2968 44496 3032
rect 44560 2968 44576 3032
rect 44640 2968 44656 3032
rect 44720 2968 44736 3032
rect 44800 2968 44816 3032
rect 44880 2968 44896 3032
rect 44960 2968 44976 3032
rect 45040 2968 45056 3032
rect 45120 2968 45136 3032
rect 45200 2968 45216 3032
rect 45280 2968 45296 3032
rect 45360 2968 45368 3032
rect 0 2952 45368 2968
rect 0 2888 8 2952
rect 72 2888 88 2952
rect 152 2888 168 2952
rect 232 2888 248 2952
rect 312 2888 328 2952
rect 392 2888 408 2952
rect 472 2888 488 2952
rect 552 2888 568 2952
rect 632 2888 648 2952
rect 712 2888 728 2952
rect 792 2888 808 2952
rect 872 2888 888 2952
rect 952 2888 968 2952
rect 1032 2888 1048 2952
rect 1112 2888 1128 2952
rect 1192 2888 1208 2952
rect 1272 2888 1288 2952
rect 1352 2888 1368 2952
rect 1432 2888 1448 2952
rect 1512 2888 1528 2952
rect 1592 2888 1608 2952
rect 1672 2888 1688 2952
rect 1752 2888 1768 2952
rect 1832 2888 1848 2952
rect 1912 2888 1928 2952
rect 1992 2888 2008 2952
rect 2072 2888 2088 2952
rect 2152 2888 2168 2952
rect 2232 2888 2248 2952
rect 2312 2888 2328 2952
rect 2392 2888 2408 2952
rect 2472 2888 2488 2952
rect 2552 2888 2568 2952
rect 2632 2888 2648 2952
rect 2712 2888 2728 2952
rect 2792 2888 2808 2952
rect 2872 2888 2888 2952
rect 2952 2888 2968 2952
rect 3032 2888 3048 2952
rect 3112 2888 3128 2952
rect 3192 2888 3208 2952
rect 3272 2888 3288 2952
rect 3352 2888 3368 2952
rect 3432 2888 3448 2952
rect 3512 2888 3528 2952
rect 3592 2888 3608 2952
rect 3672 2888 3688 2952
rect 3752 2888 3768 2952
rect 3832 2888 3848 2952
rect 3912 2888 3928 2952
rect 3992 2888 19112 2952
rect 19176 2888 19192 2952
rect 19256 2888 19272 2952
rect 19336 2888 19352 2952
rect 19416 2888 29112 2952
rect 29176 2888 29192 2952
rect 29256 2888 29272 2952
rect 29336 2888 29352 2952
rect 29416 2888 41376 2952
rect 41440 2888 41456 2952
rect 41520 2888 41536 2952
rect 41600 2888 41616 2952
rect 41680 2888 41696 2952
rect 41760 2888 41776 2952
rect 41840 2888 41856 2952
rect 41920 2888 41936 2952
rect 42000 2888 42016 2952
rect 42080 2888 42096 2952
rect 42160 2888 42176 2952
rect 42240 2888 42256 2952
rect 42320 2888 42336 2952
rect 42400 2888 42416 2952
rect 42480 2888 42496 2952
rect 42560 2888 42576 2952
rect 42640 2888 42656 2952
rect 42720 2888 42736 2952
rect 42800 2888 42816 2952
rect 42880 2888 42896 2952
rect 42960 2888 42976 2952
rect 43040 2888 43056 2952
rect 43120 2888 43136 2952
rect 43200 2888 43216 2952
rect 43280 2888 43296 2952
rect 43360 2888 43376 2952
rect 43440 2888 43456 2952
rect 43520 2888 43536 2952
rect 43600 2888 43616 2952
rect 43680 2888 43696 2952
rect 43760 2888 43776 2952
rect 43840 2888 43856 2952
rect 43920 2888 43936 2952
rect 44000 2888 44016 2952
rect 44080 2888 44096 2952
rect 44160 2888 44176 2952
rect 44240 2888 44256 2952
rect 44320 2888 44336 2952
rect 44400 2888 44416 2952
rect 44480 2888 44496 2952
rect 44560 2888 44576 2952
rect 44640 2888 44656 2952
rect 44720 2888 44736 2952
rect 44800 2888 44816 2952
rect 44880 2888 44896 2952
rect 44960 2888 44976 2952
rect 45040 2888 45056 2952
rect 45120 2888 45136 2952
rect 45200 2888 45216 2952
rect 45280 2888 45296 2952
rect 45360 2888 45368 2952
rect 0 2872 45368 2888
rect 0 2808 8 2872
rect 72 2808 88 2872
rect 152 2808 168 2872
rect 232 2808 248 2872
rect 312 2808 328 2872
rect 392 2808 408 2872
rect 472 2808 488 2872
rect 552 2808 568 2872
rect 632 2808 648 2872
rect 712 2808 728 2872
rect 792 2808 808 2872
rect 872 2808 888 2872
rect 952 2808 968 2872
rect 1032 2808 1048 2872
rect 1112 2808 1128 2872
rect 1192 2808 1208 2872
rect 1272 2808 1288 2872
rect 1352 2808 1368 2872
rect 1432 2808 1448 2872
rect 1512 2808 1528 2872
rect 1592 2808 1608 2872
rect 1672 2808 1688 2872
rect 1752 2808 1768 2872
rect 1832 2808 1848 2872
rect 1912 2808 1928 2872
rect 1992 2808 2008 2872
rect 2072 2808 2088 2872
rect 2152 2808 2168 2872
rect 2232 2808 2248 2872
rect 2312 2808 2328 2872
rect 2392 2808 2408 2872
rect 2472 2808 2488 2872
rect 2552 2808 2568 2872
rect 2632 2808 2648 2872
rect 2712 2808 2728 2872
rect 2792 2808 2808 2872
rect 2872 2808 2888 2872
rect 2952 2808 2968 2872
rect 3032 2808 3048 2872
rect 3112 2808 3128 2872
rect 3192 2808 3208 2872
rect 3272 2808 3288 2872
rect 3352 2808 3368 2872
rect 3432 2808 3448 2872
rect 3512 2808 3528 2872
rect 3592 2808 3608 2872
rect 3672 2808 3688 2872
rect 3752 2808 3768 2872
rect 3832 2808 3848 2872
rect 3912 2808 3928 2872
rect 3992 2808 19112 2872
rect 19176 2808 19192 2872
rect 19256 2808 19272 2872
rect 19336 2808 19352 2872
rect 19416 2808 29112 2872
rect 29176 2808 29192 2872
rect 29256 2808 29272 2872
rect 29336 2808 29352 2872
rect 29416 2808 41376 2872
rect 41440 2808 41456 2872
rect 41520 2808 41536 2872
rect 41600 2808 41616 2872
rect 41680 2808 41696 2872
rect 41760 2808 41776 2872
rect 41840 2808 41856 2872
rect 41920 2808 41936 2872
rect 42000 2808 42016 2872
rect 42080 2808 42096 2872
rect 42160 2808 42176 2872
rect 42240 2808 42256 2872
rect 42320 2808 42336 2872
rect 42400 2808 42416 2872
rect 42480 2808 42496 2872
rect 42560 2808 42576 2872
rect 42640 2808 42656 2872
rect 42720 2808 42736 2872
rect 42800 2808 42816 2872
rect 42880 2808 42896 2872
rect 42960 2808 42976 2872
rect 43040 2808 43056 2872
rect 43120 2808 43136 2872
rect 43200 2808 43216 2872
rect 43280 2808 43296 2872
rect 43360 2808 43376 2872
rect 43440 2808 43456 2872
rect 43520 2808 43536 2872
rect 43600 2808 43616 2872
rect 43680 2808 43696 2872
rect 43760 2808 43776 2872
rect 43840 2808 43856 2872
rect 43920 2808 43936 2872
rect 44000 2808 44016 2872
rect 44080 2808 44096 2872
rect 44160 2808 44176 2872
rect 44240 2808 44256 2872
rect 44320 2808 44336 2872
rect 44400 2808 44416 2872
rect 44480 2808 44496 2872
rect 44560 2808 44576 2872
rect 44640 2808 44656 2872
rect 44720 2808 44736 2872
rect 44800 2808 44816 2872
rect 44880 2808 44896 2872
rect 44960 2808 44976 2872
rect 45040 2808 45056 2872
rect 45120 2808 45136 2872
rect 45200 2808 45216 2872
rect 45280 2808 45296 2872
rect 45360 2808 45368 2872
rect 0 2792 45368 2808
rect 0 2728 8 2792
rect 72 2728 88 2792
rect 152 2728 168 2792
rect 232 2728 248 2792
rect 312 2728 328 2792
rect 392 2728 408 2792
rect 472 2728 488 2792
rect 552 2728 568 2792
rect 632 2728 648 2792
rect 712 2728 728 2792
rect 792 2728 808 2792
rect 872 2728 888 2792
rect 952 2728 968 2792
rect 1032 2728 1048 2792
rect 1112 2728 1128 2792
rect 1192 2728 1208 2792
rect 1272 2728 1288 2792
rect 1352 2728 1368 2792
rect 1432 2728 1448 2792
rect 1512 2728 1528 2792
rect 1592 2728 1608 2792
rect 1672 2728 1688 2792
rect 1752 2728 1768 2792
rect 1832 2728 1848 2792
rect 1912 2728 1928 2792
rect 1992 2728 2008 2792
rect 2072 2728 2088 2792
rect 2152 2728 2168 2792
rect 2232 2728 2248 2792
rect 2312 2728 2328 2792
rect 2392 2728 2408 2792
rect 2472 2728 2488 2792
rect 2552 2728 2568 2792
rect 2632 2728 2648 2792
rect 2712 2728 2728 2792
rect 2792 2728 2808 2792
rect 2872 2728 2888 2792
rect 2952 2728 2968 2792
rect 3032 2728 3048 2792
rect 3112 2728 3128 2792
rect 3192 2728 3208 2792
rect 3272 2728 3288 2792
rect 3352 2728 3368 2792
rect 3432 2728 3448 2792
rect 3512 2728 3528 2792
rect 3592 2728 3608 2792
rect 3672 2728 3688 2792
rect 3752 2728 3768 2792
rect 3832 2728 3848 2792
rect 3912 2728 3928 2792
rect 3992 2728 19112 2792
rect 19176 2728 19192 2792
rect 19256 2728 19272 2792
rect 19336 2728 19352 2792
rect 19416 2728 29112 2792
rect 29176 2728 29192 2792
rect 29256 2728 29272 2792
rect 29336 2728 29352 2792
rect 29416 2728 41376 2792
rect 41440 2728 41456 2792
rect 41520 2728 41536 2792
rect 41600 2728 41616 2792
rect 41680 2728 41696 2792
rect 41760 2728 41776 2792
rect 41840 2728 41856 2792
rect 41920 2728 41936 2792
rect 42000 2728 42016 2792
rect 42080 2728 42096 2792
rect 42160 2728 42176 2792
rect 42240 2728 42256 2792
rect 42320 2728 42336 2792
rect 42400 2728 42416 2792
rect 42480 2728 42496 2792
rect 42560 2728 42576 2792
rect 42640 2728 42656 2792
rect 42720 2728 42736 2792
rect 42800 2728 42816 2792
rect 42880 2728 42896 2792
rect 42960 2728 42976 2792
rect 43040 2728 43056 2792
rect 43120 2728 43136 2792
rect 43200 2728 43216 2792
rect 43280 2728 43296 2792
rect 43360 2728 43376 2792
rect 43440 2728 43456 2792
rect 43520 2728 43536 2792
rect 43600 2728 43616 2792
rect 43680 2728 43696 2792
rect 43760 2728 43776 2792
rect 43840 2728 43856 2792
rect 43920 2728 43936 2792
rect 44000 2728 44016 2792
rect 44080 2728 44096 2792
rect 44160 2728 44176 2792
rect 44240 2728 44256 2792
rect 44320 2728 44336 2792
rect 44400 2728 44416 2792
rect 44480 2728 44496 2792
rect 44560 2728 44576 2792
rect 44640 2728 44656 2792
rect 44720 2728 44736 2792
rect 44800 2728 44816 2792
rect 44880 2728 44896 2792
rect 44960 2728 44976 2792
rect 45040 2728 45056 2792
rect 45120 2728 45136 2792
rect 45200 2728 45216 2792
rect 45280 2728 45296 2792
rect 45360 2728 45368 2792
rect 0 2712 45368 2728
rect 0 2648 8 2712
rect 72 2648 88 2712
rect 152 2648 168 2712
rect 232 2648 248 2712
rect 312 2648 328 2712
rect 392 2648 408 2712
rect 472 2648 488 2712
rect 552 2648 568 2712
rect 632 2648 648 2712
rect 712 2648 728 2712
rect 792 2648 808 2712
rect 872 2648 888 2712
rect 952 2648 968 2712
rect 1032 2648 1048 2712
rect 1112 2648 1128 2712
rect 1192 2648 1208 2712
rect 1272 2648 1288 2712
rect 1352 2648 1368 2712
rect 1432 2648 1448 2712
rect 1512 2648 1528 2712
rect 1592 2648 1608 2712
rect 1672 2648 1688 2712
rect 1752 2648 1768 2712
rect 1832 2648 1848 2712
rect 1912 2648 1928 2712
rect 1992 2648 2008 2712
rect 2072 2648 2088 2712
rect 2152 2648 2168 2712
rect 2232 2648 2248 2712
rect 2312 2648 2328 2712
rect 2392 2648 2408 2712
rect 2472 2648 2488 2712
rect 2552 2648 2568 2712
rect 2632 2648 2648 2712
rect 2712 2648 2728 2712
rect 2792 2648 2808 2712
rect 2872 2648 2888 2712
rect 2952 2648 2968 2712
rect 3032 2648 3048 2712
rect 3112 2648 3128 2712
rect 3192 2648 3208 2712
rect 3272 2648 3288 2712
rect 3352 2648 3368 2712
rect 3432 2648 3448 2712
rect 3512 2648 3528 2712
rect 3592 2648 3608 2712
rect 3672 2648 3688 2712
rect 3752 2648 3768 2712
rect 3832 2648 3848 2712
rect 3912 2648 3928 2712
rect 3992 2648 19112 2712
rect 19176 2648 19192 2712
rect 19256 2648 19272 2712
rect 19336 2648 19352 2712
rect 19416 2648 29112 2712
rect 29176 2648 29192 2712
rect 29256 2648 29272 2712
rect 29336 2648 29352 2712
rect 29416 2648 41376 2712
rect 41440 2648 41456 2712
rect 41520 2648 41536 2712
rect 41600 2648 41616 2712
rect 41680 2648 41696 2712
rect 41760 2648 41776 2712
rect 41840 2648 41856 2712
rect 41920 2648 41936 2712
rect 42000 2648 42016 2712
rect 42080 2648 42096 2712
rect 42160 2648 42176 2712
rect 42240 2648 42256 2712
rect 42320 2648 42336 2712
rect 42400 2648 42416 2712
rect 42480 2648 42496 2712
rect 42560 2648 42576 2712
rect 42640 2648 42656 2712
rect 42720 2648 42736 2712
rect 42800 2648 42816 2712
rect 42880 2648 42896 2712
rect 42960 2648 42976 2712
rect 43040 2648 43056 2712
rect 43120 2648 43136 2712
rect 43200 2648 43216 2712
rect 43280 2648 43296 2712
rect 43360 2648 43376 2712
rect 43440 2648 43456 2712
rect 43520 2648 43536 2712
rect 43600 2648 43616 2712
rect 43680 2648 43696 2712
rect 43760 2648 43776 2712
rect 43840 2648 43856 2712
rect 43920 2648 43936 2712
rect 44000 2648 44016 2712
rect 44080 2648 44096 2712
rect 44160 2648 44176 2712
rect 44240 2648 44256 2712
rect 44320 2648 44336 2712
rect 44400 2648 44416 2712
rect 44480 2648 44496 2712
rect 44560 2648 44576 2712
rect 44640 2648 44656 2712
rect 44720 2648 44736 2712
rect 44800 2648 44816 2712
rect 44880 2648 44896 2712
rect 44960 2648 44976 2712
rect 45040 2648 45056 2712
rect 45120 2648 45136 2712
rect 45200 2648 45216 2712
rect 45280 2648 45296 2712
rect 45360 2648 45368 2712
rect 0 2632 45368 2648
rect 0 2568 8 2632
rect 72 2568 88 2632
rect 152 2568 168 2632
rect 232 2568 248 2632
rect 312 2568 328 2632
rect 392 2568 408 2632
rect 472 2568 488 2632
rect 552 2568 568 2632
rect 632 2568 648 2632
rect 712 2568 728 2632
rect 792 2568 808 2632
rect 872 2568 888 2632
rect 952 2568 968 2632
rect 1032 2568 1048 2632
rect 1112 2568 1128 2632
rect 1192 2568 1208 2632
rect 1272 2568 1288 2632
rect 1352 2568 1368 2632
rect 1432 2568 1448 2632
rect 1512 2568 1528 2632
rect 1592 2568 1608 2632
rect 1672 2568 1688 2632
rect 1752 2568 1768 2632
rect 1832 2568 1848 2632
rect 1912 2568 1928 2632
rect 1992 2568 2008 2632
rect 2072 2568 2088 2632
rect 2152 2568 2168 2632
rect 2232 2568 2248 2632
rect 2312 2568 2328 2632
rect 2392 2568 2408 2632
rect 2472 2568 2488 2632
rect 2552 2568 2568 2632
rect 2632 2568 2648 2632
rect 2712 2568 2728 2632
rect 2792 2568 2808 2632
rect 2872 2568 2888 2632
rect 2952 2568 2968 2632
rect 3032 2568 3048 2632
rect 3112 2568 3128 2632
rect 3192 2568 3208 2632
rect 3272 2568 3288 2632
rect 3352 2568 3368 2632
rect 3432 2568 3448 2632
rect 3512 2568 3528 2632
rect 3592 2568 3608 2632
rect 3672 2568 3688 2632
rect 3752 2568 3768 2632
rect 3832 2568 3848 2632
rect 3912 2568 3928 2632
rect 3992 2568 19112 2632
rect 19176 2568 19192 2632
rect 19256 2568 19272 2632
rect 19336 2568 19352 2632
rect 19416 2568 29112 2632
rect 29176 2568 29192 2632
rect 29256 2568 29272 2632
rect 29336 2568 29352 2632
rect 29416 2568 41376 2632
rect 41440 2568 41456 2632
rect 41520 2568 41536 2632
rect 41600 2568 41616 2632
rect 41680 2568 41696 2632
rect 41760 2568 41776 2632
rect 41840 2568 41856 2632
rect 41920 2568 41936 2632
rect 42000 2568 42016 2632
rect 42080 2568 42096 2632
rect 42160 2568 42176 2632
rect 42240 2568 42256 2632
rect 42320 2568 42336 2632
rect 42400 2568 42416 2632
rect 42480 2568 42496 2632
rect 42560 2568 42576 2632
rect 42640 2568 42656 2632
rect 42720 2568 42736 2632
rect 42800 2568 42816 2632
rect 42880 2568 42896 2632
rect 42960 2568 42976 2632
rect 43040 2568 43056 2632
rect 43120 2568 43136 2632
rect 43200 2568 43216 2632
rect 43280 2568 43296 2632
rect 43360 2568 43376 2632
rect 43440 2568 43456 2632
rect 43520 2568 43536 2632
rect 43600 2568 43616 2632
rect 43680 2568 43696 2632
rect 43760 2568 43776 2632
rect 43840 2568 43856 2632
rect 43920 2568 43936 2632
rect 44000 2568 44016 2632
rect 44080 2568 44096 2632
rect 44160 2568 44176 2632
rect 44240 2568 44256 2632
rect 44320 2568 44336 2632
rect 44400 2568 44416 2632
rect 44480 2568 44496 2632
rect 44560 2568 44576 2632
rect 44640 2568 44656 2632
rect 44720 2568 44736 2632
rect 44800 2568 44816 2632
rect 44880 2568 44896 2632
rect 44960 2568 44976 2632
rect 45040 2568 45056 2632
rect 45120 2568 45136 2632
rect 45200 2568 45216 2632
rect 45280 2568 45296 2632
rect 45360 2568 45368 2632
rect 0 2552 45368 2568
rect 0 2488 8 2552
rect 72 2488 88 2552
rect 152 2488 168 2552
rect 232 2488 248 2552
rect 312 2488 328 2552
rect 392 2488 408 2552
rect 472 2488 488 2552
rect 552 2488 568 2552
rect 632 2488 648 2552
rect 712 2488 728 2552
rect 792 2488 808 2552
rect 872 2488 888 2552
rect 952 2488 968 2552
rect 1032 2488 1048 2552
rect 1112 2488 1128 2552
rect 1192 2488 1208 2552
rect 1272 2488 1288 2552
rect 1352 2488 1368 2552
rect 1432 2488 1448 2552
rect 1512 2488 1528 2552
rect 1592 2488 1608 2552
rect 1672 2488 1688 2552
rect 1752 2488 1768 2552
rect 1832 2488 1848 2552
rect 1912 2488 1928 2552
rect 1992 2488 2008 2552
rect 2072 2488 2088 2552
rect 2152 2488 2168 2552
rect 2232 2488 2248 2552
rect 2312 2488 2328 2552
rect 2392 2488 2408 2552
rect 2472 2488 2488 2552
rect 2552 2488 2568 2552
rect 2632 2488 2648 2552
rect 2712 2488 2728 2552
rect 2792 2488 2808 2552
rect 2872 2488 2888 2552
rect 2952 2488 2968 2552
rect 3032 2488 3048 2552
rect 3112 2488 3128 2552
rect 3192 2488 3208 2552
rect 3272 2488 3288 2552
rect 3352 2488 3368 2552
rect 3432 2488 3448 2552
rect 3512 2488 3528 2552
rect 3592 2488 3608 2552
rect 3672 2488 3688 2552
rect 3752 2488 3768 2552
rect 3832 2488 3848 2552
rect 3912 2488 3928 2552
rect 3992 2488 19112 2552
rect 19176 2488 19192 2552
rect 19256 2488 19272 2552
rect 19336 2488 19352 2552
rect 19416 2488 29112 2552
rect 29176 2488 29192 2552
rect 29256 2488 29272 2552
rect 29336 2488 29352 2552
rect 29416 2488 41376 2552
rect 41440 2488 41456 2552
rect 41520 2488 41536 2552
rect 41600 2488 41616 2552
rect 41680 2488 41696 2552
rect 41760 2488 41776 2552
rect 41840 2488 41856 2552
rect 41920 2488 41936 2552
rect 42000 2488 42016 2552
rect 42080 2488 42096 2552
rect 42160 2488 42176 2552
rect 42240 2488 42256 2552
rect 42320 2488 42336 2552
rect 42400 2488 42416 2552
rect 42480 2488 42496 2552
rect 42560 2488 42576 2552
rect 42640 2488 42656 2552
rect 42720 2488 42736 2552
rect 42800 2488 42816 2552
rect 42880 2488 42896 2552
rect 42960 2488 42976 2552
rect 43040 2488 43056 2552
rect 43120 2488 43136 2552
rect 43200 2488 43216 2552
rect 43280 2488 43296 2552
rect 43360 2488 43376 2552
rect 43440 2488 43456 2552
rect 43520 2488 43536 2552
rect 43600 2488 43616 2552
rect 43680 2488 43696 2552
rect 43760 2488 43776 2552
rect 43840 2488 43856 2552
rect 43920 2488 43936 2552
rect 44000 2488 44016 2552
rect 44080 2488 44096 2552
rect 44160 2488 44176 2552
rect 44240 2488 44256 2552
rect 44320 2488 44336 2552
rect 44400 2488 44416 2552
rect 44480 2488 44496 2552
rect 44560 2488 44576 2552
rect 44640 2488 44656 2552
rect 44720 2488 44736 2552
rect 44800 2488 44816 2552
rect 44880 2488 44896 2552
rect 44960 2488 44976 2552
rect 45040 2488 45056 2552
rect 45120 2488 45136 2552
rect 45200 2488 45216 2552
rect 45280 2488 45296 2552
rect 45360 2488 45368 2552
rect 0 2472 45368 2488
rect 0 2408 8 2472
rect 72 2408 88 2472
rect 152 2408 168 2472
rect 232 2408 248 2472
rect 312 2408 328 2472
rect 392 2408 408 2472
rect 472 2408 488 2472
rect 552 2408 568 2472
rect 632 2408 648 2472
rect 712 2408 728 2472
rect 792 2408 808 2472
rect 872 2408 888 2472
rect 952 2408 968 2472
rect 1032 2408 1048 2472
rect 1112 2408 1128 2472
rect 1192 2408 1208 2472
rect 1272 2408 1288 2472
rect 1352 2408 1368 2472
rect 1432 2408 1448 2472
rect 1512 2408 1528 2472
rect 1592 2408 1608 2472
rect 1672 2408 1688 2472
rect 1752 2408 1768 2472
rect 1832 2408 1848 2472
rect 1912 2408 1928 2472
rect 1992 2408 2008 2472
rect 2072 2408 2088 2472
rect 2152 2408 2168 2472
rect 2232 2408 2248 2472
rect 2312 2408 2328 2472
rect 2392 2408 2408 2472
rect 2472 2408 2488 2472
rect 2552 2408 2568 2472
rect 2632 2408 2648 2472
rect 2712 2408 2728 2472
rect 2792 2408 2808 2472
rect 2872 2408 2888 2472
rect 2952 2408 2968 2472
rect 3032 2408 3048 2472
rect 3112 2408 3128 2472
rect 3192 2408 3208 2472
rect 3272 2408 3288 2472
rect 3352 2408 3368 2472
rect 3432 2408 3448 2472
rect 3512 2408 3528 2472
rect 3592 2408 3608 2472
rect 3672 2408 3688 2472
rect 3752 2408 3768 2472
rect 3832 2408 3848 2472
rect 3912 2408 3928 2472
rect 3992 2408 19112 2472
rect 19176 2408 19192 2472
rect 19256 2408 19272 2472
rect 19336 2408 19352 2472
rect 19416 2408 29112 2472
rect 29176 2408 29192 2472
rect 29256 2408 29272 2472
rect 29336 2408 29352 2472
rect 29416 2408 41376 2472
rect 41440 2408 41456 2472
rect 41520 2408 41536 2472
rect 41600 2408 41616 2472
rect 41680 2408 41696 2472
rect 41760 2408 41776 2472
rect 41840 2408 41856 2472
rect 41920 2408 41936 2472
rect 42000 2408 42016 2472
rect 42080 2408 42096 2472
rect 42160 2408 42176 2472
rect 42240 2408 42256 2472
rect 42320 2408 42336 2472
rect 42400 2408 42416 2472
rect 42480 2408 42496 2472
rect 42560 2408 42576 2472
rect 42640 2408 42656 2472
rect 42720 2408 42736 2472
rect 42800 2408 42816 2472
rect 42880 2408 42896 2472
rect 42960 2408 42976 2472
rect 43040 2408 43056 2472
rect 43120 2408 43136 2472
rect 43200 2408 43216 2472
rect 43280 2408 43296 2472
rect 43360 2408 43376 2472
rect 43440 2408 43456 2472
rect 43520 2408 43536 2472
rect 43600 2408 43616 2472
rect 43680 2408 43696 2472
rect 43760 2408 43776 2472
rect 43840 2408 43856 2472
rect 43920 2408 43936 2472
rect 44000 2408 44016 2472
rect 44080 2408 44096 2472
rect 44160 2408 44176 2472
rect 44240 2408 44256 2472
rect 44320 2408 44336 2472
rect 44400 2408 44416 2472
rect 44480 2408 44496 2472
rect 44560 2408 44576 2472
rect 44640 2408 44656 2472
rect 44720 2408 44736 2472
rect 44800 2408 44816 2472
rect 44880 2408 44896 2472
rect 44960 2408 44976 2472
rect 45040 2408 45056 2472
rect 45120 2408 45136 2472
rect 45200 2408 45216 2472
rect 45280 2408 45296 2472
rect 45360 2408 45368 2472
rect 0 2392 45368 2408
rect 0 2328 8 2392
rect 72 2328 88 2392
rect 152 2328 168 2392
rect 232 2328 248 2392
rect 312 2328 328 2392
rect 392 2328 408 2392
rect 472 2328 488 2392
rect 552 2328 568 2392
rect 632 2328 648 2392
rect 712 2328 728 2392
rect 792 2328 808 2392
rect 872 2328 888 2392
rect 952 2328 968 2392
rect 1032 2328 1048 2392
rect 1112 2328 1128 2392
rect 1192 2328 1208 2392
rect 1272 2328 1288 2392
rect 1352 2328 1368 2392
rect 1432 2328 1448 2392
rect 1512 2328 1528 2392
rect 1592 2328 1608 2392
rect 1672 2328 1688 2392
rect 1752 2328 1768 2392
rect 1832 2328 1848 2392
rect 1912 2328 1928 2392
rect 1992 2328 2008 2392
rect 2072 2328 2088 2392
rect 2152 2328 2168 2392
rect 2232 2328 2248 2392
rect 2312 2328 2328 2392
rect 2392 2328 2408 2392
rect 2472 2328 2488 2392
rect 2552 2328 2568 2392
rect 2632 2328 2648 2392
rect 2712 2328 2728 2392
rect 2792 2328 2808 2392
rect 2872 2328 2888 2392
rect 2952 2328 2968 2392
rect 3032 2328 3048 2392
rect 3112 2328 3128 2392
rect 3192 2328 3208 2392
rect 3272 2328 3288 2392
rect 3352 2328 3368 2392
rect 3432 2328 3448 2392
rect 3512 2328 3528 2392
rect 3592 2328 3608 2392
rect 3672 2328 3688 2392
rect 3752 2328 3768 2392
rect 3832 2328 3848 2392
rect 3912 2328 3928 2392
rect 3992 2328 19112 2392
rect 19176 2328 19192 2392
rect 19256 2328 19272 2392
rect 19336 2328 19352 2392
rect 19416 2328 29112 2392
rect 29176 2328 29192 2392
rect 29256 2328 29272 2392
rect 29336 2328 29352 2392
rect 29416 2328 41376 2392
rect 41440 2328 41456 2392
rect 41520 2328 41536 2392
rect 41600 2328 41616 2392
rect 41680 2328 41696 2392
rect 41760 2328 41776 2392
rect 41840 2328 41856 2392
rect 41920 2328 41936 2392
rect 42000 2328 42016 2392
rect 42080 2328 42096 2392
rect 42160 2328 42176 2392
rect 42240 2328 42256 2392
rect 42320 2328 42336 2392
rect 42400 2328 42416 2392
rect 42480 2328 42496 2392
rect 42560 2328 42576 2392
rect 42640 2328 42656 2392
rect 42720 2328 42736 2392
rect 42800 2328 42816 2392
rect 42880 2328 42896 2392
rect 42960 2328 42976 2392
rect 43040 2328 43056 2392
rect 43120 2328 43136 2392
rect 43200 2328 43216 2392
rect 43280 2328 43296 2392
rect 43360 2328 43376 2392
rect 43440 2328 43456 2392
rect 43520 2328 43536 2392
rect 43600 2328 43616 2392
rect 43680 2328 43696 2392
rect 43760 2328 43776 2392
rect 43840 2328 43856 2392
rect 43920 2328 43936 2392
rect 44000 2328 44016 2392
rect 44080 2328 44096 2392
rect 44160 2328 44176 2392
rect 44240 2328 44256 2392
rect 44320 2328 44336 2392
rect 44400 2328 44416 2392
rect 44480 2328 44496 2392
rect 44560 2328 44576 2392
rect 44640 2328 44656 2392
rect 44720 2328 44736 2392
rect 44800 2328 44816 2392
rect 44880 2328 44896 2392
rect 44960 2328 44976 2392
rect 45040 2328 45056 2392
rect 45120 2328 45136 2392
rect 45200 2328 45216 2392
rect 45280 2328 45296 2392
rect 45360 2328 45368 2392
rect 0 2312 45368 2328
rect 0 2248 8 2312
rect 72 2248 88 2312
rect 152 2248 168 2312
rect 232 2248 248 2312
rect 312 2248 328 2312
rect 392 2248 408 2312
rect 472 2248 488 2312
rect 552 2248 568 2312
rect 632 2248 648 2312
rect 712 2248 728 2312
rect 792 2248 808 2312
rect 872 2248 888 2312
rect 952 2248 968 2312
rect 1032 2248 1048 2312
rect 1112 2248 1128 2312
rect 1192 2248 1208 2312
rect 1272 2248 1288 2312
rect 1352 2248 1368 2312
rect 1432 2248 1448 2312
rect 1512 2248 1528 2312
rect 1592 2248 1608 2312
rect 1672 2248 1688 2312
rect 1752 2248 1768 2312
rect 1832 2248 1848 2312
rect 1912 2248 1928 2312
rect 1992 2248 2008 2312
rect 2072 2248 2088 2312
rect 2152 2248 2168 2312
rect 2232 2248 2248 2312
rect 2312 2248 2328 2312
rect 2392 2248 2408 2312
rect 2472 2248 2488 2312
rect 2552 2248 2568 2312
rect 2632 2248 2648 2312
rect 2712 2248 2728 2312
rect 2792 2248 2808 2312
rect 2872 2248 2888 2312
rect 2952 2248 2968 2312
rect 3032 2248 3048 2312
rect 3112 2248 3128 2312
rect 3192 2248 3208 2312
rect 3272 2248 3288 2312
rect 3352 2248 3368 2312
rect 3432 2248 3448 2312
rect 3512 2248 3528 2312
rect 3592 2248 3608 2312
rect 3672 2248 3688 2312
rect 3752 2248 3768 2312
rect 3832 2248 3848 2312
rect 3912 2248 3928 2312
rect 3992 2248 19112 2312
rect 19176 2248 19192 2312
rect 19256 2248 19272 2312
rect 19336 2248 19352 2312
rect 19416 2248 29112 2312
rect 29176 2248 29192 2312
rect 29256 2248 29272 2312
rect 29336 2248 29352 2312
rect 29416 2248 41376 2312
rect 41440 2248 41456 2312
rect 41520 2248 41536 2312
rect 41600 2248 41616 2312
rect 41680 2248 41696 2312
rect 41760 2248 41776 2312
rect 41840 2248 41856 2312
rect 41920 2248 41936 2312
rect 42000 2248 42016 2312
rect 42080 2248 42096 2312
rect 42160 2248 42176 2312
rect 42240 2248 42256 2312
rect 42320 2248 42336 2312
rect 42400 2248 42416 2312
rect 42480 2248 42496 2312
rect 42560 2248 42576 2312
rect 42640 2248 42656 2312
rect 42720 2248 42736 2312
rect 42800 2248 42816 2312
rect 42880 2248 42896 2312
rect 42960 2248 42976 2312
rect 43040 2248 43056 2312
rect 43120 2248 43136 2312
rect 43200 2248 43216 2312
rect 43280 2248 43296 2312
rect 43360 2248 43376 2312
rect 43440 2248 43456 2312
rect 43520 2248 43536 2312
rect 43600 2248 43616 2312
rect 43680 2248 43696 2312
rect 43760 2248 43776 2312
rect 43840 2248 43856 2312
rect 43920 2248 43936 2312
rect 44000 2248 44016 2312
rect 44080 2248 44096 2312
rect 44160 2248 44176 2312
rect 44240 2248 44256 2312
rect 44320 2248 44336 2312
rect 44400 2248 44416 2312
rect 44480 2248 44496 2312
rect 44560 2248 44576 2312
rect 44640 2248 44656 2312
rect 44720 2248 44736 2312
rect 44800 2248 44816 2312
rect 44880 2248 44896 2312
rect 44960 2248 44976 2312
rect 45040 2248 45056 2312
rect 45120 2248 45136 2312
rect 45200 2248 45216 2312
rect 45280 2248 45296 2312
rect 45360 2248 45368 2312
rect 0 2232 45368 2248
rect 0 2168 8 2232
rect 72 2168 88 2232
rect 152 2168 168 2232
rect 232 2168 248 2232
rect 312 2168 328 2232
rect 392 2168 408 2232
rect 472 2168 488 2232
rect 552 2168 568 2232
rect 632 2168 648 2232
rect 712 2168 728 2232
rect 792 2168 808 2232
rect 872 2168 888 2232
rect 952 2168 968 2232
rect 1032 2168 1048 2232
rect 1112 2168 1128 2232
rect 1192 2168 1208 2232
rect 1272 2168 1288 2232
rect 1352 2168 1368 2232
rect 1432 2168 1448 2232
rect 1512 2168 1528 2232
rect 1592 2168 1608 2232
rect 1672 2168 1688 2232
rect 1752 2168 1768 2232
rect 1832 2168 1848 2232
rect 1912 2168 1928 2232
rect 1992 2168 2008 2232
rect 2072 2168 2088 2232
rect 2152 2168 2168 2232
rect 2232 2168 2248 2232
rect 2312 2168 2328 2232
rect 2392 2168 2408 2232
rect 2472 2168 2488 2232
rect 2552 2168 2568 2232
rect 2632 2168 2648 2232
rect 2712 2168 2728 2232
rect 2792 2168 2808 2232
rect 2872 2168 2888 2232
rect 2952 2168 2968 2232
rect 3032 2168 3048 2232
rect 3112 2168 3128 2232
rect 3192 2168 3208 2232
rect 3272 2168 3288 2232
rect 3352 2168 3368 2232
rect 3432 2168 3448 2232
rect 3512 2168 3528 2232
rect 3592 2168 3608 2232
rect 3672 2168 3688 2232
rect 3752 2168 3768 2232
rect 3832 2168 3848 2232
rect 3912 2168 3928 2232
rect 3992 2168 19112 2232
rect 19176 2168 19192 2232
rect 19256 2168 19272 2232
rect 19336 2168 19352 2232
rect 19416 2168 29112 2232
rect 29176 2168 29192 2232
rect 29256 2168 29272 2232
rect 29336 2168 29352 2232
rect 29416 2168 41376 2232
rect 41440 2168 41456 2232
rect 41520 2168 41536 2232
rect 41600 2168 41616 2232
rect 41680 2168 41696 2232
rect 41760 2168 41776 2232
rect 41840 2168 41856 2232
rect 41920 2168 41936 2232
rect 42000 2168 42016 2232
rect 42080 2168 42096 2232
rect 42160 2168 42176 2232
rect 42240 2168 42256 2232
rect 42320 2168 42336 2232
rect 42400 2168 42416 2232
rect 42480 2168 42496 2232
rect 42560 2168 42576 2232
rect 42640 2168 42656 2232
rect 42720 2168 42736 2232
rect 42800 2168 42816 2232
rect 42880 2168 42896 2232
rect 42960 2168 42976 2232
rect 43040 2168 43056 2232
rect 43120 2168 43136 2232
rect 43200 2168 43216 2232
rect 43280 2168 43296 2232
rect 43360 2168 43376 2232
rect 43440 2168 43456 2232
rect 43520 2168 43536 2232
rect 43600 2168 43616 2232
rect 43680 2168 43696 2232
rect 43760 2168 43776 2232
rect 43840 2168 43856 2232
rect 43920 2168 43936 2232
rect 44000 2168 44016 2232
rect 44080 2168 44096 2232
rect 44160 2168 44176 2232
rect 44240 2168 44256 2232
rect 44320 2168 44336 2232
rect 44400 2168 44416 2232
rect 44480 2168 44496 2232
rect 44560 2168 44576 2232
rect 44640 2168 44656 2232
rect 44720 2168 44736 2232
rect 44800 2168 44816 2232
rect 44880 2168 44896 2232
rect 44960 2168 44976 2232
rect 45040 2168 45056 2232
rect 45120 2168 45136 2232
rect 45200 2168 45216 2232
rect 45280 2168 45296 2232
rect 45360 2168 45368 2232
rect 0 2152 45368 2168
rect 0 2088 8 2152
rect 72 2088 88 2152
rect 152 2088 168 2152
rect 232 2088 248 2152
rect 312 2088 328 2152
rect 392 2088 408 2152
rect 472 2088 488 2152
rect 552 2088 568 2152
rect 632 2088 648 2152
rect 712 2088 728 2152
rect 792 2088 808 2152
rect 872 2088 888 2152
rect 952 2088 968 2152
rect 1032 2088 1048 2152
rect 1112 2088 1128 2152
rect 1192 2088 1208 2152
rect 1272 2088 1288 2152
rect 1352 2088 1368 2152
rect 1432 2088 1448 2152
rect 1512 2088 1528 2152
rect 1592 2088 1608 2152
rect 1672 2088 1688 2152
rect 1752 2088 1768 2152
rect 1832 2088 1848 2152
rect 1912 2088 1928 2152
rect 1992 2088 2008 2152
rect 2072 2088 2088 2152
rect 2152 2088 2168 2152
rect 2232 2088 2248 2152
rect 2312 2088 2328 2152
rect 2392 2088 2408 2152
rect 2472 2088 2488 2152
rect 2552 2088 2568 2152
rect 2632 2088 2648 2152
rect 2712 2088 2728 2152
rect 2792 2088 2808 2152
rect 2872 2088 2888 2152
rect 2952 2088 2968 2152
rect 3032 2088 3048 2152
rect 3112 2088 3128 2152
rect 3192 2088 3208 2152
rect 3272 2088 3288 2152
rect 3352 2088 3368 2152
rect 3432 2088 3448 2152
rect 3512 2088 3528 2152
rect 3592 2088 3608 2152
rect 3672 2088 3688 2152
rect 3752 2088 3768 2152
rect 3832 2088 3848 2152
rect 3912 2088 3928 2152
rect 3992 2088 19112 2152
rect 19176 2088 19192 2152
rect 19256 2088 19272 2152
rect 19336 2088 19352 2152
rect 19416 2088 29112 2152
rect 29176 2088 29192 2152
rect 29256 2088 29272 2152
rect 29336 2088 29352 2152
rect 29416 2088 41376 2152
rect 41440 2088 41456 2152
rect 41520 2088 41536 2152
rect 41600 2088 41616 2152
rect 41680 2088 41696 2152
rect 41760 2088 41776 2152
rect 41840 2088 41856 2152
rect 41920 2088 41936 2152
rect 42000 2088 42016 2152
rect 42080 2088 42096 2152
rect 42160 2088 42176 2152
rect 42240 2088 42256 2152
rect 42320 2088 42336 2152
rect 42400 2088 42416 2152
rect 42480 2088 42496 2152
rect 42560 2088 42576 2152
rect 42640 2088 42656 2152
rect 42720 2088 42736 2152
rect 42800 2088 42816 2152
rect 42880 2088 42896 2152
rect 42960 2088 42976 2152
rect 43040 2088 43056 2152
rect 43120 2088 43136 2152
rect 43200 2088 43216 2152
rect 43280 2088 43296 2152
rect 43360 2088 43376 2152
rect 43440 2088 43456 2152
rect 43520 2088 43536 2152
rect 43600 2088 43616 2152
rect 43680 2088 43696 2152
rect 43760 2088 43776 2152
rect 43840 2088 43856 2152
rect 43920 2088 43936 2152
rect 44000 2088 44016 2152
rect 44080 2088 44096 2152
rect 44160 2088 44176 2152
rect 44240 2088 44256 2152
rect 44320 2088 44336 2152
rect 44400 2088 44416 2152
rect 44480 2088 44496 2152
rect 44560 2088 44576 2152
rect 44640 2088 44656 2152
rect 44720 2088 44736 2152
rect 44800 2088 44816 2152
rect 44880 2088 44896 2152
rect 44960 2088 44976 2152
rect 45040 2088 45056 2152
rect 45120 2088 45136 2152
rect 45200 2088 45216 2152
rect 45280 2088 45296 2152
rect 45360 2088 45368 2152
rect 0 2072 45368 2088
rect 0 2008 8 2072
rect 72 2008 88 2072
rect 152 2008 168 2072
rect 232 2008 248 2072
rect 312 2008 328 2072
rect 392 2008 408 2072
rect 472 2008 488 2072
rect 552 2008 568 2072
rect 632 2008 648 2072
rect 712 2008 728 2072
rect 792 2008 808 2072
rect 872 2008 888 2072
rect 952 2008 968 2072
rect 1032 2008 1048 2072
rect 1112 2008 1128 2072
rect 1192 2008 1208 2072
rect 1272 2008 1288 2072
rect 1352 2008 1368 2072
rect 1432 2008 1448 2072
rect 1512 2008 1528 2072
rect 1592 2008 1608 2072
rect 1672 2008 1688 2072
rect 1752 2008 1768 2072
rect 1832 2008 1848 2072
rect 1912 2008 1928 2072
rect 1992 2008 2008 2072
rect 2072 2008 2088 2072
rect 2152 2008 2168 2072
rect 2232 2008 2248 2072
rect 2312 2008 2328 2072
rect 2392 2008 2408 2072
rect 2472 2008 2488 2072
rect 2552 2008 2568 2072
rect 2632 2008 2648 2072
rect 2712 2008 2728 2072
rect 2792 2008 2808 2072
rect 2872 2008 2888 2072
rect 2952 2008 2968 2072
rect 3032 2008 3048 2072
rect 3112 2008 3128 2072
rect 3192 2008 3208 2072
rect 3272 2008 3288 2072
rect 3352 2008 3368 2072
rect 3432 2008 3448 2072
rect 3512 2008 3528 2072
rect 3592 2008 3608 2072
rect 3672 2008 3688 2072
rect 3752 2008 3768 2072
rect 3832 2008 3848 2072
rect 3912 2008 3928 2072
rect 3992 2008 19112 2072
rect 19176 2008 19192 2072
rect 19256 2008 19272 2072
rect 19336 2008 19352 2072
rect 19416 2008 29112 2072
rect 29176 2008 29192 2072
rect 29256 2008 29272 2072
rect 29336 2008 29352 2072
rect 29416 2008 41376 2072
rect 41440 2008 41456 2072
rect 41520 2008 41536 2072
rect 41600 2008 41616 2072
rect 41680 2008 41696 2072
rect 41760 2008 41776 2072
rect 41840 2008 41856 2072
rect 41920 2008 41936 2072
rect 42000 2008 42016 2072
rect 42080 2008 42096 2072
rect 42160 2008 42176 2072
rect 42240 2008 42256 2072
rect 42320 2008 42336 2072
rect 42400 2008 42416 2072
rect 42480 2008 42496 2072
rect 42560 2008 42576 2072
rect 42640 2008 42656 2072
rect 42720 2008 42736 2072
rect 42800 2008 42816 2072
rect 42880 2008 42896 2072
rect 42960 2008 42976 2072
rect 43040 2008 43056 2072
rect 43120 2008 43136 2072
rect 43200 2008 43216 2072
rect 43280 2008 43296 2072
rect 43360 2008 43376 2072
rect 43440 2008 43456 2072
rect 43520 2008 43536 2072
rect 43600 2008 43616 2072
rect 43680 2008 43696 2072
rect 43760 2008 43776 2072
rect 43840 2008 43856 2072
rect 43920 2008 43936 2072
rect 44000 2008 44016 2072
rect 44080 2008 44096 2072
rect 44160 2008 44176 2072
rect 44240 2008 44256 2072
rect 44320 2008 44336 2072
rect 44400 2008 44416 2072
rect 44480 2008 44496 2072
rect 44560 2008 44576 2072
rect 44640 2008 44656 2072
rect 44720 2008 44736 2072
rect 44800 2008 44816 2072
rect 44880 2008 44896 2072
rect 44960 2008 44976 2072
rect 45040 2008 45056 2072
rect 45120 2008 45136 2072
rect 45200 2008 45216 2072
rect 45280 2008 45296 2072
rect 45360 2008 45368 2072
rect 0 1992 45368 2008
rect 0 1928 8 1992
rect 72 1928 88 1992
rect 152 1928 168 1992
rect 232 1928 248 1992
rect 312 1928 328 1992
rect 392 1928 408 1992
rect 472 1928 488 1992
rect 552 1928 568 1992
rect 632 1928 648 1992
rect 712 1928 728 1992
rect 792 1928 808 1992
rect 872 1928 888 1992
rect 952 1928 968 1992
rect 1032 1928 1048 1992
rect 1112 1928 1128 1992
rect 1192 1928 1208 1992
rect 1272 1928 1288 1992
rect 1352 1928 1368 1992
rect 1432 1928 1448 1992
rect 1512 1928 1528 1992
rect 1592 1928 1608 1992
rect 1672 1928 1688 1992
rect 1752 1928 1768 1992
rect 1832 1928 1848 1992
rect 1912 1928 1928 1992
rect 1992 1928 2008 1992
rect 2072 1928 2088 1992
rect 2152 1928 2168 1992
rect 2232 1928 2248 1992
rect 2312 1928 2328 1992
rect 2392 1928 2408 1992
rect 2472 1928 2488 1992
rect 2552 1928 2568 1992
rect 2632 1928 2648 1992
rect 2712 1928 2728 1992
rect 2792 1928 2808 1992
rect 2872 1928 2888 1992
rect 2952 1928 2968 1992
rect 3032 1928 3048 1992
rect 3112 1928 3128 1992
rect 3192 1928 3208 1992
rect 3272 1928 3288 1992
rect 3352 1928 3368 1992
rect 3432 1928 3448 1992
rect 3512 1928 3528 1992
rect 3592 1928 3608 1992
rect 3672 1928 3688 1992
rect 3752 1928 3768 1992
rect 3832 1928 3848 1992
rect 3912 1928 3928 1992
rect 3992 1928 19112 1992
rect 19176 1928 19192 1992
rect 19256 1928 19272 1992
rect 19336 1928 19352 1992
rect 19416 1928 29112 1992
rect 29176 1928 29192 1992
rect 29256 1928 29272 1992
rect 29336 1928 29352 1992
rect 29416 1928 41376 1992
rect 41440 1928 41456 1992
rect 41520 1928 41536 1992
rect 41600 1928 41616 1992
rect 41680 1928 41696 1992
rect 41760 1928 41776 1992
rect 41840 1928 41856 1992
rect 41920 1928 41936 1992
rect 42000 1928 42016 1992
rect 42080 1928 42096 1992
rect 42160 1928 42176 1992
rect 42240 1928 42256 1992
rect 42320 1928 42336 1992
rect 42400 1928 42416 1992
rect 42480 1928 42496 1992
rect 42560 1928 42576 1992
rect 42640 1928 42656 1992
rect 42720 1928 42736 1992
rect 42800 1928 42816 1992
rect 42880 1928 42896 1992
rect 42960 1928 42976 1992
rect 43040 1928 43056 1992
rect 43120 1928 43136 1992
rect 43200 1928 43216 1992
rect 43280 1928 43296 1992
rect 43360 1928 43376 1992
rect 43440 1928 43456 1992
rect 43520 1928 43536 1992
rect 43600 1928 43616 1992
rect 43680 1928 43696 1992
rect 43760 1928 43776 1992
rect 43840 1928 43856 1992
rect 43920 1928 43936 1992
rect 44000 1928 44016 1992
rect 44080 1928 44096 1992
rect 44160 1928 44176 1992
rect 44240 1928 44256 1992
rect 44320 1928 44336 1992
rect 44400 1928 44416 1992
rect 44480 1928 44496 1992
rect 44560 1928 44576 1992
rect 44640 1928 44656 1992
rect 44720 1928 44736 1992
rect 44800 1928 44816 1992
rect 44880 1928 44896 1992
rect 44960 1928 44976 1992
rect 45040 1928 45056 1992
rect 45120 1928 45136 1992
rect 45200 1928 45216 1992
rect 45280 1928 45296 1992
rect 45360 1928 45368 1992
rect 0 1912 45368 1928
rect 0 1848 8 1912
rect 72 1848 88 1912
rect 152 1848 168 1912
rect 232 1848 248 1912
rect 312 1848 328 1912
rect 392 1848 408 1912
rect 472 1848 488 1912
rect 552 1848 568 1912
rect 632 1848 648 1912
rect 712 1848 728 1912
rect 792 1848 808 1912
rect 872 1848 888 1912
rect 952 1848 968 1912
rect 1032 1848 1048 1912
rect 1112 1848 1128 1912
rect 1192 1848 1208 1912
rect 1272 1848 1288 1912
rect 1352 1848 1368 1912
rect 1432 1848 1448 1912
rect 1512 1848 1528 1912
rect 1592 1848 1608 1912
rect 1672 1848 1688 1912
rect 1752 1848 1768 1912
rect 1832 1848 1848 1912
rect 1912 1848 1928 1912
rect 1992 1848 2008 1912
rect 2072 1848 2088 1912
rect 2152 1848 2168 1912
rect 2232 1848 2248 1912
rect 2312 1848 2328 1912
rect 2392 1848 2408 1912
rect 2472 1848 2488 1912
rect 2552 1848 2568 1912
rect 2632 1848 2648 1912
rect 2712 1848 2728 1912
rect 2792 1848 2808 1912
rect 2872 1848 2888 1912
rect 2952 1848 2968 1912
rect 3032 1848 3048 1912
rect 3112 1848 3128 1912
rect 3192 1848 3208 1912
rect 3272 1848 3288 1912
rect 3352 1848 3368 1912
rect 3432 1848 3448 1912
rect 3512 1848 3528 1912
rect 3592 1848 3608 1912
rect 3672 1848 3688 1912
rect 3752 1848 3768 1912
rect 3832 1848 3848 1912
rect 3912 1848 3928 1912
rect 3992 1848 19112 1912
rect 19176 1848 19192 1912
rect 19256 1848 19272 1912
rect 19336 1848 19352 1912
rect 19416 1848 29112 1912
rect 29176 1848 29192 1912
rect 29256 1848 29272 1912
rect 29336 1848 29352 1912
rect 29416 1848 41376 1912
rect 41440 1848 41456 1912
rect 41520 1848 41536 1912
rect 41600 1848 41616 1912
rect 41680 1848 41696 1912
rect 41760 1848 41776 1912
rect 41840 1848 41856 1912
rect 41920 1848 41936 1912
rect 42000 1848 42016 1912
rect 42080 1848 42096 1912
rect 42160 1848 42176 1912
rect 42240 1848 42256 1912
rect 42320 1848 42336 1912
rect 42400 1848 42416 1912
rect 42480 1848 42496 1912
rect 42560 1848 42576 1912
rect 42640 1848 42656 1912
rect 42720 1848 42736 1912
rect 42800 1848 42816 1912
rect 42880 1848 42896 1912
rect 42960 1848 42976 1912
rect 43040 1848 43056 1912
rect 43120 1848 43136 1912
rect 43200 1848 43216 1912
rect 43280 1848 43296 1912
rect 43360 1848 43376 1912
rect 43440 1848 43456 1912
rect 43520 1848 43536 1912
rect 43600 1848 43616 1912
rect 43680 1848 43696 1912
rect 43760 1848 43776 1912
rect 43840 1848 43856 1912
rect 43920 1848 43936 1912
rect 44000 1848 44016 1912
rect 44080 1848 44096 1912
rect 44160 1848 44176 1912
rect 44240 1848 44256 1912
rect 44320 1848 44336 1912
rect 44400 1848 44416 1912
rect 44480 1848 44496 1912
rect 44560 1848 44576 1912
rect 44640 1848 44656 1912
rect 44720 1848 44736 1912
rect 44800 1848 44816 1912
rect 44880 1848 44896 1912
rect 44960 1848 44976 1912
rect 45040 1848 45056 1912
rect 45120 1848 45136 1912
rect 45200 1848 45216 1912
rect 45280 1848 45296 1912
rect 45360 1848 45368 1912
rect 0 1832 45368 1848
rect 0 1768 8 1832
rect 72 1768 88 1832
rect 152 1768 168 1832
rect 232 1768 248 1832
rect 312 1768 328 1832
rect 392 1768 408 1832
rect 472 1768 488 1832
rect 552 1768 568 1832
rect 632 1768 648 1832
rect 712 1768 728 1832
rect 792 1768 808 1832
rect 872 1768 888 1832
rect 952 1768 968 1832
rect 1032 1768 1048 1832
rect 1112 1768 1128 1832
rect 1192 1768 1208 1832
rect 1272 1768 1288 1832
rect 1352 1768 1368 1832
rect 1432 1768 1448 1832
rect 1512 1768 1528 1832
rect 1592 1768 1608 1832
rect 1672 1768 1688 1832
rect 1752 1768 1768 1832
rect 1832 1768 1848 1832
rect 1912 1768 1928 1832
rect 1992 1768 2008 1832
rect 2072 1768 2088 1832
rect 2152 1768 2168 1832
rect 2232 1768 2248 1832
rect 2312 1768 2328 1832
rect 2392 1768 2408 1832
rect 2472 1768 2488 1832
rect 2552 1768 2568 1832
rect 2632 1768 2648 1832
rect 2712 1768 2728 1832
rect 2792 1768 2808 1832
rect 2872 1768 2888 1832
rect 2952 1768 2968 1832
rect 3032 1768 3048 1832
rect 3112 1768 3128 1832
rect 3192 1768 3208 1832
rect 3272 1768 3288 1832
rect 3352 1768 3368 1832
rect 3432 1768 3448 1832
rect 3512 1768 3528 1832
rect 3592 1768 3608 1832
rect 3672 1768 3688 1832
rect 3752 1768 3768 1832
rect 3832 1768 3848 1832
rect 3912 1768 3928 1832
rect 3992 1768 19112 1832
rect 19176 1768 19192 1832
rect 19256 1768 19272 1832
rect 19336 1768 19352 1832
rect 19416 1768 29112 1832
rect 29176 1768 29192 1832
rect 29256 1768 29272 1832
rect 29336 1768 29352 1832
rect 29416 1768 41376 1832
rect 41440 1768 41456 1832
rect 41520 1768 41536 1832
rect 41600 1768 41616 1832
rect 41680 1768 41696 1832
rect 41760 1768 41776 1832
rect 41840 1768 41856 1832
rect 41920 1768 41936 1832
rect 42000 1768 42016 1832
rect 42080 1768 42096 1832
rect 42160 1768 42176 1832
rect 42240 1768 42256 1832
rect 42320 1768 42336 1832
rect 42400 1768 42416 1832
rect 42480 1768 42496 1832
rect 42560 1768 42576 1832
rect 42640 1768 42656 1832
rect 42720 1768 42736 1832
rect 42800 1768 42816 1832
rect 42880 1768 42896 1832
rect 42960 1768 42976 1832
rect 43040 1768 43056 1832
rect 43120 1768 43136 1832
rect 43200 1768 43216 1832
rect 43280 1768 43296 1832
rect 43360 1768 43376 1832
rect 43440 1768 43456 1832
rect 43520 1768 43536 1832
rect 43600 1768 43616 1832
rect 43680 1768 43696 1832
rect 43760 1768 43776 1832
rect 43840 1768 43856 1832
rect 43920 1768 43936 1832
rect 44000 1768 44016 1832
rect 44080 1768 44096 1832
rect 44160 1768 44176 1832
rect 44240 1768 44256 1832
rect 44320 1768 44336 1832
rect 44400 1768 44416 1832
rect 44480 1768 44496 1832
rect 44560 1768 44576 1832
rect 44640 1768 44656 1832
rect 44720 1768 44736 1832
rect 44800 1768 44816 1832
rect 44880 1768 44896 1832
rect 44960 1768 44976 1832
rect 45040 1768 45056 1832
rect 45120 1768 45136 1832
rect 45200 1768 45216 1832
rect 45280 1768 45296 1832
rect 45360 1768 45368 1832
rect 0 1752 45368 1768
rect 0 1688 8 1752
rect 72 1688 88 1752
rect 152 1688 168 1752
rect 232 1688 248 1752
rect 312 1688 328 1752
rect 392 1688 408 1752
rect 472 1688 488 1752
rect 552 1688 568 1752
rect 632 1688 648 1752
rect 712 1688 728 1752
rect 792 1688 808 1752
rect 872 1688 888 1752
rect 952 1688 968 1752
rect 1032 1688 1048 1752
rect 1112 1688 1128 1752
rect 1192 1688 1208 1752
rect 1272 1688 1288 1752
rect 1352 1688 1368 1752
rect 1432 1688 1448 1752
rect 1512 1688 1528 1752
rect 1592 1688 1608 1752
rect 1672 1688 1688 1752
rect 1752 1688 1768 1752
rect 1832 1688 1848 1752
rect 1912 1688 1928 1752
rect 1992 1688 2008 1752
rect 2072 1688 2088 1752
rect 2152 1688 2168 1752
rect 2232 1688 2248 1752
rect 2312 1688 2328 1752
rect 2392 1688 2408 1752
rect 2472 1688 2488 1752
rect 2552 1688 2568 1752
rect 2632 1688 2648 1752
rect 2712 1688 2728 1752
rect 2792 1688 2808 1752
rect 2872 1688 2888 1752
rect 2952 1688 2968 1752
rect 3032 1688 3048 1752
rect 3112 1688 3128 1752
rect 3192 1688 3208 1752
rect 3272 1688 3288 1752
rect 3352 1688 3368 1752
rect 3432 1688 3448 1752
rect 3512 1688 3528 1752
rect 3592 1688 3608 1752
rect 3672 1688 3688 1752
rect 3752 1688 3768 1752
rect 3832 1688 3848 1752
rect 3912 1688 3928 1752
rect 3992 1688 19112 1752
rect 19176 1688 19192 1752
rect 19256 1688 19272 1752
rect 19336 1688 19352 1752
rect 19416 1688 29112 1752
rect 29176 1688 29192 1752
rect 29256 1688 29272 1752
rect 29336 1688 29352 1752
rect 29416 1688 41376 1752
rect 41440 1688 41456 1752
rect 41520 1688 41536 1752
rect 41600 1688 41616 1752
rect 41680 1688 41696 1752
rect 41760 1688 41776 1752
rect 41840 1688 41856 1752
rect 41920 1688 41936 1752
rect 42000 1688 42016 1752
rect 42080 1688 42096 1752
rect 42160 1688 42176 1752
rect 42240 1688 42256 1752
rect 42320 1688 42336 1752
rect 42400 1688 42416 1752
rect 42480 1688 42496 1752
rect 42560 1688 42576 1752
rect 42640 1688 42656 1752
rect 42720 1688 42736 1752
rect 42800 1688 42816 1752
rect 42880 1688 42896 1752
rect 42960 1688 42976 1752
rect 43040 1688 43056 1752
rect 43120 1688 43136 1752
rect 43200 1688 43216 1752
rect 43280 1688 43296 1752
rect 43360 1688 43376 1752
rect 43440 1688 43456 1752
rect 43520 1688 43536 1752
rect 43600 1688 43616 1752
rect 43680 1688 43696 1752
rect 43760 1688 43776 1752
rect 43840 1688 43856 1752
rect 43920 1688 43936 1752
rect 44000 1688 44016 1752
rect 44080 1688 44096 1752
rect 44160 1688 44176 1752
rect 44240 1688 44256 1752
rect 44320 1688 44336 1752
rect 44400 1688 44416 1752
rect 44480 1688 44496 1752
rect 44560 1688 44576 1752
rect 44640 1688 44656 1752
rect 44720 1688 44736 1752
rect 44800 1688 44816 1752
rect 44880 1688 44896 1752
rect 44960 1688 44976 1752
rect 45040 1688 45056 1752
rect 45120 1688 45136 1752
rect 45200 1688 45216 1752
rect 45280 1688 45296 1752
rect 45360 1688 45368 1752
rect 0 1672 45368 1688
rect 0 1608 8 1672
rect 72 1608 88 1672
rect 152 1608 168 1672
rect 232 1608 248 1672
rect 312 1608 328 1672
rect 392 1608 408 1672
rect 472 1608 488 1672
rect 552 1608 568 1672
rect 632 1608 648 1672
rect 712 1608 728 1672
rect 792 1608 808 1672
rect 872 1608 888 1672
rect 952 1608 968 1672
rect 1032 1608 1048 1672
rect 1112 1608 1128 1672
rect 1192 1608 1208 1672
rect 1272 1608 1288 1672
rect 1352 1608 1368 1672
rect 1432 1608 1448 1672
rect 1512 1608 1528 1672
rect 1592 1608 1608 1672
rect 1672 1608 1688 1672
rect 1752 1608 1768 1672
rect 1832 1608 1848 1672
rect 1912 1608 1928 1672
rect 1992 1608 2008 1672
rect 2072 1608 2088 1672
rect 2152 1608 2168 1672
rect 2232 1608 2248 1672
rect 2312 1608 2328 1672
rect 2392 1608 2408 1672
rect 2472 1608 2488 1672
rect 2552 1608 2568 1672
rect 2632 1608 2648 1672
rect 2712 1608 2728 1672
rect 2792 1608 2808 1672
rect 2872 1608 2888 1672
rect 2952 1608 2968 1672
rect 3032 1608 3048 1672
rect 3112 1608 3128 1672
rect 3192 1608 3208 1672
rect 3272 1608 3288 1672
rect 3352 1608 3368 1672
rect 3432 1608 3448 1672
rect 3512 1608 3528 1672
rect 3592 1608 3608 1672
rect 3672 1608 3688 1672
rect 3752 1608 3768 1672
rect 3832 1608 3848 1672
rect 3912 1608 3928 1672
rect 3992 1608 19112 1672
rect 19176 1608 19192 1672
rect 19256 1608 19272 1672
rect 19336 1608 19352 1672
rect 19416 1608 29112 1672
rect 29176 1608 29192 1672
rect 29256 1608 29272 1672
rect 29336 1608 29352 1672
rect 29416 1608 41376 1672
rect 41440 1608 41456 1672
rect 41520 1608 41536 1672
rect 41600 1608 41616 1672
rect 41680 1608 41696 1672
rect 41760 1608 41776 1672
rect 41840 1608 41856 1672
rect 41920 1608 41936 1672
rect 42000 1608 42016 1672
rect 42080 1608 42096 1672
rect 42160 1608 42176 1672
rect 42240 1608 42256 1672
rect 42320 1608 42336 1672
rect 42400 1608 42416 1672
rect 42480 1608 42496 1672
rect 42560 1608 42576 1672
rect 42640 1608 42656 1672
rect 42720 1608 42736 1672
rect 42800 1608 42816 1672
rect 42880 1608 42896 1672
rect 42960 1608 42976 1672
rect 43040 1608 43056 1672
rect 43120 1608 43136 1672
rect 43200 1608 43216 1672
rect 43280 1608 43296 1672
rect 43360 1608 43376 1672
rect 43440 1608 43456 1672
rect 43520 1608 43536 1672
rect 43600 1608 43616 1672
rect 43680 1608 43696 1672
rect 43760 1608 43776 1672
rect 43840 1608 43856 1672
rect 43920 1608 43936 1672
rect 44000 1608 44016 1672
rect 44080 1608 44096 1672
rect 44160 1608 44176 1672
rect 44240 1608 44256 1672
rect 44320 1608 44336 1672
rect 44400 1608 44416 1672
rect 44480 1608 44496 1672
rect 44560 1608 44576 1672
rect 44640 1608 44656 1672
rect 44720 1608 44736 1672
rect 44800 1608 44816 1672
rect 44880 1608 44896 1672
rect 44960 1608 44976 1672
rect 45040 1608 45056 1672
rect 45120 1608 45136 1672
rect 45200 1608 45216 1672
rect 45280 1608 45296 1672
rect 45360 1608 45368 1672
rect 0 1592 45368 1608
rect 0 1528 8 1592
rect 72 1528 88 1592
rect 152 1528 168 1592
rect 232 1528 248 1592
rect 312 1528 328 1592
rect 392 1528 408 1592
rect 472 1528 488 1592
rect 552 1528 568 1592
rect 632 1528 648 1592
rect 712 1528 728 1592
rect 792 1528 808 1592
rect 872 1528 888 1592
rect 952 1528 968 1592
rect 1032 1528 1048 1592
rect 1112 1528 1128 1592
rect 1192 1528 1208 1592
rect 1272 1528 1288 1592
rect 1352 1528 1368 1592
rect 1432 1528 1448 1592
rect 1512 1528 1528 1592
rect 1592 1528 1608 1592
rect 1672 1528 1688 1592
rect 1752 1528 1768 1592
rect 1832 1528 1848 1592
rect 1912 1528 1928 1592
rect 1992 1528 2008 1592
rect 2072 1528 2088 1592
rect 2152 1528 2168 1592
rect 2232 1528 2248 1592
rect 2312 1528 2328 1592
rect 2392 1528 2408 1592
rect 2472 1528 2488 1592
rect 2552 1528 2568 1592
rect 2632 1528 2648 1592
rect 2712 1528 2728 1592
rect 2792 1528 2808 1592
rect 2872 1528 2888 1592
rect 2952 1528 2968 1592
rect 3032 1528 3048 1592
rect 3112 1528 3128 1592
rect 3192 1528 3208 1592
rect 3272 1528 3288 1592
rect 3352 1528 3368 1592
rect 3432 1528 3448 1592
rect 3512 1528 3528 1592
rect 3592 1528 3608 1592
rect 3672 1528 3688 1592
rect 3752 1528 3768 1592
rect 3832 1528 3848 1592
rect 3912 1528 3928 1592
rect 3992 1528 19112 1592
rect 19176 1528 19192 1592
rect 19256 1528 19272 1592
rect 19336 1528 19352 1592
rect 19416 1528 29112 1592
rect 29176 1528 29192 1592
rect 29256 1528 29272 1592
rect 29336 1528 29352 1592
rect 29416 1528 41376 1592
rect 41440 1528 41456 1592
rect 41520 1528 41536 1592
rect 41600 1528 41616 1592
rect 41680 1528 41696 1592
rect 41760 1528 41776 1592
rect 41840 1528 41856 1592
rect 41920 1528 41936 1592
rect 42000 1528 42016 1592
rect 42080 1528 42096 1592
rect 42160 1528 42176 1592
rect 42240 1528 42256 1592
rect 42320 1528 42336 1592
rect 42400 1528 42416 1592
rect 42480 1528 42496 1592
rect 42560 1528 42576 1592
rect 42640 1528 42656 1592
rect 42720 1528 42736 1592
rect 42800 1528 42816 1592
rect 42880 1528 42896 1592
rect 42960 1528 42976 1592
rect 43040 1528 43056 1592
rect 43120 1528 43136 1592
rect 43200 1528 43216 1592
rect 43280 1528 43296 1592
rect 43360 1528 43376 1592
rect 43440 1528 43456 1592
rect 43520 1528 43536 1592
rect 43600 1528 43616 1592
rect 43680 1528 43696 1592
rect 43760 1528 43776 1592
rect 43840 1528 43856 1592
rect 43920 1528 43936 1592
rect 44000 1528 44016 1592
rect 44080 1528 44096 1592
rect 44160 1528 44176 1592
rect 44240 1528 44256 1592
rect 44320 1528 44336 1592
rect 44400 1528 44416 1592
rect 44480 1528 44496 1592
rect 44560 1528 44576 1592
rect 44640 1528 44656 1592
rect 44720 1528 44736 1592
rect 44800 1528 44816 1592
rect 44880 1528 44896 1592
rect 44960 1528 44976 1592
rect 45040 1528 45056 1592
rect 45120 1528 45136 1592
rect 45200 1528 45216 1592
rect 45280 1528 45296 1592
rect 45360 1528 45368 1592
rect 0 1512 45368 1528
rect 0 1448 8 1512
rect 72 1448 88 1512
rect 152 1448 168 1512
rect 232 1448 248 1512
rect 312 1448 328 1512
rect 392 1448 408 1512
rect 472 1448 488 1512
rect 552 1448 568 1512
rect 632 1448 648 1512
rect 712 1448 728 1512
rect 792 1448 808 1512
rect 872 1448 888 1512
rect 952 1448 968 1512
rect 1032 1448 1048 1512
rect 1112 1448 1128 1512
rect 1192 1448 1208 1512
rect 1272 1448 1288 1512
rect 1352 1448 1368 1512
rect 1432 1448 1448 1512
rect 1512 1448 1528 1512
rect 1592 1448 1608 1512
rect 1672 1448 1688 1512
rect 1752 1448 1768 1512
rect 1832 1448 1848 1512
rect 1912 1448 1928 1512
rect 1992 1448 2008 1512
rect 2072 1448 2088 1512
rect 2152 1448 2168 1512
rect 2232 1448 2248 1512
rect 2312 1448 2328 1512
rect 2392 1448 2408 1512
rect 2472 1448 2488 1512
rect 2552 1448 2568 1512
rect 2632 1448 2648 1512
rect 2712 1448 2728 1512
rect 2792 1448 2808 1512
rect 2872 1448 2888 1512
rect 2952 1448 2968 1512
rect 3032 1448 3048 1512
rect 3112 1448 3128 1512
rect 3192 1448 3208 1512
rect 3272 1448 3288 1512
rect 3352 1448 3368 1512
rect 3432 1448 3448 1512
rect 3512 1448 3528 1512
rect 3592 1448 3608 1512
rect 3672 1448 3688 1512
rect 3752 1448 3768 1512
rect 3832 1448 3848 1512
rect 3912 1448 3928 1512
rect 3992 1448 19112 1512
rect 19176 1448 19192 1512
rect 19256 1448 19272 1512
rect 19336 1448 19352 1512
rect 19416 1448 29112 1512
rect 29176 1448 29192 1512
rect 29256 1448 29272 1512
rect 29336 1448 29352 1512
rect 29416 1448 41376 1512
rect 41440 1448 41456 1512
rect 41520 1448 41536 1512
rect 41600 1448 41616 1512
rect 41680 1448 41696 1512
rect 41760 1448 41776 1512
rect 41840 1448 41856 1512
rect 41920 1448 41936 1512
rect 42000 1448 42016 1512
rect 42080 1448 42096 1512
rect 42160 1448 42176 1512
rect 42240 1448 42256 1512
rect 42320 1448 42336 1512
rect 42400 1448 42416 1512
rect 42480 1448 42496 1512
rect 42560 1448 42576 1512
rect 42640 1448 42656 1512
rect 42720 1448 42736 1512
rect 42800 1448 42816 1512
rect 42880 1448 42896 1512
rect 42960 1448 42976 1512
rect 43040 1448 43056 1512
rect 43120 1448 43136 1512
rect 43200 1448 43216 1512
rect 43280 1448 43296 1512
rect 43360 1448 43376 1512
rect 43440 1448 43456 1512
rect 43520 1448 43536 1512
rect 43600 1448 43616 1512
rect 43680 1448 43696 1512
rect 43760 1448 43776 1512
rect 43840 1448 43856 1512
rect 43920 1448 43936 1512
rect 44000 1448 44016 1512
rect 44080 1448 44096 1512
rect 44160 1448 44176 1512
rect 44240 1448 44256 1512
rect 44320 1448 44336 1512
rect 44400 1448 44416 1512
rect 44480 1448 44496 1512
rect 44560 1448 44576 1512
rect 44640 1448 44656 1512
rect 44720 1448 44736 1512
rect 44800 1448 44816 1512
rect 44880 1448 44896 1512
rect 44960 1448 44976 1512
rect 45040 1448 45056 1512
rect 45120 1448 45136 1512
rect 45200 1448 45216 1512
rect 45280 1448 45296 1512
rect 45360 1448 45368 1512
rect 0 1432 45368 1448
rect 0 1368 8 1432
rect 72 1368 88 1432
rect 152 1368 168 1432
rect 232 1368 248 1432
rect 312 1368 328 1432
rect 392 1368 408 1432
rect 472 1368 488 1432
rect 552 1368 568 1432
rect 632 1368 648 1432
rect 712 1368 728 1432
rect 792 1368 808 1432
rect 872 1368 888 1432
rect 952 1368 968 1432
rect 1032 1368 1048 1432
rect 1112 1368 1128 1432
rect 1192 1368 1208 1432
rect 1272 1368 1288 1432
rect 1352 1368 1368 1432
rect 1432 1368 1448 1432
rect 1512 1368 1528 1432
rect 1592 1368 1608 1432
rect 1672 1368 1688 1432
rect 1752 1368 1768 1432
rect 1832 1368 1848 1432
rect 1912 1368 1928 1432
rect 1992 1368 2008 1432
rect 2072 1368 2088 1432
rect 2152 1368 2168 1432
rect 2232 1368 2248 1432
rect 2312 1368 2328 1432
rect 2392 1368 2408 1432
rect 2472 1368 2488 1432
rect 2552 1368 2568 1432
rect 2632 1368 2648 1432
rect 2712 1368 2728 1432
rect 2792 1368 2808 1432
rect 2872 1368 2888 1432
rect 2952 1368 2968 1432
rect 3032 1368 3048 1432
rect 3112 1368 3128 1432
rect 3192 1368 3208 1432
rect 3272 1368 3288 1432
rect 3352 1368 3368 1432
rect 3432 1368 3448 1432
rect 3512 1368 3528 1432
rect 3592 1368 3608 1432
rect 3672 1368 3688 1432
rect 3752 1368 3768 1432
rect 3832 1368 3848 1432
rect 3912 1368 3928 1432
rect 3992 1368 19112 1432
rect 19176 1368 19192 1432
rect 19256 1368 19272 1432
rect 19336 1368 19352 1432
rect 19416 1368 29112 1432
rect 29176 1368 29192 1432
rect 29256 1368 29272 1432
rect 29336 1368 29352 1432
rect 29416 1368 41376 1432
rect 41440 1368 41456 1432
rect 41520 1368 41536 1432
rect 41600 1368 41616 1432
rect 41680 1368 41696 1432
rect 41760 1368 41776 1432
rect 41840 1368 41856 1432
rect 41920 1368 41936 1432
rect 42000 1368 42016 1432
rect 42080 1368 42096 1432
rect 42160 1368 42176 1432
rect 42240 1368 42256 1432
rect 42320 1368 42336 1432
rect 42400 1368 42416 1432
rect 42480 1368 42496 1432
rect 42560 1368 42576 1432
rect 42640 1368 42656 1432
rect 42720 1368 42736 1432
rect 42800 1368 42816 1432
rect 42880 1368 42896 1432
rect 42960 1368 42976 1432
rect 43040 1368 43056 1432
rect 43120 1368 43136 1432
rect 43200 1368 43216 1432
rect 43280 1368 43296 1432
rect 43360 1368 43376 1432
rect 43440 1368 43456 1432
rect 43520 1368 43536 1432
rect 43600 1368 43616 1432
rect 43680 1368 43696 1432
rect 43760 1368 43776 1432
rect 43840 1368 43856 1432
rect 43920 1368 43936 1432
rect 44000 1368 44016 1432
rect 44080 1368 44096 1432
rect 44160 1368 44176 1432
rect 44240 1368 44256 1432
rect 44320 1368 44336 1432
rect 44400 1368 44416 1432
rect 44480 1368 44496 1432
rect 44560 1368 44576 1432
rect 44640 1368 44656 1432
rect 44720 1368 44736 1432
rect 44800 1368 44816 1432
rect 44880 1368 44896 1432
rect 44960 1368 44976 1432
rect 45040 1368 45056 1432
rect 45120 1368 45136 1432
rect 45200 1368 45216 1432
rect 45280 1368 45296 1432
rect 45360 1368 45368 1432
rect 0 1352 45368 1368
rect 0 1288 8 1352
rect 72 1288 88 1352
rect 152 1288 168 1352
rect 232 1288 248 1352
rect 312 1288 328 1352
rect 392 1288 408 1352
rect 472 1288 488 1352
rect 552 1288 568 1352
rect 632 1288 648 1352
rect 712 1288 728 1352
rect 792 1288 808 1352
rect 872 1288 888 1352
rect 952 1288 968 1352
rect 1032 1288 1048 1352
rect 1112 1288 1128 1352
rect 1192 1288 1208 1352
rect 1272 1288 1288 1352
rect 1352 1288 1368 1352
rect 1432 1288 1448 1352
rect 1512 1288 1528 1352
rect 1592 1288 1608 1352
rect 1672 1288 1688 1352
rect 1752 1288 1768 1352
rect 1832 1288 1848 1352
rect 1912 1288 1928 1352
rect 1992 1288 2008 1352
rect 2072 1288 2088 1352
rect 2152 1288 2168 1352
rect 2232 1288 2248 1352
rect 2312 1288 2328 1352
rect 2392 1288 2408 1352
rect 2472 1288 2488 1352
rect 2552 1288 2568 1352
rect 2632 1288 2648 1352
rect 2712 1288 2728 1352
rect 2792 1288 2808 1352
rect 2872 1288 2888 1352
rect 2952 1288 2968 1352
rect 3032 1288 3048 1352
rect 3112 1288 3128 1352
rect 3192 1288 3208 1352
rect 3272 1288 3288 1352
rect 3352 1288 3368 1352
rect 3432 1288 3448 1352
rect 3512 1288 3528 1352
rect 3592 1288 3608 1352
rect 3672 1288 3688 1352
rect 3752 1288 3768 1352
rect 3832 1288 3848 1352
rect 3912 1288 3928 1352
rect 3992 1288 19112 1352
rect 19176 1288 19192 1352
rect 19256 1288 19272 1352
rect 19336 1288 19352 1352
rect 19416 1288 29112 1352
rect 29176 1288 29192 1352
rect 29256 1288 29272 1352
rect 29336 1288 29352 1352
rect 29416 1288 41376 1352
rect 41440 1288 41456 1352
rect 41520 1288 41536 1352
rect 41600 1288 41616 1352
rect 41680 1288 41696 1352
rect 41760 1288 41776 1352
rect 41840 1288 41856 1352
rect 41920 1288 41936 1352
rect 42000 1288 42016 1352
rect 42080 1288 42096 1352
rect 42160 1288 42176 1352
rect 42240 1288 42256 1352
rect 42320 1288 42336 1352
rect 42400 1288 42416 1352
rect 42480 1288 42496 1352
rect 42560 1288 42576 1352
rect 42640 1288 42656 1352
rect 42720 1288 42736 1352
rect 42800 1288 42816 1352
rect 42880 1288 42896 1352
rect 42960 1288 42976 1352
rect 43040 1288 43056 1352
rect 43120 1288 43136 1352
rect 43200 1288 43216 1352
rect 43280 1288 43296 1352
rect 43360 1288 43376 1352
rect 43440 1288 43456 1352
rect 43520 1288 43536 1352
rect 43600 1288 43616 1352
rect 43680 1288 43696 1352
rect 43760 1288 43776 1352
rect 43840 1288 43856 1352
rect 43920 1288 43936 1352
rect 44000 1288 44016 1352
rect 44080 1288 44096 1352
rect 44160 1288 44176 1352
rect 44240 1288 44256 1352
rect 44320 1288 44336 1352
rect 44400 1288 44416 1352
rect 44480 1288 44496 1352
rect 44560 1288 44576 1352
rect 44640 1288 44656 1352
rect 44720 1288 44736 1352
rect 44800 1288 44816 1352
rect 44880 1288 44896 1352
rect 44960 1288 44976 1352
rect 45040 1288 45056 1352
rect 45120 1288 45136 1352
rect 45200 1288 45216 1352
rect 45280 1288 45296 1352
rect 45360 1288 45368 1352
rect 0 1272 45368 1288
rect 0 1208 8 1272
rect 72 1208 88 1272
rect 152 1208 168 1272
rect 232 1208 248 1272
rect 312 1208 328 1272
rect 392 1208 408 1272
rect 472 1208 488 1272
rect 552 1208 568 1272
rect 632 1208 648 1272
rect 712 1208 728 1272
rect 792 1208 808 1272
rect 872 1208 888 1272
rect 952 1208 968 1272
rect 1032 1208 1048 1272
rect 1112 1208 1128 1272
rect 1192 1208 1208 1272
rect 1272 1208 1288 1272
rect 1352 1208 1368 1272
rect 1432 1208 1448 1272
rect 1512 1208 1528 1272
rect 1592 1208 1608 1272
rect 1672 1208 1688 1272
rect 1752 1208 1768 1272
rect 1832 1208 1848 1272
rect 1912 1208 1928 1272
rect 1992 1208 2008 1272
rect 2072 1208 2088 1272
rect 2152 1208 2168 1272
rect 2232 1208 2248 1272
rect 2312 1208 2328 1272
rect 2392 1208 2408 1272
rect 2472 1208 2488 1272
rect 2552 1208 2568 1272
rect 2632 1208 2648 1272
rect 2712 1208 2728 1272
rect 2792 1208 2808 1272
rect 2872 1208 2888 1272
rect 2952 1208 2968 1272
rect 3032 1208 3048 1272
rect 3112 1208 3128 1272
rect 3192 1208 3208 1272
rect 3272 1208 3288 1272
rect 3352 1208 3368 1272
rect 3432 1208 3448 1272
rect 3512 1208 3528 1272
rect 3592 1208 3608 1272
rect 3672 1208 3688 1272
rect 3752 1208 3768 1272
rect 3832 1208 3848 1272
rect 3912 1208 3928 1272
rect 3992 1208 19112 1272
rect 19176 1208 19192 1272
rect 19256 1208 19272 1272
rect 19336 1208 19352 1272
rect 19416 1208 29112 1272
rect 29176 1208 29192 1272
rect 29256 1208 29272 1272
rect 29336 1208 29352 1272
rect 29416 1208 41376 1272
rect 41440 1208 41456 1272
rect 41520 1208 41536 1272
rect 41600 1208 41616 1272
rect 41680 1208 41696 1272
rect 41760 1208 41776 1272
rect 41840 1208 41856 1272
rect 41920 1208 41936 1272
rect 42000 1208 42016 1272
rect 42080 1208 42096 1272
rect 42160 1208 42176 1272
rect 42240 1208 42256 1272
rect 42320 1208 42336 1272
rect 42400 1208 42416 1272
rect 42480 1208 42496 1272
rect 42560 1208 42576 1272
rect 42640 1208 42656 1272
rect 42720 1208 42736 1272
rect 42800 1208 42816 1272
rect 42880 1208 42896 1272
rect 42960 1208 42976 1272
rect 43040 1208 43056 1272
rect 43120 1208 43136 1272
rect 43200 1208 43216 1272
rect 43280 1208 43296 1272
rect 43360 1208 43376 1272
rect 43440 1208 43456 1272
rect 43520 1208 43536 1272
rect 43600 1208 43616 1272
rect 43680 1208 43696 1272
rect 43760 1208 43776 1272
rect 43840 1208 43856 1272
rect 43920 1208 43936 1272
rect 44000 1208 44016 1272
rect 44080 1208 44096 1272
rect 44160 1208 44176 1272
rect 44240 1208 44256 1272
rect 44320 1208 44336 1272
rect 44400 1208 44416 1272
rect 44480 1208 44496 1272
rect 44560 1208 44576 1272
rect 44640 1208 44656 1272
rect 44720 1208 44736 1272
rect 44800 1208 44816 1272
rect 44880 1208 44896 1272
rect 44960 1208 44976 1272
rect 45040 1208 45056 1272
rect 45120 1208 45136 1272
rect 45200 1208 45216 1272
rect 45280 1208 45296 1272
rect 45360 1208 45368 1272
rect 0 1192 45368 1208
rect 0 1128 8 1192
rect 72 1128 88 1192
rect 152 1128 168 1192
rect 232 1128 248 1192
rect 312 1128 328 1192
rect 392 1128 408 1192
rect 472 1128 488 1192
rect 552 1128 568 1192
rect 632 1128 648 1192
rect 712 1128 728 1192
rect 792 1128 808 1192
rect 872 1128 888 1192
rect 952 1128 968 1192
rect 1032 1128 1048 1192
rect 1112 1128 1128 1192
rect 1192 1128 1208 1192
rect 1272 1128 1288 1192
rect 1352 1128 1368 1192
rect 1432 1128 1448 1192
rect 1512 1128 1528 1192
rect 1592 1128 1608 1192
rect 1672 1128 1688 1192
rect 1752 1128 1768 1192
rect 1832 1128 1848 1192
rect 1912 1128 1928 1192
rect 1992 1128 2008 1192
rect 2072 1128 2088 1192
rect 2152 1128 2168 1192
rect 2232 1128 2248 1192
rect 2312 1128 2328 1192
rect 2392 1128 2408 1192
rect 2472 1128 2488 1192
rect 2552 1128 2568 1192
rect 2632 1128 2648 1192
rect 2712 1128 2728 1192
rect 2792 1128 2808 1192
rect 2872 1128 2888 1192
rect 2952 1128 2968 1192
rect 3032 1128 3048 1192
rect 3112 1128 3128 1192
rect 3192 1128 3208 1192
rect 3272 1128 3288 1192
rect 3352 1128 3368 1192
rect 3432 1128 3448 1192
rect 3512 1128 3528 1192
rect 3592 1128 3608 1192
rect 3672 1128 3688 1192
rect 3752 1128 3768 1192
rect 3832 1128 3848 1192
rect 3912 1128 3928 1192
rect 3992 1128 19112 1192
rect 19176 1128 19192 1192
rect 19256 1128 19272 1192
rect 19336 1128 19352 1192
rect 19416 1128 29112 1192
rect 29176 1128 29192 1192
rect 29256 1128 29272 1192
rect 29336 1128 29352 1192
rect 29416 1128 41376 1192
rect 41440 1128 41456 1192
rect 41520 1128 41536 1192
rect 41600 1128 41616 1192
rect 41680 1128 41696 1192
rect 41760 1128 41776 1192
rect 41840 1128 41856 1192
rect 41920 1128 41936 1192
rect 42000 1128 42016 1192
rect 42080 1128 42096 1192
rect 42160 1128 42176 1192
rect 42240 1128 42256 1192
rect 42320 1128 42336 1192
rect 42400 1128 42416 1192
rect 42480 1128 42496 1192
rect 42560 1128 42576 1192
rect 42640 1128 42656 1192
rect 42720 1128 42736 1192
rect 42800 1128 42816 1192
rect 42880 1128 42896 1192
rect 42960 1128 42976 1192
rect 43040 1128 43056 1192
rect 43120 1128 43136 1192
rect 43200 1128 43216 1192
rect 43280 1128 43296 1192
rect 43360 1128 43376 1192
rect 43440 1128 43456 1192
rect 43520 1128 43536 1192
rect 43600 1128 43616 1192
rect 43680 1128 43696 1192
rect 43760 1128 43776 1192
rect 43840 1128 43856 1192
rect 43920 1128 43936 1192
rect 44000 1128 44016 1192
rect 44080 1128 44096 1192
rect 44160 1128 44176 1192
rect 44240 1128 44256 1192
rect 44320 1128 44336 1192
rect 44400 1128 44416 1192
rect 44480 1128 44496 1192
rect 44560 1128 44576 1192
rect 44640 1128 44656 1192
rect 44720 1128 44736 1192
rect 44800 1128 44816 1192
rect 44880 1128 44896 1192
rect 44960 1128 44976 1192
rect 45040 1128 45056 1192
rect 45120 1128 45136 1192
rect 45200 1128 45216 1192
rect 45280 1128 45296 1192
rect 45360 1128 45368 1192
rect 0 1112 45368 1128
rect 0 1048 8 1112
rect 72 1048 88 1112
rect 152 1048 168 1112
rect 232 1048 248 1112
rect 312 1048 328 1112
rect 392 1048 408 1112
rect 472 1048 488 1112
rect 552 1048 568 1112
rect 632 1048 648 1112
rect 712 1048 728 1112
rect 792 1048 808 1112
rect 872 1048 888 1112
rect 952 1048 968 1112
rect 1032 1048 1048 1112
rect 1112 1048 1128 1112
rect 1192 1048 1208 1112
rect 1272 1048 1288 1112
rect 1352 1048 1368 1112
rect 1432 1048 1448 1112
rect 1512 1048 1528 1112
rect 1592 1048 1608 1112
rect 1672 1048 1688 1112
rect 1752 1048 1768 1112
rect 1832 1048 1848 1112
rect 1912 1048 1928 1112
rect 1992 1048 2008 1112
rect 2072 1048 2088 1112
rect 2152 1048 2168 1112
rect 2232 1048 2248 1112
rect 2312 1048 2328 1112
rect 2392 1048 2408 1112
rect 2472 1048 2488 1112
rect 2552 1048 2568 1112
rect 2632 1048 2648 1112
rect 2712 1048 2728 1112
rect 2792 1048 2808 1112
rect 2872 1048 2888 1112
rect 2952 1048 2968 1112
rect 3032 1048 3048 1112
rect 3112 1048 3128 1112
rect 3192 1048 3208 1112
rect 3272 1048 3288 1112
rect 3352 1048 3368 1112
rect 3432 1048 3448 1112
rect 3512 1048 3528 1112
rect 3592 1048 3608 1112
rect 3672 1048 3688 1112
rect 3752 1048 3768 1112
rect 3832 1048 3848 1112
rect 3912 1048 3928 1112
rect 3992 1048 19112 1112
rect 19176 1048 19192 1112
rect 19256 1048 19272 1112
rect 19336 1048 19352 1112
rect 19416 1048 29112 1112
rect 29176 1048 29192 1112
rect 29256 1048 29272 1112
rect 29336 1048 29352 1112
rect 29416 1048 41376 1112
rect 41440 1048 41456 1112
rect 41520 1048 41536 1112
rect 41600 1048 41616 1112
rect 41680 1048 41696 1112
rect 41760 1048 41776 1112
rect 41840 1048 41856 1112
rect 41920 1048 41936 1112
rect 42000 1048 42016 1112
rect 42080 1048 42096 1112
rect 42160 1048 42176 1112
rect 42240 1048 42256 1112
rect 42320 1048 42336 1112
rect 42400 1048 42416 1112
rect 42480 1048 42496 1112
rect 42560 1048 42576 1112
rect 42640 1048 42656 1112
rect 42720 1048 42736 1112
rect 42800 1048 42816 1112
rect 42880 1048 42896 1112
rect 42960 1048 42976 1112
rect 43040 1048 43056 1112
rect 43120 1048 43136 1112
rect 43200 1048 43216 1112
rect 43280 1048 43296 1112
rect 43360 1048 43376 1112
rect 43440 1048 43456 1112
rect 43520 1048 43536 1112
rect 43600 1048 43616 1112
rect 43680 1048 43696 1112
rect 43760 1048 43776 1112
rect 43840 1048 43856 1112
rect 43920 1048 43936 1112
rect 44000 1048 44016 1112
rect 44080 1048 44096 1112
rect 44160 1048 44176 1112
rect 44240 1048 44256 1112
rect 44320 1048 44336 1112
rect 44400 1048 44416 1112
rect 44480 1048 44496 1112
rect 44560 1048 44576 1112
rect 44640 1048 44656 1112
rect 44720 1048 44736 1112
rect 44800 1048 44816 1112
rect 44880 1048 44896 1112
rect 44960 1048 44976 1112
rect 45040 1048 45056 1112
rect 45120 1048 45136 1112
rect 45200 1048 45216 1112
rect 45280 1048 45296 1112
rect 45360 1048 45368 1112
rect 0 1032 45368 1048
rect 0 968 8 1032
rect 72 968 88 1032
rect 152 968 168 1032
rect 232 968 248 1032
rect 312 968 328 1032
rect 392 968 408 1032
rect 472 968 488 1032
rect 552 968 568 1032
rect 632 968 648 1032
rect 712 968 728 1032
rect 792 968 808 1032
rect 872 968 888 1032
rect 952 968 968 1032
rect 1032 968 1048 1032
rect 1112 968 1128 1032
rect 1192 968 1208 1032
rect 1272 968 1288 1032
rect 1352 968 1368 1032
rect 1432 968 1448 1032
rect 1512 968 1528 1032
rect 1592 968 1608 1032
rect 1672 968 1688 1032
rect 1752 968 1768 1032
rect 1832 968 1848 1032
rect 1912 968 1928 1032
rect 1992 968 2008 1032
rect 2072 968 2088 1032
rect 2152 968 2168 1032
rect 2232 968 2248 1032
rect 2312 968 2328 1032
rect 2392 968 2408 1032
rect 2472 968 2488 1032
rect 2552 968 2568 1032
rect 2632 968 2648 1032
rect 2712 968 2728 1032
rect 2792 968 2808 1032
rect 2872 968 2888 1032
rect 2952 968 2968 1032
rect 3032 968 3048 1032
rect 3112 968 3128 1032
rect 3192 968 3208 1032
rect 3272 968 3288 1032
rect 3352 968 3368 1032
rect 3432 968 3448 1032
rect 3512 968 3528 1032
rect 3592 968 3608 1032
rect 3672 968 3688 1032
rect 3752 968 3768 1032
rect 3832 968 3848 1032
rect 3912 968 3928 1032
rect 3992 968 19112 1032
rect 19176 968 19192 1032
rect 19256 968 19272 1032
rect 19336 968 19352 1032
rect 19416 968 29112 1032
rect 29176 968 29192 1032
rect 29256 968 29272 1032
rect 29336 968 29352 1032
rect 29416 968 41376 1032
rect 41440 968 41456 1032
rect 41520 968 41536 1032
rect 41600 968 41616 1032
rect 41680 968 41696 1032
rect 41760 968 41776 1032
rect 41840 968 41856 1032
rect 41920 968 41936 1032
rect 42000 968 42016 1032
rect 42080 968 42096 1032
rect 42160 968 42176 1032
rect 42240 968 42256 1032
rect 42320 968 42336 1032
rect 42400 968 42416 1032
rect 42480 968 42496 1032
rect 42560 968 42576 1032
rect 42640 968 42656 1032
rect 42720 968 42736 1032
rect 42800 968 42816 1032
rect 42880 968 42896 1032
rect 42960 968 42976 1032
rect 43040 968 43056 1032
rect 43120 968 43136 1032
rect 43200 968 43216 1032
rect 43280 968 43296 1032
rect 43360 968 43376 1032
rect 43440 968 43456 1032
rect 43520 968 43536 1032
rect 43600 968 43616 1032
rect 43680 968 43696 1032
rect 43760 968 43776 1032
rect 43840 968 43856 1032
rect 43920 968 43936 1032
rect 44000 968 44016 1032
rect 44080 968 44096 1032
rect 44160 968 44176 1032
rect 44240 968 44256 1032
rect 44320 968 44336 1032
rect 44400 968 44416 1032
rect 44480 968 44496 1032
rect 44560 968 44576 1032
rect 44640 968 44656 1032
rect 44720 968 44736 1032
rect 44800 968 44816 1032
rect 44880 968 44896 1032
rect 44960 968 44976 1032
rect 45040 968 45056 1032
rect 45120 968 45136 1032
rect 45200 968 45216 1032
rect 45280 968 45296 1032
rect 45360 968 45368 1032
rect 0 952 45368 968
rect 0 888 8 952
rect 72 888 88 952
rect 152 888 168 952
rect 232 888 248 952
rect 312 888 328 952
rect 392 888 408 952
rect 472 888 488 952
rect 552 888 568 952
rect 632 888 648 952
rect 712 888 728 952
rect 792 888 808 952
rect 872 888 888 952
rect 952 888 968 952
rect 1032 888 1048 952
rect 1112 888 1128 952
rect 1192 888 1208 952
rect 1272 888 1288 952
rect 1352 888 1368 952
rect 1432 888 1448 952
rect 1512 888 1528 952
rect 1592 888 1608 952
rect 1672 888 1688 952
rect 1752 888 1768 952
rect 1832 888 1848 952
rect 1912 888 1928 952
rect 1992 888 2008 952
rect 2072 888 2088 952
rect 2152 888 2168 952
rect 2232 888 2248 952
rect 2312 888 2328 952
rect 2392 888 2408 952
rect 2472 888 2488 952
rect 2552 888 2568 952
rect 2632 888 2648 952
rect 2712 888 2728 952
rect 2792 888 2808 952
rect 2872 888 2888 952
rect 2952 888 2968 952
rect 3032 888 3048 952
rect 3112 888 3128 952
rect 3192 888 3208 952
rect 3272 888 3288 952
rect 3352 888 3368 952
rect 3432 888 3448 952
rect 3512 888 3528 952
rect 3592 888 3608 952
rect 3672 888 3688 952
rect 3752 888 3768 952
rect 3832 888 3848 952
rect 3912 888 3928 952
rect 3992 888 19112 952
rect 19176 888 19192 952
rect 19256 888 19272 952
rect 19336 888 19352 952
rect 19416 888 29112 952
rect 29176 888 29192 952
rect 29256 888 29272 952
rect 29336 888 29352 952
rect 29416 888 41376 952
rect 41440 888 41456 952
rect 41520 888 41536 952
rect 41600 888 41616 952
rect 41680 888 41696 952
rect 41760 888 41776 952
rect 41840 888 41856 952
rect 41920 888 41936 952
rect 42000 888 42016 952
rect 42080 888 42096 952
rect 42160 888 42176 952
rect 42240 888 42256 952
rect 42320 888 42336 952
rect 42400 888 42416 952
rect 42480 888 42496 952
rect 42560 888 42576 952
rect 42640 888 42656 952
rect 42720 888 42736 952
rect 42800 888 42816 952
rect 42880 888 42896 952
rect 42960 888 42976 952
rect 43040 888 43056 952
rect 43120 888 43136 952
rect 43200 888 43216 952
rect 43280 888 43296 952
rect 43360 888 43376 952
rect 43440 888 43456 952
rect 43520 888 43536 952
rect 43600 888 43616 952
rect 43680 888 43696 952
rect 43760 888 43776 952
rect 43840 888 43856 952
rect 43920 888 43936 952
rect 44000 888 44016 952
rect 44080 888 44096 952
rect 44160 888 44176 952
rect 44240 888 44256 952
rect 44320 888 44336 952
rect 44400 888 44416 952
rect 44480 888 44496 952
rect 44560 888 44576 952
rect 44640 888 44656 952
rect 44720 888 44736 952
rect 44800 888 44816 952
rect 44880 888 44896 952
rect 44960 888 44976 952
rect 45040 888 45056 952
rect 45120 888 45136 952
rect 45200 888 45216 952
rect 45280 888 45296 952
rect 45360 888 45368 952
rect 0 872 45368 888
rect 0 808 8 872
rect 72 808 88 872
rect 152 808 168 872
rect 232 808 248 872
rect 312 808 328 872
rect 392 808 408 872
rect 472 808 488 872
rect 552 808 568 872
rect 632 808 648 872
rect 712 808 728 872
rect 792 808 808 872
rect 872 808 888 872
rect 952 808 968 872
rect 1032 808 1048 872
rect 1112 808 1128 872
rect 1192 808 1208 872
rect 1272 808 1288 872
rect 1352 808 1368 872
rect 1432 808 1448 872
rect 1512 808 1528 872
rect 1592 808 1608 872
rect 1672 808 1688 872
rect 1752 808 1768 872
rect 1832 808 1848 872
rect 1912 808 1928 872
rect 1992 808 2008 872
rect 2072 808 2088 872
rect 2152 808 2168 872
rect 2232 808 2248 872
rect 2312 808 2328 872
rect 2392 808 2408 872
rect 2472 808 2488 872
rect 2552 808 2568 872
rect 2632 808 2648 872
rect 2712 808 2728 872
rect 2792 808 2808 872
rect 2872 808 2888 872
rect 2952 808 2968 872
rect 3032 808 3048 872
rect 3112 808 3128 872
rect 3192 808 3208 872
rect 3272 808 3288 872
rect 3352 808 3368 872
rect 3432 808 3448 872
rect 3512 808 3528 872
rect 3592 808 3608 872
rect 3672 808 3688 872
rect 3752 808 3768 872
rect 3832 808 3848 872
rect 3912 808 3928 872
rect 3992 808 19112 872
rect 19176 808 19192 872
rect 19256 808 19272 872
rect 19336 808 19352 872
rect 19416 808 29112 872
rect 29176 808 29192 872
rect 29256 808 29272 872
rect 29336 808 29352 872
rect 29416 808 41376 872
rect 41440 808 41456 872
rect 41520 808 41536 872
rect 41600 808 41616 872
rect 41680 808 41696 872
rect 41760 808 41776 872
rect 41840 808 41856 872
rect 41920 808 41936 872
rect 42000 808 42016 872
rect 42080 808 42096 872
rect 42160 808 42176 872
rect 42240 808 42256 872
rect 42320 808 42336 872
rect 42400 808 42416 872
rect 42480 808 42496 872
rect 42560 808 42576 872
rect 42640 808 42656 872
rect 42720 808 42736 872
rect 42800 808 42816 872
rect 42880 808 42896 872
rect 42960 808 42976 872
rect 43040 808 43056 872
rect 43120 808 43136 872
rect 43200 808 43216 872
rect 43280 808 43296 872
rect 43360 808 43376 872
rect 43440 808 43456 872
rect 43520 808 43536 872
rect 43600 808 43616 872
rect 43680 808 43696 872
rect 43760 808 43776 872
rect 43840 808 43856 872
rect 43920 808 43936 872
rect 44000 808 44016 872
rect 44080 808 44096 872
rect 44160 808 44176 872
rect 44240 808 44256 872
rect 44320 808 44336 872
rect 44400 808 44416 872
rect 44480 808 44496 872
rect 44560 808 44576 872
rect 44640 808 44656 872
rect 44720 808 44736 872
rect 44800 808 44816 872
rect 44880 808 44896 872
rect 44960 808 44976 872
rect 45040 808 45056 872
rect 45120 808 45136 872
rect 45200 808 45216 872
rect 45280 808 45296 872
rect 45360 808 45368 872
rect 0 792 45368 808
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 808 792
rect 872 728 888 792
rect 952 728 968 792
rect 1032 728 1048 792
rect 1112 728 1128 792
rect 1192 728 1208 792
rect 1272 728 1288 792
rect 1352 728 1368 792
rect 1432 728 1448 792
rect 1512 728 1528 792
rect 1592 728 1608 792
rect 1672 728 1688 792
rect 1752 728 1768 792
rect 1832 728 1848 792
rect 1912 728 1928 792
rect 1992 728 2008 792
rect 2072 728 2088 792
rect 2152 728 2168 792
rect 2232 728 2248 792
rect 2312 728 2328 792
rect 2392 728 2408 792
rect 2472 728 2488 792
rect 2552 728 2568 792
rect 2632 728 2648 792
rect 2712 728 2728 792
rect 2792 728 2808 792
rect 2872 728 2888 792
rect 2952 728 2968 792
rect 3032 728 3048 792
rect 3112 728 3128 792
rect 3192 728 3208 792
rect 3272 728 3288 792
rect 3352 728 3368 792
rect 3432 728 3448 792
rect 3512 728 3528 792
rect 3592 728 3608 792
rect 3672 728 3688 792
rect 3752 728 3768 792
rect 3832 728 3848 792
rect 3912 728 3928 792
rect 3992 728 19112 792
rect 19176 728 19192 792
rect 19256 728 19272 792
rect 19336 728 19352 792
rect 19416 728 29112 792
rect 29176 728 29192 792
rect 29256 728 29272 792
rect 29336 728 29352 792
rect 29416 728 41376 792
rect 41440 728 41456 792
rect 41520 728 41536 792
rect 41600 728 41616 792
rect 41680 728 41696 792
rect 41760 728 41776 792
rect 41840 728 41856 792
rect 41920 728 41936 792
rect 42000 728 42016 792
rect 42080 728 42096 792
rect 42160 728 42176 792
rect 42240 728 42256 792
rect 42320 728 42336 792
rect 42400 728 42416 792
rect 42480 728 42496 792
rect 42560 728 42576 792
rect 42640 728 42656 792
rect 42720 728 42736 792
rect 42800 728 42816 792
rect 42880 728 42896 792
rect 42960 728 42976 792
rect 43040 728 43056 792
rect 43120 728 43136 792
rect 43200 728 43216 792
rect 43280 728 43296 792
rect 43360 728 43376 792
rect 43440 728 43456 792
rect 43520 728 43536 792
rect 43600 728 43616 792
rect 43680 728 43696 792
rect 43760 728 43776 792
rect 43840 728 43856 792
rect 43920 728 43936 792
rect 44000 728 44016 792
rect 44080 728 44096 792
rect 44160 728 44176 792
rect 44240 728 44256 792
rect 44320 728 44336 792
rect 44400 728 44416 792
rect 44480 728 44496 792
rect 44560 728 44576 792
rect 44640 728 44656 792
rect 44720 728 44736 792
rect 44800 728 44816 792
rect 44880 728 44896 792
rect 44960 728 44976 792
rect 45040 728 45056 792
rect 45120 728 45136 792
rect 45200 728 45216 792
rect 45280 728 45296 792
rect 45360 728 45368 792
rect 0 712 45368 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 808 712
rect 872 648 888 712
rect 952 648 968 712
rect 1032 648 1048 712
rect 1112 648 1128 712
rect 1192 648 1208 712
rect 1272 648 1288 712
rect 1352 648 1368 712
rect 1432 648 1448 712
rect 1512 648 1528 712
rect 1592 648 1608 712
rect 1672 648 1688 712
rect 1752 648 1768 712
rect 1832 648 1848 712
rect 1912 648 1928 712
rect 1992 648 2008 712
rect 2072 648 2088 712
rect 2152 648 2168 712
rect 2232 648 2248 712
rect 2312 648 2328 712
rect 2392 648 2408 712
rect 2472 648 2488 712
rect 2552 648 2568 712
rect 2632 648 2648 712
rect 2712 648 2728 712
rect 2792 648 2808 712
rect 2872 648 2888 712
rect 2952 648 2968 712
rect 3032 648 3048 712
rect 3112 648 3128 712
rect 3192 648 3208 712
rect 3272 648 3288 712
rect 3352 648 3368 712
rect 3432 648 3448 712
rect 3512 648 3528 712
rect 3592 648 3608 712
rect 3672 648 3688 712
rect 3752 648 3768 712
rect 3832 648 3848 712
rect 3912 648 3928 712
rect 3992 648 19112 712
rect 19176 648 19192 712
rect 19256 648 19272 712
rect 19336 648 19352 712
rect 19416 648 29112 712
rect 29176 648 29192 712
rect 29256 648 29272 712
rect 29336 648 29352 712
rect 29416 648 41376 712
rect 41440 648 41456 712
rect 41520 648 41536 712
rect 41600 648 41616 712
rect 41680 648 41696 712
rect 41760 648 41776 712
rect 41840 648 41856 712
rect 41920 648 41936 712
rect 42000 648 42016 712
rect 42080 648 42096 712
rect 42160 648 42176 712
rect 42240 648 42256 712
rect 42320 648 42336 712
rect 42400 648 42416 712
rect 42480 648 42496 712
rect 42560 648 42576 712
rect 42640 648 42656 712
rect 42720 648 42736 712
rect 42800 648 42816 712
rect 42880 648 42896 712
rect 42960 648 42976 712
rect 43040 648 43056 712
rect 43120 648 43136 712
rect 43200 648 43216 712
rect 43280 648 43296 712
rect 43360 648 43376 712
rect 43440 648 43456 712
rect 43520 648 43536 712
rect 43600 648 43616 712
rect 43680 648 43696 712
rect 43760 648 43776 712
rect 43840 648 43856 712
rect 43920 648 43936 712
rect 44000 648 44016 712
rect 44080 648 44096 712
rect 44160 648 44176 712
rect 44240 648 44256 712
rect 44320 648 44336 712
rect 44400 648 44416 712
rect 44480 648 44496 712
rect 44560 648 44576 712
rect 44640 648 44656 712
rect 44720 648 44736 712
rect 44800 648 44816 712
rect 44880 648 44896 712
rect 44960 648 44976 712
rect 45040 648 45056 712
rect 45120 648 45136 712
rect 45200 648 45216 712
rect 45280 648 45296 712
rect 45360 648 45368 712
rect 0 632 45368 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 808 632
rect 872 568 888 632
rect 952 568 968 632
rect 1032 568 1048 632
rect 1112 568 1128 632
rect 1192 568 1208 632
rect 1272 568 1288 632
rect 1352 568 1368 632
rect 1432 568 1448 632
rect 1512 568 1528 632
rect 1592 568 1608 632
rect 1672 568 1688 632
rect 1752 568 1768 632
rect 1832 568 1848 632
rect 1912 568 1928 632
rect 1992 568 2008 632
rect 2072 568 2088 632
rect 2152 568 2168 632
rect 2232 568 2248 632
rect 2312 568 2328 632
rect 2392 568 2408 632
rect 2472 568 2488 632
rect 2552 568 2568 632
rect 2632 568 2648 632
rect 2712 568 2728 632
rect 2792 568 2808 632
rect 2872 568 2888 632
rect 2952 568 2968 632
rect 3032 568 3048 632
rect 3112 568 3128 632
rect 3192 568 3208 632
rect 3272 568 3288 632
rect 3352 568 3368 632
rect 3432 568 3448 632
rect 3512 568 3528 632
rect 3592 568 3608 632
rect 3672 568 3688 632
rect 3752 568 3768 632
rect 3832 568 3848 632
rect 3912 568 3928 632
rect 3992 568 19112 632
rect 19176 568 19192 632
rect 19256 568 19272 632
rect 19336 568 19352 632
rect 19416 568 29112 632
rect 29176 568 29192 632
rect 29256 568 29272 632
rect 29336 568 29352 632
rect 29416 568 41376 632
rect 41440 568 41456 632
rect 41520 568 41536 632
rect 41600 568 41616 632
rect 41680 568 41696 632
rect 41760 568 41776 632
rect 41840 568 41856 632
rect 41920 568 41936 632
rect 42000 568 42016 632
rect 42080 568 42096 632
rect 42160 568 42176 632
rect 42240 568 42256 632
rect 42320 568 42336 632
rect 42400 568 42416 632
rect 42480 568 42496 632
rect 42560 568 42576 632
rect 42640 568 42656 632
rect 42720 568 42736 632
rect 42800 568 42816 632
rect 42880 568 42896 632
rect 42960 568 42976 632
rect 43040 568 43056 632
rect 43120 568 43136 632
rect 43200 568 43216 632
rect 43280 568 43296 632
rect 43360 568 43376 632
rect 43440 568 43456 632
rect 43520 568 43536 632
rect 43600 568 43616 632
rect 43680 568 43696 632
rect 43760 568 43776 632
rect 43840 568 43856 632
rect 43920 568 43936 632
rect 44000 568 44016 632
rect 44080 568 44096 632
rect 44160 568 44176 632
rect 44240 568 44256 632
rect 44320 568 44336 632
rect 44400 568 44416 632
rect 44480 568 44496 632
rect 44560 568 44576 632
rect 44640 568 44656 632
rect 44720 568 44736 632
rect 44800 568 44816 632
rect 44880 568 44896 632
rect 44960 568 44976 632
rect 45040 568 45056 632
rect 45120 568 45136 632
rect 45200 568 45216 632
rect 45280 568 45296 632
rect 45360 568 45368 632
rect 0 552 45368 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 808 552
rect 872 488 888 552
rect 952 488 968 552
rect 1032 488 1048 552
rect 1112 488 1128 552
rect 1192 488 1208 552
rect 1272 488 1288 552
rect 1352 488 1368 552
rect 1432 488 1448 552
rect 1512 488 1528 552
rect 1592 488 1608 552
rect 1672 488 1688 552
rect 1752 488 1768 552
rect 1832 488 1848 552
rect 1912 488 1928 552
rect 1992 488 2008 552
rect 2072 488 2088 552
rect 2152 488 2168 552
rect 2232 488 2248 552
rect 2312 488 2328 552
rect 2392 488 2408 552
rect 2472 488 2488 552
rect 2552 488 2568 552
rect 2632 488 2648 552
rect 2712 488 2728 552
rect 2792 488 2808 552
rect 2872 488 2888 552
rect 2952 488 2968 552
rect 3032 488 3048 552
rect 3112 488 3128 552
rect 3192 488 3208 552
rect 3272 488 3288 552
rect 3352 488 3368 552
rect 3432 488 3448 552
rect 3512 488 3528 552
rect 3592 488 3608 552
rect 3672 488 3688 552
rect 3752 488 3768 552
rect 3832 488 3848 552
rect 3912 488 3928 552
rect 3992 488 19112 552
rect 19176 488 19192 552
rect 19256 488 19272 552
rect 19336 488 19352 552
rect 19416 488 29112 552
rect 29176 488 29192 552
rect 29256 488 29272 552
rect 29336 488 29352 552
rect 29416 488 41376 552
rect 41440 488 41456 552
rect 41520 488 41536 552
rect 41600 488 41616 552
rect 41680 488 41696 552
rect 41760 488 41776 552
rect 41840 488 41856 552
rect 41920 488 41936 552
rect 42000 488 42016 552
rect 42080 488 42096 552
rect 42160 488 42176 552
rect 42240 488 42256 552
rect 42320 488 42336 552
rect 42400 488 42416 552
rect 42480 488 42496 552
rect 42560 488 42576 552
rect 42640 488 42656 552
rect 42720 488 42736 552
rect 42800 488 42816 552
rect 42880 488 42896 552
rect 42960 488 42976 552
rect 43040 488 43056 552
rect 43120 488 43136 552
rect 43200 488 43216 552
rect 43280 488 43296 552
rect 43360 488 43376 552
rect 43440 488 43456 552
rect 43520 488 43536 552
rect 43600 488 43616 552
rect 43680 488 43696 552
rect 43760 488 43776 552
rect 43840 488 43856 552
rect 43920 488 43936 552
rect 44000 488 44016 552
rect 44080 488 44096 552
rect 44160 488 44176 552
rect 44240 488 44256 552
rect 44320 488 44336 552
rect 44400 488 44416 552
rect 44480 488 44496 552
rect 44560 488 44576 552
rect 44640 488 44656 552
rect 44720 488 44736 552
rect 44800 488 44816 552
rect 44880 488 44896 552
rect 44960 488 44976 552
rect 45040 488 45056 552
rect 45120 488 45136 552
rect 45200 488 45216 552
rect 45280 488 45296 552
rect 45360 488 45368 552
rect 0 472 45368 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 808 472
rect 872 408 888 472
rect 952 408 968 472
rect 1032 408 1048 472
rect 1112 408 1128 472
rect 1192 408 1208 472
rect 1272 408 1288 472
rect 1352 408 1368 472
rect 1432 408 1448 472
rect 1512 408 1528 472
rect 1592 408 1608 472
rect 1672 408 1688 472
rect 1752 408 1768 472
rect 1832 408 1848 472
rect 1912 408 1928 472
rect 1992 408 2008 472
rect 2072 408 2088 472
rect 2152 408 2168 472
rect 2232 408 2248 472
rect 2312 408 2328 472
rect 2392 408 2408 472
rect 2472 408 2488 472
rect 2552 408 2568 472
rect 2632 408 2648 472
rect 2712 408 2728 472
rect 2792 408 2808 472
rect 2872 408 2888 472
rect 2952 408 2968 472
rect 3032 408 3048 472
rect 3112 408 3128 472
rect 3192 408 3208 472
rect 3272 408 3288 472
rect 3352 408 3368 472
rect 3432 408 3448 472
rect 3512 408 3528 472
rect 3592 408 3608 472
rect 3672 408 3688 472
rect 3752 408 3768 472
rect 3832 408 3848 472
rect 3912 408 3928 472
rect 3992 408 19112 472
rect 19176 408 19192 472
rect 19256 408 19272 472
rect 19336 408 19352 472
rect 19416 408 29112 472
rect 29176 408 29192 472
rect 29256 408 29272 472
rect 29336 408 29352 472
rect 29416 408 41376 472
rect 41440 408 41456 472
rect 41520 408 41536 472
rect 41600 408 41616 472
rect 41680 408 41696 472
rect 41760 408 41776 472
rect 41840 408 41856 472
rect 41920 408 41936 472
rect 42000 408 42016 472
rect 42080 408 42096 472
rect 42160 408 42176 472
rect 42240 408 42256 472
rect 42320 408 42336 472
rect 42400 408 42416 472
rect 42480 408 42496 472
rect 42560 408 42576 472
rect 42640 408 42656 472
rect 42720 408 42736 472
rect 42800 408 42816 472
rect 42880 408 42896 472
rect 42960 408 42976 472
rect 43040 408 43056 472
rect 43120 408 43136 472
rect 43200 408 43216 472
rect 43280 408 43296 472
rect 43360 408 43376 472
rect 43440 408 43456 472
rect 43520 408 43536 472
rect 43600 408 43616 472
rect 43680 408 43696 472
rect 43760 408 43776 472
rect 43840 408 43856 472
rect 43920 408 43936 472
rect 44000 408 44016 472
rect 44080 408 44096 472
rect 44160 408 44176 472
rect 44240 408 44256 472
rect 44320 408 44336 472
rect 44400 408 44416 472
rect 44480 408 44496 472
rect 44560 408 44576 472
rect 44640 408 44656 472
rect 44720 408 44736 472
rect 44800 408 44816 472
rect 44880 408 44896 472
rect 44960 408 44976 472
rect 45040 408 45056 472
rect 45120 408 45136 472
rect 45200 408 45216 472
rect 45280 408 45296 472
rect 45360 408 45368 472
rect 0 392 45368 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 808 392
rect 872 328 888 392
rect 952 328 968 392
rect 1032 328 1048 392
rect 1112 328 1128 392
rect 1192 328 1208 392
rect 1272 328 1288 392
rect 1352 328 1368 392
rect 1432 328 1448 392
rect 1512 328 1528 392
rect 1592 328 1608 392
rect 1672 328 1688 392
rect 1752 328 1768 392
rect 1832 328 1848 392
rect 1912 328 1928 392
rect 1992 328 2008 392
rect 2072 328 2088 392
rect 2152 328 2168 392
rect 2232 328 2248 392
rect 2312 328 2328 392
rect 2392 328 2408 392
rect 2472 328 2488 392
rect 2552 328 2568 392
rect 2632 328 2648 392
rect 2712 328 2728 392
rect 2792 328 2808 392
rect 2872 328 2888 392
rect 2952 328 2968 392
rect 3032 328 3048 392
rect 3112 328 3128 392
rect 3192 328 3208 392
rect 3272 328 3288 392
rect 3352 328 3368 392
rect 3432 328 3448 392
rect 3512 328 3528 392
rect 3592 328 3608 392
rect 3672 328 3688 392
rect 3752 328 3768 392
rect 3832 328 3848 392
rect 3912 328 3928 392
rect 3992 328 19112 392
rect 19176 328 19192 392
rect 19256 328 19272 392
rect 19336 328 19352 392
rect 19416 328 29112 392
rect 29176 328 29192 392
rect 29256 328 29272 392
rect 29336 328 29352 392
rect 29416 328 41376 392
rect 41440 328 41456 392
rect 41520 328 41536 392
rect 41600 328 41616 392
rect 41680 328 41696 392
rect 41760 328 41776 392
rect 41840 328 41856 392
rect 41920 328 41936 392
rect 42000 328 42016 392
rect 42080 328 42096 392
rect 42160 328 42176 392
rect 42240 328 42256 392
rect 42320 328 42336 392
rect 42400 328 42416 392
rect 42480 328 42496 392
rect 42560 328 42576 392
rect 42640 328 42656 392
rect 42720 328 42736 392
rect 42800 328 42816 392
rect 42880 328 42896 392
rect 42960 328 42976 392
rect 43040 328 43056 392
rect 43120 328 43136 392
rect 43200 328 43216 392
rect 43280 328 43296 392
rect 43360 328 43376 392
rect 43440 328 43456 392
rect 43520 328 43536 392
rect 43600 328 43616 392
rect 43680 328 43696 392
rect 43760 328 43776 392
rect 43840 328 43856 392
rect 43920 328 43936 392
rect 44000 328 44016 392
rect 44080 328 44096 392
rect 44160 328 44176 392
rect 44240 328 44256 392
rect 44320 328 44336 392
rect 44400 328 44416 392
rect 44480 328 44496 392
rect 44560 328 44576 392
rect 44640 328 44656 392
rect 44720 328 44736 392
rect 44800 328 44816 392
rect 44880 328 44896 392
rect 44960 328 44976 392
rect 45040 328 45056 392
rect 45120 328 45136 392
rect 45200 328 45216 392
rect 45280 328 45296 392
rect 45360 328 45368 392
rect 0 312 45368 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 808 312
rect 872 248 888 312
rect 952 248 968 312
rect 1032 248 1048 312
rect 1112 248 1128 312
rect 1192 248 1208 312
rect 1272 248 1288 312
rect 1352 248 1368 312
rect 1432 248 1448 312
rect 1512 248 1528 312
rect 1592 248 1608 312
rect 1672 248 1688 312
rect 1752 248 1768 312
rect 1832 248 1848 312
rect 1912 248 1928 312
rect 1992 248 2008 312
rect 2072 248 2088 312
rect 2152 248 2168 312
rect 2232 248 2248 312
rect 2312 248 2328 312
rect 2392 248 2408 312
rect 2472 248 2488 312
rect 2552 248 2568 312
rect 2632 248 2648 312
rect 2712 248 2728 312
rect 2792 248 2808 312
rect 2872 248 2888 312
rect 2952 248 2968 312
rect 3032 248 3048 312
rect 3112 248 3128 312
rect 3192 248 3208 312
rect 3272 248 3288 312
rect 3352 248 3368 312
rect 3432 248 3448 312
rect 3512 248 3528 312
rect 3592 248 3608 312
rect 3672 248 3688 312
rect 3752 248 3768 312
rect 3832 248 3848 312
rect 3912 248 3928 312
rect 3992 248 19112 312
rect 19176 248 19192 312
rect 19256 248 19272 312
rect 19336 248 19352 312
rect 19416 248 29112 312
rect 29176 248 29192 312
rect 29256 248 29272 312
rect 29336 248 29352 312
rect 29416 248 41376 312
rect 41440 248 41456 312
rect 41520 248 41536 312
rect 41600 248 41616 312
rect 41680 248 41696 312
rect 41760 248 41776 312
rect 41840 248 41856 312
rect 41920 248 41936 312
rect 42000 248 42016 312
rect 42080 248 42096 312
rect 42160 248 42176 312
rect 42240 248 42256 312
rect 42320 248 42336 312
rect 42400 248 42416 312
rect 42480 248 42496 312
rect 42560 248 42576 312
rect 42640 248 42656 312
rect 42720 248 42736 312
rect 42800 248 42816 312
rect 42880 248 42896 312
rect 42960 248 42976 312
rect 43040 248 43056 312
rect 43120 248 43136 312
rect 43200 248 43216 312
rect 43280 248 43296 312
rect 43360 248 43376 312
rect 43440 248 43456 312
rect 43520 248 43536 312
rect 43600 248 43616 312
rect 43680 248 43696 312
rect 43760 248 43776 312
rect 43840 248 43856 312
rect 43920 248 43936 312
rect 44000 248 44016 312
rect 44080 248 44096 312
rect 44160 248 44176 312
rect 44240 248 44256 312
rect 44320 248 44336 312
rect 44400 248 44416 312
rect 44480 248 44496 312
rect 44560 248 44576 312
rect 44640 248 44656 312
rect 44720 248 44736 312
rect 44800 248 44816 312
rect 44880 248 44896 312
rect 44960 248 44976 312
rect 45040 248 45056 312
rect 45120 248 45136 312
rect 45200 248 45216 312
rect 45280 248 45296 312
rect 45360 248 45368 312
rect 0 232 45368 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 808 232
rect 872 168 888 232
rect 952 168 968 232
rect 1032 168 1048 232
rect 1112 168 1128 232
rect 1192 168 1208 232
rect 1272 168 1288 232
rect 1352 168 1368 232
rect 1432 168 1448 232
rect 1512 168 1528 232
rect 1592 168 1608 232
rect 1672 168 1688 232
rect 1752 168 1768 232
rect 1832 168 1848 232
rect 1912 168 1928 232
rect 1992 168 2008 232
rect 2072 168 2088 232
rect 2152 168 2168 232
rect 2232 168 2248 232
rect 2312 168 2328 232
rect 2392 168 2408 232
rect 2472 168 2488 232
rect 2552 168 2568 232
rect 2632 168 2648 232
rect 2712 168 2728 232
rect 2792 168 2808 232
rect 2872 168 2888 232
rect 2952 168 2968 232
rect 3032 168 3048 232
rect 3112 168 3128 232
rect 3192 168 3208 232
rect 3272 168 3288 232
rect 3352 168 3368 232
rect 3432 168 3448 232
rect 3512 168 3528 232
rect 3592 168 3608 232
rect 3672 168 3688 232
rect 3752 168 3768 232
rect 3832 168 3848 232
rect 3912 168 3928 232
rect 3992 168 19112 232
rect 19176 168 19192 232
rect 19256 168 19272 232
rect 19336 168 19352 232
rect 19416 168 29112 232
rect 29176 168 29192 232
rect 29256 168 29272 232
rect 29336 168 29352 232
rect 29416 168 41376 232
rect 41440 168 41456 232
rect 41520 168 41536 232
rect 41600 168 41616 232
rect 41680 168 41696 232
rect 41760 168 41776 232
rect 41840 168 41856 232
rect 41920 168 41936 232
rect 42000 168 42016 232
rect 42080 168 42096 232
rect 42160 168 42176 232
rect 42240 168 42256 232
rect 42320 168 42336 232
rect 42400 168 42416 232
rect 42480 168 42496 232
rect 42560 168 42576 232
rect 42640 168 42656 232
rect 42720 168 42736 232
rect 42800 168 42816 232
rect 42880 168 42896 232
rect 42960 168 42976 232
rect 43040 168 43056 232
rect 43120 168 43136 232
rect 43200 168 43216 232
rect 43280 168 43296 232
rect 43360 168 43376 232
rect 43440 168 43456 232
rect 43520 168 43536 232
rect 43600 168 43616 232
rect 43680 168 43696 232
rect 43760 168 43776 232
rect 43840 168 43856 232
rect 43920 168 43936 232
rect 44000 168 44016 232
rect 44080 168 44096 232
rect 44160 168 44176 232
rect 44240 168 44256 232
rect 44320 168 44336 232
rect 44400 168 44416 232
rect 44480 168 44496 232
rect 44560 168 44576 232
rect 44640 168 44656 232
rect 44720 168 44736 232
rect 44800 168 44816 232
rect 44880 168 44896 232
rect 44960 168 44976 232
rect 45040 168 45056 232
rect 45120 168 45136 232
rect 45200 168 45216 232
rect 45280 168 45296 232
rect 45360 168 45368 232
rect 0 152 45368 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 808 152
rect 872 88 888 152
rect 952 88 968 152
rect 1032 88 1048 152
rect 1112 88 1128 152
rect 1192 88 1208 152
rect 1272 88 1288 152
rect 1352 88 1368 152
rect 1432 88 1448 152
rect 1512 88 1528 152
rect 1592 88 1608 152
rect 1672 88 1688 152
rect 1752 88 1768 152
rect 1832 88 1848 152
rect 1912 88 1928 152
rect 1992 88 2008 152
rect 2072 88 2088 152
rect 2152 88 2168 152
rect 2232 88 2248 152
rect 2312 88 2328 152
rect 2392 88 2408 152
rect 2472 88 2488 152
rect 2552 88 2568 152
rect 2632 88 2648 152
rect 2712 88 2728 152
rect 2792 88 2808 152
rect 2872 88 2888 152
rect 2952 88 2968 152
rect 3032 88 3048 152
rect 3112 88 3128 152
rect 3192 88 3208 152
rect 3272 88 3288 152
rect 3352 88 3368 152
rect 3432 88 3448 152
rect 3512 88 3528 152
rect 3592 88 3608 152
rect 3672 88 3688 152
rect 3752 88 3768 152
rect 3832 88 3848 152
rect 3912 88 3928 152
rect 3992 88 19112 152
rect 19176 88 19192 152
rect 19256 88 19272 152
rect 19336 88 19352 152
rect 19416 88 29112 152
rect 29176 88 29192 152
rect 29256 88 29272 152
rect 29336 88 29352 152
rect 29416 88 41376 152
rect 41440 88 41456 152
rect 41520 88 41536 152
rect 41600 88 41616 152
rect 41680 88 41696 152
rect 41760 88 41776 152
rect 41840 88 41856 152
rect 41920 88 41936 152
rect 42000 88 42016 152
rect 42080 88 42096 152
rect 42160 88 42176 152
rect 42240 88 42256 152
rect 42320 88 42336 152
rect 42400 88 42416 152
rect 42480 88 42496 152
rect 42560 88 42576 152
rect 42640 88 42656 152
rect 42720 88 42736 152
rect 42800 88 42816 152
rect 42880 88 42896 152
rect 42960 88 42976 152
rect 43040 88 43056 152
rect 43120 88 43136 152
rect 43200 88 43216 152
rect 43280 88 43296 152
rect 43360 88 43376 152
rect 43440 88 43456 152
rect 43520 88 43536 152
rect 43600 88 43616 152
rect 43680 88 43696 152
rect 43760 88 43776 152
rect 43840 88 43856 152
rect 43920 88 43936 152
rect 44000 88 44016 152
rect 44080 88 44096 152
rect 44160 88 44176 152
rect 44240 88 44256 152
rect 44320 88 44336 152
rect 44400 88 44416 152
rect 44480 88 44496 152
rect 44560 88 44576 152
rect 44640 88 44656 152
rect 44720 88 44736 152
rect 44800 88 44816 152
rect 44880 88 44896 152
rect 44960 88 44976 152
rect 45040 88 45056 152
rect 45120 88 45136 152
rect 45200 88 45216 152
rect 45280 88 45296 152
rect 45360 88 45368 152
rect 0 72 45368 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 808 72
rect 872 8 888 72
rect 952 8 968 72
rect 1032 8 1048 72
rect 1112 8 1128 72
rect 1192 8 1208 72
rect 1272 8 1288 72
rect 1352 8 1368 72
rect 1432 8 1448 72
rect 1512 8 1528 72
rect 1592 8 1608 72
rect 1672 8 1688 72
rect 1752 8 1768 72
rect 1832 8 1848 72
rect 1912 8 1928 72
rect 1992 8 2008 72
rect 2072 8 2088 72
rect 2152 8 2168 72
rect 2232 8 2248 72
rect 2312 8 2328 72
rect 2392 8 2408 72
rect 2472 8 2488 72
rect 2552 8 2568 72
rect 2632 8 2648 72
rect 2712 8 2728 72
rect 2792 8 2808 72
rect 2872 8 2888 72
rect 2952 8 2968 72
rect 3032 8 3048 72
rect 3112 8 3128 72
rect 3192 8 3208 72
rect 3272 8 3288 72
rect 3352 8 3368 72
rect 3432 8 3448 72
rect 3512 8 3528 72
rect 3592 8 3608 72
rect 3672 8 3688 72
rect 3752 8 3768 72
rect 3832 8 3848 72
rect 3912 8 3928 72
rect 3992 8 19112 72
rect 19176 8 19192 72
rect 19256 8 19272 72
rect 19336 8 19352 72
rect 19416 8 29112 72
rect 29176 8 29192 72
rect 29256 8 29272 72
rect 29336 8 29352 72
rect 29416 8 41376 72
rect 41440 8 41456 72
rect 41520 8 41536 72
rect 41600 8 41616 72
rect 41680 8 41696 72
rect 41760 8 41776 72
rect 41840 8 41856 72
rect 41920 8 41936 72
rect 42000 8 42016 72
rect 42080 8 42096 72
rect 42160 8 42176 72
rect 42240 8 42256 72
rect 42320 8 42336 72
rect 42400 8 42416 72
rect 42480 8 42496 72
rect 42560 8 42576 72
rect 42640 8 42656 72
rect 42720 8 42736 72
rect 42800 8 42816 72
rect 42880 8 42896 72
rect 42960 8 42976 72
rect 43040 8 43056 72
rect 43120 8 43136 72
rect 43200 8 43216 72
rect 43280 8 43296 72
rect 43360 8 43376 72
rect 43440 8 43456 72
rect 43520 8 43536 72
rect 43600 8 43616 72
rect 43680 8 43696 72
rect 43760 8 43776 72
rect 43840 8 43856 72
rect 43920 8 43936 72
rect 44000 8 44016 72
rect 44080 8 44096 72
rect 44160 8 44176 72
rect 44240 8 44256 72
rect 44320 8 44336 72
rect 44400 8 44416 72
rect 44480 8 44496 72
rect 44560 8 44576 72
rect 44640 8 44656 72
rect 44720 8 44736 72
rect 44800 8 44816 72
rect 44880 8 44896 72
rect 44960 8 44976 72
rect 45040 8 45056 72
rect 45120 8 45136 72
rect 45200 8 45216 72
rect 45280 8 45296 72
rect 45360 8 45368 72
rect 0 0 45368 8
<< via3 >>
rect 8 45320 72 45384
rect 88 45320 152 45384
rect 168 45320 232 45384
rect 248 45320 312 45384
rect 328 45320 392 45384
rect 408 45320 472 45384
rect 488 45320 552 45384
rect 568 45320 632 45384
rect 648 45320 712 45384
rect 728 45320 792 45384
rect 808 45320 872 45384
rect 888 45320 952 45384
rect 968 45320 1032 45384
rect 1048 45320 1112 45384
rect 1128 45320 1192 45384
rect 1208 45320 1272 45384
rect 1288 45320 1352 45384
rect 1368 45320 1432 45384
rect 1448 45320 1512 45384
rect 1528 45320 1592 45384
rect 1608 45320 1672 45384
rect 1688 45320 1752 45384
rect 1768 45320 1832 45384
rect 1848 45320 1912 45384
rect 1928 45320 1992 45384
rect 2008 45320 2072 45384
rect 2088 45320 2152 45384
rect 2168 45320 2232 45384
rect 2248 45320 2312 45384
rect 2328 45320 2392 45384
rect 2408 45320 2472 45384
rect 2488 45320 2552 45384
rect 2568 45320 2632 45384
rect 2648 45320 2712 45384
rect 2728 45320 2792 45384
rect 2808 45320 2872 45384
rect 2888 45320 2952 45384
rect 2968 45320 3032 45384
rect 3048 45320 3112 45384
rect 3128 45320 3192 45384
rect 3208 45320 3272 45384
rect 3288 45320 3352 45384
rect 3368 45320 3432 45384
rect 3448 45320 3512 45384
rect 3528 45320 3592 45384
rect 3608 45320 3672 45384
rect 3688 45320 3752 45384
rect 3768 45320 3832 45384
rect 3848 45320 3912 45384
rect 3928 45320 3992 45384
rect 19112 45320 19176 45384
rect 19192 45320 19256 45384
rect 19272 45320 19336 45384
rect 19352 45320 19416 45384
rect 29112 45320 29176 45384
rect 29192 45320 29256 45384
rect 29272 45320 29336 45384
rect 29352 45320 29416 45384
rect 41376 45320 41440 45384
rect 41456 45320 41520 45384
rect 41536 45320 41600 45384
rect 41616 45320 41680 45384
rect 41696 45320 41760 45384
rect 41776 45320 41840 45384
rect 41856 45320 41920 45384
rect 41936 45320 42000 45384
rect 42016 45320 42080 45384
rect 42096 45320 42160 45384
rect 42176 45320 42240 45384
rect 42256 45320 42320 45384
rect 42336 45320 42400 45384
rect 42416 45320 42480 45384
rect 42496 45320 42560 45384
rect 42576 45320 42640 45384
rect 42656 45320 42720 45384
rect 42736 45320 42800 45384
rect 42816 45320 42880 45384
rect 42896 45320 42960 45384
rect 42976 45320 43040 45384
rect 43056 45320 43120 45384
rect 43136 45320 43200 45384
rect 43216 45320 43280 45384
rect 43296 45320 43360 45384
rect 43376 45320 43440 45384
rect 43456 45320 43520 45384
rect 43536 45320 43600 45384
rect 43616 45320 43680 45384
rect 43696 45320 43760 45384
rect 43776 45320 43840 45384
rect 43856 45320 43920 45384
rect 43936 45320 44000 45384
rect 44016 45320 44080 45384
rect 44096 45320 44160 45384
rect 44176 45320 44240 45384
rect 44256 45320 44320 45384
rect 44336 45320 44400 45384
rect 44416 45320 44480 45384
rect 44496 45320 44560 45384
rect 44576 45320 44640 45384
rect 44656 45320 44720 45384
rect 44736 45320 44800 45384
rect 44816 45320 44880 45384
rect 44896 45320 44960 45384
rect 44976 45320 45040 45384
rect 45056 45320 45120 45384
rect 45136 45320 45200 45384
rect 45216 45320 45280 45384
rect 45296 45320 45360 45384
rect 8 45240 72 45304
rect 88 45240 152 45304
rect 168 45240 232 45304
rect 248 45240 312 45304
rect 328 45240 392 45304
rect 408 45240 472 45304
rect 488 45240 552 45304
rect 568 45240 632 45304
rect 648 45240 712 45304
rect 728 45240 792 45304
rect 808 45240 872 45304
rect 888 45240 952 45304
rect 968 45240 1032 45304
rect 1048 45240 1112 45304
rect 1128 45240 1192 45304
rect 1208 45240 1272 45304
rect 1288 45240 1352 45304
rect 1368 45240 1432 45304
rect 1448 45240 1512 45304
rect 1528 45240 1592 45304
rect 1608 45240 1672 45304
rect 1688 45240 1752 45304
rect 1768 45240 1832 45304
rect 1848 45240 1912 45304
rect 1928 45240 1992 45304
rect 2008 45240 2072 45304
rect 2088 45240 2152 45304
rect 2168 45240 2232 45304
rect 2248 45240 2312 45304
rect 2328 45240 2392 45304
rect 2408 45240 2472 45304
rect 2488 45240 2552 45304
rect 2568 45240 2632 45304
rect 2648 45240 2712 45304
rect 2728 45240 2792 45304
rect 2808 45240 2872 45304
rect 2888 45240 2952 45304
rect 2968 45240 3032 45304
rect 3048 45240 3112 45304
rect 3128 45240 3192 45304
rect 3208 45240 3272 45304
rect 3288 45240 3352 45304
rect 3368 45240 3432 45304
rect 3448 45240 3512 45304
rect 3528 45240 3592 45304
rect 3608 45240 3672 45304
rect 3688 45240 3752 45304
rect 3768 45240 3832 45304
rect 3848 45240 3912 45304
rect 3928 45240 3992 45304
rect 19112 45240 19176 45304
rect 19192 45240 19256 45304
rect 19272 45240 19336 45304
rect 19352 45240 19416 45304
rect 29112 45240 29176 45304
rect 29192 45240 29256 45304
rect 29272 45240 29336 45304
rect 29352 45240 29416 45304
rect 41376 45240 41440 45304
rect 41456 45240 41520 45304
rect 41536 45240 41600 45304
rect 41616 45240 41680 45304
rect 41696 45240 41760 45304
rect 41776 45240 41840 45304
rect 41856 45240 41920 45304
rect 41936 45240 42000 45304
rect 42016 45240 42080 45304
rect 42096 45240 42160 45304
rect 42176 45240 42240 45304
rect 42256 45240 42320 45304
rect 42336 45240 42400 45304
rect 42416 45240 42480 45304
rect 42496 45240 42560 45304
rect 42576 45240 42640 45304
rect 42656 45240 42720 45304
rect 42736 45240 42800 45304
rect 42816 45240 42880 45304
rect 42896 45240 42960 45304
rect 42976 45240 43040 45304
rect 43056 45240 43120 45304
rect 43136 45240 43200 45304
rect 43216 45240 43280 45304
rect 43296 45240 43360 45304
rect 43376 45240 43440 45304
rect 43456 45240 43520 45304
rect 43536 45240 43600 45304
rect 43616 45240 43680 45304
rect 43696 45240 43760 45304
rect 43776 45240 43840 45304
rect 43856 45240 43920 45304
rect 43936 45240 44000 45304
rect 44016 45240 44080 45304
rect 44096 45240 44160 45304
rect 44176 45240 44240 45304
rect 44256 45240 44320 45304
rect 44336 45240 44400 45304
rect 44416 45240 44480 45304
rect 44496 45240 44560 45304
rect 44576 45240 44640 45304
rect 44656 45240 44720 45304
rect 44736 45240 44800 45304
rect 44816 45240 44880 45304
rect 44896 45240 44960 45304
rect 44976 45240 45040 45304
rect 45056 45240 45120 45304
rect 45136 45240 45200 45304
rect 45216 45240 45280 45304
rect 45296 45240 45360 45304
rect 8 45160 72 45224
rect 88 45160 152 45224
rect 168 45160 232 45224
rect 248 45160 312 45224
rect 328 45160 392 45224
rect 408 45160 472 45224
rect 488 45160 552 45224
rect 568 45160 632 45224
rect 648 45160 712 45224
rect 728 45160 792 45224
rect 808 45160 872 45224
rect 888 45160 952 45224
rect 968 45160 1032 45224
rect 1048 45160 1112 45224
rect 1128 45160 1192 45224
rect 1208 45160 1272 45224
rect 1288 45160 1352 45224
rect 1368 45160 1432 45224
rect 1448 45160 1512 45224
rect 1528 45160 1592 45224
rect 1608 45160 1672 45224
rect 1688 45160 1752 45224
rect 1768 45160 1832 45224
rect 1848 45160 1912 45224
rect 1928 45160 1992 45224
rect 2008 45160 2072 45224
rect 2088 45160 2152 45224
rect 2168 45160 2232 45224
rect 2248 45160 2312 45224
rect 2328 45160 2392 45224
rect 2408 45160 2472 45224
rect 2488 45160 2552 45224
rect 2568 45160 2632 45224
rect 2648 45160 2712 45224
rect 2728 45160 2792 45224
rect 2808 45160 2872 45224
rect 2888 45160 2952 45224
rect 2968 45160 3032 45224
rect 3048 45160 3112 45224
rect 3128 45160 3192 45224
rect 3208 45160 3272 45224
rect 3288 45160 3352 45224
rect 3368 45160 3432 45224
rect 3448 45160 3512 45224
rect 3528 45160 3592 45224
rect 3608 45160 3672 45224
rect 3688 45160 3752 45224
rect 3768 45160 3832 45224
rect 3848 45160 3912 45224
rect 3928 45160 3992 45224
rect 19112 45160 19176 45224
rect 19192 45160 19256 45224
rect 19272 45160 19336 45224
rect 19352 45160 19416 45224
rect 29112 45160 29176 45224
rect 29192 45160 29256 45224
rect 29272 45160 29336 45224
rect 29352 45160 29416 45224
rect 41376 45160 41440 45224
rect 41456 45160 41520 45224
rect 41536 45160 41600 45224
rect 41616 45160 41680 45224
rect 41696 45160 41760 45224
rect 41776 45160 41840 45224
rect 41856 45160 41920 45224
rect 41936 45160 42000 45224
rect 42016 45160 42080 45224
rect 42096 45160 42160 45224
rect 42176 45160 42240 45224
rect 42256 45160 42320 45224
rect 42336 45160 42400 45224
rect 42416 45160 42480 45224
rect 42496 45160 42560 45224
rect 42576 45160 42640 45224
rect 42656 45160 42720 45224
rect 42736 45160 42800 45224
rect 42816 45160 42880 45224
rect 42896 45160 42960 45224
rect 42976 45160 43040 45224
rect 43056 45160 43120 45224
rect 43136 45160 43200 45224
rect 43216 45160 43280 45224
rect 43296 45160 43360 45224
rect 43376 45160 43440 45224
rect 43456 45160 43520 45224
rect 43536 45160 43600 45224
rect 43616 45160 43680 45224
rect 43696 45160 43760 45224
rect 43776 45160 43840 45224
rect 43856 45160 43920 45224
rect 43936 45160 44000 45224
rect 44016 45160 44080 45224
rect 44096 45160 44160 45224
rect 44176 45160 44240 45224
rect 44256 45160 44320 45224
rect 44336 45160 44400 45224
rect 44416 45160 44480 45224
rect 44496 45160 44560 45224
rect 44576 45160 44640 45224
rect 44656 45160 44720 45224
rect 44736 45160 44800 45224
rect 44816 45160 44880 45224
rect 44896 45160 44960 45224
rect 44976 45160 45040 45224
rect 45056 45160 45120 45224
rect 45136 45160 45200 45224
rect 45216 45160 45280 45224
rect 45296 45160 45360 45224
rect 8 45080 72 45144
rect 88 45080 152 45144
rect 168 45080 232 45144
rect 248 45080 312 45144
rect 328 45080 392 45144
rect 408 45080 472 45144
rect 488 45080 552 45144
rect 568 45080 632 45144
rect 648 45080 712 45144
rect 728 45080 792 45144
rect 808 45080 872 45144
rect 888 45080 952 45144
rect 968 45080 1032 45144
rect 1048 45080 1112 45144
rect 1128 45080 1192 45144
rect 1208 45080 1272 45144
rect 1288 45080 1352 45144
rect 1368 45080 1432 45144
rect 1448 45080 1512 45144
rect 1528 45080 1592 45144
rect 1608 45080 1672 45144
rect 1688 45080 1752 45144
rect 1768 45080 1832 45144
rect 1848 45080 1912 45144
rect 1928 45080 1992 45144
rect 2008 45080 2072 45144
rect 2088 45080 2152 45144
rect 2168 45080 2232 45144
rect 2248 45080 2312 45144
rect 2328 45080 2392 45144
rect 2408 45080 2472 45144
rect 2488 45080 2552 45144
rect 2568 45080 2632 45144
rect 2648 45080 2712 45144
rect 2728 45080 2792 45144
rect 2808 45080 2872 45144
rect 2888 45080 2952 45144
rect 2968 45080 3032 45144
rect 3048 45080 3112 45144
rect 3128 45080 3192 45144
rect 3208 45080 3272 45144
rect 3288 45080 3352 45144
rect 3368 45080 3432 45144
rect 3448 45080 3512 45144
rect 3528 45080 3592 45144
rect 3608 45080 3672 45144
rect 3688 45080 3752 45144
rect 3768 45080 3832 45144
rect 3848 45080 3912 45144
rect 3928 45080 3992 45144
rect 19112 45080 19176 45144
rect 19192 45080 19256 45144
rect 19272 45080 19336 45144
rect 19352 45080 19416 45144
rect 29112 45080 29176 45144
rect 29192 45080 29256 45144
rect 29272 45080 29336 45144
rect 29352 45080 29416 45144
rect 41376 45080 41440 45144
rect 41456 45080 41520 45144
rect 41536 45080 41600 45144
rect 41616 45080 41680 45144
rect 41696 45080 41760 45144
rect 41776 45080 41840 45144
rect 41856 45080 41920 45144
rect 41936 45080 42000 45144
rect 42016 45080 42080 45144
rect 42096 45080 42160 45144
rect 42176 45080 42240 45144
rect 42256 45080 42320 45144
rect 42336 45080 42400 45144
rect 42416 45080 42480 45144
rect 42496 45080 42560 45144
rect 42576 45080 42640 45144
rect 42656 45080 42720 45144
rect 42736 45080 42800 45144
rect 42816 45080 42880 45144
rect 42896 45080 42960 45144
rect 42976 45080 43040 45144
rect 43056 45080 43120 45144
rect 43136 45080 43200 45144
rect 43216 45080 43280 45144
rect 43296 45080 43360 45144
rect 43376 45080 43440 45144
rect 43456 45080 43520 45144
rect 43536 45080 43600 45144
rect 43616 45080 43680 45144
rect 43696 45080 43760 45144
rect 43776 45080 43840 45144
rect 43856 45080 43920 45144
rect 43936 45080 44000 45144
rect 44016 45080 44080 45144
rect 44096 45080 44160 45144
rect 44176 45080 44240 45144
rect 44256 45080 44320 45144
rect 44336 45080 44400 45144
rect 44416 45080 44480 45144
rect 44496 45080 44560 45144
rect 44576 45080 44640 45144
rect 44656 45080 44720 45144
rect 44736 45080 44800 45144
rect 44816 45080 44880 45144
rect 44896 45080 44960 45144
rect 44976 45080 45040 45144
rect 45056 45080 45120 45144
rect 45136 45080 45200 45144
rect 45216 45080 45280 45144
rect 45296 45080 45360 45144
rect 8 45000 72 45064
rect 88 45000 152 45064
rect 168 45000 232 45064
rect 248 45000 312 45064
rect 328 45000 392 45064
rect 408 45000 472 45064
rect 488 45000 552 45064
rect 568 45000 632 45064
rect 648 45000 712 45064
rect 728 45000 792 45064
rect 808 45000 872 45064
rect 888 45000 952 45064
rect 968 45000 1032 45064
rect 1048 45000 1112 45064
rect 1128 45000 1192 45064
rect 1208 45000 1272 45064
rect 1288 45000 1352 45064
rect 1368 45000 1432 45064
rect 1448 45000 1512 45064
rect 1528 45000 1592 45064
rect 1608 45000 1672 45064
rect 1688 45000 1752 45064
rect 1768 45000 1832 45064
rect 1848 45000 1912 45064
rect 1928 45000 1992 45064
rect 2008 45000 2072 45064
rect 2088 45000 2152 45064
rect 2168 45000 2232 45064
rect 2248 45000 2312 45064
rect 2328 45000 2392 45064
rect 2408 45000 2472 45064
rect 2488 45000 2552 45064
rect 2568 45000 2632 45064
rect 2648 45000 2712 45064
rect 2728 45000 2792 45064
rect 2808 45000 2872 45064
rect 2888 45000 2952 45064
rect 2968 45000 3032 45064
rect 3048 45000 3112 45064
rect 3128 45000 3192 45064
rect 3208 45000 3272 45064
rect 3288 45000 3352 45064
rect 3368 45000 3432 45064
rect 3448 45000 3512 45064
rect 3528 45000 3592 45064
rect 3608 45000 3672 45064
rect 3688 45000 3752 45064
rect 3768 45000 3832 45064
rect 3848 45000 3912 45064
rect 3928 45000 3992 45064
rect 19112 45000 19176 45064
rect 19192 45000 19256 45064
rect 19272 45000 19336 45064
rect 19352 45000 19416 45064
rect 29112 45000 29176 45064
rect 29192 45000 29256 45064
rect 29272 45000 29336 45064
rect 29352 45000 29416 45064
rect 41376 45000 41440 45064
rect 41456 45000 41520 45064
rect 41536 45000 41600 45064
rect 41616 45000 41680 45064
rect 41696 45000 41760 45064
rect 41776 45000 41840 45064
rect 41856 45000 41920 45064
rect 41936 45000 42000 45064
rect 42016 45000 42080 45064
rect 42096 45000 42160 45064
rect 42176 45000 42240 45064
rect 42256 45000 42320 45064
rect 42336 45000 42400 45064
rect 42416 45000 42480 45064
rect 42496 45000 42560 45064
rect 42576 45000 42640 45064
rect 42656 45000 42720 45064
rect 42736 45000 42800 45064
rect 42816 45000 42880 45064
rect 42896 45000 42960 45064
rect 42976 45000 43040 45064
rect 43056 45000 43120 45064
rect 43136 45000 43200 45064
rect 43216 45000 43280 45064
rect 43296 45000 43360 45064
rect 43376 45000 43440 45064
rect 43456 45000 43520 45064
rect 43536 45000 43600 45064
rect 43616 45000 43680 45064
rect 43696 45000 43760 45064
rect 43776 45000 43840 45064
rect 43856 45000 43920 45064
rect 43936 45000 44000 45064
rect 44016 45000 44080 45064
rect 44096 45000 44160 45064
rect 44176 45000 44240 45064
rect 44256 45000 44320 45064
rect 44336 45000 44400 45064
rect 44416 45000 44480 45064
rect 44496 45000 44560 45064
rect 44576 45000 44640 45064
rect 44656 45000 44720 45064
rect 44736 45000 44800 45064
rect 44816 45000 44880 45064
rect 44896 45000 44960 45064
rect 44976 45000 45040 45064
rect 45056 45000 45120 45064
rect 45136 45000 45200 45064
rect 45216 45000 45280 45064
rect 45296 45000 45360 45064
rect 8 44920 72 44984
rect 88 44920 152 44984
rect 168 44920 232 44984
rect 248 44920 312 44984
rect 328 44920 392 44984
rect 408 44920 472 44984
rect 488 44920 552 44984
rect 568 44920 632 44984
rect 648 44920 712 44984
rect 728 44920 792 44984
rect 808 44920 872 44984
rect 888 44920 952 44984
rect 968 44920 1032 44984
rect 1048 44920 1112 44984
rect 1128 44920 1192 44984
rect 1208 44920 1272 44984
rect 1288 44920 1352 44984
rect 1368 44920 1432 44984
rect 1448 44920 1512 44984
rect 1528 44920 1592 44984
rect 1608 44920 1672 44984
rect 1688 44920 1752 44984
rect 1768 44920 1832 44984
rect 1848 44920 1912 44984
rect 1928 44920 1992 44984
rect 2008 44920 2072 44984
rect 2088 44920 2152 44984
rect 2168 44920 2232 44984
rect 2248 44920 2312 44984
rect 2328 44920 2392 44984
rect 2408 44920 2472 44984
rect 2488 44920 2552 44984
rect 2568 44920 2632 44984
rect 2648 44920 2712 44984
rect 2728 44920 2792 44984
rect 2808 44920 2872 44984
rect 2888 44920 2952 44984
rect 2968 44920 3032 44984
rect 3048 44920 3112 44984
rect 3128 44920 3192 44984
rect 3208 44920 3272 44984
rect 3288 44920 3352 44984
rect 3368 44920 3432 44984
rect 3448 44920 3512 44984
rect 3528 44920 3592 44984
rect 3608 44920 3672 44984
rect 3688 44920 3752 44984
rect 3768 44920 3832 44984
rect 3848 44920 3912 44984
rect 3928 44920 3992 44984
rect 19112 44920 19176 44984
rect 19192 44920 19256 44984
rect 19272 44920 19336 44984
rect 19352 44920 19416 44984
rect 29112 44920 29176 44984
rect 29192 44920 29256 44984
rect 29272 44920 29336 44984
rect 29352 44920 29416 44984
rect 41376 44920 41440 44984
rect 41456 44920 41520 44984
rect 41536 44920 41600 44984
rect 41616 44920 41680 44984
rect 41696 44920 41760 44984
rect 41776 44920 41840 44984
rect 41856 44920 41920 44984
rect 41936 44920 42000 44984
rect 42016 44920 42080 44984
rect 42096 44920 42160 44984
rect 42176 44920 42240 44984
rect 42256 44920 42320 44984
rect 42336 44920 42400 44984
rect 42416 44920 42480 44984
rect 42496 44920 42560 44984
rect 42576 44920 42640 44984
rect 42656 44920 42720 44984
rect 42736 44920 42800 44984
rect 42816 44920 42880 44984
rect 42896 44920 42960 44984
rect 42976 44920 43040 44984
rect 43056 44920 43120 44984
rect 43136 44920 43200 44984
rect 43216 44920 43280 44984
rect 43296 44920 43360 44984
rect 43376 44920 43440 44984
rect 43456 44920 43520 44984
rect 43536 44920 43600 44984
rect 43616 44920 43680 44984
rect 43696 44920 43760 44984
rect 43776 44920 43840 44984
rect 43856 44920 43920 44984
rect 43936 44920 44000 44984
rect 44016 44920 44080 44984
rect 44096 44920 44160 44984
rect 44176 44920 44240 44984
rect 44256 44920 44320 44984
rect 44336 44920 44400 44984
rect 44416 44920 44480 44984
rect 44496 44920 44560 44984
rect 44576 44920 44640 44984
rect 44656 44920 44720 44984
rect 44736 44920 44800 44984
rect 44816 44920 44880 44984
rect 44896 44920 44960 44984
rect 44976 44920 45040 44984
rect 45056 44920 45120 44984
rect 45136 44920 45200 44984
rect 45216 44920 45280 44984
rect 45296 44920 45360 44984
rect 8 44840 72 44904
rect 88 44840 152 44904
rect 168 44840 232 44904
rect 248 44840 312 44904
rect 328 44840 392 44904
rect 408 44840 472 44904
rect 488 44840 552 44904
rect 568 44840 632 44904
rect 648 44840 712 44904
rect 728 44840 792 44904
rect 808 44840 872 44904
rect 888 44840 952 44904
rect 968 44840 1032 44904
rect 1048 44840 1112 44904
rect 1128 44840 1192 44904
rect 1208 44840 1272 44904
rect 1288 44840 1352 44904
rect 1368 44840 1432 44904
rect 1448 44840 1512 44904
rect 1528 44840 1592 44904
rect 1608 44840 1672 44904
rect 1688 44840 1752 44904
rect 1768 44840 1832 44904
rect 1848 44840 1912 44904
rect 1928 44840 1992 44904
rect 2008 44840 2072 44904
rect 2088 44840 2152 44904
rect 2168 44840 2232 44904
rect 2248 44840 2312 44904
rect 2328 44840 2392 44904
rect 2408 44840 2472 44904
rect 2488 44840 2552 44904
rect 2568 44840 2632 44904
rect 2648 44840 2712 44904
rect 2728 44840 2792 44904
rect 2808 44840 2872 44904
rect 2888 44840 2952 44904
rect 2968 44840 3032 44904
rect 3048 44840 3112 44904
rect 3128 44840 3192 44904
rect 3208 44840 3272 44904
rect 3288 44840 3352 44904
rect 3368 44840 3432 44904
rect 3448 44840 3512 44904
rect 3528 44840 3592 44904
rect 3608 44840 3672 44904
rect 3688 44840 3752 44904
rect 3768 44840 3832 44904
rect 3848 44840 3912 44904
rect 3928 44840 3992 44904
rect 19112 44840 19176 44904
rect 19192 44840 19256 44904
rect 19272 44840 19336 44904
rect 19352 44840 19416 44904
rect 29112 44840 29176 44904
rect 29192 44840 29256 44904
rect 29272 44840 29336 44904
rect 29352 44840 29416 44904
rect 41376 44840 41440 44904
rect 41456 44840 41520 44904
rect 41536 44840 41600 44904
rect 41616 44840 41680 44904
rect 41696 44840 41760 44904
rect 41776 44840 41840 44904
rect 41856 44840 41920 44904
rect 41936 44840 42000 44904
rect 42016 44840 42080 44904
rect 42096 44840 42160 44904
rect 42176 44840 42240 44904
rect 42256 44840 42320 44904
rect 42336 44840 42400 44904
rect 42416 44840 42480 44904
rect 42496 44840 42560 44904
rect 42576 44840 42640 44904
rect 42656 44840 42720 44904
rect 42736 44840 42800 44904
rect 42816 44840 42880 44904
rect 42896 44840 42960 44904
rect 42976 44840 43040 44904
rect 43056 44840 43120 44904
rect 43136 44840 43200 44904
rect 43216 44840 43280 44904
rect 43296 44840 43360 44904
rect 43376 44840 43440 44904
rect 43456 44840 43520 44904
rect 43536 44840 43600 44904
rect 43616 44840 43680 44904
rect 43696 44840 43760 44904
rect 43776 44840 43840 44904
rect 43856 44840 43920 44904
rect 43936 44840 44000 44904
rect 44016 44840 44080 44904
rect 44096 44840 44160 44904
rect 44176 44840 44240 44904
rect 44256 44840 44320 44904
rect 44336 44840 44400 44904
rect 44416 44840 44480 44904
rect 44496 44840 44560 44904
rect 44576 44840 44640 44904
rect 44656 44840 44720 44904
rect 44736 44840 44800 44904
rect 44816 44840 44880 44904
rect 44896 44840 44960 44904
rect 44976 44840 45040 44904
rect 45056 44840 45120 44904
rect 45136 44840 45200 44904
rect 45216 44840 45280 44904
rect 45296 44840 45360 44904
rect 8 44760 72 44824
rect 88 44760 152 44824
rect 168 44760 232 44824
rect 248 44760 312 44824
rect 328 44760 392 44824
rect 408 44760 472 44824
rect 488 44760 552 44824
rect 568 44760 632 44824
rect 648 44760 712 44824
rect 728 44760 792 44824
rect 808 44760 872 44824
rect 888 44760 952 44824
rect 968 44760 1032 44824
rect 1048 44760 1112 44824
rect 1128 44760 1192 44824
rect 1208 44760 1272 44824
rect 1288 44760 1352 44824
rect 1368 44760 1432 44824
rect 1448 44760 1512 44824
rect 1528 44760 1592 44824
rect 1608 44760 1672 44824
rect 1688 44760 1752 44824
rect 1768 44760 1832 44824
rect 1848 44760 1912 44824
rect 1928 44760 1992 44824
rect 2008 44760 2072 44824
rect 2088 44760 2152 44824
rect 2168 44760 2232 44824
rect 2248 44760 2312 44824
rect 2328 44760 2392 44824
rect 2408 44760 2472 44824
rect 2488 44760 2552 44824
rect 2568 44760 2632 44824
rect 2648 44760 2712 44824
rect 2728 44760 2792 44824
rect 2808 44760 2872 44824
rect 2888 44760 2952 44824
rect 2968 44760 3032 44824
rect 3048 44760 3112 44824
rect 3128 44760 3192 44824
rect 3208 44760 3272 44824
rect 3288 44760 3352 44824
rect 3368 44760 3432 44824
rect 3448 44760 3512 44824
rect 3528 44760 3592 44824
rect 3608 44760 3672 44824
rect 3688 44760 3752 44824
rect 3768 44760 3832 44824
rect 3848 44760 3912 44824
rect 3928 44760 3992 44824
rect 19112 44760 19176 44824
rect 19192 44760 19256 44824
rect 19272 44760 19336 44824
rect 19352 44760 19416 44824
rect 29112 44760 29176 44824
rect 29192 44760 29256 44824
rect 29272 44760 29336 44824
rect 29352 44760 29416 44824
rect 41376 44760 41440 44824
rect 41456 44760 41520 44824
rect 41536 44760 41600 44824
rect 41616 44760 41680 44824
rect 41696 44760 41760 44824
rect 41776 44760 41840 44824
rect 41856 44760 41920 44824
rect 41936 44760 42000 44824
rect 42016 44760 42080 44824
rect 42096 44760 42160 44824
rect 42176 44760 42240 44824
rect 42256 44760 42320 44824
rect 42336 44760 42400 44824
rect 42416 44760 42480 44824
rect 42496 44760 42560 44824
rect 42576 44760 42640 44824
rect 42656 44760 42720 44824
rect 42736 44760 42800 44824
rect 42816 44760 42880 44824
rect 42896 44760 42960 44824
rect 42976 44760 43040 44824
rect 43056 44760 43120 44824
rect 43136 44760 43200 44824
rect 43216 44760 43280 44824
rect 43296 44760 43360 44824
rect 43376 44760 43440 44824
rect 43456 44760 43520 44824
rect 43536 44760 43600 44824
rect 43616 44760 43680 44824
rect 43696 44760 43760 44824
rect 43776 44760 43840 44824
rect 43856 44760 43920 44824
rect 43936 44760 44000 44824
rect 44016 44760 44080 44824
rect 44096 44760 44160 44824
rect 44176 44760 44240 44824
rect 44256 44760 44320 44824
rect 44336 44760 44400 44824
rect 44416 44760 44480 44824
rect 44496 44760 44560 44824
rect 44576 44760 44640 44824
rect 44656 44760 44720 44824
rect 44736 44760 44800 44824
rect 44816 44760 44880 44824
rect 44896 44760 44960 44824
rect 44976 44760 45040 44824
rect 45056 44760 45120 44824
rect 45136 44760 45200 44824
rect 45216 44760 45280 44824
rect 45296 44760 45360 44824
rect 8 44680 72 44744
rect 88 44680 152 44744
rect 168 44680 232 44744
rect 248 44680 312 44744
rect 328 44680 392 44744
rect 408 44680 472 44744
rect 488 44680 552 44744
rect 568 44680 632 44744
rect 648 44680 712 44744
rect 728 44680 792 44744
rect 808 44680 872 44744
rect 888 44680 952 44744
rect 968 44680 1032 44744
rect 1048 44680 1112 44744
rect 1128 44680 1192 44744
rect 1208 44680 1272 44744
rect 1288 44680 1352 44744
rect 1368 44680 1432 44744
rect 1448 44680 1512 44744
rect 1528 44680 1592 44744
rect 1608 44680 1672 44744
rect 1688 44680 1752 44744
rect 1768 44680 1832 44744
rect 1848 44680 1912 44744
rect 1928 44680 1992 44744
rect 2008 44680 2072 44744
rect 2088 44680 2152 44744
rect 2168 44680 2232 44744
rect 2248 44680 2312 44744
rect 2328 44680 2392 44744
rect 2408 44680 2472 44744
rect 2488 44680 2552 44744
rect 2568 44680 2632 44744
rect 2648 44680 2712 44744
rect 2728 44680 2792 44744
rect 2808 44680 2872 44744
rect 2888 44680 2952 44744
rect 2968 44680 3032 44744
rect 3048 44680 3112 44744
rect 3128 44680 3192 44744
rect 3208 44680 3272 44744
rect 3288 44680 3352 44744
rect 3368 44680 3432 44744
rect 3448 44680 3512 44744
rect 3528 44680 3592 44744
rect 3608 44680 3672 44744
rect 3688 44680 3752 44744
rect 3768 44680 3832 44744
rect 3848 44680 3912 44744
rect 3928 44680 3992 44744
rect 19112 44680 19176 44744
rect 19192 44680 19256 44744
rect 19272 44680 19336 44744
rect 19352 44680 19416 44744
rect 29112 44680 29176 44744
rect 29192 44680 29256 44744
rect 29272 44680 29336 44744
rect 29352 44680 29416 44744
rect 41376 44680 41440 44744
rect 41456 44680 41520 44744
rect 41536 44680 41600 44744
rect 41616 44680 41680 44744
rect 41696 44680 41760 44744
rect 41776 44680 41840 44744
rect 41856 44680 41920 44744
rect 41936 44680 42000 44744
rect 42016 44680 42080 44744
rect 42096 44680 42160 44744
rect 42176 44680 42240 44744
rect 42256 44680 42320 44744
rect 42336 44680 42400 44744
rect 42416 44680 42480 44744
rect 42496 44680 42560 44744
rect 42576 44680 42640 44744
rect 42656 44680 42720 44744
rect 42736 44680 42800 44744
rect 42816 44680 42880 44744
rect 42896 44680 42960 44744
rect 42976 44680 43040 44744
rect 43056 44680 43120 44744
rect 43136 44680 43200 44744
rect 43216 44680 43280 44744
rect 43296 44680 43360 44744
rect 43376 44680 43440 44744
rect 43456 44680 43520 44744
rect 43536 44680 43600 44744
rect 43616 44680 43680 44744
rect 43696 44680 43760 44744
rect 43776 44680 43840 44744
rect 43856 44680 43920 44744
rect 43936 44680 44000 44744
rect 44016 44680 44080 44744
rect 44096 44680 44160 44744
rect 44176 44680 44240 44744
rect 44256 44680 44320 44744
rect 44336 44680 44400 44744
rect 44416 44680 44480 44744
rect 44496 44680 44560 44744
rect 44576 44680 44640 44744
rect 44656 44680 44720 44744
rect 44736 44680 44800 44744
rect 44816 44680 44880 44744
rect 44896 44680 44960 44744
rect 44976 44680 45040 44744
rect 45056 44680 45120 44744
rect 45136 44680 45200 44744
rect 45216 44680 45280 44744
rect 45296 44680 45360 44744
rect 8 44600 72 44664
rect 88 44600 152 44664
rect 168 44600 232 44664
rect 248 44600 312 44664
rect 328 44600 392 44664
rect 408 44600 472 44664
rect 488 44600 552 44664
rect 568 44600 632 44664
rect 648 44600 712 44664
rect 728 44600 792 44664
rect 808 44600 872 44664
rect 888 44600 952 44664
rect 968 44600 1032 44664
rect 1048 44600 1112 44664
rect 1128 44600 1192 44664
rect 1208 44600 1272 44664
rect 1288 44600 1352 44664
rect 1368 44600 1432 44664
rect 1448 44600 1512 44664
rect 1528 44600 1592 44664
rect 1608 44600 1672 44664
rect 1688 44600 1752 44664
rect 1768 44600 1832 44664
rect 1848 44600 1912 44664
rect 1928 44600 1992 44664
rect 2008 44600 2072 44664
rect 2088 44600 2152 44664
rect 2168 44600 2232 44664
rect 2248 44600 2312 44664
rect 2328 44600 2392 44664
rect 2408 44600 2472 44664
rect 2488 44600 2552 44664
rect 2568 44600 2632 44664
rect 2648 44600 2712 44664
rect 2728 44600 2792 44664
rect 2808 44600 2872 44664
rect 2888 44600 2952 44664
rect 2968 44600 3032 44664
rect 3048 44600 3112 44664
rect 3128 44600 3192 44664
rect 3208 44600 3272 44664
rect 3288 44600 3352 44664
rect 3368 44600 3432 44664
rect 3448 44600 3512 44664
rect 3528 44600 3592 44664
rect 3608 44600 3672 44664
rect 3688 44600 3752 44664
rect 3768 44600 3832 44664
rect 3848 44600 3912 44664
rect 3928 44600 3992 44664
rect 19112 44600 19176 44664
rect 19192 44600 19256 44664
rect 19272 44600 19336 44664
rect 19352 44600 19416 44664
rect 29112 44600 29176 44664
rect 29192 44600 29256 44664
rect 29272 44600 29336 44664
rect 29352 44600 29416 44664
rect 41376 44600 41440 44664
rect 41456 44600 41520 44664
rect 41536 44600 41600 44664
rect 41616 44600 41680 44664
rect 41696 44600 41760 44664
rect 41776 44600 41840 44664
rect 41856 44600 41920 44664
rect 41936 44600 42000 44664
rect 42016 44600 42080 44664
rect 42096 44600 42160 44664
rect 42176 44600 42240 44664
rect 42256 44600 42320 44664
rect 42336 44600 42400 44664
rect 42416 44600 42480 44664
rect 42496 44600 42560 44664
rect 42576 44600 42640 44664
rect 42656 44600 42720 44664
rect 42736 44600 42800 44664
rect 42816 44600 42880 44664
rect 42896 44600 42960 44664
rect 42976 44600 43040 44664
rect 43056 44600 43120 44664
rect 43136 44600 43200 44664
rect 43216 44600 43280 44664
rect 43296 44600 43360 44664
rect 43376 44600 43440 44664
rect 43456 44600 43520 44664
rect 43536 44600 43600 44664
rect 43616 44600 43680 44664
rect 43696 44600 43760 44664
rect 43776 44600 43840 44664
rect 43856 44600 43920 44664
rect 43936 44600 44000 44664
rect 44016 44600 44080 44664
rect 44096 44600 44160 44664
rect 44176 44600 44240 44664
rect 44256 44600 44320 44664
rect 44336 44600 44400 44664
rect 44416 44600 44480 44664
rect 44496 44600 44560 44664
rect 44576 44600 44640 44664
rect 44656 44600 44720 44664
rect 44736 44600 44800 44664
rect 44816 44600 44880 44664
rect 44896 44600 44960 44664
rect 44976 44600 45040 44664
rect 45056 44600 45120 44664
rect 45136 44600 45200 44664
rect 45216 44600 45280 44664
rect 45296 44600 45360 44664
rect 8 44520 72 44584
rect 88 44520 152 44584
rect 168 44520 232 44584
rect 248 44520 312 44584
rect 328 44520 392 44584
rect 408 44520 472 44584
rect 488 44520 552 44584
rect 568 44520 632 44584
rect 648 44520 712 44584
rect 728 44520 792 44584
rect 808 44520 872 44584
rect 888 44520 952 44584
rect 968 44520 1032 44584
rect 1048 44520 1112 44584
rect 1128 44520 1192 44584
rect 1208 44520 1272 44584
rect 1288 44520 1352 44584
rect 1368 44520 1432 44584
rect 1448 44520 1512 44584
rect 1528 44520 1592 44584
rect 1608 44520 1672 44584
rect 1688 44520 1752 44584
rect 1768 44520 1832 44584
rect 1848 44520 1912 44584
rect 1928 44520 1992 44584
rect 2008 44520 2072 44584
rect 2088 44520 2152 44584
rect 2168 44520 2232 44584
rect 2248 44520 2312 44584
rect 2328 44520 2392 44584
rect 2408 44520 2472 44584
rect 2488 44520 2552 44584
rect 2568 44520 2632 44584
rect 2648 44520 2712 44584
rect 2728 44520 2792 44584
rect 2808 44520 2872 44584
rect 2888 44520 2952 44584
rect 2968 44520 3032 44584
rect 3048 44520 3112 44584
rect 3128 44520 3192 44584
rect 3208 44520 3272 44584
rect 3288 44520 3352 44584
rect 3368 44520 3432 44584
rect 3448 44520 3512 44584
rect 3528 44520 3592 44584
rect 3608 44520 3672 44584
rect 3688 44520 3752 44584
rect 3768 44520 3832 44584
rect 3848 44520 3912 44584
rect 3928 44520 3992 44584
rect 19112 44520 19176 44584
rect 19192 44520 19256 44584
rect 19272 44520 19336 44584
rect 19352 44520 19416 44584
rect 29112 44520 29176 44584
rect 29192 44520 29256 44584
rect 29272 44520 29336 44584
rect 29352 44520 29416 44584
rect 41376 44520 41440 44584
rect 41456 44520 41520 44584
rect 41536 44520 41600 44584
rect 41616 44520 41680 44584
rect 41696 44520 41760 44584
rect 41776 44520 41840 44584
rect 41856 44520 41920 44584
rect 41936 44520 42000 44584
rect 42016 44520 42080 44584
rect 42096 44520 42160 44584
rect 42176 44520 42240 44584
rect 42256 44520 42320 44584
rect 42336 44520 42400 44584
rect 42416 44520 42480 44584
rect 42496 44520 42560 44584
rect 42576 44520 42640 44584
rect 42656 44520 42720 44584
rect 42736 44520 42800 44584
rect 42816 44520 42880 44584
rect 42896 44520 42960 44584
rect 42976 44520 43040 44584
rect 43056 44520 43120 44584
rect 43136 44520 43200 44584
rect 43216 44520 43280 44584
rect 43296 44520 43360 44584
rect 43376 44520 43440 44584
rect 43456 44520 43520 44584
rect 43536 44520 43600 44584
rect 43616 44520 43680 44584
rect 43696 44520 43760 44584
rect 43776 44520 43840 44584
rect 43856 44520 43920 44584
rect 43936 44520 44000 44584
rect 44016 44520 44080 44584
rect 44096 44520 44160 44584
rect 44176 44520 44240 44584
rect 44256 44520 44320 44584
rect 44336 44520 44400 44584
rect 44416 44520 44480 44584
rect 44496 44520 44560 44584
rect 44576 44520 44640 44584
rect 44656 44520 44720 44584
rect 44736 44520 44800 44584
rect 44816 44520 44880 44584
rect 44896 44520 44960 44584
rect 44976 44520 45040 44584
rect 45056 44520 45120 44584
rect 45136 44520 45200 44584
rect 45216 44520 45280 44584
rect 45296 44520 45360 44584
rect 8 44440 72 44504
rect 88 44440 152 44504
rect 168 44440 232 44504
rect 248 44440 312 44504
rect 328 44440 392 44504
rect 408 44440 472 44504
rect 488 44440 552 44504
rect 568 44440 632 44504
rect 648 44440 712 44504
rect 728 44440 792 44504
rect 808 44440 872 44504
rect 888 44440 952 44504
rect 968 44440 1032 44504
rect 1048 44440 1112 44504
rect 1128 44440 1192 44504
rect 1208 44440 1272 44504
rect 1288 44440 1352 44504
rect 1368 44440 1432 44504
rect 1448 44440 1512 44504
rect 1528 44440 1592 44504
rect 1608 44440 1672 44504
rect 1688 44440 1752 44504
rect 1768 44440 1832 44504
rect 1848 44440 1912 44504
rect 1928 44440 1992 44504
rect 2008 44440 2072 44504
rect 2088 44440 2152 44504
rect 2168 44440 2232 44504
rect 2248 44440 2312 44504
rect 2328 44440 2392 44504
rect 2408 44440 2472 44504
rect 2488 44440 2552 44504
rect 2568 44440 2632 44504
rect 2648 44440 2712 44504
rect 2728 44440 2792 44504
rect 2808 44440 2872 44504
rect 2888 44440 2952 44504
rect 2968 44440 3032 44504
rect 3048 44440 3112 44504
rect 3128 44440 3192 44504
rect 3208 44440 3272 44504
rect 3288 44440 3352 44504
rect 3368 44440 3432 44504
rect 3448 44440 3512 44504
rect 3528 44440 3592 44504
rect 3608 44440 3672 44504
rect 3688 44440 3752 44504
rect 3768 44440 3832 44504
rect 3848 44440 3912 44504
rect 3928 44440 3992 44504
rect 19112 44440 19176 44504
rect 19192 44440 19256 44504
rect 19272 44440 19336 44504
rect 19352 44440 19416 44504
rect 29112 44440 29176 44504
rect 29192 44440 29256 44504
rect 29272 44440 29336 44504
rect 29352 44440 29416 44504
rect 41376 44440 41440 44504
rect 41456 44440 41520 44504
rect 41536 44440 41600 44504
rect 41616 44440 41680 44504
rect 41696 44440 41760 44504
rect 41776 44440 41840 44504
rect 41856 44440 41920 44504
rect 41936 44440 42000 44504
rect 42016 44440 42080 44504
rect 42096 44440 42160 44504
rect 42176 44440 42240 44504
rect 42256 44440 42320 44504
rect 42336 44440 42400 44504
rect 42416 44440 42480 44504
rect 42496 44440 42560 44504
rect 42576 44440 42640 44504
rect 42656 44440 42720 44504
rect 42736 44440 42800 44504
rect 42816 44440 42880 44504
rect 42896 44440 42960 44504
rect 42976 44440 43040 44504
rect 43056 44440 43120 44504
rect 43136 44440 43200 44504
rect 43216 44440 43280 44504
rect 43296 44440 43360 44504
rect 43376 44440 43440 44504
rect 43456 44440 43520 44504
rect 43536 44440 43600 44504
rect 43616 44440 43680 44504
rect 43696 44440 43760 44504
rect 43776 44440 43840 44504
rect 43856 44440 43920 44504
rect 43936 44440 44000 44504
rect 44016 44440 44080 44504
rect 44096 44440 44160 44504
rect 44176 44440 44240 44504
rect 44256 44440 44320 44504
rect 44336 44440 44400 44504
rect 44416 44440 44480 44504
rect 44496 44440 44560 44504
rect 44576 44440 44640 44504
rect 44656 44440 44720 44504
rect 44736 44440 44800 44504
rect 44816 44440 44880 44504
rect 44896 44440 44960 44504
rect 44976 44440 45040 44504
rect 45056 44440 45120 44504
rect 45136 44440 45200 44504
rect 45216 44440 45280 44504
rect 45296 44440 45360 44504
rect 8 44360 72 44424
rect 88 44360 152 44424
rect 168 44360 232 44424
rect 248 44360 312 44424
rect 328 44360 392 44424
rect 408 44360 472 44424
rect 488 44360 552 44424
rect 568 44360 632 44424
rect 648 44360 712 44424
rect 728 44360 792 44424
rect 808 44360 872 44424
rect 888 44360 952 44424
rect 968 44360 1032 44424
rect 1048 44360 1112 44424
rect 1128 44360 1192 44424
rect 1208 44360 1272 44424
rect 1288 44360 1352 44424
rect 1368 44360 1432 44424
rect 1448 44360 1512 44424
rect 1528 44360 1592 44424
rect 1608 44360 1672 44424
rect 1688 44360 1752 44424
rect 1768 44360 1832 44424
rect 1848 44360 1912 44424
rect 1928 44360 1992 44424
rect 2008 44360 2072 44424
rect 2088 44360 2152 44424
rect 2168 44360 2232 44424
rect 2248 44360 2312 44424
rect 2328 44360 2392 44424
rect 2408 44360 2472 44424
rect 2488 44360 2552 44424
rect 2568 44360 2632 44424
rect 2648 44360 2712 44424
rect 2728 44360 2792 44424
rect 2808 44360 2872 44424
rect 2888 44360 2952 44424
rect 2968 44360 3032 44424
rect 3048 44360 3112 44424
rect 3128 44360 3192 44424
rect 3208 44360 3272 44424
rect 3288 44360 3352 44424
rect 3368 44360 3432 44424
rect 3448 44360 3512 44424
rect 3528 44360 3592 44424
rect 3608 44360 3672 44424
rect 3688 44360 3752 44424
rect 3768 44360 3832 44424
rect 3848 44360 3912 44424
rect 3928 44360 3992 44424
rect 19112 44360 19176 44424
rect 19192 44360 19256 44424
rect 19272 44360 19336 44424
rect 19352 44360 19416 44424
rect 29112 44360 29176 44424
rect 29192 44360 29256 44424
rect 29272 44360 29336 44424
rect 29352 44360 29416 44424
rect 41376 44360 41440 44424
rect 41456 44360 41520 44424
rect 41536 44360 41600 44424
rect 41616 44360 41680 44424
rect 41696 44360 41760 44424
rect 41776 44360 41840 44424
rect 41856 44360 41920 44424
rect 41936 44360 42000 44424
rect 42016 44360 42080 44424
rect 42096 44360 42160 44424
rect 42176 44360 42240 44424
rect 42256 44360 42320 44424
rect 42336 44360 42400 44424
rect 42416 44360 42480 44424
rect 42496 44360 42560 44424
rect 42576 44360 42640 44424
rect 42656 44360 42720 44424
rect 42736 44360 42800 44424
rect 42816 44360 42880 44424
rect 42896 44360 42960 44424
rect 42976 44360 43040 44424
rect 43056 44360 43120 44424
rect 43136 44360 43200 44424
rect 43216 44360 43280 44424
rect 43296 44360 43360 44424
rect 43376 44360 43440 44424
rect 43456 44360 43520 44424
rect 43536 44360 43600 44424
rect 43616 44360 43680 44424
rect 43696 44360 43760 44424
rect 43776 44360 43840 44424
rect 43856 44360 43920 44424
rect 43936 44360 44000 44424
rect 44016 44360 44080 44424
rect 44096 44360 44160 44424
rect 44176 44360 44240 44424
rect 44256 44360 44320 44424
rect 44336 44360 44400 44424
rect 44416 44360 44480 44424
rect 44496 44360 44560 44424
rect 44576 44360 44640 44424
rect 44656 44360 44720 44424
rect 44736 44360 44800 44424
rect 44816 44360 44880 44424
rect 44896 44360 44960 44424
rect 44976 44360 45040 44424
rect 45056 44360 45120 44424
rect 45136 44360 45200 44424
rect 45216 44360 45280 44424
rect 45296 44360 45360 44424
rect 8 44280 72 44344
rect 88 44280 152 44344
rect 168 44280 232 44344
rect 248 44280 312 44344
rect 328 44280 392 44344
rect 408 44280 472 44344
rect 488 44280 552 44344
rect 568 44280 632 44344
rect 648 44280 712 44344
rect 728 44280 792 44344
rect 808 44280 872 44344
rect 888 44280 952 44344
rect 968 44280 1032 44344
rect 1048 44280 1112 44344
rect 1128 44280 1192 44344
rect 1208 44280 1272 44344
rect 1288 44280 1352 44344
rect 1368 44280 1432 44344
rect 1448 44280 1512 44344
rect 1528 44280 1592 44344
rect 1608 44280 1672 44344
rect 1688 44280 1752 44344
rect 1768 44280 1832 44344
rect 1848 44280 1912 44344
rect 1928 44280 1992 44344
rect 2008 44280 2072 44344
rect 2088 44280 2152 44344
rect 2168 44280 2232 44344
rect 2248 44280 2312 44344
rect 2328 44280 2392 44344
rect 2408 44280 2472 44344
rect 2488 44280 2552 44344
rect 2568 44280 2632 44344
rect 2648 44280 2712 44344
rect 2728 44280 2792 44344
rect 2808 44280 2872 44344
rect 2888 44280 2952 44344
rect 2968 44280 3032 44344
rect 3048 44280 3112 44344
rect 3128 44280 3192 44344
rect 3208 44280 3272 44344
rect 3288 44280 3352 44344
rect 3368 44280 3432 44344
rect 3448 44280 3512 44344
rect 3528 44280 3592 44344
rect 3608 44280 3672 44344
rect 3688 44280 3752 44344
rect 3768 44280 3832 44344
rect 3848 44280 3912 44344
rect 3928 44280 3992 44344
rect 19112 44280 19176 44344
rect 19192 44280 19256 44344
rect 19272 44280 19336 44344
rect 19352 44280 19416 44344
rect 29112 44280 29176 44344
rect 29192 44280 29256 44344
rect 29272 44280 29336 44344
rect 29352 44280 29416 44344
rect 41376 44280 41440 44344
rect 41456 44280 41520 44344
rect 41536 44280 41600 44344
rect 41616 44280 41680 44344
rect 41696 44280 41760 44344
rect 41776 44280 41840 44344
rect 41856 44280 41920 44344
rect 41936 44280 42000 44344
rect 42016 44280 42080 44344
rect 42096 44280 42160 44344
rect 42176 44280 42240 44344
rect 42256 44280 42320 44344
rect 42336 44280 42400 44344
rect 42416 44280 42480 44344
rect 42496 44280 42560 44344
rect 42576 44280 42640 44344
rect 42656 44280 42720 44344
rect 42736 44280 42800 44344
rect 42816 44280 42880 44344
rect 42896 44280 42960 44344
rect 42976 44280 43040 44344
rect 43056 44280 43120 44344
rect 43136 44280 43200 44344
rect 43216 44280 43280 44344
rect 43296 44280 43360 44344
rect 43376 44280 43440 44344
rect 43456 44280 43520 44344
rect 43536 44280 43600 44344
rect 43616 44280 43680 44344
rect 43696 44280 43760 44344
rect 43776 44280 43840 44344
rect 43856 44280 43920 44344
rect 43936 44280 44000 44344
rect 44016 44280 44080 44344
rect 44096 44280 44160 44344
rect 44176 44280 44240 44344
rect 44256 44280 44320 44344
rect 44336 44280 44400 44344
rect 44416 44280 44480 44344
rect 44496 44280 44560 44344
rect 44576 44280 44640 44344
rect 44656 44280 44720 44344
rect 44736 44280 44800 44344
rect 44816 44280 44880 44344
rect 44896 44280 44960 44344
rect 44976 44280 45040 44344
rect 45056 44280 45120 44344
rect 45136 44280 45200 44344
rect 45216 44280 45280 44344
rect 45296 44280 45360 44344
rect 8 44200 72 44264
rect 88 44200 152 44264
rect 168 44200 232 44264
rect 248 44200 312 44264
rect 328 44200 392 44264
rect 408 44200 472 44264
rect 488 44200 552 44264
rect 568 44200 632 44264
rect 648 44200 712 44264
rect 728 44200 792 44264
rect 808 44200 872 44264
rect 888 44200 952 44264
rect 968 44200 1032 44264
rect 1048 44200 1112 44264
rect 1128 44200 1192 44264
rect 1208 44200 1272 44264
rect 1288 44200 1352 44264
rect 1368 44200 1432 44264
rect 1448 44200 1512 44264
rect 1528 44200 1592 44264
rect 1608 44200 1672 44264
rect 1688 44200 1752 44264
rect 1768 44200 1832 44264
rect 1848 44200 1912 44264
rect 1928 44200 1992 44264
rect 2008 44200 2072 44264
rect 2088 44200 2152 44264
rect 2168 44200 2232 44264
rect 2248 44200 2312 44264
rect 2328 44200 2392 44264
rect 2408 44200 2472 44264
rect 2488 44200 2552 44264
rect 2568 44200 2632 44264
rect 2648 44200 2712 44264
rect 2728 44200 2792 44264
rect 2808 44200 2872 44264
rect 2888 44200 2952 44264
rect 2968 44200 3032 44264
rect 3048 44200 3112 44264
rect 3128 44200 3192 44264
rect 3208 44200 3272 44264
rect 3288 44200 3352 44264
rect 3368 44200 3432 44264
rect 3448 44200 3512 44264
rect 3528 44200 3592 44264
rect 3608 44200 3672 44264
rect 3688 44200 3752 44264
rect 3768 44200 3832 44264
rect 3848 44200 3912 44264
rect 3928 44200 3992 44264
rect 19112 44200 19176 44264
rect 19192 44200 19256 44264
rect 19272 44200 19336 44264
rect 19352 44200 19416 44264
rect 29112 44200 29176 44264
rect 29192 44200 29256 44264
rect 29272 44200 29336 44264
rect 29352 44200 29416 44264
rect 41376 44200 41440 44264
rect 41456 44200 41520 44264
rect 41536 44200 41600 44264
rect 41616 44200 41680 44264
rect 41696 44200 41760 44264
rect 41776 44200 41840 44264
rect 41856 44200 41920 44264
rect 41936 44200 42000 44264
rect 42016 44200 42080 44264
rect 42096 44200 42160 44264
rect 42176 44200 42240 44264
rect 42256 44200 42320 44264
rect 42336 44200 42400 44264
rect 42416 44200 42480 44264
rect 42496 44200 42560 44264
rect 42576 44200 42640 44264
rect 42656 44200 42720 44264
rect 42736 44200 42800 44264
rect 42816 44200 42880 44264
rect 42896 44200 42960 44264
rect 42976 44200 43040 44264
rect 43056 44200 43120 44264
rect 43136 44200 43200 44264
rect 43216 44200 43280 44264
rect 43296 44200 43360 44264
rect 43376 44200 43440 44264
rect 43456 44200 43520 44264
rect 43536 44200 43600 44264
rect 43616 44200 43680 44264
rect 43696 44200 43760 44264
rect 43776 44200 43840 44264
rect 43856 44200 43920 44264
rect 43936 44200 44000 44264
rect 44016 44200 44080 44264
rect 44096 44200 44160 44264
rect 44176 44200 44240 44264
rect 44256 44200 44320 44264
rect 44336 44200 44400 44264
rect 44416 44200 44480 44264
rect 44496 44200 44560 44264
rect 44576 44200 44640 44264
rect 44656 44200 44720 44264
rect 44736 44200 44800 44264
rect 44816 44200 44880 44264
rect 44896 44200 44960 44264
rect 44976 44200 45040 44264
rect 45056 44200 45120 44264
rect 45136 44200 45200 44264
rect 45216 44200 45280 44264
rect 45296 44200 45360 44264
rect 8 44120 72 44184
rect 88 44120 152 44184
rect 168 44120 232 44184
rect 248 44120 312 44184
rect 328 44120 392 44184
rect 408 44120 472 44184
rect 488 44120 552 44184
rect 568 44120 632 44184
rect 648 44120 712 44184
rect 728 44120 792 44184
rect 808 44120 872 44184
rect 888 44120 952 44184
rect 968 44120 1032 44184
rect 1048 44120 1112 44184
rect 1128 44120 1192 44184
rect 1208 44120 1272 44184
rect 1288 44120 1352 44184
rect 1368 44120 1432 44184
rect 1448 44120 1512 44184
rect 1528 44120 1592 44184
rect 1608 44120 1672 44184
rect 1688 44120 1752 44184
rect 1768 44120 1832 44184
rect 1848 44120 1912 44184
rect 1928 44120 1992 44184
rect 2008 44120 2072 44184
rect 2088 44120 2152 44184
rect 2168 44120 2232 44184
rect 2248 44120 2312 44184
rect 2328 44120 2392 44184
rect 2408 44120 2472 44184
rect 2488 44120 2552 44184
rect 2568 44120 2632 44184
rect 2648 44120 2712 44184
rect 2728 44120 2792 44184
rect 2808 44120 2872 44184
rect 2888 44120 2952 44184
rect 2968 44120 3032 44184
rect 3048 44120 3112 44184
rect 3128 44120 3192 44184
rect 3208 44120 3272 44184
rect 3288 44120 3352 44184
rect 3368 44120 3432 44184
rect 3448 44120 3512 44184
rect 3528 44120 3592 44184
rect 3608 44120 3672 44184
rect 3688 44120 3752 44184
rect 3768 44120 3832 44184
rect 3848 44120 3912 44184
rect 3928 44120 3992 44184
rect 19112 44120 19176 44184
rect 19192 44120 19256 44184
rect 19272 44120 19336 44184
rect 19352 44120 19416 44184
rect 29112 44120 29176 44184
rect 29192 44120 29256 44184
rect 29272 44120 29336 44184
rect 29352 44120 29416 44184
rect 41376 44120 41440 44184
rect 41456 44120 41520 44184
rect 41536 44120 41600 44184
rect 41616 44120 41680 44184
rect 41696 44120 41760 44184
rect 41776 44120 41840 44184
rect 41856 44120 41920 44184
rect 41936 44120 42000 44184
rect 42016 44120 42080 44184
rect 42096 44120 42160 44184
rect 42176 44120 42240 44184
rect 42256 44120 42320 44184
rect 42336 44120 42400 44184
rect 42416 44120 42480 44184
rect 42496 44120 42560 44184
rect 42576 44120 42640 44184
rect 42656 44120 42720 44184
rect 42736 44120 42800 44184
rect 42816 44120 42880 44184
rect 42896 44120 42960 44184
rect 42976 44120 43040 44184
rect 43056 44120 43120 44184
rect 43136 44120 43200 44184
rect 43216 44120 43280 44184
rect 43296 44120 43360 44184
rect 43376 44120 43440 44184
rect 43456 44120 43520 44184
rect 43536 44120 43600 44184
rect 43616 44120 43680 44184
rect 43696 44120 43760 44184
rect 43776 44120 43840 44184
rect 43856 44120 43920 44184
rect 43936 44120 44000 44184
rect 44016 44120 44080 44184
rect 44096 44120 44160 44184
rect 44176 44120 44240 44184
rect 44256 44120 44320 44184
rect 44336 44120 44400 44184
rect 44416 44120 44480 44184
rect 44496 44120 44560 44184
rect 44576 44120 44640 44184
rect 44656 44120 44720 44184
rect 44736 44120 44800 44184
rect 44816 44120 44880 44184
rect 44896 44120 44960 44184
rect 44976 44120 45040 44184
rect 45056 44120 45120 44184
rect 45136 44120 45200 44184
rect 45216 44120 45280 44184
rect 45296 44120 45360 44184
rect 8 44040 72 44104
rect 88 44040 152 44104
rect 168 44040 232 44104
rect 248 44040 312 44104
rect 328 44040 392 44104
rect 408 44040 472 44104
rect 488 44040 552 44104
rect 568 44040 632 44104
rect 648 44040 712 44104
rect 728 44040 792 44104
rect 808 44040 872 44104
rect 888 44040 952 44104
rect 968 44040 1032 44104
rect 1048 44040 1112 44104
rect 1128 44040 1192 44104
rect 1208 44040 1272 44104
rect 1288 44040 1352 44104
rect 1368 44040 1432 44104
rect 1448 44040 1512 44104
rect 1528 44040 1592 44104
rect 1608 44040 1672 44104
rect 1688 44040 1752 44104
rect 1768 44040 1832 44104
rect 1848 44040 1912 44104
rect 1928 44040 1992 44104
rect 2008 44040 2072 44104
rect 2088 44040 2152 44104
rect 2168 44040 2232 44104
rect 2248 44040 2312 44104
rect 2328 44040 2392 44104
rect 2408 44040 2472 44104
rect 2488 44040 2552 44104
rect 2568 44040 2632 44104
rect 2648 44040 2712 44104
rect 2728 44040 2792 44104
rect 2808 44040 2872 44104
rect 2888 44040 2952 44104
rect 2968 44040 3032 44104
rect 3048 44040 3112 44104
rect 3128 44040 3192 44104
rect 3208 44040 3272 44104
rect 3288 44040 3352 44104
rect 3368 44040 3432 44104
rect 3448 44040 3512 44104
rect 3528 44040 3592 44104
rect 3608 44040 3672 44104
rect 3688 44040 3752 44104
rect 3768 44040 3832 44104
rect 3848 44040 3912 44104
rect 3928 44040 3992 44104
rect 19112 44040 19176 44104
rect 19192 44040 19256 44104
rect 19272 44040 19336 44104
rect 19352 44040 19416 44104
rect 29112 44040 29176 44104
rect 29192 44040 29256 44104
rect 29272 44040 29336 44104
rect 29352 44040 29416 44104
rect 41376 44040 41440 44104
rect 41456 44040 41520 44104
rect 41536 44040 41600 44104
rect 41616 44040 41680 44104
rect 41696 44040 41760 44104
rect 41776 44040 41840 44104
rect 41856 44040 41920 44104
rect 41936 44040 42000 44104
rect 42016 44040 42080 44104
rect 42096 44040 42160 44104
rect 42176 44040 42240 44104
rect 42256 44040 42320 44104
rect 42336 44040 42400 44104
rect 42416 44040 42480 44104
rect 42496 44040 42560 44104
rect 42576 44040 42640 44104
rect 42656 44040 42720 44104
rect 42736 44040 42800 44104
rect 42816 44040 42880 44104
rect 42896 44040 42960 44104
rect 42976 44040 43040 44104
rect 43056 44040 43120 44104
rect 43136 44040 43200 44104
rect 43216 44040 43280 44104
rect 43296 44040 43360 44104
rect 43376 44040 43440 44104
rect 43456 44040 43520 44104
rect 43536 44040 43600 44104
rect 43616 44040 43680 44104
rect 43696 44040 43760 44104
rect 43776 44040 43840 44104
rect 43856 44040 43920 44104
rect 43936 44040 44000 44104
rect 44016 44040 44080 44104
rect 44096 44040 44160 44104
rect 44176 44040 44240 44104
rect 44256 44040 44320 44104
rect 44336 44040 44400 44104
rect 44416 44040 44480 44104
rect 44496 44040 44560 44104
rect 44576 44040 44640 44104
rect 44656 44040 44720 44104
rect 44736 44040 44800 44104
rect 44816 44040 44880 44104
rect 44896 44040 44960 44104
rect 44976 44040 45040 44104
rect 45056 44040 45120 44104
rect 45136 44040 45200 44104
rect 45216 44040 45280 44104
rect 45296 44040 45360 44104
rect 8 43960 72 44024
rect 88 43960 152 44024
rect 168 43960 232 44024
rect 248 43960 312 44024
rect 328 43960 392 44024
rect 408 43960 472 44024
rect 488 43960 552 44024
rect 568 43960 632 44024
rect 648 43960 712 44024
rect 728 43960 792 44024
rect 808 43960 872 44024
rect 888 43960 952 44024
rect 968 43960 1032 44024
rect 1048 43960 1112 44024
rect 1128 43960 1192 44024
rect 1208 43960 1272 44024
rect 1288 43960 1352 44024
rect 1368 43960 1432 44024
rect 1448 43960 1512 44024
rect 1528 43960 1592 44024
rect 1608 43960 1672 44024
rect 1688 43960 1752 44024
rect 1768 43960 1832 44024
rect 1848 43960 1912 44024
rect 1928 43960 1992 44024
rect 2008 43960 2072 44024
rect 2088 43960 2152 44024
rect 2168 43960 2232 44024
rect 2248 43960 2312 44024
rect 2328 43960 2392 44024
rect 2408 43960 2472 44024
rect 2488 43960 2552 44024
rect 2568 43960 2632 44024
rect 2648 43960 2712 44024
rect 2728 43960 2792 44024
rect 2808 43960 2872 44024
rect 2888 43960 2952 44024
rect 2968 43960 3032 44024
rect 3048 43960 3112 44024
rect 3128 43960 3192 44024
rect 3208 43960 3272 44024
rect 3288 43960 3352 44024
rect 3368 43960 3432 44024
rect 3448 43960 3512 44024
rect 3528 43960 3592 44024
rect 3608 43960 3672 44024
rect 3688 43960 3752 44024
rect 3768 43960 3832 44024
rect 3848 43960 3912 44024
rect 3928 43960 3992 44024
rect 19112 43960 19176 44024
rect 19192 43960 19256 44024
rect 19272 43960 19336 44024
rect 19352 43960 19416 44024
rect 29112 43960 29176 44024
rect 29192 43960 29256 44024
rect 29272 43960 29336 44024
rect 29352 43960 29416 44024
rect 41376 43960 41440 44024
rect 41456 43960 41520 44024
rect 41536 43960 41600 44024
rect 41616 43960 41680 44024
rect 41696 43960 41760 44024
rect 41776 43960 41840 44024
rect 41856 43960 41920 44024
rect 41936 43960 42000 44024
rect 42016 43960 42080 44024
rect 42096 43960 42160 44024
rect 42176 43960 42240 44024
rect 42256 43960 42320 44024
rect 42336 43960 42400 44024
rect 42416 43960 42480 44024
rect 42496 43960 42560 44024
rect 42576 43960 42640 44024
rect 42656 43960 42720 44024
rect 42736 43960 42800 44024
rect 42816 43960 42880 44024
rect 42896 43960 42960 44024
rect 42976 43960 43040 44024
rect 43056 43960 43120 44024
rect 43136 43960 43200 44024
rect 43216 43960 43280 44024
rect 43296 43960 43360 44024
rect 43376 43960 43440 44024
rect 43456 43960 43520 44024
rect 43536 43960 43600 44024
rect 43616 43960 43680 44024
rect 43696 43960 43760 44024
rect 43776 43960 43840 44024
rect 43856 43960 43920 44024
rect 43936 43960 44000 44024
rect 44016 43960 44080 44024
rect 44096 43960 44160 44024
rect 44176 43960 44240 44024
rect 44256 43960 44320 44024
rect 44336 43960 44400 44024
rect 44416 43960 44480 44024
rect 44496 43960 44560 44024
rect 44576 43960 44640 44024
rect 44656 43960 44720 44024
rect 44736 43960 44800 44024
rect 44816 43960 44880 44024
rect 44896 43960 44960 44024
rect 44976 43960 45040 44024
rect 45056 43960 45120 44024
rect 45136 43960 45200 44024
rect 45216 43960 45280 44024
rect 45296 43960 45360 44024
rect 8 43880 72 43944
rect 88 43880 152 43944
rect 168 43880 232 43944
rect 248 43880 312 43944
rect 328 43880 392 43944
rect 408 43880 472 43944
rect 488 43880 552 43944
rect 568 43880 632 43944
rect 648 43880 712 43944
rect 728 43880 792 43944
rect 808 43880 872 43944
rect 888 43880 952 43944
rect 968 43880 1032 43944
rect 1048 43880 1112 43944
rect 1128 43880 1192 43944
rect 1208 43880 1272 43944
rect 1288 43880 1352 43944
rect 1368 43880 1432 43944
rect 1448 43880 1512 43944
rect 1528 43880 1592 43944
rect 1608 43880 1672 43944
rect 1688 43880 1752 43944
rect 1768 43880 1832 43944
rect 1848 43880 1912 43944
rect 1928 43880 1992 43944
rect 2008 43880 2072 43944
rect 2088 43880 2152 43944
rect 2168 43880 2232 43944
rect 2248 43880 2312 43944
rect 2328 43880 2392 43944
rect 2408 43880 2472 43944
rect 2488 43880 2552 43944
rect 2568 43880 2632 43944
rect 2648 43880 2712 43944
rect 2728 43880 2792 43944
rect 2808 43880 2872 43944
rect 2888 43880 2952 43944
rect 2968 43880 3032 43944
rect 3048 43880 3112 43944
rect 3128 43880 3192 43944
rect 3208 43880 3272 43944
rect 3288 43880 3352 43944
rect 3368 43880 3432 43944
rect 3448 43880 3512 43944
rect 3528 43880 3592 43944
rect 3608 43880 3672 43944
rect 3688 43880 3752 43944
rect 3768 43880 3832 43944
rect 3848 43880 3912 43944
rect 3928 43880 3992 43944
rect 19112 43880 19176 43944
rect 19192 43880 19256 43944
rect 19272 43880 19336 43944
rect 19352 43880 19416 43944
rect 29112 43880 29176 43944
rect 29192 43880 29256 43944
rect 29272 43880 29336 43944
rect 29352 43880 29416 43944
rect 41376 43880 41440 43944
rect 41456 43880 41520 43944
rect 41536 43880 41600 43944
rect 41616 43880 41680 43944
rect 41696 43880 41760 43944
rect 41776 43880 41840 43944
rect 41856 43880 41920 43944
rect 41936 43880 42000 43944
rect 42016 43880 42080 43944
rect 42096 43880 42160 43944
rect 42176 43880 42240 43944
rect 42256 43880 42320 43944
rect 42336 43880 42400 43944
rect 42416 43880 42480 43944
rect 42496 43880 42560 43944
rect 42576 43880 42640 43944
rect 42656 43880 42720 43944
rect 42736 43880 42800 43944
rect 42816 43880 42880 43944
rect 42896 43880 42960 43944
rect 42976 43880 43040 43944
rect 43056 43880 43120 43944
rect 43136 43880 43200 43944
rect 43216 43880 43280 43944
rect 43296 43880 43360 43944
rect 43376 43880 43440 43944
rect 43456 43880 43520 43944
rect 43536 43880 43600 43944
rect 43616 43880 43680 43944
rect 43696 43880 43760 43944
rect 43776 43880 43840 43944
rect 43856 43880 43920 43944
rect 43936 43880 44000 43944
rect 44016 43880 44080 43944
rect 44096 43880 44160 43944
rect 44176 43880 44240 43944
rect 44256 43880 44320 43944
rect 44336 43880 44400 43944
rect 44416 43880 44480 43944
rect 44496 43880 44560 43944
rect 44576 43880 44640 43944
rect 44656 43880 44720 43944
rect 44736 43880 44800 43944
rect 44816 43880 44880 43944
rect 44896 43880 44960 43944
rect 44976 43880 45040 43944
rect 45056 43880 45120 43944
rect 45136 43880 45200 43944
rect 45216 43880 45280 43944
rect 45296 43880 45360 43944
rect 8 43800 72 43864
rect 88 43800 152 43864
rect 168 43800 232 43864
rect 248 43800 312 43864
rect 328 43800 392 43864
rect 408 43800 472 43864
rect 488 43800 552 43864
rect 568 43800 632 43864
rect 648 43800 712 43864
rect 728 43800 792 43864
rect 808 43800 872 43864
rect 888 43800 952 43864
rect 968 43800 1032 43864
rect 1048 43800 1112 43864
rect 1128 43800 1192 43864
rect 1208 43800 1272 43864
rect 1288 43800 1352 43864
rect 1368 43800 1432 43864
rect 1448 43800 1512 43864
rect 1528 43800 1592 43864
rect 1608 43800 1672 43864
rect 1688 43800 1752 43864
rect 1768 43800 1832 43864
rect 1848 43800 1912 43864
rect 1928 43800 1992 43864
rect 2008 43800 2072 43864
rect 2088 43800 2152 43864
rect 2168 43800 2232 43864
rect 2248 43800 2312 43864
rect 2328 43800 2392 43864
rect 2408 43800 2472 43864
rect 2488 43800 2552 43864
rect 2568 43800 2632 43864
rect 2648 43800 2712 43864
rect 2728 43800 2792 43864
rect 2808 43800 2872 43864
rect 2888 43800 2952 43864
rect 2968 43800 3032 43864
rect 3048 43800 3112 43864
rect 3128 43800 3192 43864
rect 3208 43800 3272 43864
rect 3288 43800 3352 43864
rect 3368 43800 3432 43864
rect 3448 43800 3512 43864
rect 3528 43800 3592 43864
rect 3608 43800 3672 43864
rect 3688 43800 3752 43864
rect 3768 43800 3832 43864
rect 3848 43800 3912 43864
rect 3928 43800 3992 43864
rect 19112 43800 19176 43864
rect 19192 43800 19256 43864
rect 19272 43800 19336 43864
rect 19352 43800 19416 43864
rect 29112 43800 29176 43864
rect 29192 43800 29256 43864
rect 29272 43800 29336 43864
rect 29352 43800 29416 43864
rect 41376 43800 41440 43864
rect 41456 43800 41520 43864
rect 41536 43800 41600 43864
rect 41616 43800 41680 43864
rect 41696 43800 41760 43864
rect 41776 43800 41840 43864
rect 41856 43800 41920 43864
rect 41936 43800 42000 43864
rect 42016 43800 42080 43864
rect 42096 43800 42160 43864
rect 42176 43800 42240 43864
rect 42256 43800 42320 43864
rect 42336 43800 42400 43864
rect 42416 43800 42480 43864
rect 42496 43800 42560 43864
rect 42576 43800 42640 43864
rect 42656 43800 42720 43864
rect 42736 43800 42800 43864
rect 42816 43800 42880 43864
rect 42896 43800 42960 43864
rect 42976 43800 43040 43864
rect 43056 43800 43120 43864
rect 43136 43800 43200 43864
rect 43216 43800 43280 43864
rect 43296 43800 43360 43864
rect 43376 43800 43440 43864
rect 43456 43800 43520 43864
rect 43536 43800 43600 43864
rect 43616 43800 43680 43864
rect 43696 43800 43760 43864
rect 43776 43800 43840 43864
rect 43856 43800 43920 43864
rect 43936 43800 44000 43864
rect 44016 43800 44080 43864
rect 44096 43800 44160 43864
rect 44176 43800 44240 43864
rect 44256 43800 44320 43864
rect 44336 43800 44400 43864
rect 44416 43800 44480 43864
rect 44496 43800 44560 43864
rect 44576 43800 44640 43864
rect 44656 43800 44720 43864
rect 44736 43800 44800 43864
rect 44816 43800 44880 43864
rect 44896 43800 44960 43864
rect 44976 43800 45040 43864
rect 45056 43800 45120 43864
rect 45136 43800 45200 43864
rect 45216 43800 45280 43864
rect 45296 43800 45360 43864
rect 8 43720 72 43784
rect 88 43720 152 43784
rect 168 43720 232 43784
rect 248 43720 312 43784
rect 328 43720 392 43784
rect 408 43720 472 43784
rect 488 43720 552 43784
rect 568 43720 632 43784
rect 648 43720 712 43784
rect 728 43720 792 43784
rect 808 43720 872 43784
rect 888 43720 952 43784
rect 968 43720 1032 43784
rect 1048 43720 1112 43784
rect 1128 43720 1192 43784
rect 1208 43720 1272 43784
rect 1288 43720 1352 43784
rect 1368 43720 1432 43784
rect 1448 43720 1512 43784
rect 1528 43720 1592 43784
rect 1608 43720 1672 43784
rect 1688 43720 1752 43784
rect 1768 43720 1832 43784
rect 1848 43720 1912 43784
rect 1928 43720 1992 43784
rect 2008 43720 2072 43784
rect 2088 43720 2152 43784
rect 2168 43720 2232 43784
rect 2248 43720 2312 43784
rect 2328 43720 2392 43784
rect 2408 43720 2472 43784
rect 2488 43720 2552 43784
rect 2568 43720 2632 43784
rect 2648 43720 2712 43784
rect 2728 43720 2792 43784
rect 2808 43720 2872 43784
rect 2888 43720 2952 43784
rect 2968 43720 3032 43784
rect 3048 43720 3112 43784
rect 3128 43720 3192 43784
rect 3208 43720 3272 43784
rect 3288 43720 3352 43784
rect 3368 43720 3432 43784
rect 3448 43720 3512 43784
rect 3528 43720 3592 43784
rect 3608 43720 3672 43784
rect 3688 43720 3752 43784
rect 3768 43720 3832 43784
rect 3848 43720 3912 43784
rect 3928 43720 3992 43784
rect 19112 43720 19176 43784
rect 19192 43720 19256 43784
rect 19272 43720 19336 43784
rect 19352 43720 19416 43784
rect 29112 43720 29176 43784
rect 29192 43720 29256 43784
rect 29272 43720 29336 43784
rect 29352 43720 29416 43784
rect 41376 43720 41440 43784
rect 41456 43720 41520 43784
rect 41536 43720 41600 43784
rect 41616 43720 41680 43784
rect 41696 43720 41760 43784
rect 41776 43720 41840 43784
rect 41856 43720 41920 43784
rect 41936 43720 42000 43784
rect 42016 43720 42080 43784
rect 42096 43720 42160 43784
rect 42176 43720 42240 43784
rect 42256 43720 42320 43784
rect 42336 43720 42400 43784
rect 42416 43720 42480 43784
rect 42496 43720 42560 43784
rect 42576 43720 42640 43784
rect 42656 43720 42720 43784
rect 42736 43720 42800 43784
rect 42816 43720 42880 43784
rect 42896 43720 42960 43784
rect 42976 43720 43040 43784
rect 43056 43720 43120 43784
rect 43136 43720 43200 43784
rect 43216 43720 43280 43784
rect 43296 43720 43360 43784
rect 43376 43720 43440 43784
rect 43456 43720 43520 43784
rect 43536 43720 43600 43784
rect 43616 43720 43680 43784
rect 43696 43720 43760 43784
rect 43776 43720 43840 43784
rect 43856 43720 43920 43784
rect 43936 43720 44000 43784
rect 44016 43720 44080 43784
rect 44096 43720 44160 43784
rect 44176 43720 44240 43784
rect 44256 43720 44320 43784
rect 44336 43720 44400 43784
rect 44416 43720 44480 43784
rect 44496 43720 44560 43784
rect 44576 43720 44640 43784
rect 44656 43720 44720 43784
rect 44736 43720 44800 43784
rect 44816 43720 44880 43784
rect 44896 43720 44960 43784
rect 44976 43720 45040 43784
rect 45056 43720 45120 43784
rect 45136 43720 45200 43784
rect 45216 43720 45280 43784
rect 45296 43720 45360 43784
rect 8 43640 72 43704
rect 88 43640 152 43704
rect 168 43640 232 43704
rect 248 43640 312 43704
rect 328 43640 392 43704
rect 408 43640 472 43704
rect 488 43640 552 43704
rect 568 43640 632 43704
rect 648 43640 712 43704
rect 728 43640 792 43704
rect 808 43640 872 43704
rect 888 43640 952 43704
rect 968 43640 1032 43704
rect 1048 43640 1112 43704
rect 1128 43640 1192 43704
rect 1208 43640 1272 43704
rect 1288 43640 1352 43704
rect 1368 43640 1432 43704
rect 1448 43640 1512 43704
rect 1528 43640 1592 43704
rect 1608 43640 1672 43704
rect 1688 43640 1752 43704
rect 1768 43640 1832 43704
rect 1848 43640 1912 43704
rect 1928 43640 1992 43704
rect 2008 43640 2072 43704
rect 2088 43640 2152 43704
rect 2168 43640 2232 43704
rect 2248 43640 2312 43704
rect 2328 43640 2392 43704
rect 2408 43640 2472 43704
rect 2488 43640 2552 43704
rect 2568 43640 2632 43704
rect 2648 43640 2712 43704
rect 2728 43640 2792 43704
rect 2808 43640 2872 43704
rect 2888 43640 2952 43704
rect 2968 43640 3032 43704
rect 3048 43640 3112 43704
rect 3128 43640 3192 43704
rect 3208 43640 3272 43704
rect 3288 43640 3352 43704
rect 3368 43640 3432 43704
rect 3448 43640 3512 43704
rect 3528 43640 3592 43704
rect 3608 43640 3672 43704
rect 3688 43640 3752 43704
rect 3768 43640 3832 43704
rect 3848 43640 3912 43704
rect 3928 43640 3992 43704
rect 19112 43640 19176 43704
rect 19192 43640 19256 43704
rect 19272 43640 19336 43704
rect 19352 43640 19416 43704
rect 29112 43640 29176 43704
rect 29192 43640 29256 43704
rect 29272 43640 29336 43704
rect 29352 43640 29416 43704
rect 41376 43640 41440 43704
rect 41456 43640 41520 43704
rect 41536 43640 41600 43704
rect 41616 43640 41680 43704
rect 41696 43640 41760 43704
rect 41776 43640 41840 43704
rect 41856 43640 41920 43704
rect 41936 43640 42000 43704
rect 42016 43640 42080 43704
rect 42096 43640 42160 43704
rect 42176 43640 42240 43704
rect 42256 43640 42320 43704
rect 42336 43640 42400 43704
rect 42416 43640 42480 43704
rect 42496 43640 42560 43704
rect 42576 43640 42640 43704
rect 42656 43640 42720 43704
rect 42736 43640 42800 43704
rect 42816 43640 42880 43704
rect 42896 43640 42960 43704
rect 42976 43640 43040 43704
rect 43056 43640 43120 43704
rect 43136 43640 43200 43704
rect 43216 43640 43280 43704
rect 43296 43640 43360 43704
rect 43376 43640 43440 43704
rect 43456 43640 43520 43704
rect 43536 43640 43600 43704
rect 43616 43640 43680 43704
rect 43696 43640 43760 43704
rect 43776 43640 43840 43704
rect 43856 43640 43920 43704
rect 43936 43640 44000 43704
rect 44016 43640 44080 43704
rect 44096 43640 44160 43704
rect 44176 43640 44240 43704
rect 44256 43640 44320 43704
rect 44336 43640 44400 43704
rect 44416 43640 44480 43704
rect 44496 43640 44560 43704
rect 44576 43640 44640 43704
rect 44656 43640 44720 43704
rect 44736 43640 44800 43704
rect 44816 43640 44880 43704
rect 44896 43640 44960 43704
rect 44976 43640 45040 43704
rect 45056 43640 45120 43704
rect 45136 43640 45200 43704
rect 45216 43640 45280 43704
rect 45296 43640 45360 43704
rect 8 43560 72 43624
rect 88 43560 152 43624
rect 168 43560 232 43624
rect 248 43560 312 43624
rect 328 43560 392 43624
rect 408 43560 472 43624
rect 488 43560 552 43624
rect 568 43560 632 43624
rect 648 43560 712 43624
rect 728 43560 792 43624
rect 808 43560 872 43624
rect 888 43560 952 43624
rect 968 43560 1032 43624
rect 1048 43560 1112 43624
rect 1128 43560 1192 43624
rect 1208 43560 1272 43624
rect 1288 43560 1352 43624
rect 1368 43560 1432 43624
rect 1448 43560 1512 43624
rect 1528 43560 1592 43624
rect 1608 43560 1672 43624
rect 1688 43560 1752 43624
rect 1768 43560 1832 43624
rect 1848 43560 1912 43624
rect 1928 43560 1992 43624
rect 2008 43560 2072 43624
rect 2088 43560 2152 43624
rect 2168 43560 2232 43624
rect 2248 43560 2312 43624
rect 2328 43560 2392 43624
rect 2408 43560 2472 43624
rect 2488 43560 2552 43624
rect 2568 43560 2632 43624
rect 2648 43560 2712 43624
rect 2728 43560 2792 43624
rect 2808 43560 2872 43624
rect 2888 43560 2952 43624
rect 2968 43560 3032 43624
rect 3048 43560 3112 43624
rect 3128 43560 3192 43624
rect 3208 43560 3272 43624
rect 3288 43560 3352 43624
rect 3368 43560 3432 43624
rect 3448 43560 3512 43624
rect 3528 43560 3592 43624
rect 3608 43560 3672 43624
rect 3688 43560 3752 43624
rect 3768 43560 3832 43624
rect 3848 43560 3912 43624
rect 3928 43560 3992 43624
rect 19112 43560 19176 43624
rect 19192 43560 19256 43624
rect 19272 43560 19336 43624
rect 19352 43560 19416 43624
rect 29112 43560 29176 43624
rect 29192 43560 29256 43624
rect 29272 43560 29336 43624
rect 29352 43560 29416 43624
rect 41376 43560 41440 43624
rect 41456 43560 41520 43624
rect 41536 43560 41600 43624
rect 41616 43560 41680 43624
rect 41696 43560 41760 43624
rect 41776 43560 41840 43624
rect 41856 43560 41920 43624
rect 41936 43560 42000 43624
rect 42016 43560 42080 43624
rect 42096 43560 42160 43624
rect 42176 43560 42240 43624
rect 42256 43560 42320 43624
rect 42336 43560 42400 43624
rect 42416 43560 42480 43624
rect 42496 43560 42560 43624
rect 42576 43560 42640 43624
rect 42656 43560 42720 43624
rect 42736 43560 42800 43624
rect 42816 43560 42880 43624
rect 42896 43560 42960 43624
rect 42976 43560 43040 43624
rect 43056 43560 43120 43624
rect 43136 43560 43200 43624
rect 43216 43560 43280 43624
rect 43296 43560 43360 43624
rect 43376 43560 43440 43624
rect 43456 43560 43520 43624
rect 43536 43560 43600 43624
rect 43616 43560 43680 43624
rect 43696 43560 43760 43624
rect 43776 43560 43840 43624
rect 43856 43560 43920 43624
rect 43936 43560 44000 43624
rect 44016 43560 44080 43624
rect 44096 43560 44160 43624
rect 44176 43560 44240 43624
rect 44256 43560 44320 43624
rect 44336 43560 44400 43624
rect 44416 43560 44480 43624
rect 44496 43560 44560 43624
rect 44576 43560 44640 43624
rect 44656 43560 44720 43624
rect 44736 43560 44800 43624
rect 44816 43560 44880 43624
rect 44896 43560 44960 43624
rect 44976 43560 45040 43624
rect 45056 43560 45120 43624
rect 45136 43560 45200 43624
rect 45216 43560 45280 43624
rect 45296 43560 45360 43624
rect 8 43480 72 43544
rect 88 43480 152 43544
rect 168 43480 232 43544
rect 248 43480 312 43544
rect 328 43480 392 43544
rect 408 43480 472 43544
rect 488 43480 552 43544
rect 568 43480 632 43544
rect 648 43480 712 43544
rect 728 43480 792 43544
rect 808 43480 872 43544
rect 888 43480 952 43544
rect 968 43480 1032 43544
rect 1048 43480 1112 43544
rect 1128 43480 1192 43544
rect 1208 43480 1272 43544
rect 1288 43480 1352 43544
rect 1368 43480 1432 43544
rect 1448 43480 1512 43544
rect 1528 43480 1592 43544
rect 1608 43480 1672 43544
rect 1688 43480 1752 43544
rect 1768 43480 1832 43544
rect 1848 43480 1912 43544
rect 1928 43480 1992 43544
rect 2008 43480 2072 43544
rect 2088 43480 2152 43544
rect 2168 43480 2232 43544
rect 2248 43480 2312 43544
rect 2328 43480 2392 43544
rect 2408 43480 2472 43544
rect 2488 43480 2552 43544
rect 2568 43480 2632 43544
rect 2648 43480 2712 43544
rect 2728 43480 2792 43544
rect 2808 43480 2872 43544
rect 2888 43480 2952 43544
rect 2968 43480 3032 43544
rect 3048 43480 3112 43544
rect 3128 43480 3192 43544
rect 3208 43480 3272 43544
rect 3288 43480 3352 43544
rect 3368 43480 3432 43544
rect 3448 43480 3512 43544
rect 3528 43480 3592 43544
rect 3608 43480 3672 43544
rect 3688 43480 3752 43544
rect 3768 43480 3832 43544
rect 3848 43480 3912 43544
rect 3928 43480 3992 43544
rect 19112 43480 19176 43544
rect 19192 43480 19256 43544
rect 19272 43480 19336 43544
rect 19352 43480 19416 43544
rect 29112 43480 29176 43544
rect 29192 43480 29256 43544
rect 29272 43480 29336 43544
rect 29352 43480 29416 43544
rect 41376 43480 41440 43544
rect 41456 43480 41520 43544
rect 41536 43480 41600 43544
rect 41616 43480 41680 43544
rect 41696 43480 41760 43544
rect 41776 43480 41840 43544
rect 41856 43480 41920 43544
rect 41936 43480 42000 43544
rect 42016 43480 42080 43544
rect 42096 43480 42160 43544
rect 42176 43480 42240 43544
rect 42256 43480 42320 43544
rect 42336 43480 42400 43544
rect 42416 43480 42480 43544
rect 42496 43480 42560 43544
rect 42576 43480 42640 43544
rect 42656 43480 42720 43544
rect 42736 43480 42800 43544
rect 42816 43480 42880 43544
rect 42896 43480 42960 43544
rect 42976 43480 43040 43544
rect 43056 43480 43120 43544
rect 43136 43480 43200 43544
rect 43216 43480 43280 43544
rect 43296 43480 43360 43544
rect 43376 43480 43440 43544
rect 43456 43480 43520 43544
rect 43536 43480 43600 43544
rect 43616 43480 43680 43544
rect 43696 43480 43760 43544
rect 43776 43480 43840 43544
rect 43856 43480 43920 43544
rect 43936 43480 44000 43544
rect 44016 43480 44080 43544
rect 44096 43480 44160 43544
rect 44176 43480 44240 43544
rect 44256 43480 44320 43544
rect 44336 43480 44400 43544
rect 44416 43480 44480 43544
rect 44496 43480 44560 43544
rect 44576 43480 44640 43544
rect 44656 43480 44720 43544
rect 44736 43480 44800 43544
rect 44816 43480 44880 43544
rect 44896 43480 44960 43544
rect 44976 43480 45040 43544
rect 45056 43480 45120 43544
rect 45136 43480 45200 43544
rect 45216 43480 45280 43544
rect 45296 43480 45360 43544
rect 8 43400 72 43464
rect 88 43400 152 43464
rect 168 43400 232 43464
rect 248 43400 312 43464
rect 328 43400 392 43464
rect 408 43400 472 43464
rect 488 43400 552 43464
rect 568 43400 632 43464
rect 648 43400 712 43464
rect 728 43400 792 43464
rect 808 43400 872 43464
rect 888 43400 952 43464
rect 968 43400 1032 43464
rect 1048 43400 1112 43464
rect 1128 43400 1192 43464
rect 1208 43400 1272 43464
rect 1288 43400 1352 43464
rect 1368 43400 1432 43464
rect 1448 43400 1512 43464
rect 1528 43400 1592 43464
rect 1608 43400 1672 43464
rect 1688 43400 1752 43464
rect 1768 43400 1832 43464
rect 1848 43400 1912 43464
rect 1928 43400 1992 43464
rect 2008 43400 2072 43464
rect 2088 43400 2152 43464
rect 2168 43400 2232 43464
rect 2248 43400 2312 43464
rect 2328 43400 2392 43464
rect 2408 43400 2472 43464
rect 2488 43400 2552 43464
rect 2568 43400 2632 43464
rect 2648 43400 2712 43464
rect 2728 43400 2792 43464
rect 2808 43400 2872 43464
rect 2888 43400 2952 43464
rect 2968 43400 3032 43464
rect 3048 43400 3112 43464
rect 3128 43400 3192 43464
rect 3208 43400 3272 43464
rect 3288 43400 3352 43464
rect 3368 43400 3432 43464
rect 3448 43400 3512 43464
rect 3528 43400 3592 43464
rect 3608 43400 3672 43464
rect 3688 43400 3752 43464
rect 3768 43400 3832 43464
rect 3848 43400 3912 43464
rect 3928 43400 3992 43464
rect 19112 43400 19176 43464
rect 19192 43400 19256 43464
rect 19272 43400 19336 43464
rect 19352 43400 19416 43464
rect 29112 43400 29176 43464
rect 29192 43400 29256 43464
rect 29272 43400 29336 43464
rect 29352 43400 29416 43464
rect 41376 43400 41440 43464
rect 41456 43400 41520 43464
rect 41536 43400 41600 43464
rect 41616 43400 41680 43464
rect 41696 43400 41760 43464
rect 41776 43400 41840 43464
rect 41856 43400 41920 43464
rect 41936 43400 42000 43464
rect 42016 43400 42080 43464
rect 42096 43400 42160 43464
rect 42176 43400 42240 43464
rect 42256 43400 42320 43464
rect 42336 43400 42400 43464
rect 42416 43400 42480 43464
rect 42496 43400 42560 43464
rect 42576 43400 42640 43464
rect 42656 43400 42720 43464
rect 42736 43400 42800 43464
rect 42816 43400 42880 43464
rect 42896 43400 42960 43464
rect 42976 43400 43040 43464
rect 43056 43400 43120 43464
rect 43136 43400 43200 43464
rect 43216 43400 43280 43464
rect 43296 43400 43360 43464
rect 43376 43400 43440 43464
rect 43456 43400 43520 43464
rect 43536 43400 43600 43464
rect 43616 43400 43680 43464
rect 43696 43400 43760 43464
rect 43776 43400 43840 43464
rect 43856 43400 43920 43464
rect 43936 43400 44000 43464
rect 44016 43400 44080 43464
rect 44096 43400 44160 43464
rect 44176 43400 44240 43464
rect 44256 43400 44320 43464
rect 44336 43400 44400 43464
rect 44416 43400 44480 43464
rect 44496 43400 44560 43464
rect 44576 43400 44640 43464
rect 44656 43400 44720 43464
rect 44736 43400 44800 43464
rect 44816 43400 44880 43464
rect 44896 43400 44960 43464
rect 44976 43400 45040 43464
rect 45056 43400 45120 43464
rect 45136 43400 45200 43464
rect 45216 43400 45280 43464
rect 45296 43400 45360 43464
rect 8 43320 72 43384
rect 88 43320 152 43384
rect 168 43320 232 43384
rect 248 43320 312 43384
rect 328 43320 392 43384
rect 408 43320 472 43384
rect 488 43320 552 43384
rect 568 43320 632 43384
rect 648 43320 712 43384
rect 728 43320 792 43384
rect 808 43320 872 43384
rect 888 43320 952 43384
rect 968 43320 1032 43384
rect 1048 43320 1112 43384
rect 1128 43320 1192 43384
rect 1208 43320 1272 43384
rect 1288 43320 1352 43384
rect 1368 43320 1432 43384
rect 1448 43320 1512 43384
rect 1528 43320 1592 43384
rect 1608 43320 1672 43384
rect 1688 43320 1752 43384
rect 1768 43320 1832 43384
rect 1848 43320 1912 43384
rect 1928 43320 1992 43384
rect 2008 43320 2072 43384
rect 2088 43320 2152 43384
rect 2168 43320 2232 43384
rect 2248 43320 2312 43384
rect 2328 43320 2392 43384
rect 2408 43320 2472 43384
rect 2488 43320 2552 43384
rect 2568 43320 2632 43384
rect 2648 43320 2712 43384
rect 2728 43320 2792 43384
rect 2808 43320 2872 43384
rect 2888 43320 2952 43384
rect 2968 43320 3032 43384
rect 3048 43320 3112 43384
rect 3128 43320 3192 43384
rect 3208 43320 3272 43384
rect 3288 43320 3352 43384
rect 3368 43320 3432 43384
rect 3448 43320 3512 43384
rect 3528 43320 3592 43384
rect 3608 43320 3672 43384
rect 3688 43320 3752 43384
rect 3768 43320 3832 43384
rect 3848 43320 3912 43384
rect 3928 43320 3992 43384
rect 19112 43320 19176 43384
rect 19192 43320 19256 43384
rect 19272 43320 19336 43384
rect 19352 43320 19416 43384
rect 29112 43320 29176 43384
rect 29192 43320 29256 43384
rect 29272 43320 29336 43384
rect 29352 43320 29416 43384
rect 41376 43320 41440 43384
rect 41456 43320 41520 43384
rect 41536 43320 41600 43384
rect 41616 43320 41680 43384
rect 41696 43320 41760 43384
rect 41776 43320 41840 43384
rect 41856 43320 41920 43384
rect 41936 43320 42000 43384
rect 42016 43320 42080 43384
rect 42096 43320 42160 43384
rect 42176 43320 42240 43384
rect 42256 43320 42320 43384
rect 42336 43320 42400 43384
rect 42416 43320 42480 43384
rect 42496 43320 42560 43384
rect 42576 43320 42640 43384
rect 42656 43320 42720 43384
rect 42736 43320 42800 43384
rect 42816 43320 42880 43384
rect 42896 43320 42960 43384
rect 42976 43320 43040 43384
rect 43056 43320 43120 43384
rect 43136 43320 43200 43384
rect 43216 43320 43280 43384
rect 43296 43320 43360 43384
rect 43376 43320 43440 43384
rect 43456 43320 43520 43384
rect 43536 43320 43600 43384
rect 43616 43320 43680 43384
rect 43696 43320 43760 43384
rect 43776 43320 43840 43384
rect 43856 43320 43920 43384
rect 43936 43320 44000 43384
rect 44016 43320 44080 43384
rect 44096 43320 44160 43384
rect 44176 43320 44240 43384
rect 44256 43320 44320 43384
rect 44336 43320 44400 43384
rect 44416 43320 44480 43384
rect 44496 43320 44560 43384
rect 44576 43320 44640 43384
rect 44656 43320 44720 43384
rect 44736 43320 44800 43384
rect 44816 43320 44880 43384
rect 44896 43320 44960 43384
rect 44976 43320 45040 43384
rect 45056 43320 45120 43384
rect 45136 43320 45200 43384
rect 45216 43320 45280 43384
rect 45296 43320 45360 43384
rect 8 43240 72 43304
rect 88 43240 152 43304
rect 168 43240 232 43304
rect 248 43240 312 43304
rect 328 43240 392 43304
rect 408 43240 472 43304
rect 488 43240 552 43304
rect 568 43240 632 43304
rect 648 43240 712 43304
rect 728 43240 792 43304
rect 808 43240 872 43304
rect 888 43240 952 43304
rect 968 43240 1032 43304
rect 1048 43240 1112 43304
rect 1128 43240 1192 43304
rect 1208 43240 1272 43304
rect 1288 43240 1352 43304
rect 1368 43240 1432 43304
rect 1448 43240 1512 43304
rect 1528 43240 1592 43304
rect 1608 43240 1672 43304
rect 1688 43240 1752 43304
rect 1768 43240 1832 43304
rect 1848 43240 1912 43304
rect 1928 43240 1992 43304
rect 2008 43240 2072 43304
rect 2088 43240 2152 43304
rect 2168 43240 2232 43304
rect 2248 43240 2312 43304
rect 2328 43240 2392 43304
rect 2408 43240 2472 43304
rect 2488 43240 2552 43304
rect 2568 43240 2632 43304
rect 2648 43240 2712 43304
rect 2728 43240 2792 43304
rect 2808 43240 2872 43304
rect 2888 43240 2952 43304
rect 2968 43240 3032 43304
rect 3048 43240 3112 43304
rect 3128 43240 3192 43304
rect 3208 43240 3272 43304
rect 3288 43240 3352 43304
rect 3368 43240 3432 43304
rect 3448 43240 3512 43304
rect 3528 43240 3592 43304
rect 3608 43240 3672 43304
rect 3688 43240 3752 43304
rect 3768 43240 3832 43304
rect 3848 43240 3912 43304
rect 3928 43240 3992 43304
rect 19112 43240 19176 43304
rect 19192 43240 19256 43304
rect 19272 43240 19336 43304
rect 19352 43240 19416 43304
rect 29112 43240 29176 43304
rect 29192 43240 29256 43304
rect 29272 43240 29336 43304
rect 29352 43240 29416 43304
rect 41376 43240 41440 43304
rect 41456 43240 41520 43304
rect 41536 43240 41600 43304
rect 41616 43240 41680 43304
rect 41696 43240 41760 43304
rect 41776 43240 41840 43304
rect 41856 43240 41920 43304
rect 41936 43240 42000 43304
rect 42016 43240 42080 43304
rect 42096 43240 42160 43304
rect 42176 43240 42240 43304
rect 42256 43240 42320 43304
rect 42336 43240 42400 43304
rect 42416 43240 42480 43304
rect 42496 43240 42560 43304
rect 42576 43240 42640 43304
rect 42656 43240 42720 43304
rect 42736 43240 42800 43304
rect 42816 43240 42880 43304
rect 42896 43240 42960 43304
rect 42976 43240 43040 43304
rect 43056 43240 43120 43304
rect 43136 43240 43200 43304
rect 43216 43240 43280 43304
rect 43296 43240 43360 43304
rect 43376 43240 43440 43304
rect 43456 43240 43520 43304
rect 43536 43240 43600 43304
rect 43616 43240 43680 43304
rect 43696 43240 43760 43304
rect 43776 43240 43840 43304
rect 43856 43240 43920 43304
rect 43936 43240 44000 43304
rect 44016 43240 44080 43304
rect 44096 43240 44160 43304
rect 44176 43240 44240 43304
rect 44256 43240 44320 43304
rect 44336 43240 44400 43304
rect 44416 43240 44480 43304
rect 44496 43240 44560 43304
rect 44576 43240 44640 43304
rect 44656 43240 44720 43304
rect 44736 43240 44800 43304
rect 44816 43240 44880 43304
rect 44896 43240 44960 43304
rect 44976 43240 45040 43304
rect 45056 43240 45120 43304
rect 45136 43240 45200 43304
rect 45216 43240 45280 43304
rect 45296 43240 45360 43304
rect 8 43160 72 43224
rect 88 43160 152 43224
rect 168 43160 232 43224
rect 248 43160 312 43224
rect 328 43160 392 43224
rect 408 43160 472 43224
rect 488 43160 552 43224
rect 568 43160 632 43224
rect 648 43160 712 43224
rect 728 43160 792 43224
rect 808 43160 872 43224
rect 888 43160 952 43224
rect 968 43160 1032 43224
rect 1048 43160 1112 43224
rect 1128 43160 1192 43224
rect 1208 43160 1272 43224
rect 1288 43160 1352 43224
rect 1368 43160 1432 43224
rect 1448 43160 1512 43224
rect 1528 43160 1592 43224
rect 1608 43160 1672 43224
rect 1688 43160 1752 43224
rect 1768 43160 1832 43224
rect 1848 43160 1912 43224
rect 1928 43160 1992 43224
rect 2008 43160 2072 43224
rect 2088 43160 2152 43224
rect 2168 43160 2232 43224
rect 2248 43160 2312 43224
rect 2328 43160 2392 43224
rect 2408 43160 2472 43224
rect 2488 43160 2552 43224
rect 2568 43160 2632 43224
rect 2648 43160 2712 43224
rect 2728 43160 2792 43224
rect 2808 43160 2872 43224
rect 2888 43160 2952 43224
rect 2968 43160 3032 43224
rect 3048 43160 3112 43224
rect 3128 43160 3192 43224
rect 3208 43160 3272 43224
rect 3288 43160 3352 43224
rect 3368 43160 3432 43224
rect 3448 43160 3512 43224
rect 3528 43160 3592 43224
rect 3608 43160 3672 43224
rect 3688 43160 3752 43224
rect 3768 43160 3832 43224
rect 3848 43160 3912 43224
rect 3928 43160 3992 43224
rect 19112 43160 19176 43224
rect 19192 43160 19256 43224
rect 19272 43160 19336 43224
rect 19352 43160 19416 43224
rect 29112 43160 29176 43224
rect 29192 43160 29256 43224
rect 29272 43160 29336 43224
rect 29352 43160 29416 43224
rect 41376 43160 41440 43224
rect 41456 43160 41520 43224
rect 41536 43160 41600 43224
rect 41616 43160 41680 43224
rect 41696 43160 41760 43224
rect 41776 43160 41840 43224
rect 41856 43160 41920 43224
rect 41936 43160 42000 43224
rect 42016 43160 42080 43224
rect 42096 43160 42160 43224
rect 42176 43160 42240 43224
rect 42256 43160 42320 43224
rect 42336 43160 42400 43224
rect 42416 43160 42480 43224
rect 42496 43160 42560 43224
rect 42576 43160 42640 43224
rect 42656 43160 42720 43224
rect 42736 43160 42800 43224
rect 42816 43160 42880 43224
rect 42896 43160 42960 43224
rect 42976 43160 43040 43224
rect 43056 43160 43120 43224
rect 43136 43160 43200 43224
rect 43216 43160 43280 43224
rect 43296 43160 43360 43224
rect 43376 43160 43440 43224
rect 43456 43160 43520 43224
rect 43536 43160 43600 43224
rect 43616 43160 43680 43224
rect 43696 43160 43760 43224
rect 43776 43160 43840 43224
rect 43856 43160 43920 43224
rect 43936 43160 44000 43224
rect 44016 43160 44080 43224
rect 44096 43160 44160 43224
rect 44176 43160 44240 43224
rect 44256 43160 44320 43224
rect 44336 43160 44400 43224
rect 44416 43160 44480 43224
rect 44496 43160 44560 43224
rect 44576 43160 44640 43224
rect 44656 43160 44720 43224
rect 44736 43160 44800 43224
rect 44816 43160 44880 43224
rect 44896 43160 44960 43224
rect 44976 43160 45040 43224
rect 45056 43160 45120 43224
rect 45136 43160 45200 43224
rect 45216 43160 45280 43224
rect 45296 43160 45360 43224
rect 8 43080 72 43144
rect 88 43080 152 43144
rect 168 43080 232 43144
rect 248 43080 312 43144
rect 328 43080 392 43144
rect 408 43080 472 43144
rect 488 43080 552 43144
rect 568 43080 632 43144
rect 648 43080 712 43144
rect 728 43080 792 43144
rect 808 43080 872 43144
rect 888 43080 952 43144
rect 968 43080 1032 43144
rect 1048 43080 1112 43144
rect 1128 43080 1192 43144
rect 1208 43080 1272 43144
rect 1288 43080 1352 43144
rect 1368 43080 1432 43144
rect 1448 43080 1512 43144
rect 1528 43080 1592 43144
rect 1608 43080 1672 43144
rect 1688 43080 1752 43144
rect 1768 43080 1832 43144
rect 1848 43080 1912 43144
rect 1928 43080 1992 43144
rect 2008 43080 2072 43144
rect 2088 43080 2152 43144
rect 2168 43080 2232 43144
rect 2248 43080 2312 43144
rect 2328 43080 2392 43144
rect 2408 43080 2472 43144
rect 2488 43080 2552 43144
rect 2568 43080 2632 43144
rect 2648 43080 2712 43144
rect 2728 43080 2792 43144
rect 2808 43080 2872 43144
rect 2888 43080 2952 43144
rect 2968 43080 3032 43144
rect 3048 43080 3112 43144
rect 3128 43080 3192 43144
rect 3208 43080 3272 43144
rect 3288 43080 3352 43144
rect 3368 43080 3432 43144
rect 3448 43080 3512 43144
rect 3528 43080 3592 43144
rect 3608 43080 3672 43144
rect 3688 43080 3752 43144
rect 3768 43080 3832 43144
rect 3848 43080 3912 43144
rect 3928 43080 3992 43144
rect 19112 43080 19176 43144
rect 19192 43080 19256 43144
rect 19272 43080 19336 43144
rect 19352 43080 19416 43144
rect 29112 43080 29176 43144
rect 29192 43080 29256 43144
rect 29272 43080 29336 43144
rect 29352 43080 29416 43144
rect 41376 43080 41440 43144
rect 41456 43080 41520 43144
rect 41536 43080 41600 43144
rect 41616 43080 41680 43144
rect 41696 43080 41760 43144
rect 41776 43080 41840 43144
rect 41856 43080 41920 43144
rect 41936 43080 42000 43144
rect 42016 43080 42080 43144
rect 42096 43080 42160 43144
rect 42176 43080 42240 43144
rect 42256 43080 42320 43144
rect 42336 43080 42400 43144
rect 42416 43080 42480 43144
rect 42496 43080 42560 43144
rect 42576 43080 42640 43144
rect 42656 43080 42720 43144
rect 42736 43080 42800 43144
rect 42816 43080 42880 43144
rect 42896 43080 42960 43144
rect 42976 43080 43040 43144
rect 43056 43080 43120 43144
rect 43136 43080 43200 43144
rect 43216 43080 43280 43144
rect 43296 43080 43360 43144
rect 43376 43080 43440 43144
rect 43456 43080 43520 43144
rect 43536 43080 43600 43144
rect 43616 43080 43680 43144
rect 43696 43080 43760 43144
rect 43776 43080 43840 43144
rect 43856 43080 43920 43144
rect 43936 43080 44000 43144
rect 44016 43080 44080 43144
rect 44096 43080 44160 43144
rect 44176 43080 44240 43144
rect 44256 43080 44320 43144
rect 44336 43080 44400 43144
rect 44416 43080 44480 43144
rect 44496 43080 44560 43144
rect 44576 43080 44640 43144
rect 44656 43080 44720 43144
rect 44736 43080 44800 43144
rect 44816 43080 44880 43144
rect 44896 43080 44960 43144
rect 44976 43080 45040 43144
rect 45056 43080 45120 43144
rect 45136 43080 45200 43144
rect 45216 43080 45280 43144
rect 45296 43080 45360 43144
rect 8 43000 72 43064
rect 88 43000 152 43064
rect 168 43000 232 43064
rect 248 43000 312 43064
rect 328 43000 392 43064
rect 408 43000 472 43064
rect 488 43000 552 43064
rect 568 43000 632 43064
rect 648 43000 712 43064
rect 728 43000 792 43064
rect 808 43000 872 43064
rect 888 43000 952 43064
rect 968 43000 1032 43064
rect 1048 43000 1112 43064
rect 1128 43000 1192 43064
rect 1208 43000 1272 43064
rect 1288 43000 1352 43064
rect 1368 43000 1432 43064
rect 1448 43000 1512 43064
rect 1528 43000 1592 43064
rect 1608 43000 1672 43064
rect 1688 43000 1752 43064
rect 1768 43000 1832 43064
rect 1848 43000 1912 43064
rect 1928 43000 1992 43064
rect 2008 43000 2072 43064
rect 2088 43000 2152 43064
rect 2168 43000 2232 43064
rect 2248 43000 2312 43064
rect 2328 43000 2392 43064
rect 2408 43000 2472 43064
rect 2488 43000 2552 43064
rect 2568 43000 2632 43064
rect 2648 43000 2712 43064
rect 2728 43000 2792 43064
rect 2808 43000 2872 43064
rect 2888 43000 2952 43064
rect 2968 43000 3032 43064
rect 3048 43000 3112 43064
rect 3128 43000 3192 43064
rect 3208 43000 3272 43064
rect 3288 43000 3352 43064
rect 3368 43000 3432 43064
rect 3448 43000 3512 43064
rect 3528 43000 3592 43064
rect 3608 43000 3672 43064
rect 3688 43000 3752 43064
rect 3768 43000 3832 43064
rect 3848 43000 3912 43064
rect 3928 43000 3992 43064
rect 19112 43000 19176 43064
rect 19192 43000 19256 43064
rect 19272 43000 19336 43064
rect 19352 43000 19416 43064
rect 29112 43000 29176 43064
rect 29192 43000 29256 43064
rect 29272 43000 29336 43064
rect 29352 43000 29416 43064
rect 41376 43000 41440 43064
rect 41456 43000 41520 43064
rect 41536 43000 41600 43064
rect 41616 43000 41680 43064
rect 41696 43000 41760 43064
rect 41776 43000 41840 43064
rect 41856 43000 41920 43064
rect 41936 43000 42000 43064
rect 42016 43000 42080 43064
rect 42096 43000 42160 43064
rect 42176 43000 42240 43064
rect 42256 43000 42320 43064
rect 42336 43000 42400 43064
rect 42416 43000 42480 43064
rect 42496 43000 42560 43064
rect 42576 43000 42640 43064
rect 42656 43000 42720 43064
rect 42736 43000 42800 43064
rect 42816 43000 42880 43064
rect 42896 43000 42960 43064
rect 42976 43000 43040 43064
rect 43056 43000 43120 43064
rect 43136 43000 43200 43064
rect 43216 43000 43280 43064
rect 43296 43000 43360 43064
rect 43376 43000 43440 43064
rect 43456 43000 43520 43064
rect 43536 43000 43600 43064
rect 43616 43000 43680 43064
rect 43696 43000 43760 43064
rect 43776 43000 43840 43064
rect 43856 43000 43920 43064
rect 43936 43000 44000 43064
rect 44016 43000 44080 43064
rect 44096 43000 44160 43064
rect 44176 43000 44240 43064
rect 44256 43000 44320 43064
rect 44336 43000 44400 43064
rect 44416 43000 44480 43064
rect 44496 43000 44560 43064
rect 44576 43000 44640 43064
rect 44656 43000 44720 43064
rect 44736 43000 44800 43064
rect 44816 43000 44880 43064
rect 44896 43000 44960 43064
rect 44976 43000 45040 43064
rect 45056 43000 45120 43064
rect 45136 43000 45200 43064
rect 45216 43000 45280 43064
rect 45296 43000 45360 43064
rect 8 42920 72 42984
rect 88 42920 152 42984
rect 168 42920 232 42984
rect 248 42920 312 42984
rect 328 42920 392 42984
rect 408 42920 472 42984
rect 488 42920 552 42984
rect 568 42920 632 42984
rect 648 42920 712 42984
rect 728 42920 792 42984
rect 808 42920 872 42984
rect 888 42920 952 42984
rect 968 42920 1032 42984
rect 1048 42920 1112 42984
rect 1128 42920 1192 42984
rect 1208 42920 1272 42984
rect 1288 42920 1352 42984
rect 1368 42920 1432 42984
rect 1448 42920 1512 42984
rect 1528 42920 1592 42984
rect 1608 42920 1672 42984
rect 1688 42920 1752 42984
rect 1768 42920 1832 42984
rect 1848 42920 1912 42984
rect 1928 42920 1992 42984
rect 2008 42920 2072 42984
rect 2088 42920 2152 42984
rect 2168 42920 2232 42984
rect 2248 42920 2312 42984
rect 2328 42920 2392 42984
rect 2408 42920 2472 42984
rect 2488 42920 2552 42984
rect 2568 42920 2632 42984
rect 2648 42920 2712 42984
rect 2728 42920 2792 42984
rect 2808 42920 2872 42984
rect 2888 42920 2952 42984
rect 2968 42920 3032 42984
rect 3048 42920 3112 42984
rect 3128 42920 3192 42984
rect 3208 42920 3272 42984
rect 3288 42920 3352 42984
rect 3368 42920 3432 42984
rect 3448 42920 3512 42984
rect 3528 42920 3592 42984
rect 3608 42920 3672 42984
rect 3688 42920 3752 42984
rect 3768 42920 3832 42984
rect 3848 42920 3912 42984
rect 3928 42920 3992 42984
rect 19112 42920 19176 42984
rect 19192 42920 19256 42984
rect 19272 42920 19336 42984
rect 19352 42920 19416 42984
rect 29112 42920 29176 42984
rect 29192 42920 29256 42984
rect 29272 42920 29336 42984
rect 29352 42920 29416 42984
rect 41376 42920 41440 42984
rect 41456 42920 41520 42984
rect 41536 42920 41600 42984
rect 41616 42920 41680 42984
rect 41696 42920 41760 42984
rect 41776 42920 41840 42984
rect 41856 42920 41920 42984
rect 41936 42920 42000 42984
rect 42016 42920 42080 42984
rect 42096 42920 42160 42984
rect 42176 42920 42240 42984
rect 42256 42920 42320 42984
rect 42336 42920 42400 42984
rect 42416 42920 42480 42984
rect 42496 42920 42560 42984
rect 42576 42920 42640 42984
rect 42656 42920 42720 42984
rect 42736 42920 42800 42984
rect 42816 42920 42880 42984
rect 42896 42920 42960 42984
rect 42976 42920 43040 42984
rect 43056 42920 43120 42984
rect 43136 42920 43200 42984
rect 43216 42920 43280 42984
rect 43296 42920 43360 42984
rect 43376 42920 43440 42984
rect 43456 42920 43520 42984
rect 43536 42920 43600 42984
rect 43616 42920 43680 42984
rect 43696 42920 43760 42984
rect 43776 42920 43840 42984
rect 43856 42920 43920 42984
rect 43936 42920 44000 42984
rect 44016 42920 44080 42984
rect 44096 42920 44160 42984
rect 44176 42920 44240 42984
rect 44256 42920 44320 42984
rect 44336 42920 44400 42984
rect 44416 42920 44480 42984
rect 44496 42920 44560 42984
rect 44576 42920 44640 42984
rect 44656 42920 44720 42984
rect 44736 42920 44800 42984
rect 44816 42920 44880 42984
rect 44896 42920 44960 42984
rect 44976 42920 45040 42984
rect 45056 42920 45120 42984
rect 45136 42920 45200 42984
rect 45216 42920 45280 42984
rect 45296 42920 45360 42984
rect 8 42840 72 42904
rect 88 42840 152 42904
rect 168 42840 232 42904
rect 248 42840 312 42904
rect 328 42840 392 42904
rect 408 42840 472 42904
rect 488 42840 552 42904
rect 568 42840 632 42904
rect 648 42840 712 42904
rect 728 42840 792 42904
rect 808 42840 872 42904
rect 888 42840 952 42904
rect 968 42840 1032 42904
rect 1048 42840 1112 42904
rect 1128 42840 1192 42904
rect 1208 42840 1272 42904
rect 1288 42840 1352 42904
rect 1368 42840 1432 42904
rect 1448 42840 1512 42904
rect 1528 42840 1592 42904
rect 1608 42840 1672 42904
rect 1688 42840 1752 42904
rect 1768 42840 1832 42904
rect 1848 42840 1912 42904
rect 1928 42840 1992 42904
rect 2008 42840 2072 42904
rect 2088 42840 2152 42904
rect 2168 42840 2232 42904
rect 2248 42840 2312 42904
rect 2328 42840 2392 42904
rect 2408 42840 2472 42904
rect 2488 42840 2552 42904
rect 2568 42840 2632 42904
rect 2648 42840 2712 42904
rect 2728 42840 2792 42904
rect 2808 42840 2872 42904
rect 2888 42840 2952 42904
rect 2968 42840 3032 42904
rect 3048 42840 3112 42904
rect 3128 42840 3192 42904
rect 3208 42840 3272 42904
rect 3288 42840 3352 42904
rect 3368 42840 3432 42904
rect 3448 42840 3512 42904
rect 3528 42840 3592 42904
rect 3608 42840 3672 42904
rect 3688 42840 3752 42904
rect 3768 42840 3832 42904
rect 3848 42840 3912 42904
rect 3928 42840 3992 42904
rect 19112 42840 19176 42904
rect 19192 42840 19256 42904
rect 19272 42840 19336 42904
rect 19352 42840 19416 42904
rect 29112 42840 29176 42904
rect 29192 42840 29256 42904
rect 29272 42840 29336 42904
rect 29352 42840 29416 42904
rect 41376 42840 41440 42904
rect 41456 42840 41520 42904
rect 41536 42840 41600 42904
rect 41616 42840 41680 42904
rect 41696 42840 41760 42904
rect 41776 42840 41840 42904
rect 41856 42840 41920 42904
rect 41936 42840 42000 42904
rect 42016 42840 42080 42904
rect 42096 42840 42160 42904
rect 42176 42840 42240 42904
rect 42256 42840 42320 42904
rect 42336 42840 42400 42904
rect 42416 42840 42480 42904
rect 42496 42840 42560 42904
rect 42576 42840 42640 42904
rect 42656 42840 42720 42904
rect 42736 42840 42800 42904
rect 42816 42840 42880 42904
rect 42896 42840 42960 42904
rect 42976 42840 43040 42904
rect 43056 42840 43120 42904
rect 43136 42840 43200 42904
rect 43216 42840 43280 42904
rect 43296 42840 43360 42904
rect 43376 42840 43440 42904
rect 43456 42840 43520 42904
rect 43536 42840 43600 42904
rect 43616 42840 43680 42904
rect 43696 42840 43760 42904
rect 43776 42840 43840 42904
rect 43856 42840 43920 42904
rect 43936 42840 44000 42904
rect 44016 42840 44080 42904
rect 44096 42840 44160 42904
rect 44176 42840 44240 42904
rect 44256 42840 44320 42904
rect 44336 42840 44400 42904
rect 44416 42840 44480 42904
rect 44496 42840 44560 42904
rect 44576 42840 44640 42904
rect 44656 42840 44720 42904
rect 44736 42840 44800 42904
rect 44816 42840 44880 42904
rect 44896 42840 44960 42904
rect 44976 42840 45040 42904
rect 45056 42840 45120 42904
rect 45136 42840 45200 42904
rect 45216 42840 45280 42904
rect 45296 42840 45360 42904
rect 8 42760 72 42824
rect 88 42760 152 42824
rect 168 42760 232 42824
rect 248 42760 312 42824
rect 328 42760 392 42824
rect 408 42760 472 42824
rect 488 42760 552 42824
rect 568 42760 632 42824
rect 648 42760 712 42824
rect 728 42760 792 42824
rect 808 42760 872 42824
rect 888 42760 952 42824
rect 968 42760 1032 42824
rect 1048 42760 1112 42824
rect 1128 42760 1192 42824
rect 1208 42760 1272 42824
rect 1288 42760 1352 42824
rect 1368 42760 1432 42824
rect 1448 42760 1512 42824
rect 1528 42760 1592 42824
rect 1608 42760 1672 42824
rect 1688 42760 1752 42824
rect 1768 42760 1832 42824
rect 1848 42760 1912 42824
rect 1928 42760 1992 42824
rect 2008 42760 2072 42824
rect 2088 42760 2152 42824
rect 2168 42760 2232 42824
rect 2248 42760 2312 42824
rect 2328 42760 2392 42824
rect 2408 42760 2472 42824
rect 2488 42760 2552 42824
rect 2568 42760 2632 42824
rect 2648 42760 2712 42824
rect 2728 42760 2792 42824
rect 2808 42760 2872 42824
rect 2888 42760 2952 42824
rect 2968 42760 3032 42824
rect 3048 42760 3112 42824
rect 3128 42760 3192 42824
rect 3208 42760 3272 42824
rect 3288 42760 3352 42824
rect 3368 42760 3432 42824
rect 3448 42760 3512 42824
rect 3528 42760 3592 42824
rect 3608 42760 3672 42824
rect 3688 42760 3752 42824
rect 3768 42760 3832 42824
rect 3848 42760 3912 42824
rect 3928 42760 3992 42824
rect 19112 42760 19176 42824
rect 19192 42760 19256 42824
rect 19272 42760 19336 42824
rect 19352 42760 19416 42824
rect 29112 42760 29176 42824
rect 29192 42760 29256 42824
rect 29272 42760 29336 42824
rect 29352 42760 29416 42824
rect 41376 42760 41440 42824
rect 41456 42760 41520 42824
rect 41536 42760 41600 42824
rect 41616 42760 41680 42824
rect 41696 42760 41760 42824
rect 41776 42760 41840 42824
rect 41856 42760 41920 42824
rect 41936 42760 42000 42824
rect 42016 42760 42080 42824
rect 42096 42760 42160 42824
rect 42176 42760 42240 42824
rect 42256 42760 42320 42824
rect 42336 42760 42400 42824
rect 42416 42760 42480 42824
rect 42496 42760 42560 42824
rect 42576 42760 42640 42824
rect 42656 42760 42720 42824
rect 42736 42760 42800 42824
rect 42816 42760 42880 42824
rect 42896 42760 42960 42824
rect 42976 42760 43040 42824
rect 43056 42760 43120 42824
rect 43136 42760 43200 42824
rect 43216 42760 43280 42824
rect 43296 42760 43360 42824
rect 43376 42760 43440 42824
rect 43456 42760 43520 42824
rect 43536 42760 43600 42824
rect 43616 42760 43680 42824
rect 43696 42760 43760 42824
rect 43776 42760 43840 42824
rect 43856 42760 43920 42824
rect 43936 42760 44000 42824
rect 44016 42760 44080 42824
rect 44096 42760 44160 42824
rect 44176 42760 44240 42824
rect 44256 42760 44320 42824
rect 44336 42760 44400 42824
rect 44416 42760 44480 42824
rect 44496 42760 44560 42824
rect 44576 42760 44640 42824
rect 44656 42760 44720 42824
rect 44736 42760 44800 42824
rect 44816 42760 44880 42824
rect 44896 42760 44960 42824
rect 44976 42760 45040 42824
rect 45056 42760 45120 42824
rect 45136 42760 45200 42824
rect 45216 42760 45280 42824
rect 45296 42760 45360 42824
rect 8 42680 72 42744
rect 88 42680 152 42744
rect 168 42680 232 42744
rect 248 42680 312 42744
rect 328 42680 392 42744
rect 408 42680 472 42744
rect 488 42680 552 42744
rect 568 42680 632 42744
rect 648 42680 712 42744
rect 728 42680 792 42744
rect 808 42680 872 42744
rect 888 42680 952 42744
rect 968 42680 1032 42744
rect 1048 42680 1112 42744
rect 1128 42680 1192 42744
rect 1208 42680 1272 42744
rect 1288 42680 1352 42744
rect 1368 42680 1432 42744
rect 1448 42680 1512 42744
rect 1528 42680 1592 42744
rect 1608 42680 1672 42744
rect 1688 42680 1752 42744
rect 1768 42680 1832 42744
rect 1848 42680 1912 42744
rect 1928 42680 1992 42744
rect 2008 42680 2072 42744
rect 2088 42680 2152 42744
rect 2168 42680 2232 42744
rect 2248 42680 2312 42744
rect 2328 42680 2392 42744
rect 2408 42680 2472 42744
rect 2488 42680 2552 42744
rect 2568 42680 2632 42744
rect 2648 42680 2712 42744
rect 2728 42680 2792 42744
rect 2808 42680 2872 42744
rect 2888 42680 2952 42744
rect 2968 42680 3032 42744
rect 3048 42680 3112 42744
rect 3128 42680 3192 42744
rect 3208 42680 3272 42744
rect 3288 42680 3352 42744
rect 3368 42680 3432 42744
rect 3448 42680 3512 42744
rect 3528 42680 3592 42744
rect 3608 42680 3672 42744
rect 3688 42680 3752 42744
rect 3768 42680 3832 42744
rect 3848 42680 3912 42744
rect 3928 42680 3992 42744
rect 19112 42680 19176 42744
rect 19192 42680 19256 42744
rect 19272 42680 19336 42744
rect 19352 42680 19416 42744
rect 29112 42680 29176 42744
rect 29192 42680 29256 42744
rect 29272 42680 29336 42744
rect 29352 42680 29416 42744
rect 41376 42680 41440 42744
rect 41456 42680 41520 42744
rect 41536 42680 41600 42744
rect 41616 42680 41680 42744
rect 41696 42680 41760 42744
rect 41776 42680 41840 42744
rect 41856 42680 41920 42744
rect 41936 42680 42000 42744
rect 42016 42680 42080 42744
rect 42096 42680 42160 42744
rect 42176 42680 42240 42744
rect 42256 42680 42320 42744
rect 42336 42680 42400 42744
rect 42416 42680 42480 42744
rect 42496 42680 42560 42744
rect 42576 42680 42640 42744
rect 42656 42680 42720 42744
rect 42736 42680 42800 42744
rect 42816 42680 42880 42744
rect 42896 42680 42960 42744
rect 42976 42680 43040 42744
rect 43056 42680 43120 42744
rect 43136 42680 43200 42744
rect 43216 42680 43280 42744
rect 43296 42680 43360 42744
rect 43376 42680 43440 42744
rect 43456 42680 43520 42744
rect 43536 42680 43600 42744
rect 43616 42680 43680 42744
rect 43696 42680 43760 42744
rect 43776 42680 43840 42744
rect 43856 42680 43920 42744
rect 43936 42680 44000 42744
rect 44016 42680 44080 42744
rect 44096 42680 44160 42744
rect 44176 42680 44240 42744
rect 44256 42680 44320 42744
rect 44336 42680 44400 42744
rect 44416 42680 44480 42744
rect 44496 42680 44560 42744
rect 44576 42680 44640 42744
rect 44656 42680 44720 42744
rect 44736 42680 44800 42744
rect 44816 42680 44880 42744
rect 44896 42680 44960 42744
rect 44976 42680 45040 42744
rect 45056 42680 45120 42744
rect 45136 42680 45200 42744
rect 45216 42680 45280 42744
rect 45296 42680 45360 42744
rect 8 42600 72 42664
rect 88 42600 152 42664
rect 168 42600 232 42664
rect 248 42600 312 42664
rect 328 42600 392 42664
rect 408 42600 472 42664
rect 488 42600 552 42664
rect 568 42600 632 42664
rect 648 42600 712 42664
rect 728 42600 792 42664
rect 808 42600 872 42664
rect 888 42600 952 42664
rect 968 42600 1032 42664
rect 1048 42600 1112 42664
rect 1128 42600 1192 42664
rect 1208 42600 1272 42664
rect 1288 42600 1352 42664
rect 1368 42600 1432 42664
rect 1448 42600 1512 42664
rect 1528 42600 1592 42664
rect 1608 42600 1672 42664
rect 1688 42600 1752 42664
rect 1768 42600 1832 42664
rect 1848 42600 1912 42664
rect 1928 42600 1992 42664
rect 2008 42600 2072 42664
rect 2088 42600 2152 42664
rect 2168 42600 2232 42664
rect 2248 42600 2312 42664
rect 2328 42600 2392 42664
rect 2408 42600 2472 42664
rect 2488 42600 2552 42664
rect 2568 42600 2632 42664
rect 2648 42600 2712 42664
rect 2728 42600 2792 42664
rect 2808 42600 2872 42664
rect 2888 42600 2952 42664
rect 2968 42600 3032 42664
rect 3048 42600 3112 42664
rect 3128 42600 3192 42664
rect 3208 42600 3272 42664
rect 3288 42600 3352 42664
rect 3368 42600 3432 42664
rect 3448 42600 3512 42664
rect 3528 42600 3592 42664
rect 3608 42600 3672 42664
rect 3688 42600 3752 42664
rect 3768 42600 3832 42664
rect 3848 42600 3912 42664
rect 3928 42600 3992 42664
rect 19112 42600 19176 42664
rect 19192 42600 19256 42664
rect 19272 42600 19336 42664
rect 19352 42600 19416 42664
rect 29112 42600 29176 42664
rect 29192 42600 29256 42664
rect 29272 42600 29336 42664
rect 29352 42600 29416 42664
rect 41376 42600 41440 42664
rect 41456 42600 41520 42664
rect 41536 42600 41600 42664
rect 41616 42600 41680 42664
rect 41696 42600 41760 42664
rect 41776 42600 41840 42664
rect 41856 42600 41920 42664
rect 41936 42600 42000 42664
rect 42016 42600 42080 42664
rect 42096 42600 42160 42664
rect 42176 42600 42240 42664
rect 42256 42600 42320 42664
rect 42336 42600 42400 42664
rect 42416 42600 42480 42664
rect 42496 42600 42560 42664
rect 42576 42600 42640 42664
rect 42656 42600 42720 42664
rect 42736 42600 42800 42664
rect 42816 42600 42880 42664
rect 42896 42600 42960 42664
rect 42976 42600 43040 42664
rect 43056 42600 43120 42664
rect 43136 42600 43200 42664
rect 43216 42600 43280 42664
rect 43296 42600 43360 42664
rect 43376 42600 43440 42664
rect 43456 42600 43520 42664
rect 43536 42600 43600 42664
rect 43616 42600 43680 42664
rect 43696 42600 43760 42664
rect 43776 42600 43840 42664
rect 43856 42600 43920 42664
rect 43936 42600 44000 42664
rect 44016 42600 44080 42664
rect 44096 42600 44160 42664
rect 44176 42600 44240 42664
rect 44256 42600 44320 42664
rect 44336 42600 44400 42664
rect 44416 42600 44480 42664
rect 44496 42600 44560 42664
rect 44576 42600 44640 42664
rect 44656 42600 44720 42664
rect 44736 42600 44800 42664
rect 44816 42600 44880 42664
rect 44896 42600 44960 42664
rect 44976 42600 45040 42664
rect 45056 42600 45120 42664
rect 45136 42600 45200 42664
rect 45216 42600 45280 42664
rect 45296 42600 45360 42664
rect 8 42520 72 42584
rect 88 42520 152 42584
rect 168 42520 232 42584
rect 248 42520 312 42584
rect 328 42520 392 42584
rect 408 42520 472 42584
rect 488 42520 552 42584
rect 568 42520 632 42584
rect 648 42520 712 42584
rect 728 42520 792 42584
rect 808 42520 872 42584
rect 888 42520 952 42584
rect 968 42520 1032 42584
rect 1048 42520 1112 42584
rect 1128 42520 1192 42584
rect 1208 42520 1272 42584
rect 1288 42520 1352 42584
rect 1368 42520 1432 42584
rect 1448 42520 1512 42584
rect 1528 42520 1592 42584
rect 1608 42520 1672 42584
rect 1688 42520 1752 42584
rect 1768 42520 1832 42584
rect 1848 42520 1912 42584
rect 1928 42520 1992 42584
rect 2008 42520 2072 42584
rect 2088 42520 2152 42584
rect 2168 42520 2232 42584
rect 2248 42520 2312 42584
rect 2328 42520 2392 42584
rect 2408 42520 2472 42584
rect 2488 42520 2552 42584
rect 2568 42520 2632 42584
rect 2648 42520 2712 42584
rect 2728 42520 2792 42584
rect 2808 42520 2872 42584
rect 2888 42520 2952 42584
rect 2968 42520 3032 42584
rect 3048 42520 3112 42584
rect 3128 42520 3192 42584
rect 3208 42520 3272 42584
rect 3288 42520 3352 42584
rect 3368 42520 3432 42584
rect 3448 42520 3512 42584
rect 3528 42520 3592 42584
rect 3608 42520 3672 42584
rect 3688 42520 3752 42584
rect 3768 42520 3832 42584
rect 3848 42520 3912 42584
rect 3928 42520 3992 42584
rect 19112 42520 19176 42584
rect 19192 42520 19256 42584
rect 19272 42520 19336 42584
rect 19352 42520 19416 42584
rect 29112 42520 29176 42584
rect 29192 42520 29256 42584
rect 29272 42520 29336 42584
rect 29352 42520 29416 42584
rect 41376 42520 41440 42584
rect 41456 42520 41520 42584
rect 41536 42520 41600 42584
rect 41616 42520 41680 42584
rect 41696 42520 41760 42584
rect 41776 42520 41840 42584
rect 41856 42520 41920 42584
rect 41936 42520 42000 42584
rect 42016 42520 42080 42584
rect 42096 42520 42160 42584
rect 42176 42520 42240 42584
rect 42256 42520 42320 42584
rect 42336 42520 42400 42584
rect 42416 42520 42480 42584
rect 42496 42520 42560 42584
rect 42576 42520 42640 42584
rect 42656 42520 42720 42584
rect 42736 42520 42800 42584
rect 42816 42520 42880 42584
rect 42896 42520 42960 42584
rect 42976 42520 43040 42584
rect 43056 42520 43120 42584
rect 43136 42520 43200 42584
rect 43216 42520 43280 42584
rect 43296 42520 43360 42584
rect 43376 42520 43440 42584
rect 43456 42520 43520 42584
rect 43536 42520 43600 42584
rect 43616 42520 43680 42584
rect 43696 42520 43760 42584
rect 43776 42520 43840 42584
rect 43856 42520 43920 42584
rect 43936 42520 44000 42584
rect 44016 42520 44080 42584
rect 44096 42520 44160 42584
rect 44176 42520 44240 42584
rect 44256 42520 44320 42584
rect 44336 42520 44400 42584
rect 44416 42520 44480 42584
rect 44496 42520 44560 42584
rect 44576 42520 44640 42584
rect 44656 42520 44720 42584
rect 44736 42520 44800 42584
rect 44816 42520 44880 42584
rect 44896 42520 44960 42584
rect 44976 42520 45040 42584
rect 45056 42520 45120 42584
rect 45136 42520 45200 42584
rect 45216 42520 45280 42584
rect 45296 42520 45360 42584
rect 8 42440 72 42504
rect 88 42440 152 42504
rect 168 42440 232 42504
rect 248 42440 312 42504
rect 328 42440 392 42504
rect 408 42440 472 42504
rect 488 42440 552 42504
rect 568 42440 632 42504
rect 648 42440 712 42504
rect 728 42440 792 42504
rect 808 42440 872 42504
rect 888 42440 952 42504
rect 968 42440 1032 42504
rect 1048 42440 1112 42504
rect 1128 42440 1192 42504
rect 1208 42440 1272 42504
rect 1288 42440 1352 42504
rect 1368 42440 1432 42504
rect 1448 42440 1512 42504
rect 1528 42440 1592 42504
rect 1608 42440 1672 42504
rect 1688 42440 1752 42504
rect 1768 42440 1832 42504
rect 1848 42440 1912 42504
rect 1928 42440 1992 42504
rect 2008 42440 2072 42504
rect 2088 42440 2152 42504
rect 2168 42440 2232 42504
rect 2248 42440 2312 42504
rect 2328 42440 2392 42504
rect 2408 42440 2472 42504
rect 2488 42440 2552 42504
rect 2568 42440 2632 42504
rect 2648 42440 2712 42504
rect 2728 42440 2792 42504
rect 2808 42440 2872 42504
rect 2888 42440 2952 42504
rect 2968 42440 3032 42504
rect 3048 42440 3112 42504
rect 3128 42440 3192 42504
rect 3208 42440 3272 42504
rect 3288 42440 3352 42504
rect 3368 42440 3432 42504
rect 3448 42440 3512 42504
rect 3528 42440 3592 42504
rect 3608 42440 3672 42504
rect 3688 42440 3752 42504
rect 3768 42440 3832 42504
rect 3848 42440 3912 42504
rect 3928 42440 3992 42504
rect 19112 42440 19176 42504
rect 19192 42440 19256 42504
rect 19272 42440 19336 42504
rect 19352 42440 19416 42504
rect 29112 42440 29176 42504
rect 29192 42440 29256 42504
rect 29272 42440 29336 42504
rect 29352 42440 29416 42504
rect 41376 42440 41440 42504
rect 41456 42440 41520 42504
rect 41536 42440 41600 42504
rect 41616 42440 41680 42504
rect 41696 42440 41760 42504
rect 41776 42440 41840 42504
rect 41856 42440 41920 42504
rect 41936 42440 42000 42504
rect 42016 42440 42080 42504
rect 42096 42440 42160 42504
rect 42176 42440 42240 42504
rect 42256 42440 42320 42504
rect 42336 42440 42400 42504
rect 42416 42440 42480 42504
rect 42496 42440 42560 42504
rect 42576 42440 42640 42504
rect 42656 42440 42720 42504
rect 42736 42440 42800 42504
rect 42816 42440 42880 42504
rect 42896 42440 42960 42504
rect 42976 42440 43040 42504
rect 43056 42440 43120 42504
rect 43136 42440 43200 42504
rect 43216 42440 43280 42504
rect 43296 42440 43360 42504
rect 43376 42440 43440 42504
rect 43456 42440 43520 42504
rect 43536 42440 43600 42504
rect 43616 42440 43680 42504
rect 43696 42440 43760 42504
rect 43776 42440 43840 42504
rect 43856 42440 43920 42504
rect 43936 42440 44000 42504
rect 44016 42440 44080 42504
rect 44096 42440 44160 42504
rect 44176 42440 44240 42504
rect 44256 42440 44320 42504
rect 44336 42440 44400 42504
rect 44416 42440 44480 42504
rect 44496 42440 44560 42504
rect 44576 42440 44640 42504
rect 44656 42440 44720 42504
rect 44736 42440 44800 42504
rect 44816 42440 44880 42504
rect 44896 42440 44960 42504
rect 44976 42440 45040 42504
rect 45056 42440 45120 42504
rect 45136 42440 45200 42504
rect 45216 42440 45280 42504
rect 45296 42440 45360 42504
rect 8 42360 72 42424
rect 88 42360 152 42424
rect 168 42360 232 42424
rect 248 42360 312 42424
rect 328 42360 392 42424
rect 408 42360 472 42424
rect 488 42360 552 42424
rect 568 42360 632 42424
rect 648 42360 712 42424
rect 728 42360 792 42424
rect 808 42360 872 42424
rect 888 42360 952 42424
rect 968 42360 1032 42424
rect 1048 42360 1112 42424
rect 1128 42360 1192 42424
rect 1208 42360 1272 42424
rect 1288 42360 1352 42424
rect 1368 42360 1432 42424
rect 1448 42360 1512 42424
rect 1528 42360 1592 42424
rect 1608 42360 1672 42424
rect 1688 42360 1752 42424
rect 1768 42360 1832 42424
rect 1848 42360 1912 42424
rect 1928 42360 1992 42424
rect 2008 42360 2072 42424
rect 2088 42360 2152 42424
rect 2168 42360 2232 42424
rect 2248 42360 2312 42424
rect 2328 42360 2392 42424
rect 2408 42360 2472 42424
rect 2488 42360 2552 42424
rect 2568 42360 2632 42424
rect 2648 42360 2712 42424
rect 2728 42360 2792 42424
rect 2808 42360 2872 42424
rect 2888 42360 2952 42424
rect 2968 42360 3032 42424
rect 3048 42360 3112 42424
rect 3128 42360 3192 42424
rect 3208 42360 3272 42424
rect 3288 42360 3352 42424
rect 3368 42360 3432 42424
rect 3448 42360 3512 42424
rect 3528 42360 3592 42424
rect 3608 42360 3672 42424
rect 3688 42360 3752 42424
rect 3768 42360 3832 42424
rect 3848 42360 3912 42424
rect 3928 42360 3992 42424
rect 19112 42360 19176 42424
rect 19192 42360 19256 42424
rect 19272 42360 19336 42424
rect 19352 42360 19416 42424
rect 29112 42360 29176 42424
rect 29192 42360 29256 42424
rect 29272 42360 29336 42424
rect 29352 42360 29416 42424
rect 41376 42360 41440 42424
rect 41456 42360 41520 42424
rect 41536 42360 41600 42424
rect 41616 42360 41680 42424
rect 41696 42360 41760 42424
rect 41776 42360 41840 42424
rect 41856 42360 41920 42424
rect 41936 42360 42000 42424
rect 42016 42360 42080 42424
rect 42096 42360 42160 42424
rect 42176 42360 42240 42424
rect 42256 42360 42320 42424
rect 42336 42360 42400 42424
rect 42416 42360 42480 42424
rect 42496 42360 42560 42424
rect 42576 42360 42640 42424
rect 42656 42360 42720 42424
rect 42736 42360 42800 42424
rect 42816 42360 42880 42424
rect 42896 42360 42960 42424
rect 42976 42360 43040 42424
rect 43056 42360 43120 42424
rect 43136 42360 43200 42424
rect 43216 42360 43280 42424
rect 43296 42360 43360 42424
rect 43376 42360 43440 42424
rect 43456 42360 43520 42424
rect 43536 42360 43600 42424
rect 43616 42360 43680 42424
rect 43696 42360 43760 42424
rect 43776 42360 43840 42424
rect 43856 42360 43920 42424
rect 43936 42360 44000 42424
rect 44016 42360 44080 42424
rect 44096 42360 44160 42424
rect 44176 42360 44240 42424
rect 44256 42360 44320 42424
rect 44336 42360 44400 42424
rect 44416 42360 44480 42424
rect 44496 42360 44560 42424
rect 44576 42360 44640 42424
rect 44656 42360 44720 42424
rect 44736 42360 44800 42424
rect 44816 42360 44880 42424
rect 44896 42360 44960 42424
rect 44976 42360 45040 42424
rect 45056 42360 45120 42424
rect 45136 42360 45200 42424
rect 45216 42360 45280 42424
rect 45296 42360 45360 42424
rect 8 42280 72 42344
rect 88 42280 152 42344
rect 168 42280 232 42344
rect 248 42280 312 42344
rect 328 42280 392 42344
rect 408 42280 472 42344
rect 488 42280 552 42344
rect 568 42280 632 42344
rect 648 42280 712 42344
rect 728 42280 792 42344
rect 808 42280 872 42344
rect 888 42280 952 42344
rect 968 42280 1032 42344
rect 1048 42280 1112 42344
rect 1128 42280 1192 42344
rect 1208 42280 1272 42344
rect 1288 42280 1352 42344
rect 1368 42280 1432 42344
rect 1448 42280 1512 42344
rect 1528 42280 1592 42344
rect 1608 42280 1672 42344
rect 1688 42280 1752 42344
rect 1768 42280 1832 42344
rect 1848 42280 1912 42344
rect 1928 42280 1992 42344
rect 2008 42280 2072 42344
rect 2088 42280 2152 42344
rect 2168 42280 2232 42344
rect 2248 42280 2312 42344
rect 2328 42280 2392 42344
rect 2408 42280 2472 42344
rect 2488 42280 2552 42344
rect 2568 42280 2632 42344
rect 2648 42280 2712 42344
rect 2728 42280 2792 42344
rect 2808 42280 2872 42344
rect 2888 42280 2952 42344
rect 2968 42280 3032 42344
rect 3048 42280 3112 42344
rect 3128 42280 3192 42344
rect 3208 42280 3272 42344
rect 3288 42280 3352 42344
rect 3368 42280 3432 42344
rect 3448 42280 3512 42344
rect 3528 42280 3592 42344
rect 3608 42280 3672 42344
rect 3688 42280 3752 42344
rect 3768 42280 3832 42344
rect 3848 42280 3912 42344
rect 3928 42280 3992 42344
rect 19112 42280 19176 42344
rect 19192 42280 19256 42344
rect 19272 42280 19336 42344
rect 19352 42280 19416 42344
rect 29112 42280 29176 42344
rect 29192 42280 29256 42344
rect 29272 42280 29336 42344
rect 29352 42280 29416 42344
rect 41376 42280 41440 42344
rect 41456 42280 41520 42344
rect 41536 42280 41600 42344
rect 41616 42280 41680 42344
rect 41696 42280 41760 42344
rect 41776 42280 41840 42344
rect 41856 42280 41920 42344
rect 41936 42280 42000 42344
rect 42016 42280 42080 42344
rect 42096 42280 42160 42344
rect 42176 42280 42240 42344
rect 42256 42280 42320 42344
rect 42336 42280 42400 42344
rect 42416 42280 42480 42344
rect 42496 42280 42560 42344
rect 42576 42280 42640 42344
rect 42656 42280 42720 42344
rect 42736 42280 42800 42344
rect 42816 42280 42880 42344
rect 42896 42280 42960 42344
rect 42976 42280 43040 42344
rect 43056 42280 43120 42344
rect 43136 42280 43200 42344
rect 43216 42280 43280 42344
rect 43296 42280 43360 42344
rect 43376 42280 43440 42344
rect 43456 42280 43520 42344
rect 43536 42280 43600 42344
rect 43616 42280 43680 42344
rect 43696 42280 43760 42344
rect 43776 42280 43840 42344
rect 43856 42280 43920 42344
rect 43936 42280 44000 42344
rect 44016 42280 44080 42344
rect 44096 42280 44160 42344
rect 44176 42280 44240 42344
rect 44256 42280 44320 42344
rect 44336 42280 44400 42344
rect 44416 42280 44480 42344
rect 44496 42280 44560 42344
rect 44576 42280 44640 42344
rect 44656 42280 44720 42344
rect 44736 42280 44800 42344
rect 44816 42280 44880 42344
rect 44896 42280 44960 42344
rect 44976 42280 45040 42344
rect 45056 42280 45120 42344
rect 45136 42280 45200 42344
rect 45216 42280 45280 42344
rect 45296 42280 45360 42344
rect 8 42200 72 42264
rect 88 42200 152 42264
rect 168 42200 232 42264
rect 248 42200 312 42264
rect 328 42200 392 42264
rect 408 42200 472 42264
rect 488 42200 552 42264
rect 568 42200 632 42264
rect 648 42200 712 42264
rect 728 42200 792 42264
rect 808 42200 872 42264
rect 888 42200 952 42264
rect 968 42200 1032 42264
rect 1048 42200 1112 42264
rect 1128 42200 1192 42264
rect 1208 42200 1272 42264
rect 1288 42200 1352 42264
rect 1368 42200 1432 42264
rect 1448 42200 1512 42264
rect 1528 42200 1592 42264
rect 1608 42200 1672 42264
rect 1688 42200 1752 42264
rect 1768 42200 1832 42264
rect 1848 42200 1912 42264
rect 1928 42200 1992 42264
rect 2008 42200 2072 42264
rect 2088 42200 2152 42264
rect 2168 42200 2232 42264
rect 2248 42200 2312 42264
rect 2328 42200 2392 42264
rect 2408 42200 2472 42264
rect 2488 42200 2552 42264
rect 2568 42200 2632 42264
rect 2648 42200 2712 42264
rect 2728 42200 2792 42264
rect 2808 42200 2872 42264
rect 2888 42200 2952 42264
rect 2968 42200 3032 42264
rect 3048 42200 3112 42264
rect 3128 42200 3192 42264
rect 3208 42200 3272 42264
rect 3288 42200 3352 42264
rect 3368 42200 3432 42264
rect 3448 42200 3512 42264
rect 3528 42200 3592 42264
rect 3608 42200 3672 42264
rect 3688 42200 3752 42264
rect 3768 42200 3832 42264
rect 3848 42200 3912 42264
rect 3928 42200 3992 42264
rect 19112 42200 19176 42264
rect 19192 42200 19256 42264
rect 19272 42200 19336 42264
rect 19352 42200 19416 42264
rect 29112 42200 29176 42264
rect 29192 42200 29256 42264
rect 29272 42200 29336 42264
rect 29352 42200 29416 42264
rect 41376 42200 41440 42264
rect 41456 42200 41520 42264
rect 41536 42200 41600 42264
rect 41616 42200 41680 42264
rect 41696 42200 41760 42264
rect 41776 42200 41840 42264
rect 41856 42200 41920 42264
rect 41936 42200 42000 42264
rect 42016 42200 42080 42264
rect 42096 42200 42160 42264
rect 42176 42200 42240 42264
rect 42256 42200 42320 42264
rect 42336 42200 42400 42264
rect 42416 42200 42480 42264
rect 42496 42200 42560 42264
rect 42576 42200 42640 42264
rect 42656 42200 42720 42264
rect 42736 42200 42800 42264
rect 42816 42200 42880 42264
rect 42896 42200 42960 42264
rect 42976 42200 43040 42264
rect 43056 42200 43120 42264
rect 43136 42200 43200 42264
rect 43216 42200 43280 42264
rect 43296 42200 43360 42264
rect 43376 42200 43440 42264
rect 43456 42200 43520 42264
rect 43536 42200 43600 42264
rect 43616 42200 43680 42264
rect 43696 42200 43760 42264
rect 43776 42200 43840 42264
rect 43856 42200 43920 42264
rect 43936 42200 44000 42264
rect 44016 42200 44080 42264
rect 44096 42200 44160 42264
rect 44176 42200 44240 42264
rect 44256 42200 44320 42264
rect 44336 42200 44400 42264
rect 44416 42200 44480 42264
rect 44496 42200 44560 42264
rect 44576 42200 44640 42264
rect 44656 42200 44720 42264
rect 44736 42200 44800 42264
rect 44816 42200 44880 42264
rect 44896 42200 44960 42264
rect 44976 42200 45040 42264
rect 45056 42200 45120 42264
rect 45136 42200 45200 42264
rect 45216 42200 45280 42264
rect 45296 42200 45360 42264
rect 8 42120 72 42184
rect 88 42120 152 42184
rect 168 42120 232 42184
rect 248 42120 312 42184
rect 328 42120 392 42184
rect 408 42120 472 42184
rect 488 42120 552 42184
rect 568 42120 632 42184
rect 648 42120 712 42184
rect 728 42120 792 42184
rect 808 42120 872 42184
rect 888 42120 952 42184
rect 968 42120 1032 42184
rect 1048 42120 1112 42184
rect 1128 42120 1192 42184
rect 1208 42120 1272 42184
rect 1288 42120 1352 42184
rect 1368 42120 1432 42184
rect 1448 42120 1512 42184
rect 1528 42120 1592 42184
rect 1608 42120 1672 42184
rect 1688 42120 1752 42184
rect 1768 42120 1832 42184
rect 1848 42120 1912 42184
rect 1928 42120 1992 42184
rect 2008 42120 2072 42184
rect 2088 42120 2152 42184
rect 2168 42120 2232 42184
rect 2248 42120 2312 42184
rect 2328 42120 2392 42184
rect 2408 42120 2472 42184
rect 2488 42120 2552 42184
rect 2568 42120 2632 42184
rect 2648 42120 2712 42184
rect 2728 42120 2792 42184
rect 2808 42120 2872 42184
rect 2888 42120 2952 42184
rect 2968 42120 3032 42184
rect 3048 42120 3112 42184
rect 3128 42120 3192 42184
rect 3208 42120 3272 42184
rect 3288 42120 3352 42184
rect 3368 42120 3432 42184
rect 3448 42120 3512 42184
rect 3528 42120 3592 42184
rect 3608 42120 3672 42184
rect 3688 42120 3752 42184
rect 3768 42120 3832 42184
rect 3848 42120 3912 42184
rect 3928 42120 3992 42184
rect 19112 42120 19176 42184
rect 19192 42120 19256 42184
rect 19272 42120 19336 42184
rect 19352 42120 19416 42184
rect 29112 42120 29176 42184
rect 29192 42120 29256 42184
rect 29272 42120 29336 42184
rect 29352 42120 29416 42184
rect 41376 42120 41440 42184
rect 41456 42120 41520 42184
rect 41536 42120 41600 42184
rect 41616 42120 41680 42184
rect 41696 42120 41760 42184
rect 41776 42120 41840 42184
rect 41856 42120 41920 42184
rect 41936 42120 42000 42184
rect 42016 42120 42080 42184
rect 42096 42120 42160 42184
rect 42176 42120 42240 42184
rect 42256 42120 42320 42184
rect 42336 42120 42400 42184
rect 42416 42120 42480 42184
rect 42496 42120 42560 42184
rect 42576 42120 42640 42184
rect 42656 42120 42720 42184
rect 42736 42120 42800 42184
rect 42816 42120 42880 42184
rect 42896 42120 42960 42184
rect 42976 42120 43040 42184
rect 43056 42120 43120 42184
rect 43136 42120 43200 42184
rect 43216 42120 43280 42184
rect 43296 42120 43360 42184
rect 43376 42120 43440 42184
rect 43456 42120 43520 42184
rect 43536 42120 43600 42184
rect 43616 42120 43680 42184
rect 43696 42120 43760 42184
rect 43776 42120 43840 42184
rect 43856 42120 43920 42184
rect 43936 42120 44000 42184
rect 44016 42120 44080 42184
rect 44096 42120 44160 42184
rect 44176 42120 44240 42184
rect 44256 42120 44320 42184
rect 44336 42120 44400 42184
rect 44416 42120 44480 42184
rect 44496 42120 44560 42184
rect 44576 42120 44640 42184
rect 44656 42120 44720 42184
rect 44736 42120 44800 42184
rect 44816 42120 44880 42184
rect 44896 42120 44960 42184
rect 44976 42120 45040 42184
rect 45056 42120 45120 42184
rect 45136 42120 45200 42184
rect 45216 42120 45280 42184
rect 45296 42120 45360 42184
rect 8 42040 72 42104
rect 88 42040 152 42104
rect 168 42040 232 42104
rect 248 42040 312 42104
rect 328 42040 392 42104
rect 408 42040 472 42104
rect 488 42040 552 42104
rect 568 42040 632 42104
rect 648 42040 712 42104
rect 728 42040 792 42104
rect 808 42040 872 42104
rect 888 42040 952 42104
rect 968 42040 1032 42104
rect 1048 42040 1112 42104
rect 1128 42040 1192 42104
rect 1208 42040 1272 42104
rect 1288 42040 1352 42104
rect 1368 42040 1432 42104
rect 1448 42040 1512 42104
rect 1528 42040 1592 42104
rect 1608 42040 1672 42104
rect 1688 42040 1752 42104
rect 1768 42040 1832 42104
rect 1848 42040 1912 42104
rect 1928 42040 1992 42104
rect 2008 42040 2072 42104
rect 2088 42040 2152 42104
rect 2168 42040 2232 42104
rect 2248 42040 2312 42104
rect 2328 42040 2392 42104
rect 2408 42040 2472 42104
rect 2488 42040 2552 42104
rect 2568 42040 2632 42104
rect 2648 42040 2712 42104
rect 2728 42040 2792 42104
rect 2808 42040 2872 42104
rect 2888 42040 2952 42104
rect 2968 42040 3032 42104
rect 3048 42040 3112 42104
rect 3128 42040 3192 42104
rect 3208 42040 3272 42104
rect 3288 42040 3352 42104
rect 3368 42040 3432 42104
rect 3448 42040 3512 42104
rect 3528 42040 3592 42104
rect 3608 42040 3672 42104
rect 3688 42040 3752 42104
rect 3768 42040 3832 42104
rect 3848 42040 3912 42104
rect 3928 42040 3992 42104
rect 19112 42040 19176 42104
rect 19192 42040 19256 42104
rect 19272 42040 19336 42104
rect 19352 42040 19416 42104
rect 29112 42040 29176 42104
rect 29192 42040 29256 42104
rect 29272 42040 29336 42104
rect 29352 42040 29416 42104
rect 41376 42040 41440 42104
rect 41456 42040 41520 42104
rect 41536 42040 41600 42104
rect 41616 42040 41680 42104
rect 41696 42040 41760 42104
rect 41776 42040 41840 42104
rect 41856 42040 41920 42104
rect 41936 42040 42000 42104
rect 42016 42040 42080 42104
rect 42096 42040 42160 42104
rect 42176 42040 42240 42104
rect 42256 42040 42320 42104
rect 42336 42040 42400 42104
rect 42416 42040 42480 42104
rect 42496 42040 42560 42104
rect 42576 42040 42640 42104
rect 42656 42040 42720 42104
rect 42736 42040 42800 42104
rect 42816 42040 42880 42104
rect 42896 42040 42960 42104
rect 42976 42040 43040 42104
rect 43056 42040 43120 42104
rect 43136 42040 43200 42104
rect 43216 42040 43280 42104
rect 43296 42040 43360 42104
rect 43376 42040 43440 42104
rect 43456 42040 43520 42104
rect 43536 42040 43600 42104
rect 43616 42040 43680 42104
rect 43696 42040 43760 42104
rect 43776 42040 43840 42104
rect 43856 42040 43920 42104
rect 43936 42040 44000 42104
rect 44016 42040 44080 42104
rect 44096 42040 44160 42104
rect 44176 42040 44240 42104
rect 44256 42040 44320 42104
rect 44336 42040 44400 42104
rect 44416 42040 44480 42104
rect 44496 42040 44560 42104
rect 44576 42040 44640 42104
rect 44656 42040 44720 42104
rect 44736 42040 44800 42104
rect 44816 42040 44880 42104
rect 44896 42040 44960 42104
rect 44976 42040 45040 42104
rect 45056 42040 45120 42104
rect 45136 42040 45200 42104
rect 45216 42040 45280 42104
rect 45296 42040 45360 42104
rect 8 41960 72 42024
rect 88 41960 152 42024
rect 168 41960 232 42024
rect 248 41960 312 42024
rect 328 41960 392 42024
rect 408 41960 472 42024
rect 488 41960 552 42024
rect 568 41960 632 42024
rect 648 41960 712 42024
rect 728 41960 792 42024
rect 808 41960 872 42024
rect 888 41960 952 42024
rect 968 41960 1032 42024
rect 1048 41960 1112 42024
rect 1128 41960 1192 42024
rect 1208 41960 1272 42024
rect 1288 41960 1352 42024
rect 1368 41960 1432 42024
rect 1448 41960 1512 42024
rect 1528 41960 1592 42024
rect 1608 41960 1672 42024
rect 1688 41960 1752 42024
rect 1768 41960 1832 42024
rect 1848 41960 1912 42024
rect 1928 41960 1992 42024
rect 2008 41960 2072 42024
rect 2088 41960 2152 42024
rect 2168 41960 2232 42024
rect 2248 41960 2312 42024
rect 2328 41960 2392 42024
rect 2408 41960 2472 42024
rect 2488 41960 2552 42024
rect 2568 41960 2632 42024
rect 2648 41960 2712 42024
rect 2728 41960 2792 42024
rect 2808 41960 2872 42024
rect 2888 41960 2952 42024
rect 2968 41960 3032 42024
rect 3048 41960 3112 42024
rect 3128 41960 3192 42024
rect 3208 41960 3272 42024
rect 3288 41960 3352 42024
rect 3368 41960 3432 42024
rect 3448 41960 3512 42024
rect 3528 41960 3592 42024
rect 3608 41960 3672 42024
rect 3688 41960 3752 42024
rect 3768 41960 3832 42024
rect 3848 41960 3912 42024
rect 3928 41960 3992 42024
rect 19112 41960 19176 42024
rect 19192 41960 19256 42024
rect 19272 41960 19336 42024
rect 19352 41960 19416 42024
rect 29112 41960 29176 42024
rect 29192 41960 29256 42024
rect 29272 41960 29336 42024
rect 29352 41960 29416 42024
rect 41376 41960 41440 42024
rect 41456 41960 41520 42024
rect 41536 41960 41600 42024
rect 41616 41960 41680 42024
rect 41696 41960 41760 42024
rect 41776 41960 41840 42024
rect 41856 41960 41920 42024
rect 41936 41960 42000 42024
rect 42016 41960 42080 42024
rect 42096 41960 42160 42024
rect 42176 41960 42240 42024
rect 42256 41960 42320 42024
rect 42336 41960 42400 42024
rect 42416 41960 42480 42024
rect 42496 41960 42560 42024
rect 42576 41960 42640 42024
rect 42656 41960 42720 42024
rect 42736 41960 42800 42024
rect 42816 41960 42880 42024
rect 42896 41960 42960 42024
rect 42976 41960 43040 42024
rect 43056 41960 43120 42024
rect 43136 41960 43200 42024
rect 43216 41960 43280 42024
rect 43296 41960 43360 42024
rect 43376 41960 43440 42024
rect 43456 41960 43520 42024
rect 43536 41960 43600 42024
rect 43616 41960 43680 42024
rect 43696 41960 43760 42024
rect 43776 41960 43840 42024
rect 43856 41960 43920 42024
rect 43936 41960 44000 42024
rect 44016 41960 44080 42024
rect 44096 41960 44160 42024
rect 44176 41960 44240 42024
rect 44256 41960 44320 42024
rect 44336 41960 44400 42024
rect 44416 41960 44480 42024
rect 44496 41960 44560 42024
rect 44576 41960 44640 42024
rect 44656 41960 44720 42024
rect 44736 41960 44800 42024
rect 44816 41960 44880 42024
rect 44896 41960 44960 42024
rect 44976 41960 45040 42024
rect 45056 41960 45120 42024
rect 45136 41960 45200 42024
rect 45216 41960 45280 42024
rect 45296 41960 45360 42024
rect 8 41880 72 41944
rect 88 41880 152 41944
rect 168 41880 232 41944
rect 248 41880 312 41944
rect 328 41880 392 41944
rect 408 41880 472 41944
rect 488 41880 552 41944
rect 568 41880 632 41944
rect 648 41880 712 41944
rect 728 41880 792 41944
rect 808 41880 872 41944
rect 888 41880 952 41944
rect 968 41880 1032 41944
rect 1048 41880 1112 41944
rect 1128 41880 1192 41944
rect 1208 41880 1272 41944
rect 1288 41880 1352 41944
rect 1368 41880 1432 41944
rect 1448 41880 1512 41944
rect 1528 41880 1592 41944
rect 1608 41880 1672 41944
rect 1688 41880 1752 41944
rect 1768 41880 1832 41944
rect 1848 41880 1912 41944
rect 1928 41880 1992 41944
rect 2008 41880 2072 41944
rect 2088 41880 2152 41944
rect 2168 41880 2232 41944
rect 2248 41880 2312 41944
rect 2328 41880 2392 41944
rect 2408 41880 2472 41944
rect 2488 41880 2552 41944
rect 2568 41880 2632 41944
rect 2648 41880 2712 41944
rect 2728 41880 2792 41944
rect 2808 41880 2872 41944
rect 2888 41880 2952 41944
rect 2968 41880 3032 41944
rect 3048 41880 3112 41944
rect 3128 41880 3192 41944
rect 3208 41880 3272 41944
rect 3288 41880 3352 41944
rect 3368 41880 3432 41944
rect 3448 41880 3512 41944
rect 3528 41880 3592 41944
rect 3608 41880 3672 41944
rect 3688 41880 3752 41944
rect 3768 41880 3832 41944
rect 3848 41880 3912 41944
rect 3928 41880 3992 41944
rect 19112 41880 19176 41944
rect 19192 41880 19256 41944
rect 19272 41880 19336 41944
rect 19352 41880 19416 41944
rect 29112 41880 29176 41944
rect 29192 41880 29256 41944
rect 29272 41880 29336 41944
rect 29352 41880 29416 41944
rect 41376 41880 41440 41944
rect 41456 41880 41520 41944
rect 41536 41880 41600 41944
rect 41616 41880 41680 41944
rect 41696 41880 41760 41944
rect 41776 41880 41840 41944
rect 41856 41880 41920 41944
rect 41936 41880 42000 41944
rect 42016 41880 42080 41944
rect 42096 41880 42160 41944
rect 42176 41880 42240 41944
rect 42256 41880 42320 41944
rect 42336 41880 42400 41944
rect 42416 41880 42480 41944
rect 42496 41880 42560 41944
rect 42576 41880 42640 41944
rect 42656 41880 42720 41944
rect 42736 41880 42800 41944
rect 42816 41880 42880 41944
rect 42896 41880 42960 41944
rect 42976 41880 43040 41944
rect 43056 41880 43120 41944
rect 43136 41880 43200 41944
rect 43216 41880 43280 41944
rect 43296 41880 43360 41944
rect 43376 41880 43440 41944
rect 43456 41880 43520 41944
rect 43536 41880 43600 41944
rect 43616 41880 43680 41944
rect 43696 41880 43760 41944
rect 43776 41880 43840 41944
rect 43856 41880 43920 41944
rect 43936 41880 44000 41944
rect 44016 41880 44080 41944
rect 44096 41880 44160 41944
rect 44176 41880 44240 41944
rect 44256 41880 44320 41944
rect 44336 41880 44400 41944
rect 44416 41880 44480 41944
rect 44496 41880 44560 41944
rect 44576 41880 44640 41944
rect 44656 41880 44720 41944
rect 44736 41880 44800 41944
rect 44816 41880 44880 41944
rect 44896 41880 44960 41944
rect 44976 41880 45040 41944
rect 45056 41880 45120 41944
rect 45136 41880 45200 41944
rect 45216 41880 45280 41944
rect 45296 41880 45360 41944
rect 8 41800 72 41864
rect 88 41800 152 41864
rect 168 41800 232 41864
rect 248 41800 312 41864
rect 328 41800 392 41864
rect 408 41800 472 41864
rect 488 41800 552 41864
rect 568 41800 632 41864
rect 648 41800 712 41864
rect 728 41800 792 41864
rect 808 41800 872 41864
rect 888 41800 952 41864
rect 968 41800 1032 41864
rect 1048 41800 1112 41864
rect 1128 41800 1192 41864
rect 1208 41800 1272 41864
rect 1288 41800 1352 41864
rect 1368 41800 1432 41864
rect 1448 41800 1512 41864
rect 1528 41800 1592 41864
rect 1608 41800 1672 41864
rect 1688 41800 1752 41864
rect 1768 41800 1832 41864
rect 1848 41800 1912 41864
rect 1928 41800 1992 41864
rect 2008 41800 2072 41864
rect 2088 41800 2152 41864
rect 2168 41800 2232 41864
rect 2248 41800 2312 41864
rect 2328 41800 2392 41864
rect 2408 41800 2472 41864
rect 2488 41800 2552 41864
rect 2568 41800 2632 41864
rect 2648 41800 2712 41864
rect 2728 41800 2792 41864
rect 2808 41800 2872 41864
rect 2888 41800 2952 41864
rect 2968 41800 3032 41864
rect 3048 41800 3112 41864
rect 3128 41800 3192 41864
rect 3208 41800 3272 41864
rect 3288 41800 3352 41864
rect 3368 41800 3432 41864
rect 3448 41800 3512 41864
rect 3528 41800 3592 41864
rect 3608 41800 3672 41864
rect 3688 41800 3752 41864
rect 3768 41800 3832 41864
rect 3848 41800 3912 41864
rect 3928 41800 3992 41864
rect 19112 41800 19176 41864
rect 19192 41800 19256 41864
rect 19272 41800 19336 41864
rect 19352 41800 19416 41864
rect 29112 41800 29176 41864
rect 29192 41800 29256 41864
rect 29272 41800 29336 41864
rect 29352 41800 29416 41864
rect 41376 41800 41440 41864
rect 41456 41800 41520 41864
rect 41536 41800 41600 41864
rect 41616 41800 41680 41864
rect 41696 41800 41760 41864
rect 41776 41800 41840 41864
rect 41856 41800 41920 41864
rect 41936 41800 42000 41864
rect 42016 41800 42080 41864
rect 42096 41800 42160 41864
rect 42176 41800 42240 41864
rect 42256 41800 42320 41864
rect 42336 41800 42400 41864
rect 42416 41800 42480 41864
rect 42496 41800 42560 41864
rect 42576 41800 42640 41864
rect 42656 41800 42720 41864
rect 42736 41800 42800 41864
rect 42816 41800 42880 41864
rect 42896 41800 42960 41864
rect 42976 41800 43040 41864
rect 43056 41800 43120 41864
rect 43136 41800 43200 41864
rect 43216 41800 43280 41864
rect 43296 41800 43360 41864
rect 43376 41800 43440 41864
rect 43456 41800 43520 41864
rect 43536 41800 43600 41864
rect 43616 41800 43680 41864
rect 43696 41800 43760 41864
rect 43776 41800 43840 41864
rect 43856 41800 43920 41864
rect 43936 41800 44000 41864
rect 44016 41800 44080 41864
rect 44096 41800 44160 41864
rect 44176 41800 44240 41864
rect 44256 41800 44320 41864
rect 44336 41800 44400 41864
rect 44416 41800 44480 41864
rect 44496 41800 44560 41864
rect 44576 41800 44640 41864
rect 44656 41800 44720 41864
rect 44736 41800 44800 41864
rect 44816 41800 44880 41864
rect 44896 41800 44960 41864
rect 44976 41800 45040 41864
rect 45056 41800 45120 41864
rect 45136 41800 45200 41864
rect 45216 41800 45280 41864
rect 45296 41800 45360 41864
rect 8 41720 72 41784
rect 88 41720 152 41784
rect 168 41720 232 41784
rect 248 41720 312 41784
rect 328 41720 392 41784
rect 408 41720 472 41784
rect 488 41720 552 41784
rect 568 41720 632 41784
rect 648 41720 712 41784
rect 728 41720 792 41784
rect 808 41720 872 41784
rect 888 41720 952 41784
rect 968 41720 1032 41784
rect 1048 41720 1112 41784
rect 1128 41720 1192 41784
rect 1208 41720 1272 41784
rect 1288 41720 1352 41784
rect 1368 41720 1432 41784
rect 1448 41720 1512 41784
rect 1528 41720 1592 41784
rect 1608 41720 1672 41784
rect 1688 41720 1752 41784
rect 1768 41720 1832 41784
rect 1848 41720 1912 41784
rect 1928 41720 1992 41784
rect 2008 41720 2072 41784
rect 2088 41720 2152 41784
rect 2168 41720 2232 41784
rect 2248 41720 2312 41784
rect 2328 41720 2392 41784
rect 2408 41720 2472 41784
rect 2488 41720 2552 41784
rect 2568 41720 2632 41784
rect 2648 41720 2712 41784
rect 2728 41720 2792 41784
rect 2808 41720 2872 41784
rect 2888 41720 2952 41784
rect 2968 41720 3032 41784
rect 3048 41720 3112 41784
rect 3128 41720 3192 41784
rect 3208 41720 3272 41784
rect 3288 41720 3352 41784
rect 3368 41720 3432 41784
rect 3448 41720 3512 41784
rect 3528 41720 3592 41784
rect 3608 41720 3672 41784
rect 3688 41720 3752 41784
rect 3768 41720 3832 41784
rect 3848 41720 3912 41784
rect 3928 41720 3992 41784
rect 19112 41720 19176 41784
rect 19192 41720 19256 41784
rect 19272 41720 19336 41784
rect 19352 41720 19416 41784
rect 29112 41720 29176 41784
rect 29192 41720 29256 41784
rect 29272 41720 29336 41784
rect 29352 41720 29416 41784
rect 41376 41720 41440 41784
rect 41456 41720 41520 41784
rect 41536 41720 41600 41784
rect 41616 41720 41680 41784
rect 41696 41720 41760 41784
rect 41776 41720 41840 41784
rect 41856 41720 41920 41784
rect 41936 41720 42000 41784
rect 42016 41720 42080 41784
rect 42096 41720 42160 41784
rect 42176 41720 42240 41784
rect 42256 41720 42320 41784
rect 42336 41720 42400 41784
rect 42416 41720 42480 41784
rect 42496 41720 42560 41784
rect 42576 41720 42640 41784
rect 42656 41720 42720 41784
rect 42736 41720 42800 41784
rect 42816 41720 42880 41784
rect 42896 41720 42960 41784
rect 42976 41720 43040 41784
rect 43056 41720 43120 41784
rect 43136 41720 43200 41784
rect 43216 41720 43280 41784
rect 43296 41720 43360 41784
rect 43376 41720 43440 41784
rect 43456 41720 43520 41784
rect 43536 41720 43600 41784
rect 43616 41720 43680 41784
rect 43696 41720 43760 41784
rect 43776 41720 43840 41784
rect 43856 41720 43920 41784
rect 43936 41720 44000 41784
rect 44016 41720 44080 41784
rect 44096 41720 44160 41784
rect 44176 41720 44240 41784
rect 44256 41720 44320 41784
rect 44336 41720 44400 41784
rect 44416 41720 44480 41784
rect 44496 41720 44560 41784
rect 44576 41720 44640 41784
rect 44656 41720 44720 41784
rect 44736 41720 44800 41784
rect 44816 41720 44880 41784
rect 44896 41720 44960 41784
rect 44976 41720 45040 41784
rect 45056 41720 45120 41784
rect 45136 41720 45200 41784
rect 45216 41720 45280 41784
rect 45296 41720 45360 41784
rect 8 41640 72 41704
rect 88 41640 152 41704
rect 168 41640 232 41704
rect 248 41640 312 41704
rect 328 41640 392 41704
rect 408 41640 472 41704
rect 488 41640 552 41704
rect 568 41640 632 41704
rect 648 41640 712 41704
rect 728 41640 792 41704
rect 808 41640 872 41704
rect 888 41640 952 41704
rect 968 41640 1032 41704
rect 1048 41640 1112 41704
rect 1128 41640 1192 41704
rect 1208 41640 1272 41704
rect 1288 41640 1352 41704
rect 1368 41640 1432 41704
rect 1448 41640 1512 41704
rect 1528 41640 1592 41704
rect 1608 41640 1672 41704
rect 1688 41640 1752 41704
rect 1768 41640 1832 41704
rect 1848 41640 1912 41704
rect 1928 41640 1992 41704
rect 2008 41640 2072 41704
rect 2088 41640 2152 41704
rect 2168 41640 2232 41704
rect 2248 41640 2312 41704
rect 2328 41640 2392 41704
rect 2408 41640 2472 41704
rect 2488 41640 2552 41704
rect 2568 41640 2632 41704
rect 2648 41640 2712 41704
rect 2728 41640 2792 41704
rect 2808 41640 2872 41704
rect 2888 41640 2952 41704
rect 2968 41640 3032 41704
rect 3048 41640 3112 41704
rect 3128 41640 3192 41704
rect 3208 41640 3272 41704
rect 3288 41640 3352 41704
rect 3368 41640 3432 41704
rect 3448 41640 3512 41704
rect 3528 41640 3592 41704
rect 3608 41640 3672 41704
rect 3688 41640 3752 41704
rect 3768 41640 3832 41704
rect 3848 41640 3912 41704
rect 3928 41640 3992 41704
rect 19112 41640 19176 41704
rect 19192 41640 19256 41704
rect 19272 41640 19336 41704
rect 19352 41640 19416 41704
rect 29112 41640 29176 41704
rect 29192 41640 29256 41704
rect 29272 41640 29336 41704
rect 29352 41640 29416 41704
rect 41376 41640 41440 41704
rect 41456 41640 41520 41704
rect 41536 41640 41600 41704
rect 41616 41640 41680 41704
rect 41696 41640 41760 41704
rect 41776 41640 41840 41704
rect 41856 41640 41920 41704
rect 41936 41640 42000 41704
rect 42016 41640 42080 41704
rect 42096 41640 42160 41704
rect 42176 41640 42240 41704
rect 42256 41640 42320 41704
rect 42336 41640 42400 41704
rect 42416 41640 42480 41704
rect 42496 41640 42560 41704
rect 42576 41640 42640 41704
rect 42656 41640 42720 41704
rect 42736 41640 42800 41704
rect 42816 41640 42880 41704
rect 42896 41640 42960 41704
rect 42976 41640 43040 41704
rect 43056 41640 43120 41704
rect 43136 41640 43200 41704
rect 43216 41640 43280 41704
rect 43296 41640 43360 41704
rect 43376 41640 43440 41704
rect 43456 41640 43520 41704
rect 43536 41640 43600 41704
rect 43616 41640 43680 41704
rect 43696 41640 43760 41704
rect 43776 41640 43840 41704
rect 43856 41640 43920 41704
rect 43936 41640 44000 41704
rect 44016 41640 44080 41704
rect 44096 41640 44160 41704
rect 44176 41640 44240 41704
rect 44256 41640 44320 41704
rect 44336 41640 44400 41704
rect 44416 41640 44480 41704
rect 44496 41640 44560 41704
rect 44576 41640 44640 41704
rect 44656 41640 44720 41704
rect 44736 41640 44800 41704
rect 44816 41640 44880 41704
rect 44896 41640 44960 41704
rect 44976 41640 45040 41704
rect 45056 41640 45120 41704
rect 45136 41640 45200 41704
rect 45216 41640 45280 41704
rect 45296 41640 45360 41704
rect 8 41560 72 41624
rect 88 41560 152 41624
rect 168 41560 232 41624
rect 248 41560 312 41624
rect 328 41560 392 41624
rect 408 41560 472 41624
rect 488 41560 552 41624
rect 568 41560 632 41624
rect 648 41560 712 41624
rect 728 41560 792 41624
rect 808 41560 872 41624
rect 888 41560 952 41624
rect 968 41560 1032 41624
rect 1048 41560 1112 41624
rect 1128 41560 1192 41624
rect 1208 41560 1272 41624
rect 1288 41560 1352 41624
rect 1368 41560 1432 41624
rect 1448 41560 1512 41624
rect 1528 41560 1592 41624
rect 1608 41560 1672 41624
rect 1688 41560 1752 41624
rect 1768 41560 1832 41624
rect 1848 41560 1912 41624
rect 1928 41560 1992 41624
rect 2008 41560 2072 41624
rect 2088 41560 2152 41624
rect 2168 41560 2232 41624
rect 2248 41560 2312 41624
rect 2328 41560 2392 41624
rect 2408 41560 2472 41624
rect 2488 41560 2552 41624
rect 2568 41560 2632 41624
rect 2648 41560 2712 41624
rect 2728 41560 2792 41624
rect 2808 41560 2872 41624
rect 2888 41560 2952 41624
rect 2968 41560 3032 41624
rect 3048 41560 3112 41624
rect 3128 41560 3192 41624
rect 3208 41560 3272 41624
rect 3288 41560 3352 41624
rect 3368 41560 3432 41624
rect 3448 41560 3512 41624
rect 3528 41560 3592 41624
rect 3608 41560 3672 41624
rect 3688 41560 3752 41624
rect 3768 41560 3832 41624
rect 3848 41560 3912 41624
rect 3928 41560 3992 41624
rect 19112 41560 19176 41624
rect 19192 41560 19256 41624
rect 19272 41560 19336 41624
rect 19352 41560 19416 41624
rect 29112 41560 29176 41624
rect 29192 41560 29256 41624
rect 29272 41560 29336 41624
rect 29352 41560 29416 41624
rect 41376 41560 41440 41624
rect 41456 41560 41520 41624
rect 41536 41560 41600 41624
rect 41616 41560 41680 41624
rect 41696 41560 41760 41624
rect 41776 41560 41840 41624
rect 41856 41560 41920 41624
rect 41936 41560 42000 41624
rect 42016 41560 42080 41624
rect 42096 41560 42160 41624
rect 42176 41560 42240 41624
rect 42256 41560 42320 41624
rect 42336 41560 42400 41624
rect 42416 41560 42480 41624
rect 42496 41560 42560 41624
rect 42576 41560 42640 41624
rect 42656 41560 42720 41624
rect 42736 41560 42800 41624
rect 42816 41560 42880 41624
rect 42896 41560 42960 41624
rect 42976 41560 43040 41624
rect 43056 41560 43120 41624
rect 43136 41560 43200 41624
rect 43216 41560 43280 41624
rect 43296 41560 43360 41624
rect 43376 41560 43440 41624
rect 43456 41560 43520 41624
rect 43536 41560 43600 41624
rect 43616 41560 43680 41624
rect 43696 41560 43760 41624
rect 43776 41560 43840 41624
rect 43856 41560 43920 41624
rect 43936 41560 44000 41624
rect 44016 41560 44080 41624
rect 44096 41560 44160 41624
rect 44176 41560 44240 41624
rect 44256 41560 44320 41624
rect 44336 41560 44400 41624
rect 44416 41560 44480 41624
rect 44496 41560 44560 41624
rect 44576 41560 44640 41624
rect 44656 41560 44720 41624
rect 44736 41560 44800 41624
rect 44816 41560 44880 41624
rect 44896 41560 44960 41624
rect 44976 41560 45040 41624
rect 45056 41560 45120 41624
rect 45136 41560 45200 41624
rect 45216 41560 45280 41624
rect 45296 41560 45360 41624
rect 8 41480 72 41544
rect 88 41480 152 41544
rect 168 41480 232 41544
rect 248 41480 312 41544
rect 328 41480 392 41544
rect 408 41480 472 41544
rect 488 41480 552 41544
rect 568 41480 632 41544
rect 648 41480 712 41544
rect 728 41480 792 41544
rect 808 41480 872 41544
rect 888 41480 952 41544
rect 968 41480 1032 41544
rect 1048 41480 1112 41544
rect 1128 41480 1192 41544
rect 1208 41480 1272 41544
rect 1288 41480 1352 41544
rect 1368 41480 1432 41544
rect 1448 41480 1512 41544
rect 1528 41480 1592 41544
rect 1608 41480 1672 41544
rect 1688 41480 1752 41544
rect 1768 41480 1832 41544
rect 1848 41480 1912 41544
rect 1928 41480 1992 41544
rect 2008 41480 2072 41544
rect 2088 41480 2152 41544
rect 2168 41480 2232 41544
rect 2248 41480 2312 41544
rect 2328 41480 2392 41544
rect 2408 41480 2472 41544
rect 2488 41480 2552 41544
rect 2568 41480 2632 41544
rect 2648 41480 2712 41544
rect 2728 41480 2792 41544
rect 2808 41480 2872 41544
rect 2888 41480 2952 41544
rect 2968 41480 3032 41544
rect 3048 41480 3112 41544
rect 3128 41480 3192 41544
rect 3208 41480 3272 41544
rect 3288 41480 3352 41544
rect 3368 41480 3432 41544
rect 3448 41480 3512 41544
rect 3528 41480 3592 41544
rect 3608 41480 3672 41544
rect 3688 41480 3752 41544
rect 3768 41480 3832 41544
rect 3848 41480 3912 41544
rect 3928 41480 3992 41544
rect 19112 41480 19176 41544
rect 19192 41480 19256 41544
rect 19272 41480 19336 41544
rect 19352 41480 19416 41544
rect 29112 41480 29176 41544
rect 29192 41480 29256 41544
rect 29272 41480 29336 41544
rect 29352 41480 29416 41544
rect 41376 41480 41440 41544
rect 41456 41480 41520 41544
rect 41536 41480 41600 41544
rect 41616 41480 41680 41544
rect 41696 41480 41760 41544
rect 41776 41480 41840 41544
rect 41856 41480 41920 41544
rect 41936 41480 42000 41544
rect 42016 41480 42080 41544
rect 42096 41480 42160 41544
rect 42176 41480 42240 41544
rect 42256 41480 42320 41544
rect 42336 41480 42400 41544
rect 42416 41480 42480 41544
rect 42496 41480 42560 41544
rect 42576 41480 42640 41544
rect 42656 41480 42720 41544
rect 42736 41480 42800 41544
rect 42816 41480 42880 41544
rect 42896 41480 42960 41544
rect 42976 41480 43040 41544
rect 43056 41480 43120 41544
rect 43136 41480 43200 41544
rect 43216 41480 43280 41544
rect 43296 41480 43360 41544
rect 43376 41480 43440 41544
rect 43456 41480 43520 41544
rect 43536 41480 43600 41544
rect 43616 41480 43680 41544
rect 43696 41480 43760 41544
rect 43776 41480 43840 41544
rect 43856 41480 43920 41544
rect 43936 41480 44000 41544
rect 44016 41480 44080 41544
rect 44096 41480 44160 41544
rect 44176 41480 44240 41544
rect 44256 41480 44320 41544
rect 44336 41480 44400 41544
rect 44416 41480 44480 41544
rect 44496 41480 44560 41544
rect 44576 41480 44640 41544
rect 44656 41480 44720 41544
rect 44736 41480 44800 41544
rect 44816 41480 44880 41544
rect 44896 41480 44960 41544
rect 44976 41480 45040 41544
rect 45056 41480 45120 41544
rect 45136 41480 45200 41544
rect 45216 41480 45280 41544
rect 45296 41480 45360 41544
rect 8 41400 72 41464
rect 88 41400 152 41464
rect 168 41400 232 41464
rect 248 41400 312 41464
rect 328 41400 392 41464
rect 408 41400 472 41464
rect 488 41400 552 41464
rect 568 41400 632 41464
rect 648 41400 712 41464
rect 728 41400 792 41464
rect 808 41400 872 41464
rect 888 41400 952 41464
rect 968 41400 1032 41464
rect 1048 41400 1112 41464
rect 1128 41400 1192 41464
rect 1208 41400 1272 41464
rect 1288 41400 1352 41464
rect 1368 41400 1432 41464
rect 1448 41400 1512 41464
rect 1528 41400 1592 41464
rect 1608 41400 1672 41464
rect 1688 41400 1752 41464
rect 1768 41400 1832 41464
rect 1848 41400 1912 41464
rect 1928 41400 1992 41464
rect 2008 41400 2072 41464
rect 2088 41400 2152 41464
rect 2168 41400 2232 41464
rect 2248 41400 2312 41464
rect 2328 41400 2392 41464
rect 2408 41400 2472 41464
rect 2488 41400 2552 41464
rect 2568 41400 2632 41464
rect 2648 41400 2712 41464
rect 2728 41400 2792 41464
rect 2808 41400 2872 41464
rect 2888 41400 2952 41464
rect 2968 41400 3032 41464
rect 3048 41400 3112 41464
rect 3128 41400 3192 41464
rect 3208 41400 3272 41464
rect 3288 41400 3352 41464
rect 3368 41400 3432 41464
rect 3448 41400 3512 41464
rect 3528 41400 3592 41464
rect 3608 41400 3672 41464
rect 3688 41400 3752 41464
rect 3768 41400 3832 41464
rect 3848 41400 3912 41464
rect 3928 41400 3992 41464
rect 19112 41400 19176 41464
rect 19192 41400 19256 41464
rect 19272 41400 19336 41464
rect 19352 41400 19416 41464
rect 29112 41400 29176 41464
rect 29192 41400 29256 41464
rect 29272 41400 29336 41464
rect 29352 41400 29416 41464
rect 41376 41400 41440 41464
rect 41456 41400 41520 41464
rect 41536 41400 41600 41464
rect 41616 41400 41680 41464
rect 41696 41400 41760 41464
rect 41776 41400 41840 41464
rect 41856 41400 41920 41464
rect 41936 41400 42000 41464
rect 42016 41400 42080 41464
rect 42096 41400 42160 41464
rect 42176 41400 42240 41464
rect 42256 41400 42320 41464
rect 42336 41400 42400 41464
rect 42416 41400 42480 41464
rect 42496 41400 42560 41464
rect 42576 41400 42640 41464
rect 42656 41400 42720 41464
rect 42736 41400 42800 41464
rect 42816 41400 42880 41464
rect 42896 41400 42960 41464
rect 42976 41400 43040 41464
rect 43056 41400 43120 41464
rect 43136 41400 43200 41464
rect 43216 41400 43280 41464
rect 43296 41400 43360 41464
rect 43376 41400 43440 41464
rect 43456 41400 43520 41464
rect 43536 41400 43600 41464
rect 43616 41400 43680 41464
rect 43696 41400 43760 41464
rect 43776 41400 43840 41464
rect 43856 41400 43920 41464
rect 43936 41400 44000 41464
rect 44016 41400 44080 41464
rect 44096 41400 44160 41464
rect 44176 41400 44240 41464
rect 44256 41400 44320 41464
rect 44336 41400 44400 41464
rect 44416 41400 44480 41464
rect 44496 41400 44560 41464
rect 44576 41400 44640 41464
rect 44656 41400 44720 41464
rect 44736 41400 44800 41464
rect 44816 41400 44880 41464
rect 44896 41400 44960 41464
rect 44976 41400 45040 41464
rect 45056 41400 45120 41464
rect 45136 41400 45200 41464
rect 45216 41400 45280 41464
rect 45296 41400 45360 41464
rect 5008 40320 5072 40384
rect 5088 40320 5152 40384
rect 5168 40320 5232 40384
rect 5248 40320 5312 40384
rect 5328 40320 5392 40384
rect 5408 40320 5472 40384
rect 5488 40320 5552 40384
rect 5568 40320 5632 40384
rect 5648 40320 5712 40384
rect 5728 40320 5792 40384
rect 5808 40320 5872 40384
rect 5888 40320 5952 40384
rect 5968 40320 6032 40384
rect 6048 40320 6112 40384
rect 6128 40320 6192 40384
rect 6208 40320 6272 40384
rect 6288 40320 6352 40384
rect 6368 40320 6432 40384
rect 6448 40320 6512 40384
rect 6528 40320 6592 40384
rect 6608 40320 6672 40384
rect 6688 40320 6752 40384
rect 6768 40320 6832 40384
rect 6848 40320 6912 40384
rect 6928 40320 6992 40384
rect 7008 40320 7072 40384
rect 7088 40320 7152 40384
rect 7168 40320 7232 40384
rect 7248 40320 7312 40384
rect 7328 40320 7392 40384
rect 7408 40320 7472 40384
rect 7488 40320 7552 40384
rect 7568 40320 7632 40384
rect 7648 40320 7712 40384
rect 7728 40320 7792 40384
rect 7808 40320 7872 40384
rect 7888 40320 7952 40384
rect 7968 40320 8032 40384
rect 8048 40320 8112 40384
rect 8128 40320 8192 40384
rect 8208 40320 8272 40384
rect 8288 40320 8352 40384
rect 8368 40320 8432 40384
rect 8448 40320 8512 40384
rect 8528 40320 8592 40384
rect 8608 40320 8672 40384
rect 8688 40320 8752 40384
rect 8768 40320 8832 40384
rect 8848 40320 8912 40384
rect 8928 40320 8992 40384
rect 14112 40320 14176 40384
rect 14192 40320 14256 40384
rect 14272 40320 14336 40384
rect 14352 40320 14416 40384
rect 24112 40320 24176 40384
rect 24192 40320 24256 40384
rect 24272 40320 24336 40384
rect 24352 40320 24416 40384
rect 36376 40320 36440 40384
rect 36456 40320 36520 40384
rect 36536 40320 36600 40384
rect 36616 40320 36680 40384
rect 36696 40320 36760 40384
rect 36776 40320 36840 40384
rect 36856 40320 36920 40384
rect 36936 40320 37000 40384
rect 37016 40320 37080 40384
rect 37096 40320 37160 40384
rect 37176 40320 37240 40384
rect 37256 40320 37320 40384
rect 37336 40320 37400 40384
rect 37416 40320 37480 40384
rect 37496 40320 37560 40384
rect 37576 40320 37640 40384
rect 37656 40320 37720 40384
rect 37736 40320 37800 40384
rect 37816 40320 37880 40384
rect 37896 40320 37960 40384
rect 37976 40320 38040 40384
rect 38056 40320 38120 40384
rect 38136 40320 38200 40384
rect 38216 40320 38280 40384
rect 38296 40320 38360 40384
rect 38376 40320 38440 40384
rect 38456 40320 38520 40384
rect 38536 40320 38600 40384
rect 38616 40320 38680 40384
rect 38696 40320 38760 40384
rect 38776 40320 38840 40384
rect 38856 40320 38920 40384
rect 38936 40320 39000 40384
rect 39016 40320 39080 40384
rect 39096 40320 39160 40384
rect 39176 40320 39240 40384
rect 39256 40320 39320 40384
rect 39336 40320 39400 40384
rect 39416 40320 39480 40384
rect 39496 40320 39560 40384
rect 39576 40320 39640 40384
rect 39656 40320 39720 40384
rect 39736 40320 39800 40384
rect 39816 40320 39880 40384
rect 39896 40320 39960 40384
rect 39976 40320 40040 40384
rect 40056 40320 40120 40384
rect 40136 40320 40200 40384
rect 40216 40320 40280 40384
rect 40296 40320 40360 40384
rect 5008 40240 5072 40304
rect 5088 40240 5152 40304
rect 5168 40240 5232 40304
rect 5248 40240 5312 40304
rect 5328 40240 5392 40304
rect 5408 40240 5472 40304
rect 5488 40240 5552 40304
rect 5568 40240 5632 40304
rect 5648 40240 5712 40304
rect 5728 40240 5792 40304
rect 5808 40240 5872 40304
rect 5888 40240 5952 40304
rect 5968 40240 6032 40304
rect 6048 40240 6112 40304
rect 6128 40240 6192 40304
rect 6208 40240 6272 40304
rect 6288 40240 6352 40304
rect 6368 40240 6432 40304
rect 6448 40240 6512 40304
rect 6528 40240 6592 40304
rect 6608 40240 6672 40304
rect 6688 40240 6752 40304
rect 6768 40240 6832 40304
rect 6848 40240 6912 40304
rect 6928 40240 6992 40304
rect 7008 40240 7072 40304
rect 7088 40240 7152 40304
rect 7168 40240 7232 40304
rect 7248 40240 7312 40304
rect 7328 40240 7392 40304
rect 7408 40240 7472 40304
rect 7488 40240 7552 40304
rect 7568 40240 7632 40304
rect 7648 40240 7712 40304
rect 7728 40240 7792 40304
rect 7808 40240 7872 40304
rect 7888 40240 7952 40304
rect 7968 40240 8032 40304
rect 8048 40240 8112 40304
rect 8128 40240 8192 40304
rect 8208 40240 8272 40304
rect 8288 40240 8352 40304
rect 8368 40240 8432 40304
rect 8448 40240 8512 40304
rect 8528 40240 8592 40304
rect 8608 40240 8672 40304
rect 8688 40240 8752 40304
rect 8768 40240 8832 40304
rect 8848 40240 8912 40304
rect 8928 40240 8992 40304
rect 14112 40240 14176 40304
rect 14192 40240 14256 40304
rect 14272 40240 14336 40304
rect 14352 40240 14416 40304
rect 24112 40240 24176 40304
rect 24192 40240 24256 40304
rect 24272 40240 24336 40304
rect 24352 40240 24416 40304
rect 36376 40240 36440 40304
rect 36456 40240 36520 40304
rect 36536 40240 36600 40304
rect 36616 40240 36680 40304
rect 36696 40240 36760 40304
rect 36776 40240 36840 40304
rect 36856 40240 36920 40304
rect 36936 40240 37000 40304
rect 37016 40240 37080 40304
rect 37096 40240 37160 40304
rect 37176 40240 37240 40304
rect 37256 40240 37320 40304
rect 37336 40240 37400 40304
rect 37416 40240 37480 40304
rect 37496 40240 37560 40304
rect 37576 40240 37640 40304
rect 37656 40240 37720 40304
rect 37736 40240 37800 40304
rect 37816 40240 37880 40304
rect 37896 40240 37960 40304
rect 37976 40240 38040 40304
rect 38056 40240 38120 40304
rect 38136 40240 38200 40304
rect 38216 40240 38280 40304
rect 38296 40240 38360 40304
rect 38376 40240 38440 40304
rect 38456 40240 38520 40304
rect 38536 40240 38600 40304
rect 38616 40240 38680 40304
rect 38696 40240 38760 40304
rect 38776 40240 38840 40304
rect 38856 40240 38920 40304
rect 38936 40240 39000 40304
rect 39016 40240 39080 40304
rect 39096 40240 39160 40304
rect 39176 40240 39240 40304
rect 39256 40240 39320 40304
rect 39336 40240 39400 40304
rect 39416 40240 39480 40304
rect 39496 40240 39560 40304
rect 39576 40240 39640 40304
rect 39656 40240 39720 40304
rect 39736 40240 39800 40304
rect 39816 40240 39880 40304
rect 39896 40240 39960 40304
rect 39976 40240 40040 40304
rect 40056 40240 40120 40304
rect 40136 40240 40200 40304
rect 40216 40240 40280 40304
rect 40296 40240 40360 40304
rect 5008 40160 5072 40224
rect 5088 40160 5152 40224
rect 5168 40160 5232 40224
rect 5248 40160 5312 40224
rect 5328 40160 5392 40224
rect 5408 40160 5472 40224
rect 5488 40160 5552 40224
rect 5568 40160 5632 40224
rect 5648 40160 5712 40224
rect 5728 40160 5792 40224
rect 5808 40160 5872 40224
rect 5888 40160 5952 40224
rect 5968 40160 6032 40224
rect 6048 40160 6112 40224
rect 6128 40160 6192 40224
rect 6208 40160 6272 40224
rect 6288 40160 6352 40224
rect 6368 40160 6432 40224
rect 6448 40160 6512 40224
rect 6528 40160 6592 40224
rect 6608 40160 6672 40224
rect 6688 40160 6752 40224
rect 6768 40160 6832 40224
rect 6848 40160 6912 40224
rect 6928 40160 6992 40224
rect 7008 40160 7072 40224
rect 7088 40160 7152 40224
rect 7168 40160 7232 40224
rect 7248 40160 7312 40224
rect 7328 40160 7392 40224
rect 7408 40160 7472 40224
rect 7488 40160 7552 40224
rect 7568 40160 7632 40224
rect 7648 40160 7712 40224
rect 7728 40160 7792 40224
rect 7808 40160 7872 40224
rect 7888 40160 7952 40224
rect 7968 40160 8032 40224
rect 8048 40160 8112 40224
rect 8128 40160 8192 40224
rect 8208 40160 8272 40224
rect 8288 40160 8352 40224
rect 8368 40160 8432 40224
rect 8448 40160 8512 40224
rect 8528 40160 8592 40224
rect 8608 40160 8672 40224
rect 8688 40160 8752 40224
rect 8768 40160 8832 40224
rect 8848 40160 8912 40224
rect 8928 40160 8992 40224
rect 14112 40160 14176 40224
rect 14192 40160 14256 40224
rect 14272 40160 14336 40224
rect 14352 40160 14416 40224
rect 24112 40160 24176 40224
rect 24192 40160 24256 40224
rect 24272 40160 24336 40224
rect 24352 40160 24416 40224
rect 36376 40160 36440 40224
rect 36456 40160 36520 40224
rect 36536 40160 36600 40224
rect 36616 40160 36680 40224
rect 36696 40160 36760 40224
rect 36776 40160 36840 40224
rect 36856 40160 36920 40224
rect 36936 40160 37000 40224
rect 37016 40160 37080 40224
rect 37096 40160 37160 40224
rect 37176 40160 37240 40224
rect 37256 40160 37320 40224
rect 37336 40160 37400 40224
rect 37416 40160 37480 40224
rect 37496 40160 37560 40224
rect 37576 40160 37640 40224
rect 37656 40160 37720 40224
rect 37736 40160 37800 40224
rect 37816 40160 37880 40224
rect 37896 40160 37960 40224
rect 37976 40160 38040 40224
rect 38056 40160 38120 40224
rect 38136 40160 38200 40224
rect 38216 40160 38280 40224
rect 38296 40160 38360 40224
rect 38376 40160 38440 40224
rect 38456 40160 38520 40224
rect 38536 40160 38600 40224
rect 38616 40160 38680 40224
rect 38696 40160 38760 40224
rect 38776 40160 38840 40224
rect 38856 40160 38920 40224
rect 38936 40160 39000 40224
rect 39016 40160 39080 40224
rect 39096 40160 39160 40224
rect 39176 40160 39240 40224
rect 39256 40160 39320 40224
rect 39336 40160 39400 40224
rect 39416 40160 39480 40224
rect 39496 40160 39560 40224
rect 39576 40160 39640 40224
rect 39656 40160 39720 40224
rect 39736 40160 39800 40224
rect 39816 40160 39880 40224
rect 39896 40160 39960 40224
rect 39976 40160 40040 40224
rect 40056 40160 40120 40224
rect 40136 40160 40200 40224
rect 40216 40160 40280 40224
rect 40296 40160 40360 40224
rect 5008 40080 5072 40144
rect 5088 40080 5152 40144
rect 5168 40080 5232 40144
rect 5248 40080 5312 40144
rect 5328 40080 5392 40144
rect 5408 40080 5472 40144
rect 5488 40080 5552 40144
rect 5568 40080 5632 40144
rect 5648 40080 5712 40144
rect 5728 40080 5792 40144
rect 5808 40080 5872 40144
rect 5888 40080 5952 40144
rect 5968 40080 6032 40144
rect 6048 40080 6112 40144
rect 6128 40080 6192 40144
rect 6208 40080 6272 40144
rect 6288 40080 6352 40144
rect 6368 40080 6432 40144
rect 6448 40080 6512 40144
rect 6528 40080 6592 40144
rect 6608 40080 6672 40144
rect 6688 40080 6752 40144
rect 6768 40080 6832 40144
rect 6848 40080 6912 40144
rect 6928 40080 6992 40144
rect 7008 40080 7072 40144
rect 7088 40080 7152 40144
rect 7168 40080 7232 40144
rect 7248 40080 7312 40144
rect 7328 40080 7392 40144
rect 7408 40080 7472 40144
rect 7488 40080 7552 40144
rect 7568 40080 7632 40144
rect 7648 40080 7712 40144
rect 7728 40080 7792 40144
rect 7808 40080 7872 40144
rect 7888 40080 7952 40144
rect 7968 40080 8032 40144
rect 8048 40080 8112 40144
rect 8128 40080 8192 40144
rect 8208 40080 8272 40144
rect 8288 40080 8352 40144
rect 8368 40080 8432 40144
rect 8448 40080 8512 40144
rect 8528 40080 8592 40144
rect 8608 40080 8672 40144
rect 8688 40080 8752 40144
rect 8768 40080 8832 40144
rect 8848 40080 8912 40144
rect 8928 40080 8992 40144
rect 14112 40080 14176 40144
rect 14192 40080 14256 40144
rect 14272 40080 14336 40144
rect 14352 40080 14416 40144
rect 24112 40080 24176 40144
rect 24192 40080 24256 40144
rect 24272 40080 24336 40144
rect 24352 40080 24416 40144
rect 36376 40080 36440 40144
rect 36456 40080 36520 40144
rect 36536 40080 36600 40144
rect 36616 40080 36680 40144
rect 36696 40080 36760 40144
rect 36776 40080 36840 40144
rect 36856 40080 36920 40144
rect 36936 40080 37000 40144
rect 37016 40080 37080 40144
rect 37096 40080 37160 40144
rect 37176 40080 37240 40144
rect 37256 40080 37320 40144
rect 37336 40080 37400 40144
rect 37416 40080 37480 40144
rect 37496 40080 37560 40144
rect 37576 40080 37640 40144
rect 37656 40080 37720 40144
rect 37736 40080 37800 40144
rect 37816 40080 37880 40144
rect 37896 40080 37960 40144
rect 37976 40080 38040 40144
rect 38056 40080 38120 40144
rect 38136 40080 38200 40144
rect 38216 40080 38280 40144
rect 38296 40080 38360 40144
rect 38376 40080 38440 40144
rect 38456 40080 38520 40144
rect 38536 40080 38600 40144
rect 38616 40080 38680 40144
rect 38696 40080 38760 40144
rect 38776 40080 38840 40144
rect 38856 40080 38920 40144
rect 38936 40080 39000 40144
rect 39016 40080 39080 40144
rect 39096 40080 39160 40144
rect 39176 40080 39240 40144
rect 39256 40080 39320 40144
rect 39336 40080 39400 40144
rect 39416 40080 39480 40144
rect 39496 40080 39560 40144
rect 39576 40080 39640 40144
rect 39656 40080 39720 40144
rect 39736 40080 39800 40144
rect 39816 40080 39880 40144
rect 39896 40080 39960 40144
rect 39976 40080 40040 40144
rect 40056 40080 40120 40144
rect 40136 40080 40200 40144
rect 40216 40080 40280 40144
rect 40296 40080 40360 40144
rect 5008 40000 5072 40064
rect 5088 40000 5152 40064
rect 5168 40000 5232 40064
rect 5248 40000 5312 40064
rect 5328 40000 5392 40064
rect 5408 40000 5472 40064
rect 5488 40000 5552 40064
rect 5568 40000 5632 40064
rect 5648 40000 5712 40064
rect 5728 40000 5792 40064
rect 5808 40000 5872 40064
rect 5888 40000 5952 40064
rect 5968 40000 6032 40064
rect 6048 40000 6112 40064
rect 6128 40000 6192 40064
rect 6208 40000 6272 40064
rect 6288 40000 6352 40064
rect 6368 40000 6432 40064
rect 6448 40000 6512 40064
rect 6528 40000 6592 40064
rect 6608 40000 6672 40064
rect 6688 40000 6752 40064
rect 6768 40000 6832 40064
rect 6848 40000 6912 40064
rect 6928 40000 6992 40064
rect 7008 40000 7072 40064
rect 7088 40000 7152 40064
rect 7168 40000 7232 40064
rect 7248 40000 7312 40064
rect 7328 40000 7392 40064
rect 7408 40000 7472 40064
rect 7488 40000 7552 40064
rect 7568 40000 7632 40064
rect 7648 40000 7712 40064
rect 7728 40000 7792 40064
rect 7808 40000 7872 40064
rect 7888 40000 7952 40064
rect 7968 40000 8032 40064
rect 8048 40000 8112 40064
rect 8128 40000 8192 40064
rect 8208 40000 8272 40064
rect 8288 40000 8352 40064
rect 8368 40000 8432 40064
rect 8448 40000 8512 40064
rect 8528 40000 8592 40064
rect 8608 40000 8672 40064
rect 8688 40000 8752 40064
rect 8768 40000 8832 40064
rect 8848 40000 8912 40064
rect 8928 40000 8992 40064
rect 14112 40000 14176 40064
rect 14192 40000 14256 40064
rect 14272 40000 14336 40064
rect 14352 40000 14416 40064
rect 24112 40000 24176 40064
rect 24192 40000 24256 40064
rect 24272 40000 24336 40064
rect 24352 40000 24416 40064
rect 36376 40000 36440 40064
rect 36456 40000 36520 40064
rect 36536 40000 36600 40064
rect 36616 40000 36680 40064
rect 36696 40000 36760 40064
rect 36776 40000 36840 40064
rect 36856 40000 36920 40064
rect 36936 40000 37000 40064
rect 37016 40000 37080 40064
rect 37096 40000 37160 40064
rect 37176 40000 37240 40064
rect 37256 40000 37320 40064
rect 37336 40000 37400 40064
rect 37416 40000 37480 40064
rect 37496 40000 37560 40064
rect 37576 40000 37640 40064
rect 37656 40000 37720 40064
rect 37736 40000 37800 40064
rect 37816 40000 37880 40064
rect 37896 40000 37960 40064
rect 37976 40000 38040 40064
rect 38056 40000 38120 40064
rect 38136 40000 38200 40064
rect 38216 40000 38280 40064
rect 38296 40000 38360 40064
rect 38376 40000 38440 40064
rect 38456 40000 38520 40064
rect 38536 40000 38600 40064
rect 38616 40000 38680 40064
rect 38696 40000 38760 40064
rect 38776 40000 38840 40064
rect 38856 40000 38920 40064
rect 38936 40000 39000 40064
rect 39016 40000 39080 40064
rect 39096 40000 39160 40064
rect 39176 40000 39240 40064
rect 39256 40000 39320 40064
rect 39336 40000 39400 40064
rect 39416 40000 39480 40064
rect 39496 40000 39560 40064
rect 39576 40000 39640 40064
rect 39656 40000 39720 40064
rect 39736 40000 39800 40064
rect 39816 40000 39880 40064
rect 39896 40000 39960 40064
rect 39976 40000 40040 40064
rect 40056 40000 40120 40064
rect 40136 40000 40200 40064
rect 40216 40000 40280 40064
rect 40296 40000 40360 40064
rect 5008 39920 5072 39984
rect 5088 39920 5152 39984
rect 5168 39920 5232 39984
rect 5248 39920 5312 39984
rect 5328 39920 5392 39984
rect 5408 39920 5472 39984
rect 5488 39920 5552 39984
rect 5568 39920 5632 39984
rect 5648 39920 5712 39984
rect 5728 39920 5792 39984
rect 5808 39920 5872 39984
rect 5888 39920 5952 39984
rect 5968 39920 6032 39984
rect 6048 39920 6112 39984
rect 6128 39920 6192 39984
rect 6208 39920 6272 39984
rect 6288 39920 6352 39984
rect 6368 39920 6432 39984
rect 6448 39920 6512 39984
rect 6528 39920 6592 39984
rect 6608 39920 6672 39984
rect 6688 39920 6752 39984
rect 6768 39920 6832 39984
rect 6848 39920 6912 39984
rect 6928 39920 6992 39984
rect 7008 39920 7072 39984
rect 7088 39920 7152 39984
rect 7168 39920 7232 39984
rect 7248 39920 7312 39984
rect 7328 39920 7392 39984
rect 7408 39920 7472 39984
rect 7488 39920 7552 39984
rect 7568 39920 7632 39984
rect 7648 39920 7712 39984
rect 7728 39920 7792 39984
rect 7808 39920 7872 39984
rect 7888 39920 7952 39984
rect 7968 39920 8032 39984
rect 8048 39920 8112 39984
rect 8128 39920 8192 39984
rect 8208 39920 8272 39984
rect 8288 39920 8352 39984
rect 8368 39920 8432 39984
rect 8448 39920 8512 39984
rect 8528 39920 8592 39984
rect 8608 39920 8672 39984
rect 8688 39920 8752 39984
rect 8768 39920 8832 39984
rect 8848 39920 8912 39984
rect 8928 39920 8992 39984
rect 14112 39920 14176 39984
rect 14192 39920 14256 39984
rect 14272 39920 14336 39984
rect 14352 39920 14416 39984
rect 24112 39920 24176 39984
rect 24192 39920 24256 39984
rect 24272 39920 24336 39984
rect 24352 39920 24416 39984
rect 36376 39920 36440 39984
rect 36456 39920 36520 39984
rect 36536 39920 36600 39984
rect 36616 39920 36680 39984
rect 36696 39920 36760 39984
rect 36776 39920 36840 39984
rect 36856 39920 36920 39984
rect 36936 39920 37000 39984
rect 37016 39920 37080 39984
rect 37096 39920 37160 39984
rect 37176 39920 37240 39984
rect 37256 39920 37320 39984
rect 37336 39920 37400 39984
rect 37416 39920 37480 39984
rect 37496 39920 37560 39984
rect 37576 39920 37640 39984
rect 37656 39920 37720 39984
rect 37736 39920 37800 39984
rect 37816 39920 37880 39984
rect 37896 39920 37960 39984
rect 37976 39920 38040 39984
rect 38056 39920 38120 39984
rect 38136 39920 38200 39984
rect 38216 39920 38280 39984
rect 38296 39920 38360 39984
rect 38376 39920 38440 39984
rect 38456 39920 38520 39984
rect 38536 39920 38600 39984
rect 38616 39920 38680 39984
rect 38696 39920 38760 39984
rect 38776 39920 38840 39984
rect 38856 39920 38920 39984
rect 38936 39920 39000 39984
rect 39016 39920 39080 39984
rect 39096 39920 39160 39984
rect 39176 39920 39240 39984
rect 39256 39920 39320 39984
rect 39336 39920 39400 39984
rect 39416 39920 39480 39984
rect 39496 39920 39560 39984
rect 39576 39920 39640 39984
rect 39656 39920 39720 39984
rect 39736 39920 39800 39984
rect 39816 39920 39880 39984
rect 39896 39920 39960 39984
rect 39976 39920 40040 39984
rect 40056 39920 40120 39984
rect 40136 39920 40200 39984
rect 40216 39920 40280 39984
rect 40296 39920 40360 39984
rect 5008 39840 5072 39904
rect 5088 39840 5152 39904
rect 5168 39840 5232 39904
rect 5248 39840 5312 39904
rect 5328 39840 5392 39904
rect 5408 39840 5472 39904
rect 5488 39840 5552 39904
rect 5568 39840 5632 39904
rect 5648 39840 5712 39904
rect 5728 39840 5792 39904
rect 5808 39840 5872 39904
rect 5888 39840 5952 39904
rect 5968 39840 6032 39904
rect 6048 39840 6112 39904
rect 6128 39840 6192 39904
rect 6208 39840 6272 39904
rect 6288 39840 6352 39904
rect 6368 39840 6432 39904
rect 6448 39840 6512 39904
rect 6528 39840 6592 39904
rect 6608 39840 6672 39904
rect 6688 39840 6752 39904
rect 6768 39840 6832 39904
rect 6848 39840 6912 39904
rect 6928 39840 6992 39904
rect 7008 39840 7072 39904
rect 7088 39840 7152 39904
rect 7168 39840 7232 39904
rect 7248 39840 7312 39904
rect 7328 39840 7392 39904
rect 7408 39840 7472 39904
rect 7488 39840 7552 39904
rect 7568 39840 7632 39904
rect 7648 39840 7712 39904
rect 7728 39840 7792 39904
rect 7808 39840 7872 39904
rect 7888 39840 7952 39904
rect 7968 39840 8032 39904
rect 8048 39840 8112 39904
rect 8128 39840 8192 39904
rect 8208 39840 8272 39904
rect 8288 39840 8352 39904
rect 8368 39840 8432 39904
rect 8448 39840 8512 39904
rect 8528 39840 8592 39904
rect 8608 39840 8672 39904
rect 8688 39840 8752 39904
rect 8768 39840 8832 39904
rect 8848 39840 8912 39904
rect 8928 39840 8992 39904
rect 14112 39840 14176 39904
rect 14192 39840 14256 39904
rect 14272 39840 14336 39904
rect 14352 39840 14416 39904
rect 24112 39840 24176 39904
rect 24192 39840 24256 39904
rect 24272 39840 24336 39904
rect 24352 39840 24416 39904
rect 36376 39840 36440 39904
rect 36456 39840 36520 39904
rect 36536 39840 36600 39904
rect 36616 39840 36680 39904
rect 36696 39840 36760 39904
rect 36776 39840 36840 39904
rect 36856 39840 36920 39904
rect 36936 39840 37000 39904
rect 37016 39840 37080 39904
rect 37096 39840 37160 39904
rect 37176 39840 37240 39904
rect 37256 39840 37320 39904
rect 37336 39840 37400 39904
rect 37416 39840 37480 39904
rect 37496 39840 37560 39904
rect 37576 39840 37640 39904
rect 37656 39840 37720 39904
rect 37736 39840 37800 39904
rect 37816 39840 37880 39904
rect 37896 39840 37960 39904
rect 37976 39840 38040 39904
rect 38056 39840 38120 39904
rect 38136 39840 38200 39904
rect 38216 39840 38280 39904
rect 38296 39840 38360 39904
rect 38376 39840 38440 39904
rect 38456 39840 38520 39904
rect 38536 39840 38600 39904
rect 38616 39840 38680 39904
rect 38696 39840 38760 39904
rect 38776 39840 38840 39904
rect 38856 39840 38920 39904
rect 38936 39840 39000 39904
rect 39016 39840 39080 39904
rect 39096 39840 39160 39904
rect 39176 39840 39240 39904
rect 39256 39840 39320 39904
rect 39336 39840 39400 39904
rect 39416 39840 39480 39904
rect 39496 39840 39560 39904
rect 39576 39840 39640 39904
rect 39656 39840 39720 39904
rect 39736 39840 39800 39904
rect 39816 39840 39880 39904
rect 39896 39840 39960 39904
rect 39976 39840 40040 39904
rect 40056 39840 40120 39904
rect 40136 39840 40200 39904
rect 40216 39840 40280 39904
rect 40296 39840 40360 39904
rect 5008 39760 5072 39824
rect 5088 39760 5152 39824
rect 5168 39760 5232 39824
rect 5248 39760 5312 39824
rect 5328 39760 5392 39824
rect 5408 39760 5472 39824
rect 5488 39760 5552 39824
rect 5568 39760 5632 39824
rect 5648 39760 5712 39824
rect 5728 39760 5792 39824
rect 5808 39760 5872 39824
rect 5888 39760 5952 39824
rect 5968 39760 6032 39824
rect 6048 39760 6112 39824
rect 6128 39760 6192 39824
rect 6208 39760 6272 39824
rect 6288 39760 6352 39824
rect 6368 39760 6432 39824
rect 6448 39760 6512 39824
rect 6528 39760 6592 39824
rect 6608 39760 6672 39824
rect 6688 39760 6752 39824
rect 6768 39760 6832 39824
rect 6848 39760 6912 39824
rect 6928 39760 6992 39824
rect 7008 39760 7072 39824
rect 7088 39760 7152 39824
rect 7168 39760 7232 39824
rect 7248 39760 7312 39824
rect 7328 39760 7392 39824
rect 7408 39760 7472 39824
rect 7488 39760 7552 39824
rect 7568 39760 7632 39824
rect 7648 39760 7712 39824
rect 7728 39760 7792 39824
rect 7808 39760 7872 39824
rect 7888 39760 7952 39824
rect 7968 39760 8032 39824
rect 8048 39760 8112 39824
rect 8128 39760 8192 39824
rect 8208 39760 8272 39824
rect 8288 39760 8352 39824
rect 8368 39760 8432 39824
rect 8448 39760 8512 39824
rect 8528 39760 8592 39824
rect 8608 39760 8672 39824
rect 8688 39760 8752 39824
rect 8768 39760 8832 39824
rect 8848 39760 8912 39824
rect 8928 39760 8992 39824
rect 14112 39760 14176 39824
rect 14192 39760 14256 39824
rect 14272 39760 14336 39824
rect 14352 39760 14416 39824
rect 24112 39760 24176 39824
rect 24192 39760 24256 39824
rect 24272 39760 24336 39824
rect 24352 39760 24416 39824
rect 36376 39760 36440 39824
rect 36456 39760 36520 39824
rect 36536 39760 36600 39824
rect 36616 39760 36680 39824
rect 36696 39760 36760 39824
rect 36776 39760 36840 39824
rect 36856 39760 36920 39824
rect 36936 39760 37000 39824
rect 37016 39760 37080 39824
rect 37096 39760 37160 39824
rect 37176 39760 37240 39824
rect 37256 39760 37320 39824
rect 37336 39760 37400 39824
rect 37416 39760 37480 39824
rect 37496 39760 37560 39824
rect 37576 39760 37640 39824
rect 37656 39760 37720 39824
rect 37736 39760 37800 39824
rect 37816 39760 37880 39824
rect 37896 39760 37960 39824
rect 37976 39760 38040 39824
rect 38056 39760 38120 39824
rect 38136 39760 38200 39824
rect 38216 39760 38280 39824
rect 38296 39760 38360 39824
rect 38376 39760 38440 39824
rect 38456 39760 38520 39824
rect 38536 39760 38600 39824
rect 38616 39760 38680 39824
rect 38696 39760 38760 39824
rect 38776 39760 38840 39824
rect 38856 39760 38920 39824
rect 38936 39760 39000 39824
rect 39016 39760 39080 39824
rect 39096 39760 39160 39824
rect 39176 39760 39240 39824
rect 39256 39760 39320 39824
rect 39336 39760 39400 39824
rect 39416 39760 39480 39824
rect 39496 39760 39560 39824
rect 39576 39760 39640 39824
rect 39656 39760 39720 39824
rect 39736 39760 39800 39824
rect 39816 39760 39880 39824
rect 39896 39760 39960 39824
rect 39976 39760 40040 39824
rect 40056 39760 40120 39824
rect 40136 39760 40200 39824
rect 40216 39760 40280 39824
rect 40296 39760 40360 39824
rect 5008 39680 5072 39744
rect 5088 39680 5152 39744
rect 5168 39680 5232 39744
rect 5248 39680 5312 39744
rect 5328 39680 5392 39744
rect 5408 39680 5472 39744
rect 5488 39680 5552 39744
rect 5568 39680 5632 39744
rect 5648 39680 5712 39744
rect 5728 39680 5792 39744
rect 5808 39680 5872 39744
rect 5888 39680 5952 39744
rect 5968 39680 6032 39744
rect 6048 39680 6112 39744
rect 6128 39680 6192 39744
rect 6208 39680 6272 39744
rect 6288 39680 6352 39744
rect 6368 39680 6432 39744
rect 6448 39680 6512 39744
rect 6528 39680 6592 39744
rect 6608 39680 6672 39744
rect 6688 39680 6752 39744
rect 6768 39680 6832 39744
rect 6848 39680 6912 39744
rect 6928 39680 6992 39744
rect 7008 39680 7072 39744
rect 7088 39680 7152 39744
rect 7168 39680 7232 39744
rect 7248 39680 7312 39744
rect 7328 39680 7392 39744
rect 7408 39680 7472 39744
rect 7488 39680 7552 39744
rect 7568 39680 7632 39744
rect 7648 39680 7712 39744
rect 7728 39680 7792 39744
rect 7808 39680 7872 39744
rect 7888 39680 7952 39744
rect 7968 39680 8032 39744
rect 8048 39680 8112 39744
rect 8128 39680 8192 39744
rect 8208 39680 8272 39744
rect 8288 39680 8352 39744
rect 8368 39680 8432 39744
rect 8448 39680 8512 39744
rect 8528 39680 8592 39744
rect 8608 39680 8672 39744
rect 8688 39680 8752 39744
rect 8768 39680 8832 39744
rect 8848 39680 8912 39744
rect 8928 39680 8992 39744
rect 14112 39680 14176 39744
rect 14192 39680 14256 39744
rect 14272 39680 14336 39744
rect 14352 39680 14416 39744
rect 24112 39680 24176 39744
rect 24192 39680 24256 39744
rect 24272 39680 24336 39744
rect 24352 39680 24416 39744
rect 36376 39680 36440 39744
rect 36456 39680 36520 39744
rect 36536 39680 36600 39744
rect 36616 39680 36680 39744
rect 36696 39680 36760 39744
rect 36776 39680 36840 39744
rect 36856 39680 36920 39744
rect 36936 39680 37000 39744
rect 37016 39680 37080 39744
rect 37096 39680 37160 39744
rect 37176 39680 37240 39744
rect 37256 39680 37320 39744
rect 37336 39680 37400 39744
rect 37416 39680 37480 39744
rect 37496 39680 37560 39744
rect 37576 39680 37640 39744
rect 37656 39680 37720 39744
rect 37736 39680 37800 39744
rect 37816 39680 37880 39744
rect 37896 39680 37960 39744
rect 37976 39680 38040 39744
rect 38056 39680 38120 39744
rect 38136 39680 38200 39744
rect 38216 39680 38280 39744
rect 38296 39680 38360 39744
rect 38376 39680 38440 39744
rect 38456 39680 38520 39744
rect 38536 39680 38600 39744
rect 38616 39680 38680 39744
rect 38696 39680 38760 39744
rect 38776 39680 38840 39744
rect 38856 39680 38920 39744
rect 38936 39680 39000 39744
rect 39016 39680 39080 39744
rect 39096 39680 39160 39744
rect 39176 39680 39240 39744
rect 39256 39680 39320 39744
rect 39336 39680 39400 39744
rect 39416 39680 39480 39744
rect 39496 39680 39560 39744
rect 39576 39680 39640 39744
rect 39656 39680 39720 39744
rect 39736 39680 39800 39744
rect 39816 39680 39880 39744
rect 39896 39680 39960 39744
rect 39976 39680 40040 39744
rect 40056 39680 40120 39744
rect 40136 39680 40200 39744
rect 40216 39680 40280 39744
rect 40296 39680 40360 39744
rect 5008 39600 5072 39664
rect 5088 39600 5152 39664
rect 5168 39600 5232 39664
rect 5248 39600 5312 39664
rect 5328 39600 5392 39664
rect 5408 39600 5472 39664
rect 5488 39600 5552 39664
rect 5568 39600 5632 39664
rect 5648 39600 5712 39664
rect 5728 39600 5792 39664
rect 5808 39600 5872 39664
rect 5888 39600 5952 39664
rect 5968 39600 6032 39664
rect 6048 39600 6112 39664
rect 6128 39600 6192 39664
rect 6208 39600 6272 39664
rect 6288 39600 6352 39664
rect 6368 39600 6432 39664
rect 6448 39600 6512 39664
rect 6528 39600 6592 39664
rect 6608 39600 6672 39664
rect 6688 39600 6752 39664
rect 6768 39600 6832 39664
rect 6848 39600 6912 39664
rect 6928 39600 6992 39664
rect 7008 39600 7072 39664
rect 7088 39600 7152 39664
rect 7168 39600 7232 39664
rect 7248 39600 7312 39664
rect 7328 39600 7392 39664
rect 7408 39600 7472 39664
rect 7488 39600 7552 39664
rect 7568 39600 7632 39664
rect 7648 39600 7712 39664
rect 7728 39600 7792 39664
rect 7808 39600 7872 39664
rect 7888 39600 7952 39664
rect 7968 39600 8032 39664
rect 8048 39600 8112 39664
rect 8128 39600 8192 39664
rect 8208 39600 8272 39664
rect 8288 39600 8352 39664
rect 8368 39600 8432 39664
rect 8448 39600 8512 39664
rect 8528 39600 8592 39664
rect 8608 39600 8672 39664
rect 8688 39600 8752 39664
rect 8768 39600 8832 39664
rect 8848 39600 8912 39664
rect 8928 39600 8992 39664
rect 14112 39600 14176 39664
rect 14192 39600 14256 39664
rect 14272 39600 14336 39664
rect 14352 39600 14416 39664
rect 24112 39600 24176 39664
rect 24192 39600 24256 39664
rect 24272 39600 24336 39664
rect 24352 39600 24416 39664
rect 36376 39600 36440 39664
rect 36456 39600 36520 39664
rect 36536 39600 36600 39664
rect 36616 39600 36680 39664
rect 36696 39600 36760 39664
rect 36776 39600 36840 39664
rect 36856 39600 36920 39664
rect 36936 39600 37000 39664
rect 37016 39600 37080 39664
rect 37096 39600 37160 39664
rect 37176 39600 37240 39664
rect 37256 39600 37320 39664
rect 37336 39600 37400 39664
rect 37416 39600 37480 39664
rect 37496 39600 37560 39664
rect 37576 39600 37640 39664
rect 37656 39600 37720 39664
rect 37736 39600 37800 39664
rect 37816 39600 37880 39664
rect 37896 39600 37960 39664
rect 37976 39600 38040 39664
rect 38056 39600 38120 39664
rect 38136 39600 38200 39664
rect 38216 39600 38280 39664
rect 38296 39600 38360 39664
rect 38376 39600 38440 39664
rect 38456 39600 38520 39664
rect 38536 39600 38600 39664
rect 38616 39600 38680 39664
rect 38696 39600 38760 39664
rect 38776 39600 38840 39664
rect 38856 39600 38920 39664
rect 38936 39600 39000 39664
rect 39016 39600 39080 39664
rect 39096 39600 39160 39664
rect 39176 39600 39240 39664
rect 39256 39600 39320 39664
rect 39336 39600 39400 39664
rect 39416 39600 39480 39664
rect 39496 39600 39560 39664
rect 39576 39600 39640 39664
rect 39656 39600 39720 39664
rect 39736 39600 39800 39664
rect 39816 39600 39880 39664
rect 39896 39600 39960 39664
rect 39976 39600 40040 39664
rect 40056 39600 40120 39664
rect 40136 39600 40200 39664
rect 40216 39600 40280 39664
rect 40296 39600 40360 39664
rect 5008 39520 5072 39584
rect 5088 39520 5152 39584
rect 5168 39520 5232 39584
rect 5248 39520 5312 39584
rect 5328 39520 5392 39584
rect 5408 39520 5472 39584
rect 5488 39520 5552 39584
rect 5568 39520 5632 39584
rect 5648 39520 5712 39584
rect 5728 39520 5792 39584
rect 5808 39520 5872 39584
rect 5888 39520 5952 39584
rect 5968 39520 6032 39584
rect 6048 39520 6112 39584
rect 6128 39520 6192 39584
rect 6208 39520 6272 39584
rect 6288 39520 6352 39584
rect 6368 39520 6432 39584
rect 6448 39520 6512 39584
rect 6528 39520 6592 39584
rect 6608 39520 6672 39584
rect 6688 39520 6752 39584
rect 6768 39520 6832 39584
rect 6848 39520 6912 39584
rect 6928 39520 6992 39584
rect 7008 39520 7072 39584
rect 7088 39520 7152 39584
rect 7168 39520 7232 39584
rect 7248 39520 7312 39584
rect 7328 39520 7392 39584
rect 7408 39520 7472 39584
rect 7488 39520 7552 39584
rect 7568 39520 7632 39584
rect 7648 39520 7712 39584
rect 7728 39520 7792 39584
rect 7808 39520 7872 39584
rect 7888 39520 7952 39584
rect 7968 39520 8032 39584
rect 8048 39520 8112 39584
rect 8128 39520 8192 39584
rect 8208 39520 8272 39584
rect 8288 39520 8352 39584
rect 8368 39520 8432 39584
rect 8448 39520 8512 39584
rect 8528 39520 8592 39584
rect 8608 39520 8672 39584
rect 8688 39520 8752 39584
rect 8768 39520 8832 39584
rect 8848 39520 8912 39584
rect 8928 39520 8992 39584
rect 14112 39520 14176 39584
rect 14192 39520 14256 39584
rect 14272 39520 14336 39584
rect 14352 39520 14416 39584
rect 24112 39520 24176 39584
rect 24192 39520 24256 39584
rect 24272 39520 24336 39584
rect 24352 39520 24416 39584
rect 36376 39520 36440 39584
rect 36456 39520 36520 39584
rect 36536 39520 36600 39584
rect 36616 39520 36680 39584
rect 36696 39520 36760 39584
rect 36776 39520 36840 39584
rect 36856 39520 36920 39584
rect 36936 39520 37000 39584
rect 37016 39520 37080 39584
rect 37096 39520 37160 39584
rect 37176 39520 37240 39584
rect 37256 39520 37320 39584
rect 37336 39520 37400 39584
rect 37416 39520 37480 39584
rect 37496 39520 37560 39584
rect 37576 39520 37640 39584
rect 37656 39520 37720 39584
rect 37736 39520 37800 39584
rect 37816 39520 37880 39584
rect 37896 39520 37960 39584
rect 37976 39520 38040 39584
rect 38056 39520 38120 39584
rect 38136 39520 38200 39584
rect 38216 39520 38280 39584
rect 38296 39520 38360 39584
rect 38376 39520 38440 39584
rect 38456 39520 38520 39584
rect 38536 39520 38600 39584
rect 38616 39520 38680 39584
rect 38696 39520 38760 39584
rect 38776 39520 38840 39584
rect 38856 39520 38920 39584
rect 38936 39520 39000 39584
rect 39016 39520 39080 39584
rect 39096 39520 39160 39584
rect 39176 39520 39240 39584
rect 39256 39520 39320 39584
rect 39336 39520 39400 39584
rect 39416 39520 39480 39584
rect 39496 39520 39560 39584
rect 39576 39520 39640 39584
rect 39656 39520 39720 39584
rect 39736 39520 39800 39584
rect 39816 39520 39880 39584
rect 39896 39520 39960 39584
rect 39976 39520 40040 39584
rect 40056 39520 40120 39584
rect 40136 39520 40200 39584
rect 40216 39520 40280 39584
rect 40296 39520 40360 39584
rect 5008 39440 5072 39504
rect 5088 39440 5152 39504
rect 5168 39440 5232 39504
rect 5248 39440 5312 39504
rect 5328 39440 5392 39504
rect 5408 39440 5472 39504
rect 5488 39440 5552 39504
rect 5568 39440 5632 39504
rect 5648 39440 5712 39504
rect 5728 39440 5792 39504
rect 5808 39440 5872 39504
rect 5888 39440 5952 39504
rect 5968 39440 6032 39504
rect 6048 39440 6112 39504
rect 6128 39440 6192 39504
rect 6208 39440 6272 39504
rect 6288 39440 6352 39504
rect 6368 39440 6432 39504
rect 6448 39440 6512 39504
rect 6528 39440 6592 39504
rect 6608 39440 6672 39504
rect 6688 39440 6752 39504
rect 6768 39440 6832 39504
rect 6848 39440 6912 39504
rect 6928 39440 6992 39504
rect 7008 39440 7072 39504
rect 7088 39440 7152 39504
rect 7168 39440 7232 39504
rect 7248 39440 7312 39504
rect 7328 39440 7392 39504
rect 7408 39440 7472 39504
rect 7488 39440 7552 39504
rect 7568 39440 7632 39504
rect 7648 39440 7712 39504
rect 7728 39440 7792 39504
rect 7808 39440 7872 39504
rect 7888 39440 7952 39504
rect 7968 39440 8032 39504
rect 8048 39440 8112 39504
rect 8128 39440 8192 39504
rect 8208 39440 8272 39504
rect 8288 39440 8352 39504
rect 8368 39440 8432 39504
rect 8448 39440 8512 39504
rect 8528 39440 8592 39504
rect 8608 39440 8672 39504
rect 8688 39440 8752 39504
rect 8768 39440 8832 39504
rect 8848 39440 8912 39504
rect 8928 39440 8992 39504
rect 14112 39440 14176 39504
rect 14192 39440 14256 39504
rect 14272 39440 14336 39504
rect 14352 39440 14416 39504
rect 24112 39440 24176 39504
rect 24192 39440 24256 39504
rect 24272 39440 24336 39504
rect 24352 39440 24416 39504
rect 36376 39440 36440 39504
rect 36456 39440 36520 39504
rect 36536 39440 36600 39504
rect 36616 39440 36680 39504
rect 36696 39440 36760 39504
rect 36776 39440 36840 39504
rect 36856 39440 36920 39504
rect 36936 39440 37000 39504
rect 37016 39440 37080 39504
rect 37096 39440 37160 39504
rect 37176 39440 37240 39504
rect 37256 39440 37320 39504
rect 37336 39440 37400 39504
rect 37416 39440 37480 39504
rect 37496 39440 37560 39504
rect 37576 39440 37640 39504
rect 37656 39440 37720 39504
rect 37736 39440 37800 39504
rect 37816 39440 37880 39504
rect 37896 39440 37960 39504
rect 37976 39440 38040 39504
rect 38056 39440 38120 39504
rect 38136 39440 38200 39504
rect 38216 39440 38280 39504
rect 38296 39440 38360 39504
rect 38376 39440 38440 39504
rect 38456 39440 38520 39504
rect 38536 39440 38600 39504
rect 38616 39440 38680 39504
rect 38696 39440 38760 39504
rect 38776 39440 38840 39504
rect 38856 39440 38920 39504
rect 38936 39440 39000 39504
rect 39016 39440 39080 39504
rect 39096 39440 39160 39504
rect 39176 39440 39240 39504
rect 39256 39440 39320 39504
rect 39336 39440 39400 39504
rect 39416 39440 39480 39504
rect 39496 39440 39560 39504
rect 39576 39440 39640 39504
rect 39656 39440 39720 39504
rect 39736 39440 39800 39504
rect 39816 39440 39880 39504
rect 39896 39440 39960 39504
rect 39976 39440 40040 39504
rect 40056 39440 40120 39504
rect 40136 39440 40200 39504
rect 40216 39440 40280 39504
rect 40296 39440 40360 39504
rect 5008 39360 5072 39424
rect 5088 39360 5152 39424
rect 5168 39360 5232 39424
rect 5248 39360 5312 39424
rect 5328 39360 5392 39424
rect 5408 39360 5472 39424
rect 5488 39360 5552 39424
rect 5568 39360 5632 39424
rect 5648 39360 5712 39424
rect 5728 39360 5792 39424
rect 5808 39360 5872 39424
rect 5888 39360 5952 39424
rect 5968 39360 6032 39424
rect 6048 39360 6112 39424
rect 6128 39360 6192 39424
rect 6208 39360 6272 39424
rect 6288 39360 6352 39424
rect 6368 39360 6432 39424
rect 6448 39360 6512 39424
rect 6528 39360 6592 39424
rect 6608 39360 6672 39424
rect 6688 39360 6752 39424
rect 6768 39360 6832 39424
rect 6848 39360 6912 39424
rect 6928 39360 6992 39424
rect 7008 39360 7072 39424
rect 7088 39360 7152 39424
rect 7168 39360 7232 39424
rect 7248 39360 7312 39424
rect 7328 39360 7392 39424
rect 7408 39360 7472 39424
rect 7488 39360 7552 39424
rect 7568 39360 7632 39424
rect 7648 39360 7712 39424
rect 7728 39360 7792 39424
rect 7808 39360 7872 39424
rect 7888 39360 7952 39424
rect 7968 39360 8032 39424
rect 8048 39360 8112 39424
rect 8128 39360 8192 39424
rect 8208 39360 8272 39424
rect 8288 39360 8352 39424
rect 8368 39360 8432 39424
rect 8448 39360 8512 39424
rect 8528 39360 8592 39424
rect 8608 39360 8672 39424
rect 8688 39360 8752 39424
rect 8768 39360 8832 39424
rect 8848 39360 8912 39424
rect 8928 39360 8992 39424
rect 14112 39360 14176 39424
rect 14192 39360 14256 39424
rect 14272 39360 14336 39424
rect 14352 39360 14416 39424
rect 24112 39360 24176 39424
rect 24192 39360 24256 39424
rect 24272 39360 24336 39424
rect 24352 39360 24416 39424
rect 36376 39360 36440 39424
rect 36456 39360 36520 39424
rect 36536 39360 36600 39424
rect 36616 39360 36680 39424
rect 36696 39360 36760 39424
rect 36776 39360 36840 39424
rect 36856 39360 36920 39424
rect 36936 39360 37000 39424
rect 37016 39360 37080 39424
rect 37096 39360 37160 39424
rect 37176 39360 37240 39424
rect 37256 39360 37320 39424
rect 37336 39360 37400 39424
rect 37416 39360 37480 39424
rect 37496 39360 37560 39424
rect 37576 39360 37640 39424
rect 37656 39360 37720 39424
rect 37736 39360 37800 39424
rect 37816 39360 37880 39424
rect 37896 39360 37960 39424
rect 37976 39360 38040 39424
rect 38056 39360 38120 39424
rect 38136 39360 38200 39424
rect 38216 39360 38280 39424
rect 38296 39360 38360 39424
rect 38376 39360 38440 39424
rect 38456 39360 38520 39424
rect 38536 39360 38600 39424
rect 38616 39360 38680 39424
rect 38696 39360 38760 39424
rect 38776 39360 38840 39424
rect 38856 39360 38920 39424
rect 38936 39360 39000 39424
rect 39016 39360 39080 39424
rect 39096 39360 39160 39424
rect 39176 39360 39240 39424
rect 39256 39360 39320 39424
rect 39336 39360 39400 39424
rect 39416 39360 39480 39424
rect 39496 39360 39560 39424
rect 39576 39360 39640 39424
rect 39656 39360 39720 39424
rect 39736 39360 39800 39424
rect 39816 39360 39880 39424
rect 39896 39360 39960 39424
rect 39976 39360 40040 39424
rect 40056 39360 40120 39424
rect 40136 39360 40200 39424
rect 40216 39360 40280 39424
rect 40296 39360 40360 39424
rect 5008 39280 5072 39344
rect 5088 39280 5152 39344
rect 5168 39280 5232 39344
rect 5248 39280 5312 39344
rect 5328 39280 5392 39344
rect 5408 39280 5472 39344
rect 5488 39280 5552 39344
rect 5568 39280 5632 39344
rect 5648 39280 5712 39344
rect 5728 39280 5792 39344
rect 5808 39280 5872 39344
rect 5888 39280 5952 39344
rect 5968 39280 6032 39344
rect 6048 39280 6112 39344
rect 6128 39280 6192 39344
rect 6208 39280 6272 39344
rect 6288 39280 6352 39344
rect 6368 39280 6432 39344
rect 6448 39280 6512 39344
rect 6528 39280 6592 39344
rect 6608 39280 6672 39344
rect 6688 39280 6752 39344
rect 6768 39280 6832 39344
rect 6848 39280 6912 39344
rect 6928 39280 6992 39344
rect 7008 39280 7072 39344
rect 7088 39280 7152 39344
rect 7168 39280 7232 39344
rect 7248 39280 7312 39344
rect 7328 39280 7392 39344
rect 7408 39280 7472 39344
rect 7488 39280 7552 39344
rect 7568 39280 7632 39344
rect 7648 39280 7712 39344
rect 7728 39280 7792 39344
rect 7808 39280 7872 39344
rect 7888 39280 7952 39344
rect 7968 39280 8032 39344
rect 8048 39280 8112 39344
rect 8128 39280 8192 39344
rect 8208 39280 8272 39344
rect 8288 39280 8352 39344
rect 8368 39280 8432 39344
rect 8448 39280 8512 39344
rect 8528 39280 8592 39344
rect 8608 39280 8672 39344
rect 8688 39280 8752 39344
rect 8768 39280 8832 39344
rect 8848 39280 8912 39344
rect 8928 39280 8992 39344
rect 14112 39280 14176 39344
rect 14192 39280 14256 39344
rect 14272 39280 14336 39344
rect 14352 39280 14416 39344
rect 24112 39280 24176 39344
rect 24192 39280 24256 39344
rect 24272 39280 24336 39344
rect 24352 39280 24416 39344
rect 36376 39280 36440 39344
rect 36456 39280 36520 39344
rect 36536 39280 36600 39344
rect 36616 39280 36680 39344
rect 36696 39280 36760 39344
rect 36776 39280 36840 39344
rect 36856 39280 36920 39344
rect 36936 39280 37000 39344
rect 37016 39280 37080 39344
rect 37096 39280 37160 39344
rect 37176 39280 37240 39344
rect 37256 39280 37320 39344
rect 37336 39280 37400 39344
rect 37416 39280 37480 39344
rect 37496 39280 37560 39344
rect 37576 39280 37640 39344
rect 37656 39280 37720 39344
rect 37736 39280 37800 39344
rect 37816 39280 37880 39344
rect 37896 39280 37960 39344
rect 37976 39280 38040 39344
rect 38056 39280 38120 39344
rect 38136 39280 38200 39344
rect 38216 39280 38280 39344
rect 38296 39280 38360 39344
rect 38376 39280 38440 39344
rect 38456 39280 38520 39344
rect 38536 39280 38600 39344
rect 38616 39280 38680 39344
rect 38696 39280 38760 39344
rect 38776 39280 38840 39344
rect 38856 39280 38920 39344
rect 38936 39280 39000 39344
rect 39016 39280 39080 39344
rect 39096 39280 39160 39344
rect 39176 39280 39240 39344
rect 39256 39280 39320 39344
rect 39336 39280 39400 39344
rect 39416 39280 39480 39344
rect 39496 39280 39560 39344
rect 39576 39280 39640 39344
rect 39656 39280 39720 39344
rect 39736 39280 39800 39344
rect 39816 39280 39880 39344
rect 39896 39280 39960 39344
rect 39976 39280 40040 39344
rect 40056 39280 40120 39344
rect 40136 39280 40200 39344
rect 40216 39280 40280 39344
rect 40296 39280 40360 39344
rect 5008 39200 5072 39264
rect 5088 39200 5152 39264
rect 5168 39200 5232 39264
rect 5248 39200 5312 39264
rect 5328 39200 5392 39264
rect 5408 39200 5472 39264
rect 5488 39200 5552 39264
rect 5568 39200 5632 39264
rect 5648 39200 5712 39264
rect 5728 39200 5792 39264
rect 5808 39200 5872 39264
rect 5888 39200 5952 39264
rect 5968 39200 6032 39264
rect 6048 39200 6112 39264
rect 6128 39200 6192 39264
rect 6208 39200 6272 39264
rect 6288 39200 6352 39264
rect 6368 39200 6432 39264
rect 6448 39200 6512 39264
rect 6528 39200 6592 39264
rect 6608 39200 6672 39264
rect 6688 39200 6752 39264
rect 6768 39200 6832 39264
rect 6848 39200 6912 39264
rect 6928 39200 6992 39264
rect 7008 39200 7072 39264
rect 7088 39200 7152 39264
rect 7168 39200 7232 39264
rect 7248 39200 7312 39264
rect 7328 39200 7392 39264
rect 7408 39200 7472 39264
rect 7488 39200 7552 39264
rect 7568 39200 7632 39264
rect 7648 39200 7712 39264
rect 7728 39200 7792 39264
rect 7808 39200 7872 39264
rect 7888 39200 7952 39264
rect 7968 39200 8032 39264
rect 8048 39200 8112 39264
rect 8128 39200 8192 39264
rect 8208 39200 8272 39264
rect 8288 39200 8352 39264
rect 8368 39200 8432 39264
rect 8448 39200 8512 39264
rect 8528 39200 8592 39264
rect 8608 39200 8672 39264
rect 8688 39200 8752 39264
rect 8768 39200 8832 39264
rect 8848 39200 8912 39264
rect 8928 39200 8992 39264
rect 14112 39200 14176 39264
rect 14192 39200 14256 39264
rect 14272 39200 14336 39264
rect 14352 39200 14416 39264
rect 24112 39200 24176 39264
rect 24192 39200 24256 39264
rect 24272 39200 24336 39264
rect 24352 39200 24416 39264
rect 36376 39200 36440 39264
rect 36456 39200 36520 39264
rect 36536 39200 36600 39264
rect 36616 39200 36680 39264
rect 36696 39200 36760 39264
rect 36776 39200 36840 39264
rect 36856 39200 36920 39264
rect 36936 39200 37000 39264
rect 37016 39200 37080 39264
rect 37096 39200 37160 39264
rect 37176 39200 37240 39264
rect 37256 39200 37320 39264
rect 37336 39200 37400 39264
rect 37416 39200 37480 39264
rect 37496 39200 37560 39264
rect 37576 39200 37640 39264
rect 37656 39200 37720 39264
rect 37736 39200 37800 39264
rect 37816 39200 37880 39264
rect 37896 39200 37960 39264
rect 37976 39200 38040 39264
rect 38056 39200 38120 39264
rect 38136 39200 38200 39264
rect 38216 39200 38280 39264
rect 38296 39200 38360 39264
rect 38376 39200 38440 39264
rect 38456 39200 38520 39264
rect 38536 39200 38600 39264
rect 38616 39200 38680 39264
rect 38696 39200 38760 39264
rect 38776 39200 38840 39264
rect 38856 39200 38920 39264
rect 38936 39200 39000 39264
rect 39016 39200 39080 39264
rect 39096 39200 39160 39264
rect 39176 39200 39240 39264
rect 39256 39200 39320 39264
rect 39336 39200 39400 39264
rect 39416 39200 39480 39264
rect 39496 39200 39560 39264
rect 39576 39200 39640 39264
rect 39656 39200 39720 39264
rect 39736 39200 39800 39264
rect 39816 39200 39880 39264
rect 39896 39200 39960 39264
rect 39976 39200 40040 39264
rect 40056 39200 40120 39264
rect 40136 39200 40200 39264
rect 40216 39200 40280 39264
rect 40296 39200 40360 39264
rect 5008 39120 5072 39184
rect 5088 39120 5152 39184
rect 5168 39120 5232 39184
rect 5248 39120 5312 39184
rect 5328 39120 5392 39184
rect 5408 39120 5472 39184
rect 5488 39120 5552 39184
rect 5568 39120 5632 39184
rect 5648 39120 5712 39184
rect 5728 39120 5792 39184
rect 5808 39120 5872 39184
rect 5888 39120 5952 39184
rect 5968 39120 6032 39184
rect 6048 39120 6112 39184
rect 6128 39120 6192 39184
rect 6208 39120 6272 39184
rect 6288 39120 6352 39184
rect 6368 39120 6432 39184
rect 6448 39120 6512 39184
rect 6528 39120 6592 39184
rect 6608 39120 6672 39184
rect 6688 39120 6752 39184
rect 6768 39120 6832 39184
rect 6848 39120 6912 39184
rect 6928 39120 6992 39184
rect 7008 39120 7072 39184
rect 7088 39120 7152 39184
rect 7168 39120 7232 39184
rect 7248 39120 7312 39184
rect 7328 39120 7392 39184
rect 7408 39120 7472 39184
rect 7488 39120 7552 39184
rect 7568 39120 7632 39184
rect 7648 39120 7712 39184
rect 7728 39120 7792 39184
rect 7808 39120 7872 39184
rect 7888 39120 7952 39184
rect 7968 39120 8032 39184
rect 8048 39120 8112 39184
rect 8128 39120 8192 39184
rect 8208 39120 8272 39184
rect 8288 39120 8352 39184
rect 8368 39120 8432 39184
rect 8448 39120 8512 39184
rect 8528 39120 8592 39184
rect 8608 39120 8672 39184
rect 8688 39120 8752 39184
rect 8768 39120 8832 39184
rect 8848 39120 8912 39184
rect 8928 39120 8992 39184
rect 14112 39120 14176 39184
rect 14192 39120 14256 39184
rect 14272 39120 14336 39184
rect 14352 39120 14416 39184
rect 24112 39120 24176 39184
rect 24192 39120 24256 39184
rect 24272 39120 24336 39184
rect 24352 39120 24416 39184
rect 36376 39120 36440 39184
rect 36456 39120 36520 39184
rect 36536 39120 36600 39184
rect 36616 39120 36680 39184
rect 36696 39120 36760 39184
rect 36776 39120 36840 39184
rect 36856 39120 36920 39184
rect 36936 39120 37000 39184
rect 37016 39120 37080 39184
rect 37096 39120 37160 39184
rect 37176 39120 37240 39184
rect 37256 39120 37320 39184
rect 37336 39120 37400 39184
rect 37416 39120 37480 39184
rect 37496 39120 37560 39184
rect 37576 39120 37640 39184
rect 37656 39120 37720 39184
rect 37736 39120 37800 39184
rect 37816 39120 37880 39184
rect 37896 39120 37960 39184
rect 37976 39120 38040 39184
rect 38056 39120 38120 39184
rect 38136 39120 38200 39184
rect 38216 39120 38280 39184
rect 38296 39120 38360 39184
rect 38376 39120 38440 39184
rect 38456 39120 38520 39184
rect 38536 39120 38600 39184
rect 38616 39120 38680 39184
rect 38696 39120 38760 39184
rect 38776 39120 38840 39184
rect 38856 39120 38920 39184
rect 38936 39120 39000 39184
rect 39016 39120 39080 39184
rect 39096 39120 39160 39184
rect 39176 39120 39240 39184
rect 39256 39120 39320 39184
rect 39336 39120 39400 39184
rect 39416 39120 39480 39184
rect 39496 39120 39560 39184
rect 39576 39120 39640 39184
rect 39656 39120 39720 39184
rect 39736 39120 39800 39184
rect 39816 39120 39880 39184
rect 39896 39120 39960 39184
rect 39976 39120 40040 39184
rect 40056 39120 40120 39184
rect 40136 39120 40200 39184
rect 40216 39120 40280 39184
rect 40296 39120 40360 39184
rect 5008 39040 5072 39104
rect 5088 39040 5152 39104
rect 5168 39040 5232 39104
rect 5248 39040 5312 39104
rect 5328 39040 5392 39104
rect 5408 39040 5472 39104
rect 5488 39040 5552 39104
rect 5568 39040 5632 39104
rect 5648 39040 5712 39104
rect 5728 39040 5792 39104
rect 5808 39040 5872 39104
rect 5888 39040 5952 39104
rect 5968 39040 6032 39104
rect 6048 39040 6112 39104
rect 6128 39040 6192 39104
rect 6208 39040 6272 39104
rect 6288 39040 6352 39104
rect 6368 39040 6432 39104
rect 6448 39040 6512 39104
rect 6528 39040 6592 39104
rect 6608 39040 6672 39104
rect 6688 39040 6752 39104
rect 6768 39040 6832 39104
rect 6848 39040 6912 39104
rect 6928 39040 6992 39104
rect 7008 39040 7072 39104
rect 7088 39040 7152 39104
rect 7168 39040 7232 39104
rect 7248 39040 7312 39104
rect 7328 39040 7392 39104
rect 7408 39040 7472 39104
rect 7488 39040 7552 39104
rect 7568 39040 7632 39104
rect 7648 39040 7712 39104
rect 7728 39040 7792 39104
rect 7808 39040 7872 39104
rect 7888 39040 7952 39104
rect 7968 39040 8032 39104
rect 8048 39040 8112 39104
rect 8128 39040 8192 39104
rect 8208 39040 8272 39104
rect 8288 39040 8352 39104
rect 8368 39040 8432 39104
rect 8448 39040 8512 39104
rect 8528 39040 8592 39104
rect 8608 39040 8672 39104
rect 8688 39040 8752 39104
rect 8768 39040 8832 39104
rect 8848 39040 8912 39104
rect 8928 39040 8992 39104
rect 14112 39040 14176 39104
rect 14192 39040 14256 39104
rect 14272 39040 14336 39104
rect 14352 39040 14416 39104
rect 24112 39040 24176 39104
rect 24192 39040 24256 39104
rect 24272 39040 24336 39104
rect 24352 39040 24416 39104
rect 36376 39040 36440 39104
rect 36456 39040 36520 39104
rect 36536 39040 36600 39104
rect 36616 39040 36680 39104
rect 36696 39040 36760 39104
rect 36776 39040 36840 39104
rect 36856 39040 36920 39104
rect 36936 39040 37000 39104
rect 37016 39040 37080 39104
rect 37096 39040 37160 39104
rect 37176 39040 37240 39104
rect 37256 39040 37320 39104
rect 37336 39040 37400 39104
rect 37416 39040 37480 39104
rect 37496 39040 37560 39104
rect 37576 39040 37640 39104
rect 37656 39040 37720 39104
rect 37736 39040 37800 39104
rect 37816 39040 37880 39104
rect 37896 39040 37960 39104
rect 37976 39040 38040 39104
rect 38056 39040 38120 39104
rect 38136 39040 38200 39104
rect 38216 39040 38280 39104
rect 38296 39040 38360 39104
rect 38376 39040 38440 39104
rect 38456 39040 38520 39104
rect 38536 39040 38600 39104
rect 38616 39040 38680 39104
rect 38696 39040 38760 39104
rect 38776 39040 38840 39104
rect 38856 39040 38920 39104
rect 38936 39040 39000 39104
rect 39016 39040 39080 39104
rect 39096 39040 39160 39104
rect 39176 39040 39240 39104
rect 39256 39040 39320 39104
rect 39336 39040 39400 39104
rect 39416 39040 39480 39104
rect 39496 39040 39560 39104
rect 39576 39040 39640 39104
rect 39656 39040 39720 39104
rect 39736 39040 39800 39104
rect 39816 39040 39880 39104
rect 39896 39040 39960 39104
rect 39976 39040 40040 39104
rect 40056 39040 40120 39104
rect 40136 39040 40200 39104
rect 40216 39040 40280 39104
rect 40296 39040 40360 39104
rect 5008 38960 5072 39024
rect 5088 38960 5152 39024
rect 5168 38960 5232 39024
rect 5248 38960 5312 39024
rect 5328 38960 5392 39024
rect 5408 38960 5472 39024
rect 5488 38960 5552 39024
rect 5568 38960 5632 39024
rect 5648 38960 5712 39024
rect 5728 38960 5792 39024
rect 5808 38960 5872 39024
rect 5888 38960 5952 39024
rect 5968 38960 6032 39024
rect 6048 38960 6112 39024
rect 6128 38960 6192 39024
rect 6208 38960 6272 39024
rect 6288 38960 6352 39024
rect 6368 38960 6432 39024
rect 6448 38960 6512 39024
rect 6528 38960 6592 39024
rect 6608 38960 6672 39024
rect 6688 38960 6752 39024
rect 6768 38960 6832 39024
rect 6848 38960 6912 39024
rect 6928 38960 6992 39024
rect 7008 38960 7072 39024
rect 7088 38960 7152 39024
rect 7168 38960 7232 39024
rect 7248 38960 7312 39024
rect 7328 38960 7392 39024
rect 7408 38960 7472 39024
rect 7488 38960 7552 39024
rect 7568 38960 7632 39024
rect 7648 38960 7712 39024
rect 7728 38960 7792 39024
rect 7808 38960 7872 39024
rect 7888 38960 7952 39024
rect 7968 38960 8032 39024
rect 8048 38960 8112 39024
rect 8128 38960 8192 39024
rect 8208 38960 8272 39024
rect 8288 38960 8352 39024
rect 8368 38960 8432 39024
rect 8448 38960 8512 39024
rect 8528 38960 8592 39024
rect 8608 38960 8672 39024
rect 8688 38960 8752 39024
rect 8768 38960 8832 39024
rect 8848 38960 8912 39024
rect 8928 38960 8992 39024
rect 14112 38960 14176 39024
rect 14192 38960 14256 39024
rect 14272 38960 14336 39024
rect 14352 38960 14416 39024
rect 24112 38960 24176 39024
rect 24192 38960 24256 39024
rect 24272 38960 24336 39024
rect 24352 38960 24416 39024
rect 36376 38960 36440 39024
rect 36456 38960 36520 39024
rect 36536 38960 36600 39024
rect 36616 38960 36680 39024
rect 36696 38960 36760 39024
rect 36776 38960 36840 39024
rect 36856 38960 36920 39024
rect 36936 38960 37000 39024
rect 37016 38960 37080 39024
rect 37096 38960 37160 39024
rect 37176 38960 37240 39024
rect 37256 38960 37320 39024
rect 37336 38960 37400 39024
rect 37416 38960 37480 39024
rect 37496 38960 37560 39024
rect 37576 38960 37640 39024
rect 37656 38960 37720 39024
rect 37736 38960 37800 39024
rect 37816 38960 37880 39024
rect 37896 38960 37960 39024
rect 37976 38960 38040 39024
rect 38056 38960 38120 39024
rect 38136 38960 38200 39024
rect 38216 38960 38280 39024
rect 38296 38960 38360 39024
rect 38376 38960 38440 39024
rect 38456 38960 38520 39024
rect 38536 38960 38600 39024
rect 38616 38960 38680 39024
rect 38696 38960 38760 39024
rect 38776 38960 38840 39024
rect 38856 38960 38920 39024
rect 38936 38960 39000 39024
rect 39016 38960 39080 39024
rect 39096 38960 39160 39024
rect 39176 38960 39240 39024
rect 39256 38960 39320 39024
rect 39336 38960 39400 39024
rect 39416 38960 39480 39024
rect 39496 38960 39560 39024
rect 39576 38960 39640 39024
rect 39656 38960 39720 39024
rect 39736 38960 39800 39024
rect 39816 38960 39880 39024
rect 39896 38960 39960 39024
rect 39976 38960 40040 39024
rect 40056 38960 40120 39024
rect 40136 38960 40200 39024
rect 40216 38960 40280 39024
rect 40296 38960 40360 39024
rect 5008 38880 5072 38944
rect 5088 38880 5152 38944
rect 5168 38880 5232 38944
rect 5248 38880 5312 38944
rect 5328 38880 5392 38944
rect 5408 38880 5472 38944
rect 5488 38880 5552 38944
rect 5568 38880 5632 38944
rect 5648 38880 5712 38944
rect 5728 38880 5792 38944
rect 5808 38880 5872 38944
rect 5888 38880 5952 38944
rect 5968 38880 6032 38944
rect 6048 38880 6112 38944
rect 6128 38880 6192 38944
rect 6208 38880 6272 38944
rect 6288 38880 6352 38944
rect 6368 38880 6432 38944
rect 6448 38880 6512 38944
rect 6528 38880 6592 38944
rect 6608 38880 6672 38944
rect 6688 38880 6752 38944
rect 6768 38880 6832 38944
rect 6848 38880 6912 38944
rect 6928 38880 6992 38944
rect 7008 38880 7072 38944
rect 7088 38880 7152 38944
rect 7168 38880 7232 38944
rect 7248 38880 7312 38944
rect 7328 38880 7392 38944
rect 7408 38880 7472 38944
rect 7488 38880 7552 38944
rect 7568 38880 7632 38944
rect 7648 38880 7712 38944
rect 7728 38880 7792 38944
rect 7808 38880 7872 38944
rect 7888 38880 7952 38944
rect 7968 38880 8032 38944
rect 8048 38880 8112 38944
rect 8128 38880 8192 38944
rect 8208 38880 8272 38944
rect 8288 38880 8352 38944
rect 8368 38880 8432 38944
rect 8448 38880 8512 38944
rect 8528 38880 8592 38944
rect 8608 38880 8672 38944
rect 8688 38880 8752 38944
rect 8768 38880 8832 38944
rect 8848 38880 8912 38944
rect 8928 38880 8992 38944
rect 14112 38880 14176 38944
rect 14192 38880 14256 38944
rect 14272 38880 14336 38944
rect 14352 38880 14416 38944
rect 24112 38880 24176 38944
rect 24192 38880 24256 38944
rect 24272 38880 24336 38944
rect 24352 38880 24416 38944
rect 36376 38880 36440 38944
rect 36456 38880 36520 38944
rect 36536 38880 36600 38944
rect 36616 38880 36680 38944
rect 36696 38880 36760 38944
rect 36776 38880 36840 38944
rect 36856 38880 36920 38944
rect 36936 38880 37000 38944
rect 37016 38880 37080 38944
rect 37096 38880 37160 38944
rect 37176 38880 37240 38944
rect 37256 38880 37320 38944
rect 37336 38880 37400 38944
rect 37416 38880 37480 38944
rect 37496 38880 37560 38944
rect 37576 38880 37640 38944
rect 37656 38880 37720 38944
rect 37736 38880 37800 38944
rect 37816 38880 37880 38944
rect 37896 38880 37960 38944
rect 37976 38880 38040 38944
rect 38056 38880 38120 38944
rect 38136 38880 38200 38944
rect 38216 38880 38280 38944
rect 38296 38880 38360 38944
rect 38376 38880 38440 38944
rect 38456 38880 38520 38944
rect 38536 38880 38600 38944
rect 38616 38880 38680 38944
rect 38696 38880 38760 38944
rect 38776 38880 38840 38944
rect 38856 38880 38920 38944
rect 38936 38880 39000 38944
rect 39016 38880 39080 38944
rect 39096 38880 39160 38944
rect 39176 38880 39240 38944
rect 39256 38880 39320 38944
rect 39336 38880 39400 38944
rect 39416 38880 39480 38944
rect 39496 38880 39560 38944
rect 39576 38880 39640 38944
rect 39656 38880 39720 38944
rect 39736 38880 39800 38944
rect 39816 38880 39880 38944
rect 39896 38880 39960 38944
rect 39976 38880 40040 38944
rect 40056 38880 40120 38944
rect 40136 38880 40200 38944
rect 40216 38880 40280 38944
rect 40296 38880 40360 38944
rect 5008 38800 5072 38864
rect 5088 38800 5152 38864
rect 5168 38800 5232 38864
rect 5248 38800 5312 38864
rect 5328 38800 5392 38864
rect 5408 38800 5472 38864
rect 5488 38800 5552 38864
rect 5568 38800 5632 38864
rect 5648 38800 5712 38864
rect 5728 38800 5792 38864
rect 5808 38800 5872 38864
rect 5888 38800 5952 38864
rect 5968 38800 6032 38864
rect 6048 38800 6112 38864
rect 6128 38800 6192 38864
rect 6208 38800 6272 38864
rect 6288 38800 6352 38864
rect 6368 38800 6432 38864
rect 6448 38800 6512 38864
rect 6528 38800 6592 38864
rect 6608 38800 6672 38864
rect 6688 38800 6752 38864
rect 6768 38800 6832 38864
rect 6848 38800 6912 38864
rect 6928 38800 6992 38864
rect 7008 38800 7072 38864
rect 7088 38800 7152 38864
rect 7168 38800 7232 38864
rect 7248 38800 7312 38864
rect 7328 38800 7392 38864
rect 7408 38800 7472 38864
rect 7488 38800 7552 38864
rect 7568 38800 7632 38864
rect 7648 38800 7712 38864
rect 7728 38800 7792 38864
rect 7808 38800 7872 38864
rect 7888 38800 7952 38864
rect 7968 38800 8032 38864
rect 8048 38800 8112 38864
rect 8128 38800 8192 38864
rect 8208 38800 8272 38864
rect 8288 38800 8352 38864
rect 8368 38800 8432 38864
rect 8448 38800 8512 38864
rect 8528 38800 8592 38864
rect 8608 38800 8672 38864
rect 8688 38800 8752 38864
rect 8768 38800 8832 38864
rect 8848 38800 8912 38864
rect 8928 38800 8992 38864
rect 14112 38800 14176 38864
rect 14192 38800 14256 38864
rect 14272 38800 14336 38864
rect 14352 38800 14416 38864
rect 24112 38800 24176 38864
rect 24192 38800 24256 38864
rect 24272 38800 24336 38864
rect 24352 38800 24416 38864
rect 36376 38800 36440 38864
rect 36456 38800 36520 38864
rect 36536 38800 36600 38864
rect 36616 38800 36680 38864
rect 36696 38800 36760 38864
rect 36776 38800 36840 38864
rect 36856 38800 36920 38864
rect 36936 38800 37000 38864
rect 37016 38800 37080 38864
rect 37096 38800 37160 38864
rect 37176 38800 37240 38864
rect 37256 38800 37320 38864
rect 37336 38800 37400 38864
rect 37416 38800 37480 38864
rect 37496 38800 37560 38864
rect 37576 38800 37640 38864
rect 37656 38800 37720 38864
rect 37736 38800 37800 38864
rect 37816 38800 37880 38864
rect 37896 38800 37960 38864
rect 37976 38800 38040 38864
rect 38056 38800 38120 38864
rect 38136 38800 38200 38864
rect 38216 38800 38280 38864
rect 38296 38800 38360 38864
rect 38376 38800 38440 38864
rect 38456 38800 38520 38864
rect 38536 38800 38600 38864
rect 38616 38800 38680 38864
rect 38696 38800 38760 38864
rect 38776 38800 38840 38864
rect 38856 38800 38920 38864
rect 38936 38800 39000 38864
rect 39016 38800 39080 38864
rect 39096 38800 39160 38864
rect 39176 38800 39240 38864
rect 39256 38800 39320 38864
rect 39336 38800 39400 38864
rect 39416 38800 39480 38864
rect 39496 38800 39560 38864
rect 39576 38800 39640 38864
rect 39656 38800 39720 38864
rect 39736 38800 39800 38864
rect 39816 38800 39880 38864
rect 39896 38800 39960 38864
rect 39976 38800 40040 38864
rect 40056 38800 40120 38864
rect 40136 38800 40200 38864
rect 40216 38800 40280 38864
rect 40296 38800 40360 38864
rect 5008 38720 5072 38784
rect 5088 38720 5152 38784
rect 5168 38720 5232 38784
rect 5248 38720 5312 38784
rect 5328 38720 5392 38784
rect 5408 38720 5472 38784
rect 5488 38720 5552 38784
rect 5568 38720 5632 38784
rect 5648 38720 5712 38784
rect 5728 38720 5792 38784
rect 5808 38720 5872 38784
rect 5888 38720 5952 38784
rect 5968 38720 6032 38784
rect 6048 38720 6112 38784
rect 6128 38720 6192 38784
rect 6208 38720 6272 38784
rect 6288 38720 6352 38784
rect 6368 38720 6432 38784
rect 6448 38720 6512 38784
rect 6528 38720 6592 38784
rect 6608 38720 6672 38784
rect 6688 38720 6752 38784
rect 6768 38720 6832 38784
rect 6848 38720 6912 38784
rect 6928 38720 6992 38784
rect 7008 38720 7072 38784
rect 7088 38720 7152 38784
rect 7168 38720 7232 38784
rect 7248 38720 7312 38784
rect 7328 38720 7392 38784
rect 7408 38720 7472 38784
rect 7488 38720 7552 38784
rect 7568 38720 7632 38784
rect 7648 38720 7712 38784
rect 7728 38720 7792 38784
rect 7808 38720 7872 38784
rect 7888 38720 7952 38784
rect 7968 38720 8032 38784
rect 8048 38720 8112 38784
rect 8128 38720 8192 38784
rect 8208 38720 8272 38784
rect 8288 38720 8352 38784
rect 8368 38720 8432 38784
rect 8448 38720 8512 38784
rect 8528 38720 8592 38784
rect 8608 38720 8672 38784
rect 8688 38720 8752 38784
rect 8768 38720 8832 38784
rect 8848 38720 8912 38784
rect 8928 38720 8992 38784
rect 14112 38720 14176 38784
rect 14192 38720 14256 38784
rect 14272 38720 14336 38784
rect 14352 38720 14416 38784
rect 24112 38720 24176 38784
rect 24192 38720 24256 38784
rect 24272 38720 24336 38784
rect 24352 38720 24416 38784
rect 36376 38720 36440 38784
rect 36456 38720 36520 38784
rect 36536 38720 36600 38784
rect 36616 38720 36680 38784
rect 36696 38720 36760 38784
rect 36776 38720 36840 38784
rect 36856 38720 36920 38784
rect 36936 38720 37000 38784
rect 37016 38720 37080 38784
rect 37096 38720 37160 38784
rect 37176 38720 37240 38784
rect 37256 38720 37320 38784
rect 37336 38720 37400 38784
rect 37416 38720 37480 38784
rect 37496 38720 37560 38784
rect 37576 38720 37640 38784
rect 37656 38720 37720 38784
rect 37736 38720 37800 38784
rect 37816 38720 37880 38784
rect 37896 38720 37960 38784
rect 37976 38720 38040 38784
rect 38056 38720 38120 38784
rect 38136 38720 38200 38784
rect 38216 38720 38280 38784
rect 38296 38720 38360 38784
rect 38376 38720 38440 38784
rect 38456 38720 38520 38784
rect 38536 38720 38600 38784
rect 38616 38720 38680 38784
rect 38696 38720 38760 38784
rect 38776 38720 38840 38784
rect 38856 38720 38920 38784
rect 38936 38720 39000 38784
rect 39016 38720 39080 38784
rect 39096 38720 39160 38784
rect 39176 38720 39240 38784
rect 39256 38720 39320 38784
rect 39336 38720 39400 38784
rect 39416 38720 39480 38784
rect 39496 38720 39560 38784
rect 39576 38720 39640 38784
rect 39656 38720 39720 38784
rect 39736 38720 39800 38784
rect 39816 38720 39880 38784
rect 39896 38720 39960 38784
rect 39976 38720 40040 38784
rect 40056 38720 40120 38784
rect 40136 38720 40200 38784
rect 40216 38720 40280 38784
rect 40296 38720 40360 38784
rect 5008 38640 5072 38704
rect 5088 38640 5152 38704
rect 5168 38640 5232 38704
rect 5248 38640 5312 38704
rect 5328 38640 5392 38704
rect 5408 38640 5472 38704
rect 5488 38640 5552 38704
rect 5568 38640 5632 38704
rect 5648 38640 5712 38704
rect 5728 38640 5792 38704
rect 5808 38640 5872 38704
rect 5888 38640 5952 38704
rect 5968 38640 6032 38704
rect 6048 38640 6112 38704
rect 6128 38640 6192 38704
rect 6208 38640 6272 38704
rect 6288 38640 6352 38704
rect 6368 38640 6432 38704
rect 6448 38640 6512 38704
rect 6528 38640 6592 38704
rect 6608 38640 6672 38704
rect 6688 38640 6752 38704
rect 6768 38640 6832 38704
rect 6848 38640 6912 38704
rect 6928 38640 6992 38704
rect 7008 38640 7072 38704
rect 7088 38640 7152 38704
rect 7168 38640 7232 38704
rect 7248 38640 7312 38704
rect 7328 38640 7392 38704
rect 7408 38640 7472 38704
rect 7488 38640 7552 38704
rect 7568 38640 7632 38704
rect 7648 38640 7712 38704
rect 7728 38640 7792 38704
rect 7808 38640 7872 38704
rect 7888 38640 7952 38704
rect 7968 38640 8032 38704
rect 8048 38640 8112 38704
rect 8128 38640 8192 38704
rect 8208 38640 8272 38704
rect 8288 38640 8352 38704
rect 8368 38640 8432 38704
rect 8448 38640 8512 38704
rect 8528 38640 8592 38704
rect 8608 38640 8672 38704
rect 8688 38640 8752 38704
rect 8768 38640 8832 38704
rect 8848 38640 8912 38704
rect 8928 38640 8992 38704
rect 14112 38640 14176 38704
rect 14192 38640 14256 38704
rect 14272 38640 14336 38704
rect 14352 38640 14416 38704
rect 24112 38640 24176 38704
rect 24192 38640 24256 38704
rect 24272 38640 24336 38704
rect 24352 38640 24416 38704
rect 36376 38640 36440 38704
rect 36456 38640 36520 38704
rect 36536 38640 36600 38704
rect 36616 38640 36680 38704
rect 36696 38640 36760 38704
rect 36776 38640 36840 38704
rect 36856 38640 36920 38704
rect 36936 38640 37000 38704
rect 37016 38640 37080 38704
rect 37096 38640 37160 38704
rect 37176 38640 37240 38704
rect 37256 38640 37320 38704
rect 37336 38640 37400 38704
rect 37416 38640 37480 38704
rect 37496 38640 37560 38704
rect 37576 38640 37640 38704
rect 37656 38640 37720 38704
rect 37736 38640 37800 38704
rect 37816 38640 37880 38704
rect 37896 38640 37960 38704
rect 37976 38640 38040 38704
rect 38056 38640 38120 38704
rect 38136 38640 38200 38704
rect 38216 38640 38280 38704
rect 38296 38640 38360 38704
rect 38376 38640 38440 38704
rect 38456 38640 38520 38704
rect 38536 38640 38600 38704
rect 38616 38640 38680 38704
rect 38696 38640 38760 38704
rect 38776 38640 38840 38704
rect 38856 38640 38920 38704
rect 38936 38640 39000 38704
rect 39016 38640 39080 38704
rect 39096 38640 39160 38704
rect 39176 38640 39240 38704
rect 39256 38640 39320 38704
rect 39336 38640 39400 38704
rect 39416 38640 39480 38704
rect 39496 38640 39560 38704
rect 39576 38640 39640 38704
rect 39656 38640 39720 38704
rect 39736 38640 39800 38704
rect 39816 38640 39880 38704
rect 39896 38640 39960 38704
rect 39976 38640 40040 38704
rect 40056 38640 40120 38704
rect 40136 38640 40200 38704
rect 40216 38640 40280 38704
rect 40296 38640 40360 38704
rect 5008 38560 5072 38624
rect 5088 38560 5152 38624
rect 5168 38560 5232 38624
rect 5248 38560 5312 38624
rect 5328 38560 5392 38624
rect 5408 38560 5472 38624
rect 5488 38560 5552 38624
rect 5568 38560 5632 38624
rect 5648 38560 5712 38624
rect 5728 38560 5792 38624
rect 5808 38560 5872 38624
rect 5888 38560 5952 38624
rect 5968 38560 6032 38624
rect 6048 38560 6112 38624
rect 6128 38560 6192 38624
rect 6208 38560 6272 38624
rect 6288 38560 6352 38624
rect 6368 38560 6432 38624
rect 6448 38560 6512 38624
rect 6528 38560 6592 38624
rect 6608 38560 6672 38624
rect 6688 38560 6752 38624
rect 6768 38560 6832 38624
rect 6848 38560 6912 38624
rect 6928 38560 6992 38624
rect 7008 38560 7072 38624
rect 7088 38560 7152 38624
rect 7168 38560 7232 38624
rect 7248 38560 7312 38624
rect 7328 38560 7392 38624
rect 7408 38560 7472 38624
rect 7488 38560 7552 38624
rect 7568 38560 7632 38624
rect 7648 38560 7712 38624
rect 7728 38560 7792 38624
rect 7808 38560 7872 38624
rect 7888 38560 7952 38624
rect 7968 38560 8032 38624
rect 8048 38560 8112 38624
rect 8128 38560 8192 38624
rect 8208 38560 8272 38624
rect 8288 38560 8352 38624
rect 8368 38560 8432 38624
rect 8448 38560 8512 38624
rect 8528 38560 8592 38624
rect 8608 38560 8672 38624
rect 8688 38560 8752 38624
rect 8768 38560 8832 38624
rect 8848 38560 8912 38624
rect 8928 38560 8992 38624
rect 14112 38560 14176 38624
rect 14192 38560 14256 38624
rect 14272 38560 14336 38624
rect 14352 38560 14416 38624
rect 24112 38560 24176 38624
rect 24192 38560 24256 38624
rect 24272 38560 24336 38624
rect 24352 38560 24416 38624
rect 36376 38560 36440 38624
rect 36456 38560 36520 38624
rect 36536 38560 36600 38624
rect 36616 38560 36680 38624
rect 36696 38560 36760 38624
rect 36776 38560 36840 38624
rect 36856 38560 36920 38624
rect 36936 38560 37000 38624
rect 37016 38560 37080 38624
rect 37096 38560 37160 38624
rect 37176 38560 37240 38624
rect 37256 38560 37320 38624
rect 37336 38560 37400 38624
rect 37416 38560 37480 38624
rect 37496 38560 37560 38624
rect 37576 38560 37640 38624
rect 37656 38560 37720 38624
rect 37736 38560 37800 38624
rect 37816 38560 37880 38624
rect 37896 38560 37960 38624
rect 37976 38560 38040 38624
rect 38056 38560 38120 38624
rect 38136 38560 38200 38624
rect 38216 38560 38280 38624
rect 38296 38560 38360 38624
rect 38376 38560 38440 38624
rect 38456 38560 38520 38624
rect 38536 38560 38600 38624
rect 38616 38560 38680 38624
rect 38696 38560 38760 38624
rect 38776 38560 38840 38624
rect 38856 38560 38920 38624
rect 38936 38560 39000 38624
rect 39016 38560 39080 38624
rect 39096 38560 39160 38624
rect 39176 38560 39240 38624
rect 39256 38560 39320 38624
rect 39336 38560 39400 38624
rect 39416 38560 39480 38624
rect 39496 38560 39560 38624
rect 39576 38560 39640 38624
rect 39656 38560 39720 38624
rect 39736 38560 39800 38624
rect 39816 38560 39880 38624
rect 39896 38560 39960 38624
rect 39976 38560 40040 38624
rect 40056 38560 40120 38624
rect 40136 38560 40200 38624
rect 40216 38560 40280 38624
rect 40296 38560 40360 38624
rect 5008 38480 5072 38544
rect 5088 38480 5152 38544
rect 5168 38480 5232 38544
rect 5248 38480 5312 38544
rect 5328 38480 5392 38544
rect 5408 38480 5472 38544
rect 5488 38480 5552 38544
rect 5568 38480 5632 38544
rect 5648 38480 5712 38544
rect 5728 38480 5792 38544
rect 5808 38480 5872 38544
rect 5888 38480 5952 38544
rect 5968 38480 6032 38544
rect 6048 38480 6112 38544
rect 6128 38480 6192 38544
rect 6208 38480 6272 38544
rect 6288 38480 6352 38544
rect 6368 38480 6432 38544
rect 6448 38480 6512 38544
rect 6528 38480 6592 38544
rect 6608 38480 6672 38544
rect 6688 38480 6752 38544
rect 6768 38480 6832 38544
rect 6848 38480 6912 38544
rect 6928 38480 6992 38544
rect 7008 38480 7072 38544
rect 7088 38480 7152 38544
rect 7168 38480 7232 38544
rect 7248 38480 7312 38544
rect 7328 38480 7392 38544
rect 7408 38480 7472 38544
rect 7488 38480 7552 38544
rect 7568 38480 7632 38544
rect 7648 38480 7712 38544
rect 7728 38480 7792 38544
rect 7808 38480 7872 38544
rect 7888 38480 7952 38544
rect 7968 38480 8032 38544
rect 8048 38480 8112 38544
rect 8128 38480 8192 38544
rect 8208 38480 8272 38544
rect 8288 38480 8352 38544
rect 8368 38480 8432 38544
rect 8448 38480 8512 38544
rect 8528 38480 8592 38544
rect 8608 38480 8672 38544
rect 8688 38480 8752 38544
rect 8768 38480 8832 38544
rect 8848 38480 8912 38544
rect 8928 38480 8992 38544
rect 14112 38480 14176 38544
rect 14192 38480 14256 38544
rect 14272 38480 14336 38544
rect 14352 38480 14416 38544
rect 24112 38480 24176 38544
rect 24192 38480 24256 38544
rect 24272 38480 24336 38544
rect 24352 38480 24416 38544
rect 36376 38480 36440 38544
rect 36456 38480 36520 38544
rect 36536 38480 36600 38544
rect 36616 38480 36680 38544
rect 36696 38480 36760 38544
rect 36776 38480 36840 38544
rect 36856 38480 36920 38544
rect 36936 38480 37000 38544
rect 37016 38480 37080 38544
rect 37096 38480 37160 38544
rect 37176 38480 37240 38544
rect 37256 38480 37320 38544
rect 37336 38480 37400 38544
rect 37416 38480 37480 38544
rect 37496 38480 37560 38544
rect 37576 38480 37640 38544
rect 37656 38480 37720 38544
rect 37736 38480 37800 38544
rect 37816 38480 37880 38544
rect 37896 38480 37960 38544
rect 37976 38480 38040 38544
rect 38056 38480 38120 38544
rect 38136 38480 38200 38544
rect 38216 38480 38280 38544
rect 38296 38480 38360 38544
rect 38376 38480 38440 38544
rect 38456 38480 38520 38544
rect 38536 38480 38600 38544
rect 38616 38480 38680 38544
rect 38696 38480 38760 38544
rect 38776 38480 38840 38544
rect 38856 38480 38920 38544
rect 38936 38480 39000 38544
rect 39016 38480 39080 38544
rect 39096 38480 39160 38544
rect 39176 38480 39240 38544
rect 39256 38480 39320 38544
rect 39336 38480 39400 38544
rect 39416 38480 39480 38544
rect 39496 38480 39560 38544
rect 39576 38480 39640 38544
rect 39656 38480 39720 38544
rect 39736 38480 39800 38544
rect 39816 38480 39880 38544
rect 39896 38480 39960 38544
rect 39976 38480 40040 38544
rect 40056 38480 40120 38544
rect 40136 38480 40200 38544
rect 40216 38480 40280 38544
rect 40296 38480 40360 38544
rect 5008 38400 5072 38464
rect 5088 38400 5152 38464
rect 5168 38400 5232 38464
rect 5248 38400 5312 38464
rect 5328 38400 5392 38464
rect 5408 38400 5472 38464
rect 5488 38400 5552 38464
rect 5568 38400 5632 38464
rect 5648 38400 5712 38464
rect 5728 38400 5792 38464
rect 5808 38400 5872 38464
rect 5888 38400 5952 38464
rect 5968 38400 6032 38464
rect 6048 38400 6112 38464
rect 6128 38400 6192 38464
rect 6208 38400 6272 38464
rect 6288 38400 6352 38464
rect 6368 38400 6432 38464
rect 6448 38400 6512 38464
rect 6528 38400 6592 38464
rect 6608 38400 6672 38464
rect 6688 38400 6752 38464
rect 6768 38400 6832 38464
rect 6848 38400 6912 38464
rect 6928 38400 6992 38464
rect 7008 38400 7072 38464
rect 7088 38400 7152 38464
rect 7168 38400 7232 38464
rect 7248 38400 7312 38464
rect 7328 38400 7392 38464
rect 7408 38400 7472 38464
rect 7488 38400 7552 38464
rect 7568 38400 7632 38464
rect 7648 38400 7712 38464
rect 7728 38400 7792 38464
rect 7808 38400 7872 38464
rect 7888 38400 7952 38464
rect 7968 38400 8032 38464
rect 8048 38400 8112 38464
rect 8128 38400 8192 38464
rect 8208 38400 8272 38464
rect 8288 38400 8352 38464
rect 8368 38400 8432 38464
rect 8448 38400 8512 38464
rect 8528 38400 8592 38464
rect 8608 38400 8672 38464
rect 8688 38400 8752 38464
rect 8768 38400 8832 38464
rect 8848 38400 8912 38464
rect 8928 38400 8992 38464
rect 14112 38400 14176 38464
rect 14192 38400 14256 38464
rect 14272 38400 14336 38464
rect 14352 38400 14416 38464
rect 24112 38400 24176 38464
rect 24192 38400 24256 38464
rect 24272 38400 24336 38464
rect 24352 38400 24416 38464
rect 36376 38400 36440 38464
rect 36456 38400 36520 38464
rect 36536 38400 36600 38464
rect 36616 38400 36680 38464
rect 36696 38400 36760 38464
rect 36776 38400 36840 38464
rect 36856 38400 36920 38464
rect 36936 38400 37000 38464
rect 37016 38400 37080 38464
rect 37096 38400 37160 38464
rect 37176 38400 37240 38464
rect 37256 38400 37320 38464
rect 37336 38400 37400 38464
rect 37416 38400 37480 38464
rect 37496 38400 37560 38464
rect 37576 38400 37640 38464
rect 37656 38400 37720 38464
rect 37736 38400 37800 38464
rect 37816 38400 37880 38464
rect 37896 38400 37960 38464
rect 37976 38400 38040 38464
rect 38056 38400 38120 38464
rect 38136 38400 38200 38464
rect 38216 38400 38280 38464
rect 38296 38400 38360 38464
rect 38376 38400 38440 38464
rect 38456 38400 38520 38464
rect 38536 38400 38600 38464
rect 38616 38400 38680 38464
rect 38696 38400 38760 38464
rect 38776 38400 38840 38464
rect 38856 38400 38920 38464
rect 38936 38400 39000 38464
rect 39016 38400 39080 38464
rect 39096 38400 39160 38464
rect 39176 38400 39240 38464
rect 39256 38400 39320 38464
rect 39336 38400 39400 38464
rect 39416 38400 39480 38464
rect 39496 38400 39560 38464
rect 39576 38400 39640 38464
rect 39656 38400 39720 38464
rect 39736 38400 39800 38464
rect 39816 38400 39880 38464
rect 39896 38400 39960 38464
rect 39976 38400 40040 38464
rect 40056 38400 40120 38464
rect 40136 38400 40200 38464
rect 40216 38400 40280 38464
rect 40296 38400 40360 38464
rect 5008 38320 5072 38384
rect 5088 38320 5152 38384
rect 5168 38320 5232 38384
rect 5248 38320 5312 38384
rect 5328 38320 5392 38384
rect 5408 38320 5472 38384
rect 5488 38320 5552 38384
rect 5568 38320 5632 38384
rect 5648 38320 5712 38384
rect 5728 38320 5792 38384
rect 5808 38320 5872 38384
rect 5888 38320 5952 38384
rect 5968 38320 6032 38384
rect 6048 38320 6112 38384
rect 6128 38320 6192 38384
rect 6208 38320 6272 38384
rect 6288 38320 6352 38384
rect 6368 38320 6432 38384
rect 6448 38320 6512 38384
rect 6528 38320 6592 38384
rect 6608 38320 6672 38384
rect 6688 38320 6752 38384
rect 6768 38320 6832 38384
rect 6848 38320 6912 38384
rect 6928 38320 6992 38384
rect 7008 38320 7072 38384
rect 7088 38320 7152 38384
rect 7168 38320 7232 38384
rect 7248 38320 7312 38384
rect 7328 38320 7392 38384
rect 7408 38320 7472 38384
rect 7488 38320 7552 38384
rect 7568 38320 7632 38384
rect 7648 38320 7712 38384
rect 7728 38320 7792 38384
rect 7808 38320 7872 38384
rect 7888 38320 7952 38384
rect 7968 38320 8032 38384
rect 8048 38320 8112 38384
rect 8128 38320 8192 38384
rect 8208 38320 8272 38384
rect 8288 38320 8352 38384
rect 8368 38320 8432 38384
rect 8448 38320 8512 38384
rect 8528 38320 8592 38384
rect 8608 38320 8672 38384
rect 8688 38320 8752 38384
rect 8768 38320 8832 38384
rect 8848 38320 8912 38384
rect 8928 38320 8992 38384
rect 14112 38320 14176 38384
rect 14192 38320 14256 38384
rect 14272 38320 14336 38384
rect 14352 38320 14416 38384
rect 24112 38320 24176 38384
rect 24192 38320 24256 38384
rect 24272 38320 24336 38384
rect 24352 38320 24416 38384
rect 36376 38320 36440 38384
rect 36456 38320 36520 38384
rect 36536 38320 36600 38384
rect 36616 38320 36680 38384
rect 36696 38320 36760 38384
rect 36776 38320 36840 38384
rect 36856 38320 36920 38384
rect 36936 38320 37000 38384
rect 37016 38320 37080 38384
rect 37096 38320 37160 38384
rect 37176 38320 37240 38384
rect 37256 38320 37320 38384
rect 37336 38320 37400 38384
rect 37416 38320 37480 38384
rect 37496 38320 37560 38384
rect 37576 38320 37640 38384
rect 37656 38320 37720 38384
rect 37736 38320 37800 38384
rect 37816 38320 37880 38384
rect 37896 38320 37960 38384
rect 37976 38320 38040 38384
rect 38056 38320 38120 38384
rect 38136 38320 38200 38384
rect 38216 38320 38280 38384
rect 38296 38320 38360 38384
rect 38376 38320 38440 38384
rect 38456 38320 38520 38384
rect 38536 38320 38600 38384
rect 38616 38320 38680 38384
rect 38696 38320 38760 38384
rect 38776 38320 38840 38384
rect 38856 38320 38920 38384
rect 38936 38320 39000 38384
rect 39016 38320 39080 38384
rect 39096 38320 39160 38384
rect 39176 38320 39240 38384
rect 39256 38320 39320 38384
rect 39336 38320 39400 38384
rect 39416 38320 39480 38384
rect 39496 38320 39560 38384
rect 39576 38320 39640 38384
rect 39656 38320 39720 38384
rect 39736 38320 39800 38384
rect 39816 38320 39880 38384
rect 39896 38320 39960 38384
rect 39976 38320 40040 38384
rect 40056 38320 40120 38384
rect 40136 38320 40200 38384
rect 40216 38320 40280 38384
rect 40296 38320 40360 38384
rect 5008 38240 5072 38304
rect 5088 38240 5152 38304
rect 5168 38240 5232 38304
rect 5248 38240 5312 38304
rect 5328 38240 5392 38304
rect 5408 38240 5472 38304
rect 5488 38240 5552 38304
rect 5568 38240 5632 38304
rect 5648 38240 5712 38304
rect 5728 38240 5792 38304
rect 5808 38240 5872 38304
rect 5888 38240 5952 38304
rect 5968 38240 6032 38304
rect 6048 38240 6112 38304
rect 6128 38240 6192 38304
rect 6208 38240 6272 38304
rect 6288 38240 6352 38304
rect 6368 38240 6432 38304
rect 6448 38240 6512 38304
rect 6528 38240 6592 38304
rect 6608 38240 6672 38304
rect 6688 38240 6752 38304
rect 6768 38240 6832 38304
rect 6848 38240 6912 38304
rect 6928 38240 6992 38304
rect 7008 38240 7072 38304
rect 7088 38240 7152 38304
rect 7168 38240 7232 38304
rect 7248 38240 7312 38304
rect 7328 38240 7392 38304
rect 7408 38240 7472 38304
rect 7488 38240 7552 38304
rect 7568 38240 7632 38304
rect 7648 38240 7712 38304
rect 7728 38240 7792 38304
rect 7808 38240 7872 38304
rect 7888 38240 7952 38304
rect 7968 38240 8032 38304
rect 8048 38240 8112 38304
rect 8128 38240 8192 38304
rect 8208 38240 8272 38304
rect 8288 38240 8352 38304
rect 8368 38240 8432 38304
rect 8448 38240 8512 38304
rect 8528 38240 8592 38304
rect 8608 38240 8672 38304
rect 8688 38240 8752 38304
rect 8768 38240 8832 38304
rect 8848 38240 8912 38304
rect 8928 38240 8992 38304
rect 14112 38240 14176 38304
rect 14192 38240 14256 38304
rect 14272 38240 14336 38304
rect 14352 38240 14416 38304
rect 24112 38240 24176 38304
rect 24192 38240 24256 38304
rect 24272 38240 24336 38304
rect 24352 38240 24416 38304
rect 36376 38240 36440 38304
rect 36456 38240 36520 38304
rect 36536 38240 36600 38304
rect 36616 38240 36680 38304
rect 36696 38240 36760 38304
rect 36776 38240 36840 38304
rect 36856 38240 36920 38304
rect 36936 38240 37000 38304
rect 37016 38240 37080 38304
rect 37096 38240 37160 38304
rect 37176 38240 37240 38304
rect 37256 38240 37320 38304
rect 37336 38240 37400 38304
rect 37416 38240 37480 38304
rect 37496 38240 37560 38304
rect 37576 38240 37640 38304
rect 37656 38240 37720 38304
rect 37736 38240 37800 38304
rect 37816 38240 37880 38304
rect 37896 38240 37960 38304
rect 37976 38240 38040 38304
rect 38056 38240 38120 38304
rect 38136 38240 38200 38304
rect 38216 38240 38280 38304
rect 38296 38240 38360 38304
rect 38376 38240 38440 38304
rect 38456 38240 38520 38304
rect 38536 38240 38600 38304
rect 38616 38240 38680 38304
rect 38696 38240 38760 38304
rect 38776 38240 38840 38304
rect 38856 38240 38920 38304
rect 38936 38240 39000 38304
rect 39016 38240 39080 38304
rect 39096 38240 39160 38304
rect 39176 38240 39240 38304
rect 39256 38240 39320 38304
rect 39336 38240 39400 38304
rect 39416 38240 39480 38304
rect 39496 38240 39560 38304
rect 39576 38240 39640 38304
rect 39656 38240 39720 38304
rect 39736 38240 39800 38304
rect 39816 38240 39880 38304
rect 39896 38240 39960 38304
rect 39976 38240 40040 38304
rect 40056 38240 40120 38304
rect 40136 38240 40200 38304
rect 40216 38240 40280 38304
rect 40296 38240 40360 38304
rect 5008 38160 5072 38224
rect 5088 38160 5152 38224
rect 5168 38160 5232 38224
rect 5248 38160 5312 38224
rect 5328 38160 5392 38224
rect 5408 38160 5472 38224
rect 5488 38160 5552 38224
rect 5568 38160 5632 38224
rect 5648 38160 5712 38224
rect 5728 38160 5792 38224
rect 5808 38160 5872 38224
rect 5888 38160 5952 38224
rect 5968 38160 6032 38224
rect 6048 38160 6112 38224
rect 6128 38160 6192 38224
rect 6208 38160 6272 38224
rect 6288 38160 6352 38224
rect 6368 38160 6432 38224
rect 6448 38160 6512 38224
rect 6528 38160 6592 38224
rect 6608 38160 6672 38224
rect 6688 38160 6752 38224
rect 6768 38160 6832 38224
rect 6848 38160 6912 38224
rect 6928 38160 6992 38224
rect 7008 38160 7072 38224
rect 7088 38160 7152 38224
rect 7168 38160 7232 38224
rect 7248 38160 7312 38224
rect 7328 38160 7392 38224
rect 7408 38160 7472 38224
rect 7488 38160 7552 38224
rect 7568 38160 7632 38224
rect 7648 38160 7712 38224
rect 7728 38160 7792 38224
rect 7808 38160 7872 38224
rect 7888 38160 7952 38224
rect 7968 38160 8032 38224
rect 8048 38160 8112 38224
rect 8128 38160 8192 38224
rect 8208 38160 8272 38224
rect 8288 38160 8352 38224
rect 8368 38160 8432 38224
rect 8448 38160 8512 38224
rect 8528 38160 8592 38224
rect 8608 38160 8672 38224
rect 8688 38160 8752 38224
rect 8768 38160 8832 38224
rect 8848 38160 8912 38224
rect 8928 38160 8992 38224
rect 14112 38160 14176 38224
rect 14192 38160 14256 38224
rect 14272 38160 14336 38224
rect 14352 38160 14416 38224
rect 24112 38160 24176 38224
rect 24192 38160 24256 38224
rect 24272 38160 24336 38224
rect 24352 38160 24416 38224
rect 36376 38160 36440 38224
rect 36456 38160 36520 38224
rect 36536 38160 36600 38224
rect 36616 38160 36680 38224
rect 36696 38160 36760 38224
rect 36776 38160 36840 38224
rect 36856 38160 36920 38224
rect 36936 38160 37000 38224
rect 37016 38160 37080 38224
rect 37096 38160 37160 38224
rect 37176 38160 37240 38224
rect 37256 38160 37320 38224
rect 37336 38160 37400 38224
rect 37416 38160 37480 38224
rect 37496 38160 37560 38224
rect 37576 38160 37640 38224
rect 37656 38160 37720 38224
rect 37736 38160 37800 38224
rect 37816 38160 37880 38224
rect 37896 38160 37960 38224
rect 37976 38160 38040 38224
rect 38056 38160 38120 38224
rect 38136 38160 38200 38224
rect 38216 38160 38280 38224
rect 38296 38160 38360 38224
rect 38376 38160 38440 38224
rect 38456 38160 38520 38224
rect 38536 38160 38600 38224
rect 38616 38160 38680 38224
rect 38696 38160 38760 38224
rect 38776 38160 38840 38224
rect 38856 38160 38920 38224
rect 38936 38160 39000 38224
rect 39016 38160 39080 38224
rect 39096 38160 39160 38224
rect 39176 38160 39240 38224
rect 39256 38160 39320 38224
rect 39336 38160 39400 38224
rect 39416 38160 39480 38224
rect 39496 38160 39560 38224
rect 39576 38160 39640 38224
rect 39656 38160 39720 38224
rect 39736 38160 39800 38224
rect 39816 38160 39880 38224
rect 39896 38160 39960 38224
rect 39976 38160 40040 38224
rect 40056 38160 40120 38224
rect 40136 38160 40200 38224
rect 40216 38160 40280 38224
rect 40296 38160 40360 38224
rect 5008 38080 5072 38144
rect 5088 38080 5152 38144
rect 5168 38080 5232 38144
rect 5248 38080 5312 38144
rect 5328 38080 5392 38144
rect 5408 38080 5472 38144
rect 5488 38080 5552 38144
rect 5568 38080 5632 38144
rect 5648 38080 5712 38144
rect 5728 38080 5792 38144
rect 5808 38080 5872 38144
rect 5888 38080 5952 38144
rect 5968 38080 6032 38144
rect 6048 38080 6112 38144
rect 6128 38080 6192 38144
rect 6208 38080 6272 38144
rect 6288 38080 6352 38144
rect 6368 38080 6432 38144
rect 6448 38080 6512 38144
rect 6528 38080 6592 38144
rect 6608 38080 6672 38144
rect 6688 38080 6752 38144
rect 6768 38080 6832 38144
rect 6848 38080 6912 38144
rect 6928 38080 6992 38144
rect 7008 38080 7072 38144
rect 7088 38080 7152 38144
rect 7168 38080 7232 38144
rect 7248 38080 7312 38144
rect 7328 38080 7392 38144
rect 7408 38080 7472 38144
rect 7488 38080 7552 38144
rect 7568 38080 7632 38144
rect 7648 38080 7712 38144
rect 7728 38080 7792 38144
rect 7808 38080 7872 38144
rect 7888 38080 7952 38144
rect 7968 38080 8032 38144
rect 8048 38080 8112 38144
rect 8128 38080 8192 38144
rect 8208 38080 8272 38144
rect 8288 38080 8352 38144
rect 8368 38080 8432 38144
rect 8448 38080 8512 38144
rect 8528 38080 8592 38144
rect 8608 38080 8672 38144
rect 8688 38080 8752 38144
rect 8768 38080 8832 38144
rect 8848 38080 8912 38144
rect 8928 38080 8992 38144
rect 14112 38080 14176 38144
rect 14192 38080 14256 38144
rect 14272 38080 14336 38144
rect 14352 38080 14416 38144
rect 24112 38080 24176 38144
rect 24192 38080 24256 38144
rect 24272 38080 24336 38144
rect 24352 38080 24416 38144
rect 36376 38080 36440 38144
rect 36456 38080 36520 38144
rect 36536 38080 36600 38144
rect 36616 38080 36680 38144
rect 36696 38080 36760 38144
rect 36776 38080 36840 38144
rect 36856 38080 36920 38144
rect 36936 38080 37000 38144
rect 37016 38080 37080 38144
rect 37096 38080 37160 38144
rect 37176 38080 37240 38144
rect 37256 38080 37320 38144
rect 37336 38080 37400 38144
rect 37416 38080 37480 38144
rect 37496 38080 37560 38144
rect 37576 38080 37640 38144
rect 37656 38080 37720 38144
rect 37736 38080 37800 38144
rect 37816 38080 37880 38144
rect 37896 38080 37960 38144
rect 37976 38080 38040 38144
rect 38056 38080 38120 38144
rect 38136 38080 38200 38144
rect 38216 38080 38280 38144
rect 38296 38080 38360 38144
rect 38376 38080 38440 38144
rect 38456 38080 38520 38144
rect 38536 38080 38600 38144
rect 38616 38080 38680 38144
rect 38696 38080 38760 38144
rect 38776 38080 38840 38144
rect 38856 38080 38920 38144
rect 38936 38080 39000 38144
rect 39016 38080 39080 38144
rect 39096 38080 39160 38144
rect 39176 38080 39240 38144
rect 39256 38080 39320 38144
rect 39336 38080 39400 38144
rect 39416 38080 39480 38144
rect 39496 38080 39560 38144
rect 39576 38080 39640 38144
rect 39656 38080 39720 38144
rect 39736 38080 39800 38144
rect 39816 38080 39880 38144
rect 39896 38080 39960 38144
rect 39976 38080 40040 38144
rect 40056 38080 40120 38144
rect 40136 38080 40200 38144
rect 40216 38080 40280 38144
rect 40296 38080 40360 38144
rect 5008 38000 5072 38064
rect 5088 38000 5152 38064
rect 5168 38000 5232 38064
rect 5248 38000 5312 38064
rect 5328 38000 5392 38064
rect 5408 38000 5472 38064
rect 5488 38000 5552 38064
rect 5568 38000 5632 38064
rect 5648 38000 5712 38064
rect 5728 38000 5792 38064
rect 5808 38000 5872 38064
rect 5888 38000 5952 38064
rect 5968 38000 6032 38064
rect 6048 38000 6112 38064
rect 6128 38000 6192 38064
rect 6208 38000 6272 38064
rect 6288 38000 6352 38064
rect 6368 38000 6432 38064
rect 6448 38000 6512 38064
rect 6528 38000 6592 38064
rect 6608 38000 6672 38064
rect 6688 38000 6752 38064
rect 6768 38000 6832 38064
rect 6848 38000 6912 38064
rect 6928 38000 6992 38064
rect 7008 38000 7072 38064
rect 7088 38000 7152 38064
rect 7168 38000 7232 38064
rect 7248 38000 7312 38064
rect 7328 38000 7392 38064
rect 7408 38000 7472 38064
rect 7488 38000 7552 38064
rect 7568 38000 7632 38064
rect 7648 38000 7712 38064
rect 7728 38000 7792 38064
rect 7808 38000 7872 38064
rect 7888 38000 7952 38064
rect 7968 38000 8032 38064
rect 8048 38000 8112 38064
rect 8128 38000 8192 38064
rect 8208 38000 8272 38064
rect 8288 38000 8352 38064
rect 8368 38000 8432 38064
rect 8448 38000 8512 38064
rect 8528 38000 8592 38064
rect 8608 38000 8672 38064
rect 8688 38000 8752 38064
rect 8768 38000 8832 38064
rect 8848 38000 8912 38064
rect 8928 38000 8992 38064
rect 14112 38000 14176 38064
rect 14192 38000 14256 38064
rect 14272 38000 14336 38064
rect 14352 38000 14416 38064
rect 24112 38000 24176 38064
rect 24192 38000 24256 38064
rect 24272 38000 24336 38064
rect 24352 38000 24416 38064
rect 36376 38000 36440 38064
rect 36456 38000 36520 38064
rect 36536 38000 36600 38064
rect 36616 38000 36680 38064
rect 36696 38000 36760 38064
rect 36776 38000 36840 38064
rect 36856 38000 36920 38064
rect 36936 38000 37000 38064
rect 37016 38000 37080 38064
rect 37096 38000 37160 38064
rect 37176 38000 37240 38064
rect 37256 38000 37320 38064
rect 37336 38000 37400 38064
rect 37416 38000 37480 38064
rect 37496 38000 37560 38064
rect 37576 38000 37640 38064
rect 37656 38000 37720 38064
rect 37736 38000 37800 38064
rect 37816 38000 37880 38064
rect 37896 38000 37960 38064
rect 37976 38000 38040 38064
rect 38056 38000 38120 38064
rect 38136 38000 38200 38064
rect 38216 38000 38280 38064
rect 38296 38000 38360 38064
rect 38376 38000 38440 38064
rect 38456 38000 38520 38064
rect 38536 38000 38600 38064
rect 38616 38000 38680 38064
rect 38696 38000 38760 38064
rect 38776 38000 38840 38064
rect 38856 38000 38920 38064
rect 38936 38000 39000 38064
rect 39016 38000 39080 38064
rect 39096 38000 39160 38064
rect 39176 38000 39240 38064
rect 39256 38000 39320 38064
rect 39336 38000 39400 38064
rect 39416 38000 39480 38064
rect 39496 38000 39560 38064
rect 39576 38000 39640 38064
rect 39656 38000 39720 38064
rect 39736 38000 39800 38064
rect 39816 38000 39880 38064
rect 39896 38000 39960 38064
rect 39976 38000 40040 38064
rect 40056 38000 40120 38064
rect 40136 38000 40200 38064
rect 40216 38000 40280 38064
rect 40296 38000 40360 38064
rect 5008 37920 5072 37984
rect 5088 37920 5152 37984
rect 5168 37920 5232 37984
rect 5248 37920 5312 37984
rect 5328 37920 5392 37984
rect 5408 37920 5472 37984
rect 5488 37920 5552 37984
rect 5568 37920 5632 37984
rect 5648 37920 5712 37984
rect 5728 37920 5792 37984
rect 5808 37920 5872 37984
rect 5888 37920 5952 37984
rect 5968 37920 6032 37984
rect 6048 37920 6112 37984
rect 6128 37920 6192 37984
rect 6208 37920 6272 37984
rect 6288 37920 6352 37984
rect 6368 37920 6432 37984
rect 6448 37920 6512 37984
rect 6528 37920 6592 37984
rect 6608 37920 6672 37984
rect 6688 37920 6752 37984
rect 6768 37920 6832 37984
rect 6848 37920 6912 37984
rect 6928 37920 6992 37984
rect 7008 37920 7072 37984
rect 7088 37920 7152 37984
rect 7168 37920 7232 37984
rect 7248 37920 7312 37984
rect 7328 37920 7392 37984
rect 7408 37920 7472 37984
rect 7488 37920 7552 37984
rect 7568 37920 7632 37984
rect 7648 37920 7712 37984
rect 7728 37920 7792 37984
rect 7808 37920 7872 37984
rect 7888 37920 7952 37984
rect 7968 37920 8032 37984
rect 8048 37920 8112 37984
rect 8128 37920 8192 37984
rect 8208 37920 8272 37984
rect 8288 37920 8352 37984
rect 8368 37920 8432 37984
rect 8448 37920 8512 37984
rect 8528 37920 8592 37984
rect 8608 37920 8672 37984
rect 8688 37920 8752 37984
rect 8768 37920 8832 37984
rect 8848 37920 8912 37984
rect 8928 37920 8992 37984
rect 14112 37920 14176 37984
rect 14192 37920 14256 37984
rect 14272 37920 14336 37984
rect 14352 37920 14416 37984
rect 24112 37920 24176 37984
rect 24192 37920 24256 37984
rect 24272 37920 24336 37984
rect 24352 37920 24416 37984
rect 36376 37920 36440 37984
rect 36456 37920 36520 37984
rect 36536 37920 36600 37984
rect 36616 37920 36680 37984
rect 36696 37920 36760 37984
rect 36776 37920 36840 37984
rect 36856 37920 36920 37984
rect 36936 37920 37000 37984
rect 37016 37920 37080 37984
rect 37096 37920 37160 37984
rect 37176 37920 37240 37984
rect 37256 37920 37320 37984
rect 37336 37920 37400 37984
rect 37416 37920 37480 37984
rect 37496 37920 37560 37984
rect 37576 37920 37640 37984
rect 37656 37920 37720 37984
rect 37736 37920 37800 37984
rect 37816 37920 37880 37984
rect 37896 37920 37960 37984
rect 37976 37920 38040 37984
rect 38056 37920 38120 37984
rect 38136 37920 38200 37984
rect 38216 37920 38280 37984
rect 38296 37920 38360 37984
rect 38376 37920 38440 37984
rect 38456 37920 38520 37984
rect 38536 37920 38600 37984
rect 38616 37920 38680 37984
rect 38696 37920 38760 37984
rect 38776 37920 38840 37984
rect 38856 37920 38920 37984
rect 38936 37920 39000 37984
rect 39016 37920 39080 37984
rect 39096 37920 39160 37984
rect 39176 37920 39240 37984
rect 39256 37920 39320 37984
rect 39336 37920 39400 37984
rect 39416 37920 39480 37984
rect 39496 37920 39560 37984
rect 39576 37920 39640 37984
rect 39656 37920 39720 37984
rect 39736 37920 39800 37984
rect 39816 37920 39880 37984
rect 39896 37920 39960 37984
rect 39976 37920 40040 37984
rect 40056 37920 40120 37984
rect 40136 37920 40200 37984
rect 40216 37920 40280 37984
rect 40296 37920 40360 37984
rect 5008 37840 5072 37904
rect 5088 37840 5152 37904
rect 5168 37840 5232 37904
rect 5248 37840 5312 37904
rect 5328 37840 5392 37904
rect 5408 37840 5472 37904
rect 5488 37840 5552 37904
rect 5568 37840 5632 37904
rect 5648 37840 5712 37904
rect 5728 37840 5792 37904
rect 5808 37840 5872 37904
rect 5888 37840 5952 37904
rect 5968 37840 6032 37904
rect 6048 37840 6112 37904
rect 6128 37840 6192 37904
rect 6208 37840 6272 37904
rect 6288 37840 6352 37904
rect 6368 37840 6432 37904
rect 6448 37840 6512 37904
rect 6528 37840 6592 37904
rect 6608 37840 6672 37904
rect 6688 37840 6752 37904
rect 6768 37840 6832 37904
rect 6848 37840 6912 37904
rect 6928 37840 6992 37904
rect 7008 37840 7072 37904
rect 7088 37840 7152 37904
rect 7168 37840 7232 37904
rect 7248 37840 7312 37904
rect 7328 37840 7392 37904
rect 7408 37840 7472 37904
rect 7488 37840 7552 37904
rect 7568 37840 7632 37904
rect 7648 37840 7712 37904
rect 7728 37840 7792 37904
rect 7808 37840 7872 37904
rect 7888 37840 7952 37904
rect 7968 37840 8032 37904
rect 8048 37840 8112 37904
rect 8128 37840 8192 37904
rect 8208 37840 8272 37904
rect 8288 37840 8352 37904
rect 8368 37840 8432 37904
rect 8448 37840 8512 37904
rect 8528 37840 8592 37904
rect 8608 37840 8672 37904
rect 8688 37840 8752 37904
rect 8768 37840 8832 37904
rect 8848 37840 8912 37904
rect 8928 37840 8992 37904
rect 14112 37840 14176 37904
rect 14192 37840 14256 37904
rect 14272 37840 14336 37904
rect 14352 37840 14416 37904
rect 24112 37840 24176 37904
rect 24192 37840 24256 37904
rect 24272 37840 24336 37904
rect 24352 37840 24416 37904
rect 36376 37840 36440 37904
rect 36456 37840 36520 37904
rect 36536 37840 36600 37904
rect 36616 37840 36680 37904
rect 36696 37840 36760 37904
rect 36776 37840 36840 37904
rect 36856 37840 36920 37904
rect 36936 37840 37000 37904
rect 37016 37840 37080 37904
rect 37096 37840 37160 37904
rect 37176 37840 37240 37904
rect 37256 37840 37320 37904
rect 37336 37840 37400 37904
rect 37416 37840 37480 37904
rect 37496 37840 37560 37904
rect 37576 37840 37640 37904
rect 37656 37840 37720 37904
rect 37736 37840 37800 37904
rect 37816 37840 37880 37904
rect 37896 37840 37960 37904
rect 37976 37840 38040 37904
rect 38056 37840 38120 37904
rect 38136 37840 38200 37904
rect 38216 37840 38280 37904
rect 38296 37840 38360 37904
rect 38376 37840 38440 37904
rect 38456 37840 38520 37904
rect 38536 37840 38600 37904
rect 38616 37840 38680 37904
rect 38696 37840 38760 37904
rect 38776 37840 38840 37904
rect 38856 37840 38920 37904
rect 38936 37840 39000 37904
rect 39016 37840 39080 37904
rect 39096 37840 39160 37904
rect 39176 37840 39240 37904
rect 39256 37840 39320 37904
rect 39336 37840 39400 37904
rect 39416 37840 39480 37904
rect 39496 37840 39560 37904
rect 39576 37840 39640 37904
rect 39656 37840 39720 37904
rect 39736 37840 39800 37904
rect 39816 37840 39880 37904
rect 39896 37840 39960 37904
rect 39976 37840 40040 37904
rect 40056 37840 40120 37904
rect 40136 37840 40200 37904
rect 40216 37840 40280 37904
rect 40296 37840 40360 37904
rect 5008 37760 5072 37824
rect 5088 37760 5152 37824
rect 5168 37760 5232 37824
rect 5248 37760 5312 37824
rect 5328 37760 5392 37824
rect 5408 37760 5472 37824
rect 5488 37760 5552 37824
rect 5568 37760 5632 37824
rect 5648 37760 5712 37824
rect 5728 37760 5792 37824
rect 5808 37760 5872 37824
rect 5888 37760 5952 37824
rect 5968 37760 6032 37824
rect 6048 37760 6112 37824
rect 6128 37760 6192 37824
rect 6208 37760 6272 37824
rect 6288 37760 6352 37824
rect 6368 37760 6432 37824
rect 6448 37760 6512 37824
rect 6528 37760 6592 37824
rect 6608 37760 6672 37824
rect 6688 37760 6752 37824
rect 6768 37760 6832 37824
rect 6848 37760 6912 37824
rect 6928 37760 6992 37824
rect 7008 37760 7072 37824
rect 7088 37760 7152 37824
rect 7168 37760 7232 37824
rect 7248 37760 7312 37824
rect 7328 37760 7392 37824
rect 7408 37760 7472 37824
rect 7488 37760 7552 37824
rect 7568 37760 7632 37824
rect 7648 37760 7712 37824
rect 7728 37760 7792 37824
rect 7808 37760 7872 37824
rect 7888 37760 7952 37824
rect 7968 37760 8032 37824
rect 8048 37760 8112 37824
rect 8128 37760 8192 37824
rect 8208 37760 8272 37824
rect 8288 37760 8352 37824
rect 8368 37760 8432 37824
rect 8448 37760 8512 37824
rect 8528 37760 8592 37824
rect 8608 37760 8672 37824
rect 8688 37760 8752 37824
rect 8768 37760 8832 37824
rect 8848 37760 8912 37824
rect 8928 37760 8992 37824
rect 14112 37760 14176 37824
rect 14192 37760 14256 37824
rect 14272 37760 14336 37824
rect 14352 37760 14416 37824
rect 24112 37760 24176 37824
rect 24192 37760 24256 37824
rect 24272 37760 24336 37824
rect 24352 37760 24416 37824
rect 36376 37760 36440 37824
rect 36456 37760 36520 37824
rect 36536 37760 36600 37824
rect 36616 37760 36680 37824
rect 36696 37760 36760 37824
rect 36776 37760 36840 37824
rect 36856 37760 36920 37824
rect 36936 37760 37000 37824
rect 37016 37760 37080 37824
rect 37096 37760 37160 37824
rect 37176 37760 37240 37824
rect 37256 37760 37320 37824
rect 37336 37760 37400 37824
rect 37416 37760 37480 37824
rect 37496 37760 37560 37824
rect 37576 37760 37640 37824
rect 37656 37760 37720 37824
rect 37736 37760 37800 37824
rect 37816 37760 37880 37824
rect 37896 37760 37960 37824
rect 37976 37760 38040 37824
rect 38056 37760 38120 37824
rect 38136 37760 38200 37824
rect 38216 37760 38280 37824
rect 38296 37760 38360 37824
rect 38376 37760 38440 37824
rect 38456 37760 38520 37824
rect 38536 37760 38600 37824
rect 38616 37760 38680 37824
rect 38696 37760 38760 37824
rect 38776 37760 38840 37824
rect 38856 37760 38920 37824
rect 38936 37760 39000 37824
rect 39016 37760 39080 37824
rect 39096 37760 39160 37824
rect 39176 37760 39240 37824
rect 39256 37760 39320 37824
rect 39336 37760 39400 37824
rect 39416 37760 39480 37824
rect 39496 37760 39560 37824
rect 39576 37760 39640 37824
rect 39656 37760 39720 37824
rect 39736 37760 39800 37824
rect 39816 37760 39880 37824
rect 39896 37760 39960 37824
rect 39976 37760 40040 37824
rect 40056 37760 40120 37824
rect 40136 37760 40200 37824
rect 40216 37760 40280 37824
rect 40296 37760 40360 37824
rect 5008 37680 5072 37744
rect 5088 37680 5152 37744
rect 5168 37680 5232 37744
rect 5248 37680 5312 37744
rect 5328 37680 5392 37744
rect 5408 37680 5472 37744
rect 5488 37680 5552 37744
rect 5568 37680 5632 37744
rect 5648 37680 5712 37744
rect 5728 37680 5792 37744
rect 5808 37680 5872 37744
rect 5888 37680 5952 37744
rect 5968 37680 6032 37744
rect 6048 37680 6112 37744
rect 6128 37680 6192 37744
rect 6208 37680 6272 37744
rect 6288 37680 6352 37744
rect 6368 37680 6432 37744
rect 6448 37680 6512 37744
rect 6528 37680 6592 37744
rect 6608 37680 6672 37744
rect 6688 37680 6752 37744
rect 6768 37680 6832 37744
rect 6848 37680 6912 37744
rect 6928 37680 6992 37744
rect 7008 37680 7072 37744
rect 7088 37680 7152 37744
rect 7168 37680 7232 37744
rect 7248 37680 7312 37744
rect 7328 37680 7392 37744
rect 7408 37680 7472 37744
rect 7488 37680 7552 37744
rect 7568 37680 7632 37744
rect 7648 37680 7712 37744
rect 7728 37680 7792 37744
rect 7808 37680 7872 37744
rect 7888 37680 7952 37744
rect 7968 37680 8032 37744
rect 8048 37680 8112 37744
rect 8128 37680 8192 37744
rect 8208 37680 8272 37744
rect 8288 37680 8352 37744
rect 8368 37680 8432 37744
rect 8448 37680 8512 37744
rect 8528 37680 8592 37744
rect 8608 37680 8672 37744
rect 8688 37680 8752 37744
rect 8768 37680 8832 37744
rect 8848 37680 8912 37744
rect 8928 37680 8992 37744
rect 14112 37680 14176 37744
rect 14192 37680 14256 37744
rect 14272 37680 14336 37744
rect 14352 37680 14416 37744
rect 24112 37680 24176 37744
rect 24192 37680 24256 37744
rect 24272 37680 24336 37744
rect 24352 37680 24416 37744
rect 36376 37680 36440 37744
rect 36456 37680 36520 37744
rect 36536 37680 36600 37744
rect 36616 37680 36680 37744
rect 36696 37680 36760 37744
rect 36776 37680 36840 37744
rect 36856 37680 36920 37744
rect 36936 37680 37000 37744
rect 37016 37680 37080 37744
rect 37096 37680 37160 37744
rect 37176 37680 37240 37744
rect 37256 37680 37320 37744
rect 37336 37680 37400 37744
rect 37416 37680 37480 37744
rect 37496 37680 37560 37744
rect 37576 37680 37640 37744
rect 37656 37680 37720 37744
rect 37736 37680 37800 37744
rect 37816 37680 37880 37744
rect 37896 37680 37960 37744
rect 37976 37680 38040 37744
rect 38056 37680 38120 37744
rect 38136 37680 38200 37744
rect 38216 37680 38280 37744
rect 38296 37680 38360 37744
rect 38376 37680 38440 37744
rect 38456 37680 38520 37744
rect 38536 37680 38600 37744
rect 38616 37680 38680 37744
rect 38696 37680 38760 37744
rect 38776 37680 38840 37744
rect 38856 37680 38920 37744
rect 38936 37680 39000 37744
rect 39016 37680 39080 37744
rect 39096 37680 39160 37744
rect 39176 37680 39240 37744
rect 39256 37680 39320 37744
rect 39336 37680 39400 37744
rect 39416 37680 39480 37744
rect 39496 37680 39560 37744
rect 39576 37680 39640 37744
rect 39656 37680 39720 37744
rect 39736 37680 39800 37744
rect 39816 37680 39880 37744
rect 39896 37680 39960 37744
rect 39976 37680 40040 37744
rect 40056 37680 40120 37744
rect 40136 37680 40200 37744
rect 40216 37680 40280 37744
rect 40296 37680 40360 37744
rect 5008 37600 5072 37664
rect 5088 37600 5152 37664
rect 5168 37600 5232 37664
rect 5248 37600 5312 37664
rect 5328 37600 5392 37664
rect 5408 37600 5472 37664
rect 5488 37600 5552 37664
rect 5568 37600 5632 37664
rect 5648 37600 5712 37664
rect 5728 37600 5792 37664
rect 5808 37600 5872 37664
rect 5888 37600 5952 37664
rect 5968 37600 6032 37664
rect 6048 37600 6112 37664
rect 6128 37600 6192 37664
rect 6208 37600 6272 37664
rect 6288 37600 6352 37664
rect 6368 37600 6432 37664
rect 6448 37600 6512 37664
rect 6528 37600 6592 37664
rect 6608 37600 6672 37664
rect 6688 37600 6752 37664
rect 6768 37600 6832 37664
rect 6848 37600 6912 37664
rect 6928 37600 6992 37664
rect 7008 37600 7072 37664
rect 7088 37600 7152 37664
rect 7168 37600 7232 37664
rect 7248 37600 7312 37664
rect 7328 37600 7392 37664
rect 7408 37600 7472 37664
rect 7488 37600 7552 37664
rect 7568 37600 7632 37664
rect 7648 37600 7712 37664
rect 7728 37600 7792 37664
rect 7808 37600 7872 37664
rect 7888 37600 7952 37664
rect 7968 37600 8032 37664
rect 8048 37600 8112 37664
rect 8128 37600 8192 37664
rect 8208 37600 8272 37664
rect 8288 37600 8352 37664
rect 8368 37600 8432 37664
rect 8448 37600 8512 37664
rect 8528 37600 8592 37664
rect 8608 37600 8672 37664
rect 8688 37600 8752 37664
rect 8768 37600 8832 37664
rect 8848 37600 8912 37664
rect 8928 37600 8992 37664
rect 14112 37600 14176 37664
rect 14192 37600 14256 37664
rect 14272 37600 14336 37664
rect 14352 37600 14416 37664
rect 24112 37600 24176 37664
rect 24192 37600 24256 37664
rect 24272 37600 24336 37664
rect 24352 37600 24416 37664
rect 36376 37600 36440 37664
rect 36456 37600 36520 37664
rect 36536 37600 36600 37664
rect 36616 37600 36680 37664
rect 36696 37600 36760 37664
rect 36776 37600 36840 37664
rect 36856 37600 36920 37664
rect 36936 37600 37000 37664
rect 37016 37600 37080 37664
rect 37096 37600 37160 37664
rect 37176 37600 37240 37664
rect 37256 37600 37320 37664
rect 37336 37600 37400 37664
rect 37416 37600 37480 37664
rect 37496 37600 37560 37664
rect 37576 37600 37640 37664
rect 37656 37600 37720 37664
rect 37736 37600 37800 37664
rect 37816 37600 37880 37664
rect 37896 37600 37960 37664
rect 37976 37600 38040 37664
rect 38056 37600 38120 37664
rect 38136 37600 38200 37664
rect 38216 37600 38280 37664
rect 38296 37600 38360 37664
rect 38376 37600 38440 37664
rect 38456 37600 38520 37664
rect 38536 37600 38600 37664
rect 38616 37600 38680 37664
rect 38696 37600 38760 37664
rect 38776 37600 38840 37664
rect 38856 37600 38920 37664
rect 38936 37600 39000 37664
rect 39016 37600 39080 37664
rect 39096 37600 39160 37664
rect 39176 37600 39240 37664
rect 39256 37600 39320 37664
rect 39336 37600 39400 37664
rect 39416 37600 39480 37664
rect 39496 37600 39560 37664
rect 39576 37600 39640 37664
rect 39656 37600 39720 37664
rect 39736 37600 39800 37664
rect 39816 37600 39880 37664
rect 39896 37600 39960 37664
rect 39976 37600 40040 37664
rect 40056 37600 40120 37664
rect 40136 37600 40200 37664
rect 40216 37600 40280 37664
rect 40296 37600 40360 37664
rect 5008 37520 5072 37584
rect 5088 37520 5152 37584
rect 5168 37520 5232 37584
rect 5248 37520 5312 37584
rect 5328 37520 5392 37584
rect 5408 37520 5472 37584
rect 5488 37520 5552 37584
rect 5568 37520 5632 37584
rect 5648 37520 5712 37584
rect 5728 37520 5792 37584
rect 5808 37520 5872 37584
rect 5888 37520 5952 37584
rect 5968 37520 6032 37584
rect 6048 37520 6112 37584
rect 6128 37520 6192 37584
rect 6208 37520 6272 37584
rect 6288 37520 6352 37584
rect 6368 37520 6432 37584
rect 6448 37520 6512 37584
rect 6528 37520 6592 37584
rect 6608 37520 6672 37584
rect 6688 37520 6752 37584
rect 6768 37520 6832 37584
rect 6848 37520 6912 37584
rect 6928 37520 6992 37584
rect 7008 37520 7072 37584
rect 7088 37520 7152 37584
rect 7168 37520 7232 37584
rect 7248 37520 7312 37584
rect 7328 37520 7392 37584
rect 7408 37520 7472 37584
rect 7488 37520 7552 37584
rect 7568 37520 7632 37584
rect 7648 37520 7712 37584
rect 7728 37520 7792 37584
rect 7808 37520 7872 37584
rect 7888 37520 7952 37584
rect 7968 37520 8032 37584
rect 8048 37520 8112 37584
rect 8128 37520 8192 37584
rect 8208 37520 8272 37584
rect 8288 37520 8352 37584
rect 8368 37520 8432 37584
rect 8448 37520 8512 37584
rect 8528 37520 8592 37584
rect 8608 37520 8672 37584
rect 8688 37520 8752 37584
rect 8768 37520 8832 37584
rect 8848 37520 8912 37584
rect 8928 37520 8992 37584
rect 14112 37520 14176 37584
rect 14192 37520 14256 37584
rect 14272 37520 14336 37584
rect 14352 37520 14416 37584
rect 24112 37520 24176 37584
rect 24192 37520 24256 37584
rect 24272 37520 24336 37584
rect 24352 37520 24416 37584
rect 36376 37520 36440 37584
rect 36456 37520 36520 37584
rect 36536 37520 36600 37584
rect 36616 37520 36680 37584
rect 36696 37520 36760 37584
rect 36776 37520 36840 37584
rect 36856 37520 36920 37584
rect 36936 37520 37000 37584
rect 37016 37520 37080 37584
rect 37096 37520 37160 37584
rect 37176 37520 37240 37584
rect 37256 37520 37320 37584
rect 37336 37520 37400 37584
rect 37416 37520 37480 37584
rect 37496 37520 37560 37584
rect 37576 37520 37640 37584
rect 37656 37520 37720 37584
rect 37736 37520 37800 37584
rect 37816 37520 37880 37584
rect 37896 37520 37960 37584
rect 37976 37520 38040 37584
rect 38056 37520 38120 37584
rect 38136 37520 38200 37584
rect 38216 37520 38280 37584
rect 38296 37520 38360 37584
rect 38376 37520 38440 37584
rect 38456 37520 38520 37584
rect 38536 37520 38600 37584
rect 38616 37520 38680 37584
rect 38696 37520 38760 37584
rect 38776 37520 38840 37584
rect 38856 37520 38920 37584
rect 38936 37520 39000 37584
rect 39016 37520 39080 37584
rect 39096 37520 39160 37584
rect 39176 37520 39240 37584
rect 39256 37520 39320 37584
rect 39336 37520 39400 37584
rect 39416 37520 39480 37584
rect 39496 37520 39560 37584
rect 39576 37520 39640 37584
rect 39656 37520 39720 37584
rect 39736 37520 39800 37584
rect 39816 37520 39880 37584
rect 39896 37520 39960 37584
rect 39976 37520 40040 37584
rect 40056 37520 40120 37584
rect 40136 37520 40200 37584
rect 40216 37520 40280 37584
rect 40296 37520 40360 37584
rect 5008 37440 5072 37504
rect 5088 37440 5152 37504
rect 5168 37440 5232 37504
rect 5248 37440 5312 37504
rect 5328 37440 5392 37504
rect 5408 37440 5472 37504
rect 5488 37440 5552 37504
rect 5568 37440 5632 37504
rect 5648 37440 5712 37504
rect 5728 37440 5792 37504
rect 5808 37440 5872 37504
rect 5888 37440 5952 37504
rect 5968 37440 6032 37504
rect 6048 37440 6112 37504
rect 6128 37440 6192 37504
rect 6208 37440 6272 37504
rect 6288 37440 6352 37504
rect 6368 37440 6432 37504
rect 6448 37440 6512 37504
rect 6528 37440 6592 37504
rect 6608 37440 6672 37504
rect 6688 37440 6752 37504
rect 6768 37440 6832 37504
rect 6848 37440 6912 37504
rect 6928 37440 6992 37504
rect 7008 37440 7072 37504
rect 7088 37440 7152 37504
rect 7168 37440 7232 37504
rect 7248 37440 7312 37504
rect 7328 37440 7392 37504
rect 7408 37440 7472 37504
rect 7488 37440 7552 37504
rect 7568 37440 7632 37504
rect 7648 37440 7712 37504
rect 7728 37440 7792 37504
rect 7808 37440 7872 37504
rect 7888 37440 7952 37504
rect 7968 37440 8032 37504
rect 8048 37440 8112 37504
rect 8128 37440 8192 37504
rect 8208 37440 8272 37504
rect 8288 37440 8352 37504
rect 8368 37440 8432 37504
rect 8448 37440 8512 37504
rect 8528 37440 8592 37504
rect 8608 37440 8672 37504
rect 8688 37440 8752 37504
rect 8768 37440 8832 37504
rect 8848 37440 8912 37504
rect 8928 37440 8992 37504
rect 14112 37440 14176 37504
rect 14192 37440 14256 37504
rect 14272 37440 14336 37504
rect 14352 37440 14416 37504
rect 24112 37440 24176 37504
rect 24192 37440 24256 37504
rect 24272 37440 24336 37504
rect 24352 37440 24416 37504
rect 36376 37440 36440 37504
rect 36456 37440 36520 37504
rect 36536 37440 36600 37504
rect 36616 37440 36680 37504
rect 36696 37440 36760 37504
rect 36776 37440 36840 37504
rect 36856 37440 36920 37504
rect 36936 37440 37000 37504
rect 37016 37440 37080 37504
rect 37096 37440 37160 37504
rect 37176 37440 37240 37504
rect 37256 37440 37320 37504
rect 37336 37440 37400 37504
rect 37416 37440 37480 37504
rect 37496 37440 37560 37504
rect 37576 37440 37640 37504
rect 37656 37440 37720 37504
rect 37736 37440 37800 37504
rect 37816 37440 37880 37504
rect 37896 37440 37960 37504
rect 37976 37440 38040 37504
rect 38056 37440 38120 37504
rect 38136 37440 38200 37504
rect 38216 37440 38280 37504
rect 38296 37440 38360 37504
rect 38376 37440 38440 37504
rect 38456 37440 38520 37504
rect 38536 37440 38600 37504
rect 38616 37440 38680 37504
rect 38696 37440 38760 37504
rect 38776 37440 38840 37504
rect 38856 37440 38920 37504
rect 38936 37440 39000 37504
rect 39016 37440 39080 37504
rect 39096 37440 39160 37504
rect 39176 37440 39240 37504
rect 39256 37440 39320 37504
rect 39336 37440 39400 37504
rect 39416 37440 39480 37504
rect 39496 37440 39560 37504
rect 39576 37440 39640 37504
rect 39656 37440 39720 37504
rect 39736 37440 39800 37504
rect 39816 37440 39880 37504
rect 39896 37440 39960 37504
rect 39976 37440 40040 37504
rect 40056 37440 40120 37504
rect 40136 37440 40200 37504
rect 40216 37440 40280 37504
rect 40296 37440 40360 37504
rect 5008 37360 5072 37424
rect 5088 37360 5152 37424
rect 5168 37360 5232 37424
rect 5248 37360 5312 37424
rect 5328 37360 5392 37424
rect 5408 37360 5472 37424
rect 5488 37360 5552 37424
rect 5568 37360 5632 37424
rect 5648 37360 5712 37424
rect 5728 37360 5792 37424
rect 5808 37360 5872 37424
rect 5888 37360 5952 37424
rect 5968 37360 6032 37424
rect 6048 37360 6112 37424
rect 6128 37360 6192 37424
rect 6208 37360 6272 37424
rect 6288 37360 6352 37424
rect 6368 37360 6432 37424
rect 6448 37360 6512 37424
rect 6528 37360 6592 37424
rect 6608 37360 6672 37424
rect 6688 37360 6752 37424
rect 6768 37360 6832 37424
rect 6848 37360 6912 37424
rect 6928 37360 6992 37424
rect 7008 37360 7072 37424
rect 7088 37360 7152 37424
rect 7168 37360 7232 37424
rect 7248 37360 7312 37424
rect 7328 37360 7392 37424
rect 7408 37360 7472 37424
rect 7488 37360 7552 37424
rect 7568 37360 7632 37424
rect 7648 37360 7712 37424
rect 7728 37360 7792 37424
rect 7808 37360 7872 37424
rect 7888 37360 7952 37424
rect 7968 37360 8032 37424
rect 8048 37360 8112 37424
rect 8128 37360 8192 37424
rect 8208 37360 8272 37424
rect 8288 37360 8352 37424
rect 8368 37360 8432 37424
rect 8448 37360 8512 37424
rect 8528 37360 8592 37424
rect 8608 37360 8672 37424
rect 8688 37360 8752 37424
rect 8768 37360 8832 37424
rect 8848 37360 8912 37424
rect 8928 37360 8992 37424
rect 14112 37360 14176 37424
rect 14192 37360 14256 37424
rect 14272 37360 14336 37424
rect 14352 37360 14416 37424
rect 24112 37360 24176 37424
rect 24192 37360 24256 37424
rect 24272 37360 24336 37424
rect 24352 37360 24416 37424
rect 36376 37360 36440 37424
rect 36456 37360 36520 37424
rect 36536 37360 36600 37424
rect 36616 37360 36680 37424
rect 36696 37360 36760 37424
rect 36776 37360 36840 37424
rect 36856 37360 36920 37424
rect 36936 37360 37000 37424
rect 37016 37360 37080 37424
rect 37096 37360 37160 37424
rect 37176 37360 37240 37424
rect 37256 37360 37320 37424
rect 37336 37360 37400 37424
rect 37416 37360 37480 37424
rect 37496 37360 37560 37424
rect 37576 37360 37640 37424
rect 37656 37360 37720 37424
rect 37736 37360 37800 37424
rect 37816 37360 37880 37424
rect 37896 37360 37960 37424
rect 37976 37360 38040 37424
rect 38056 37360 38120 37424
rect 38136 37360 38200 37424
rect 38216 37360 38280 37424
rect 38296 37360 38360 37424
rect 38376 37360 38440 37424
rect 38456 37360 38520 37424
rect 38536 37360 38600 37424
rect 38616 37360 38680 37424
rect 38696 37360 38760 37424
rect 38776 37360 38840 37424
rect 38856 37360 38920 37424
rect 38936 37360 39000 37424
rect 39016 37360 39080 37424
rect 39096 37360 39160 37424
rect 39176 37360 39240 37424
rect 39256 37360 39320 37424
rect 39336 37360 39400 37424
rect 39416 37360 39480 37424
rect 39496 37360 39560 37424
rect 39576 37360 39640 37424
rect 39656 37360 39720 37424
rect 39736 37360 39800 37424
rect 39816 37360 39880 37424
rect 39896 37360 39960 37424
rect 39976 37360 40040 37424
rect 40056 37360 40120 37424
rect 40136 37360 40200 37424
rect 40216 37360 40280 37424
rect 40296 37360 40360 37424
rect 5008 37280 5072 37344
rect 5088 37280 5152 37344
rect 5168 37280 5232 37344
rect 5248 37280 5312 37344
rect 5328 37280 5392 37344
rect 5408 37280 5472 37344
rect 5488 37280 5552 37344
rect 5568 37280 5632 37344
rect 5648 37280 5712 37344
rect 5728 37280 5792 37344
rect 5808 37280 5872 37344
rect 5888 37280 5952 37344
rect 5968 37280 6032 37344
rect 6048 37280 6112 37344
rect 6128 37280 6192 37344
rect 6208 37280 6272 37344
rect 6288 37280 6352 37344
rect 6368 37280 6432 37344
rect 6448 37280 6512 37344
rect 6528 37280 6592 37344
rect 6608 37280 6672 37344
rect 6688 37280 6752 37344
rect 6768 37280 6832 37344
rect 6848 37280 6912 37344
rect 6928 37280 6992 37344
rect 7008 37280 7072 37344
rect 7088 37280 7152 37344
rect 7168 37280 7232 37344
rect 7248 37280 7312 37344
rect 7328 37280 7392 37344
rect 7408 37280 7472 37344
rect 7488 37280 7552 37344
rect 7568 37280 7632 37344
rect 7648 37280 7712 37344
rect 7728 37280 7792 37344
rect 7808 37280 7872 37344
rect 7888 37280 7952 37344
rect 7968 37280 8032 37344
rect 8048 37280 8112 37344
rect 8128 37280 8192 37344
rect 8208 37280 8272 37344
rect 8288 37280 8352 37344
rect 8368 37280 8432 37344
rect 8448 37280 8512 37344
rect 8528 37280 8592 37344
rect 8608 37280 8672 37344
rect 8688 37280 8752 37344
rect 8768 37280 8832 37344
rect 8848 37280 8912 37344
rect 8928 37280 8992 37344
rect 14112 37280 14176 37344
rect 14192 37280 14256 37344
rect 14272 37280 14336 37344
rect 14352 37280 14416 37344
rect 24112 37280 24176 37344
rect 24192 37280 24256 37344
rect 24272 37280 24336 37344
rect 24352 37280 24416 37344
rect 36376 37280 36440 37344
rect 36456 37280 36520 37344
rect 36536 37280 36600 37344
rect 36616 37280 36680 37344
rect 36696 37280 36760 37344
rect 36776 37280 36840 37344
rect 36856 37280 36920 37344
rect 36936 37280 37000 37344
rect 37016 37280 37080 37344
rect 37096 37280 37160 37344
rect 37176 37280 37240 37344
rect 37256 37280 37320 37344
rect 37336 37280 37400 37344
rect 37416 37280 37480 37344
rect 37496 37280 37560 37344
rect 37576 37280 37640 37344
rect 37656 37280 37720 37344
rect 37736 37280 37800 37344
rect 37816 37280 37880 37344
rect 37896 37280 37960 37344
rect 37976 37280 38040 37344
rect 38056 37280 38120 37344
rect 38136 37280 38200 37344
rect 38216 37280 38280 37344
rect 38296 37280 38360 37344
rect 38376 37280 38440 37344
rect 38456 37280 38520 37344
rect 38536 37280 38600 37344
rect 38616 37280 38680 37344
rect 38696 37280 38760 37344
rect 38776 37280 38840 37344
rect 38856 37280 38920 37344
rect 38936 37280 39000 37344
rect 39016 37280 39080 37344
rect 39096 37280 39160 37344
rect 39176 37280 39240 37344
rect 39256 37280 39320 37344
rect 39336 37280 39400 37344
rect 39416 37280 39480 37344
rect 39496 37280 39560 37344
rect 39576 37280 39640 37344
rect 39656 37280 39720 37344
rect 39736 37280 39800 37344
rect 39816 37280 39880 37344
rect 39896 37280 39960 37344
rect 39976 37280 40040 37344
rect 40056 37280 40120 37344
rect 40136 37280 40200 37344
rect 40216 37280 40280 37344
rect 40296 37280 40360 37344
rect 5008 37200 5072 37264
rect 5088 37200 5152 37264
rect 5168 37200 5232 37264
rect 5248 37200 5312 37264
rect 5328 37200 5392 37264
rect 5408 37200 5472 37264
rect 5488 37200 5552 37264
rect 5568 37200 5632 37264
rect 5648 37200 5712 37264
rect 5728 37200 5792 37264
rect 5808 37200 5872 37264
rect 5888 37200 5952 37264
rect 5968 37200 6032 37264
rect 6048 37200 6112 37264
rect 6128 37200 6192 37264
rect 6208 37200 6272 37264
rect 6288 37200 6352 37264
rect 6368 37200 6432 37264
rect 6448 37200 6512 37264
rect 6528 37200 6592 37264
rect 6608 37200 6672 37264
rect 6688 37200 6752 37264
rect 6768 37200 6832 37264
rect 6848 37200 6912 37264
rect 6928 37200 6992 37264
rect 7008 37200 7072 37264
rect 7088 37200 7152 37264
rect 7168 37200 7232 37264
rect 7248 37200 7312 37264
rect 7328 37200 7392 37264
rect 7408 37200 7472 37264
rect 7488 37200 7552 37264
rect 7568 37200 7632 37264
rect 7648 37200 7712 37264
rect 7728 37200 7792 37264
rect 7808 37200 7872 37264
rect 7888 37200 7952 37264
rect 7968 37200 8032 37264
rect 8048 37200 8112 37264
rect 8128 37200 8192 37264
rect 8208 37200 8272 37264
rect 8288 37200 8352 37264
rect 8368 37200 8432 37264
rect 8448 37200 8512 37264
rect 8528 37200 8592 37264
rect 8608 37200 8672 37264
rect 8688 37200 8752 37264
rect 8768 37200 8832 37264
rect 8848 37200 8912 37264
rect 8928 37200 8992 37264
rect 14112 37200 14176 37264
rect 14192 37200 14256 37264
rect 14272 37200 14336 37264
rect 14352 37200 14416 37264
rect 24112 37200 24176 37264
rect 24192 37200 24256 37264
rect 24272 37200 24336 37264
rect 24352 37200 24416 37264
rect 36376 37200 36440 37264
rect 36456 37200 36520 37264
rect 36536 37200 36600 37264
rect 36616 37200 36680 37264
rect 36696 37200 36760 37264
rect 36776 37200 36840 37264
rect 36856 37200 36920 37264
rect 36936 37200 37000 37264
rect 37016 37200 37080 37264
rect 37096 37200 37160 37264
rect 37176 37200 37240 37264
rect 37256 37200 37320 37264
rect 37336 37200 37400 37264
rect 37416 37200 37480 37264
rect 37496 37200 37560 37264
rect 37576 37200 37640 37264
rect 37656 37200 37720 37264
rect 37736 37200 37800 37264
rect 37816 37200 37880 37264
rect 37896 37200 37960 37264
rect 37976 37200 38040 37264
rect 38056 37200 38120 37264
rect 38136 37200 38200 37264
rect 38216 37200 38280 37264
rect 38296 37200 38360 37264
rect 38376 37200 38440 37264
rect 38456 37200 38520 37264
rect 38536 37200 38600 37264
rect 38616 37200 38680 37264
rect 38696 37200 38760 37264
rect 38776 37200 38840 37264
rect 38856 37200 38920 37264
rect 38936 37200 39000 37264
rect 39016 37200 39080 37264
rect 39096 37200 39160 37264
rect 39176 37200 39240 37264
rect 39256 37200 39320 37264
rect 39336 37200 39400 37264
rect 39416 37200 39480 37264
rect 39496 37200 39560 37264
rect 39576 37200 39640 37264
rect 39656 37200 39720 37264
rect 39736 37200 39800 37264
rect 39816 37200 39880 37264
rect 39896 37200 39960 37264
rect 39976 37200 40040 37264
rect 40056 37200 40120 37264
rect 40136 37200 40200 37264
rect 40216 37200 40280 37264
rect 40296 37200 40360 37264
rect 5008 37120 5072 37184
rect 5088 37120 5152 37184
rect 5168 37120 5232 37184
rect 5248 37120 5312 37184
rect 5328 37120 5392 37184
rect 5408 37120 5472 37184
rect 5488 37120 5552 37184
rect 5568 37120 5632 37184
rect 5648 37120 5712 37184
rect 5728 37120 5792 37184
rect 5808 37120 5872 37184
rect 5888 37120 5952 37184
rect 5968 37120 6032 37184
rect 6048 37120 6112 37184
rect 6128 37120 6192 37184
rect 6208 37120 6272 37184
rect 6288 37120 6352 37184
rect 6368 37120 6432 37184
rect 6448 37120 6512 37184
rect 6528 37120 6592 37184
rect 6608 37120 6672 37184
rect 6688 37120 6752 37184
rect 6768 37120 6832 37184
rect 6848 37120 6912 37184
rect 6928 37120 6992 37184
rect 7008 37120 7072 37184
rect 7088 37120 7152 37184
rect 7168 37120 7232 37184
rect 7248 37120 7312 37184
rect 7328 37120 7392 37184
rect 7408 37120 7472 37184
rect 7488 37120 7552 37184
rect 7568 37120 7632 37184
rect 7648 37120 7712 37184
rect 7728 37120 7792 37184
rect 7808 37120 7872 37184
rect 7888 37120 7952 37184
rect 7968 37120 8032 37184
rect 8048 37120 8112 37184
rect 8128 37120 8192 37184
rect 8208 37120 8272 37184
rect 8288 37120 8352 37184
rect 8368 37120 8432 37184
rect 8448 37120 8512 37184
rect 8528 37120 8592 37184
rect 8608 37120 8672 37184
rect 8688 37120 8752 37184
rect 8768 37120 8832 37184
rect 8848 37120 8912 37184
rect 8928 37120 8992 37184
rect 14112 37120 14176 37184
rect 14192 37120 14256 37184
rect 14272 37120 14336 37184
rect 14352 37120 14416 37184
rect 24112 37120 24176 37184
rect 24192 37120 24256 37184
rect 24272 37120 24336 37184
rect 24352 37120 24416 37184
rect 36376 37120 36440 37184
rect 36456 37120 36520 37184
rect 36536 37120 36600 37184
rect 36616 37120 36680 37184
rect 36696 37120 36760 37184
rect 36776 37120 36840 37184
rect 36856 37120 36920 37184
rect 36936 37120 37000 37184
rect 37016 37120 37080 37184
rect 37096 37120 37160 37184
rect 37176 37120 37240 37184
rect 37256 37120 37320 37184
rect 37336 37120 37400 37184
rect 37416 37120 37480 37184
rect 37496 37120 37560 37184
rect 37576 37120 37640 37184
rect 37656 37120 37720 37184
rect 37736 37120 37800 37184
rect 37816 37120 37880 37184
rect 37896 37120 37960 37184
rect 37976 37120 38040 37184
rect 38056 37120 38120 37184
rect 38136 37120 38200 37184
rect 38216 37120 38280 37184
rect 38296 37120 38360 37184
rect 38376 37120 38440 37184
rect 38456 37120 38520 37184
rect 38536 37120 38600 37184
rect 38616 37120 38680 37184
rect 38696 37120 38760 37184
rect 38776 37120 38840 37184
rect 38856 37120 38920 37184
rect 38936 37120 39000 37184
rect 39016 37120 39080 37184
rect 39096 37120 39160 37184
rect 39176 37120 39240 37184
rect 39256 37120 39320 37184
rect 39336 37120 39400 37184
rect 39416 37120 39480 37184
rect 39496 37120 39560 37184
rect 39576 37120 39640 37184
rect 39656 37120 39720 37184
rect 39736 37120 39800 37184
rect 39816 37120 39880 37184
rect 39896 37120 39960 37184
rect 39976 37120 40040 37184
rect 40056 37120 40120 37184
rect 40136 37120 40200 37184
rect 40216 37120 40280 37184
rect 40296 37120 40360 37184
rect 5008 37040 5072 37104
rect 5088 37040 5152 37104
rect 5168 37040 5232 37104
rect 5248 37040 5312 37104
rect 5328 37040 5392 37104
rect 5408 37040 5472 37104
rect 5488 37040 5552 37104
rect 5568 37040 5632 37104
rect 5648 37040 5712 37104
rect 5728 37040 5792 37104
rect 5808 37040 5872 37104
rect 5888 37040 5952 37104
rect 5968 37040 6032 37104
rect 6048 37040 6112 37104
rect 6128 37040 6192 37104
rect 6208 37040 6272 37104
rect 6288 37040 6352 37104
rect 6368 37040 6432 37104
rect 6448 37040 6512 37104
rect 6528 37040 6592 37104
rect 6608 37040 6672 37104
rect 6688 37040 6752 37104
rect 6768 37040 6832 37104
rect 6848 37040 6912 37104
rect 6928 37040 6992 37104
rect 7008 37040 7072 37104
rect 7088 37040 7152 37104
rect 7168 37040 7232 37104
rect 7248 37040 7312 37104
rect 7328 37040 7392 37104
rect 7408 37040 7472 37104
rect 7488 37040 7552 37104
rect 7568 37040 7632 37104
rect 7648 37040 7712 37104
rect 7728 37040 7792 37104
rect 7808 37040 7872 37104
rect 7888 37040 7952 37104
rect 7968 37040 8032 37104
rect 8048 37040 8112 37104
rect 8128 37040 8192 37104
rect 8208 37040 8272 37104
rect 8288 37040 8352 37104
rect 8368 37040 8432 37104
rect 8448 37040 8512 37104
rect 8528 37040 8592 37104
rect 8608 37040 8672 37104
rect 8688 37040 8752 37104
rect 8768 37040 8832 37104
rect 8848 37040 8912 37104
rect 8928 37040 8992 37104
rect 14112 37040 14176 37104
rect 14192 37040 14256 37104
rect 14272 37040 14336 37104
rect 14352 37040 14416 37104
rect 24112 37040 24176 37104
rect 24192 37040 24256 37104
rect 24272 37040 24336 37104
rect 24352 37040 24416 37104
rect 36376 37040 36440 37104
rect 36456 37040 36520 37104
rect 36536 37040 36600 37104
rect 36616 37040 36680 37104
rect 36696 37040 36760 37104
rect 36776 37040 36840 37104
rect 36856 37040 36920 37104
rect 36936 37040 37000 37104
rect 37016 37040 37080 37104
rect 37096 37040 37160 37104
rect 37176 37040 37240 37104
rect 37256 37040 37320 37104
rect 37336 37040 37400 37104
rect 37416 37040 37480 37104
rect 37496 37040 37560 37104
rect 37576 37040 37640 37104
rect 37656 37040 37720 37104
rect 37736 37040 37800 37104
rect 37816 37040 37880 37104
rect 37896 37040 37960 37104
rect 37976 37040 38040 37104
rect 38056 37040 38120 37104
rect 38136 37040 38200 37104
rect 38216 37040 38280 37104
rect 38296 37040 38360 37104
rect 38376 37040 38440 37104
rect 38456 37040 38520 37104
rect 38536 37040 38600 37104
rect 38616 37040 38680 37104
rect 38696 37040 38760 37104
rect 38776 37040 38840 37104
rect 38856 37040 38920 37104
rect 38936 37040 39000 37104
rect 39016 37040 39080 37104
rect 39096 37040 39160 37104
rect 39176 37040 39240 37104
rect 39256 37040 39320 37104
rect 39336 37040 39400 37104
rect 39416 37040 39480 37104
rect 39496 37040 39560 37104
rect 39576 37040 39640 37104
rect 39656 37040 39720 37104
rect 39736 37040 39800 37104
rect 39816 37040 39880 37104
rect 39896 37040 39960 37104
rect 39976 37040 40040 37104
rect 40056 37040 40120 37104
rect 40136 37040 40200 37104
rect 40216 37040 40280 37104
rect 40296 37040 40360 37104
rect 5008 36960 5072 37024
rect 5088 36960 5152 37024
rect 5168 36960 5232 37024
rect 5248 36960 5312 37024
rect 5328 36960 5392 37024
rect 5408 36960 5472 37024
rect 5488 36960 5552 37024
rect 5568 36960 5632 37024
rect 5648 36960 5712 37024
rect 5728 36960 5792 37024
rect 5808 36960 5872 37024
rect 5888 36960 5952 37024
rect 5968 36960 6032 37024
rect 6048 36960 6112 37024
rect 6128 36960 6192 37024
rect 6208 36960 6272 37024
rect 6288 36960 6352 37024
rect 6368 36960 6432 37024
rect 6448 36960 6512 37024
rect 6528 36960 6592 37024
rect 6608 36960 6672 37024
rect 6688 36960 6752 37024
rect 6768 36960 6832 37024
rect 6848 36960 6912 37024
rect 6928 36960 6992 37024
rect 7008 36960 7072 37024
rect 7088 36960 7152 37024
rect 7168 36960 7232 37024
rect 7248 36960 7312 37024
rect 7328 36960 7392 37024
rect 7408 36960 7472 37024
rect 7488 36960 7552 37024
rect 7568 36960 7632 37024
rect 7648 36960 7712 37024
rect 7728 36960 7792 37024
rect 7808 36960 7872 37024
rect 7888 36960 7952 37024
rect 7968 36960 8032 37024
rect 8048 36960 8112 37024
rect 8128 36960 8192 37024
rect 8208 36960 8272 37024
rect 8288 36960 8352 37024
rect 8368 36960 8432 37024
rect 8448 36960 8512 37024
rect 8528 36960 8592 37024
rect 8608 36960 8672 37024
rect 8688 36960 8752 37024
rect 8768 36960 8832 37024
rect 8848 36960 8912 37024
rect 8928 36960 8992 37024
rect 14112 36960 14176 37024
rect 14192 36960 14256 37024
rect 14272 36960 14336 37024
rect 14352 36960 14416 37024
rect 24112 36960 24176 37024
rect 24192 36960 24256 37024
rect 24272 36960 24336 37024
rect 24352 36960 24416 37024
rect 36376 36960 36440 37024
rect 36456 36960 36520 37024
rect 36536 36960 36600 37024
rect 36616 36960 36680 37024
rect 36696 36960 36760 37024
rect 36776 36960 36840 37024
rect 36856 36960 36920 37024
rect 36936 36960 37000 37024
rect 37016 36960 37080 37024
rect 37096 36960 37160 37024
rect 37176 36960 37240 37024
rect 37256 36960 37320 37024
rect 37336 36960 37400 37024
rect 37416 36960 37480 37024
rect 37496 36960 37560 37024
rect 37576 36960 37640 37024
rect 37656 36960 37720 37024
rect 37736 36960 37800 37024
rect 37816 36960 37880 37024
rect 37896 36960 37960 37024
rect 37976 36960 38040 37024
rect 38056 36960 38120 37024
rect 38136 36960 38200 37024
rect 38216 36960 38280 37024
rect 38296 36960 38360 37024
rect 38376 36960 38440 37024
rect 38456 36960 38520 37024
rect 38536 36960 38600 37024
rect 38616 36960 38680 37024
rect 38696 36960 38760 37024
rect 38776 36960 38840 37024
rect 38856 36960 38920 37024
rect 38936 36960 39000 37024
rect 39016 36960 39080 37024
rect 39096 36960 39160 37024
rect 39176 36960 39240 37024
rect 39256 36960 39320 37024
rect 39336 36960 39400 37024
rect 39416 36960 39480 37024
rect 39496 36960 39560 37024
rect 39576 36960 39640 37024
rect 39656 36960 39720 37024
rect 39736 36960 39800 37024
rect 39816 36960 39880 37024
rect 39896 36960 39960 37024
rect 39976 36960 40040 37024
rect 40056 36960 40120 37024
rect 40136 36960 40200 37024
rect 40216 36960 40280 37024
rect 40296 36960 40360 37024
rect 5008 36880 5072 36944
rect 5088 36880 5152 36944
rect 5168 36880 5232 36944
rect 5248 36880 5312 36944
rect 5328 36880 5392 36944
rect 5408 36880 5472 36944
rect 5488 36880 5552 36944
rect 5568 36880 5632 36944
rect 5648 36880 5712 36944
rect 5728 36880 5792 36944
rect 5808 36880 5872 36944
rect 5888 36880 5952 36944
rect 5968 36880 6032 36944
rect 6048 36880 6112 36944
rect 6128 36880 6192 36944
rect 6208 36880 6272 36944
rect 6288 36880 6352 36944
rect 6368 36880 6432 36944
rect 6448 36880 6512 36944
rect 6528 36880 6592 36944
rect 6608 36880 6672 36944
rect 6688 36880 6752 36944
rect 6768 36880 6832 36944
rect 6848 36880 6912 36944
rect 6928 36880 6992 36944
rect 7008 36880 7072 36944
rect 7088 36880 7152 36944
rect 7168 36880 7232 36944
rect 7248 36880 7312 36944
rect 7328 36880 7392 36944
rect 7408 36880 7472 36944
rect 7488 36880 7552 36944
rect 7568 36880 7632 36944
rect 7648 36880 7712 36944
rect 7728 36880 7792 36944
rect 7808 36880 7872 36944
rect 7888 36880 7952 36944
rect 7968 36880 8032 36944
rect 8048 36880 8112 36944
rect 8128 36880 8192 36944
rect 8208 36880 8272 36944
rect 8288 36880 8352 36944
rect 8368 36880 8432 36944
rect 8448 36880 8512 36944
rect 8528 36880 8592 36944
rect 8608 36880 8672 36944
rect 8688 36880 8752 36944
rect 8768 36880 8832 36944
rect 8848 36880 8912 36944
rect 8928 36880 8992 36944
rect 14112 36880 14176 36944
rect 14192 36880 14256 36944
rect 14272 36880 14336 36944
rect 14352 36880 14416 36944
rect 24112 36880 24176 36944
rect 24192 36880 24256 36944
rect 24272 36880 24336 36944
rect 24352 36880 24416 36944
rect 36376 36880 36440 36944
rect 36456 36880 36520 36944
rect 36536 36880 36600 36944
rect 36616 36880 36680 36944
rect 36696 36880 36760 36944
rect 36776 36880 36840 36944
rect 36856 36880 36920 36944
rect 36936 36880 37000 36944
rect 37016 36880 37080 36944
rect 37096 36880 37160 36944
rect 37176 36880 37240 36944
rect 37256 36880 37320 36944
rect 37336 36880 37400 36944
rect 37416 36880 37480 36944
rect 37496 36880 37560 36944
rect 37576 36880 37640 36944
rect 37656 36880 37720 36944
rect 37736 36880 37800 36944
rect 37816 36880 37880 36944
rect 37896 36880 37960 36944
rect 37976 36880 38040 36944
rect 38056 36880 38120 36944
rect 38136 36880 38200 36944
rect 38216 36880 38280 36944
rect 38296 36880 38360 36944
rect 38376 36880 38440 36944
rect 38456 36880 38520 36944
rect 38536 36880 38600 36944
rect 38616 36880 38680 36944
rect 38696 36880 38760 36944
rect 38776 36880 38840 36944
rect 38856 36880 38920 36944
rect 38936 36880 39000 36944
rect 39016 36880 39080 36944
rect 39096 36880 39160 36944
rect 39176 36880 39240 36944
rect 39256 36880 39320 36944
rect 39336 36880 39400 36944
rect 39416 36880 39480 36944
rect 39496 36880 39560 36944
rect 39576 36880 39640 36944
rect 39656 36880 39720 36944
rect 39736 36880 39800 36944
rect 39816 36880 39880 36944
rect 39896 36880 39960 36944
rect 39976 36880 40040 36944
rect 40056 36880 40120 36944
rect 40136 36880 40200 36944
rect 40216 36880 40280 36944
rect 40296 36880 40360 36944
rect 5008 36800 5072 36864
rect 5088 36800 5152 36864
rect 5168 36800 5232 36864
rect 5248 36800 5312 36864
rect 5328 36800 5392 36864
rect 5408 36800 5472 36864
rect 5488 36800 5552 36864
rect 5568 36800 5632 36864
rect 5648 36800 5712 36864
rect 5728 36800 5792 36864
rect 5808 36800 5872 36864
rect 5888 36800 5952 36864
rect 5968 36800 6032 36864
rect 6048 36800 6112 36864
rect 6128 36800 6192 36864
rect 6208 36800 6272 36864
rect 6288 36800 6352 36864
rect 6368 36800 6432 36864
rect 6448 36800 6512 36864
rect 6528 36800 6592 36864
rect 6608 36800 6672 36864
rect 6688 36800 6752 36864
rect 6768 36800 6832 36864
rect 6848 36800 6912 36864
rect 6928 36800 6992 36864
rect 7008 36800 7072 36864
rect 7088 36800 7152 36864
rect 7168 36800 7232 36864
rect 7248 36800 7312 36864
rect 7328 36800 7392 36864
rect 7408 36800 7472 36864
rect 7488 36800 7552 36864
rect 7568 36800 7632 36864
rect 7648 36800 7712 36864
rect 7728 36800 7792 36864
rect 7808 36800 7872 36864
rect 7888 36800 7952 36864
rect 7968 36800 8032 36864
rect 8048 36800 8112 36864
rect 8128 36800 8192 36864
rect 8208 36800 8272 36864
rect 8288 36800 8352 36864
rect 8368 36800 8432 36864
rect 8448 36800 8512 36864
rect 8528 36800 8592 36864
rect 8608 36800 8672 36864
rect 8688 36800 8752 36864
rect 8768 36800 8832 36864
rect 8848 36800 8912 36864
rect 8928 36800 8992 36864
rect 14112 36800 14176 36864
rect 14192 36800 14256 36864
rect 14272 36800 14336 36864
rect 14352 36800 14416 36864
rect 24112 36800 24176 36864
rect 24192 36800 24256 36864
rect 24272 36800 24336 36864
rect 24352 36800 24416 36864
rect 36376 36800 36440 36864
rect 36456 36800 36520 36864
rect 36536 36800 36600 36864
rect 36616 36800 36680 36864
rect 36696 36800 36760 36864
rect 36776 36800 36840 36864
rect 36856 36800 36920 36864
rect 36936 36800 37000 36864
rect 37016 36800 37080 36864
rect 37096 36800 37160 36864
rect 37176 36800 37240 36864
rect 37256 36800 37320 36864
rect 37336 36800 37400 36864
rect 37416 36800 37480 36864
rect 37496 36800 37560 36864
rect 37576 36800 37640 36864
rect 37656 36800 37720 36864
rect 37736 36800 37800 36864
rect 37816 36800 37880 36864
rect 37896 36800 37960 36864
rect 37976 36800 38040 36864
rect 38056 36800 38120 36864
rect 38136 36800 38200 36864
rect 38216 36800 38280 36864
rect 38296 36800 38360 36864
rect 38376 36800 38440 36864
rect 38456 36800 38520 36864
rect 38536 36800 38600 36864
rect 38616 36800 38680 36864
rect 38696 36800 38760 36864
rect 38776 36800 38840 36864
rect 38856 36800 38920 36864
rect 38936 36800 39000 36864
rect 39016 36800 39080 36864
rect 39096 36800 39160 36864
rect 39176 36800 39240 36864
rect 39256 36800 39320 36864
rect 39336 36800 39400 36864
rect 39416 36800 39480 36864
rect 39496 36800 39560 36864
rect 39576 36800 39640 36864
rect 39656 36800 39720 36864
rect 39736 36800 39800 36864
rect 39816 36800 39880 36864
rect 39896 36800 39960 36864
rect 39976 36800 40040 36864
rect 40056 36800 40120 36864
rect 40136 36800 40200 36864
rect 40216 36800 40280 36864
rect 40296 36800 40360 36864
rect 5008 36720 5072 36784
rect 5088 36720 5152 36784
rect 5168 36720 5232 36784
rect 5248 36720 5312 36784
rect 5328 36720 5392 36784
rect 5408 36720 5472 36784
rect 5488 36720 5552 36784
rect 5568 36720 5632 36784
rect 5648 36720 5712 36784
rect 5728 36720 5792 36784
rect 5808 36720 5872 36784
rect 5888 36720 5952 36784
rect 5968 36720 6032 36784
rect 6048 36720 6112 36784
rect 6128 36720 6192 36784
rect 6208 36720 6272 36784
rect 6288 36720 6352 36784
rect 6368 36720 6432 36784
rect 6448 36720 6512 36784
rect 6528 36720 6592 36784
rect 6608 36720 6672 36784
rect 6688 36720 6752 36784
rect 6768 36720 6832 36784
rect 6848 36720 6912 36784
rect 6928 36720 6992 36784
rect 7008 36720 7072 36784
rect 7088 36720 7152 36784
rect 7168 36720 7232 36784
rect 7248 36720 7312 36784
rect 7328 36720 7392 36784
rect 7408 36720 7472 36784
rect 7488 36720 7552 36784
rect 7568 36720 7632 36784
rect 7648 36720 7712 36784
rect 7728 36720 7792 36784
rect 7808 36720 7872 36784
rect 7888 36720 7952 36784
rect 7968 36720 8032 36784
rect 8048 36720 8112 36784
rect 8128 36720 8192 36784
rect 8208 36720 8272 36784
rect 8288 36720 8352 36784
rect 8368 36720 8432 36784
rect 8448 36720 8512 36784
rect 8528 36720 8592 36784
rect 8608 36720 8672 36784
rect 8688 36720 8752 36784
rect 8768 36720 8832 36784
rect 8848 36720 8912 36784
rect 8928 36720 8992 36784
rect 14112 36720 14176 36784
rect 14192 36720 14256 36784
rect 14272 36720 14336 36784
rect 14352 36720 14416 36784
rect 24112 36720 24176 36784
rect 24192 36720 24256 36784
rect 24272 36720 24336 36784
rect 24352 36720 24416 36784
rect 36376 36720 36440 36784
rect 36456 36720 36520 36784
rect 36536 36720 36600 36784
rect 36616 36720 36680 36784
rect 36696 36720 36760 36784
rect 36776 36720 36840 36784
rect 36856 36720 36920 36784
rect 36936 36720 37000 36784
rect 37016 36720 37080 36784
rect 37096 36720 37160 36784
rect 37176 36720 37240 36784
rect 37256 36720 37320 36784
rect 37336 36720 37400 36784
rect 37416 36720 37480 36784
rect 37496 36720 37560 36784
rect 37576 36720 37640 36784
rect 37656 36720 37720 36784
rect 37736 36720 37800 36784
rect 37816 36720 37880 36784
rect 37896 36720 37960 36784
rect 37976 36720 38040 36784
rect 38056 36720 38120 36784
rect 38136 36720 38200 36784
rect 38216 36720 38280 36784
rect 38296 36720 38360 36784
rect 38376 36720 38440 36784
rect 38456 36720 38520 36784
rect 38536 36720 38600 36784
rect 38616 36720 38680 36784
rect 38696 36720 38760 36784
rect 38776 36720 38840 36784
rect 38856 36720 38920 36784
rect 38936 36720 39000 36784
rect 39016 36720 39080 36784
rect 39096 36720 39160 36784
rect 39176 36720 39240 36784
rect 39256 36720 39320 36784
rect 39336 36720 39400 36784
rect 39416 36720 39480 36784
rect 39496 36720 39560 36784
rect 39576 36720 39640 36784
rect 39656 36720 39720 36784
rect 39736 36720 39800 36784
rect 39816 36720 39880 36784
rect 39896 36720 39960 36784
rect 39976 36720 40040 36784
rect 40056 36720 40120 36784
rect 40136 36720 40200 36784
rect 40216 36720 40280 36784
rect 40296 36720 40360 36784
rect 5008 36640 5072 36704
rect 5088 36640 5152 36704
rect 5168 36640 5232 36704
rect 5248 36640 5312 36704
rect 5328 36640 5392 36704
rect 5408 36640 5472 36704
rect 5488 36640 5552 36704
rect 5568 36640 5632 36704
rect 5648 36640 5712 36704
rect 5728 36640 5792 36704
rect 5808 36640 5872 36704
rect 5888 36640 5952 36704
rect 5968 36640 6032 36704
rect 6048 36640 6112 36704
rect 6128 36640 6192 36704
rect 6208 36640 6272 36704
rect 6288 36640 6352 36704
rect 6368 36640 6432 36704
rect 6448 36640 6512 36704
rect 6528 36640 6592 36704
rect 6608 36640 6672 36704
rect 6688 36640 6752 36704
rect 6768 36640 6832 36704
rect 6848 36640 6912 36704
rect 6928 36640 6992 36704
rect 7008 36640 7072 36704
rect 7088 36640 7152 36704
rect 7168 36640 7232 36704
rect 7248 36640 7312 36704
rect 7328 36640 7392 36704
rect 7408 36640 7472 36704
rect 7488 36640 7552 36704
rect 7568 36640 7632 36704
rect 7648 36640 7712 36704
rect 7728 36640 7792 36704
rect 7808 36640 7872 36704
rect 7888 36640 7952 36704
rect 7968 36640 8032 36704
rect 8048 36640 8112 36704
rect 8128 36640 8192 36704
rect 8208 36640 8272 36704
rect 8288 36640 8352 36704
rect 8368 36640 8432 36704
rect 8448 36640 8512 36704
rect 8528 36640 8592 36704
rect 8608 36640 8672 36704
rect 8688 36640 8752 36704
rect 8768 36640 8832 36704
rect 8848 36640 8912 36704
rect 8928 36640 8992 36704
rect 14112 36640 14176 36704
rect 14192 36640 14256 36704
rect 14272 36640 14336 36704
rect 14352 36640 14416 36704
rect 24112 36640 24176 36704
rect 24192 36640 24256 36704
rect 24272 36640 24336 36704
rect 24352 36640 24416 36704
rect 36376 36640 36440 36704
rect 36456 36640 36520 36704
rect 36536 36640 36600 36704
rect 36616 36640 36680 36704
rect 36696 36640 36760 36704
rect 36776 36640 36840 36704
rect 36856 36640 36920 36704
rect 36936 36640 37000 36704
rect 37016 36640 37080 36704
rect 37096 36640 37160 36704
rect 37176 36640 37240 36704
rect 37256 36640 37320 36704
rect 37336 36640 37400 36704
rect 37416 36640 37480 36704
rect 37496 36640 37560 36704
rect 37576 36640 37640 36704
rect 37656 36640 37720 36704
rect 37736 36640 37800 36704
rect 37816 36640 37880 36704
rect 37896 36640 37960 36704
rect 37976 36640 38040 36704
rect 38056 36640 38120 36704
rect 38136 36640 38200 36704
rect 38216 36640 38280 36704
rect 38296 36640 38360 36704
rect 38376 36640 38440 36704
rect 38456 36640 38520 36704
rect 38536 36640 38600 36704
rect 38616 36640 38680 36704
rect 38696 36640 38760 36704
rect 38776 36640 38840 36704
rect 38856 36640 38920 36704
rect 38936 36640 39000 36704
rect 39016 36640 39080 36704
rect 39096 36640 39160 36704
rect 39176 36640 39240 36704
rect 39256 36640 39320 36704
rect 39336 36640 39400 36704
rect 39416 36640 39480 36704
rect 39496 36640 39560 36704
rect 39576 36640 39640 36704
rect 39656 36640 39720 36704
rect 39736 36640 39800 36704
rect 39816 36640 39880 36704
rect 39896 36640 39960 36704
rect 39976 36640 40040 36704
rect 40056 36640 40120 36704
rect 40136 36640 40200 36704
rect 40216 36640 40280 36704
rect 40296 36640 40360 36704
rect 5008 36560 5072 36624
rect 5088 36560 5152 36624
rect 5168 36560 5232 36624
rect 5248 36560 5312 36624
rect 5328 36560 5392 36624
rect 5408 36560 5472 36624
rect 5488 36560 5552 36624
rect 5568 36560 5632 36624
rect 5648 36560 5712 36624
rect 5728 36560 5792 36624
rect 5808 36560 5872 36624
rect 5888 36560 5952 36624
rect 5968 36560 6032 36624
rect 6048 36560 6112 36624
rect 6128 36560 6192 36624
rect 6208 36560 6272 36624
rect 6288 36560 6352 36624
rect 6368 36560 6432 36624
rect 6448 36560 6512 36624
rect 6528 36560 6592 36624
rect 6608 36560 6672 36624
rect 6688 36560 6752 36624
rect 6768 36560 6832 36624
rect 6848 36560 6912 36624
rect 6928 36560 6992 36624
rect 7008 36560 7072 36624
rect 7088 36560 7152 36624
rect 7168 36560 7232 36624
rect 7248 36560 7312 36624
rect 7328 36560 7392 36624
rect 7408 36560 7472 36624
rect 7488 36560 7552 36624
rect 7568 36560 7632 36624
rect 7648 36560 7712 36624
rect 7728 36560 7792 36624
rect 7808 36560 7872 36624
rect 7888 36560 7952 36624
rect 7968 36560 8032 36624
rect 8048 36560 8112 36624
rect 8128 36560 8192 36624
rect 8208 36560 8272 36624
rect 8288 36560 8352 36624
rect 8368 36560 8432 36624
rect 8448 36560 8512 36624
rect 8528 36560 8592 36624
rect 8608 36560 8672 36624
rect 8688 36560 8752 36624
rect 8768 36560 8832 36624
rect 8848 36560 8912 36624
rect 8928 36560 8992 36624
rect 14112 36560 14176 36624
rect 14192 36560 14256 36624
rect 14272 36560 14336 36624
rect 14352 36560 14416 36624
rect 24112 36560 24176 36624
rect 24192 36560 24256 36624
rect 24272 36560 24336 36624
rect 24352 36560 24416 36624
rect 36376 36560 36440 36624
rect 36456 36560 36520 36624
rect 36536 36560 36600 36624
rect 36616 36560 36680 36624
rect 36696 36560 36760 36624
rect 36776 36560 36840 36624
rect 36856 36560 36920 36624
rect 36936 36560 37000 36624
rect 37016 36560 37080 36624
rect 37096 36560 37160 36624
rect 37176 36560 37240 36624
rect 37256 36560 37320 36624
rect 37336 36560 37400 36624
rect 37416 36560 37480 36624
rect 37496 36560 37560 36624
rect 37576 36560 37640 36624
rect 37656 36560 37720 36624
rect 37736 36560 37800 36624
rect 37816 36560 37880 36624
rect 37896 36560 37960 36624
rect 37976 36560 38040 36624
rect 38056 36560 38120 36624
rect 38136 36560 38200 36624
rect 38216 36560 38280 36624
rect 38296 36560 38360 36624
rect 38376 36560 38440 36624
rect 38456 36560 38520 36624
rect 38536 36560 38600 36624
rect 38616 36560 38680 36624
rect 38696 36560 38760 36624
rect 38776 36560 38840 36624
rect 38856 36560 38920 36624
rect 38936 36560 39000 36624
rect 39016 36560 39080 36624
rect 39096 36560 39160 36624
rect 39176 36560 39240 36624
rect 39256 36560 39320 36624
rect 39336 36560 39400 36624
rect 39416 36560 39480 36624
rect 39496 36560 39560 36624
rect 39576 36560 39640 36624
rect 39656 36560 39720 36624
rect 39736 36560 39800 36624
rect 39816 36560 39880 36624
rect 39896 36560 39960 36624
rect 39976 36560 40040 36624
rect 40056 36560 40120 36624
rect 40136 36560 40200 36624
rect 40216 36560 40280 36624
rect 40296 36560 40360 36624
rect 5008 36480 5072 36544
rect 5088 36480 5152 36544
rect 5168 36480 5232 36544
rect 5248 36480 5312 36544
rect 5328 36480 5392 36544
rect 5408 36480 5472 36544
rect 5488 36480 5552 36544
rect 5568 36480 5632 36544
rect 5648 36480 5712 36544
rect 5728 36480 5792 36544
rect 5808 36480 5872 36544
rect 5888 36480 5952 36544
rect 5968 36480 6032 36544
rect 6048 36480 6112 36544
rect 6128 36480 6192 36544
rect 6208 36480 6272 36544
rect 6288 36480 6352 36544
rect 6368 36480 6432 36544
rect 6448 36480 6512 36544
rect 6528 36480 6592 36544
rect 6608 36480 6672 36544
rect 6688 36480 6752 36544
rect 6768 36480 6832 36544
rect 6848 36480 6912 36544
rect 6928 36480 6992 36544
rect 7008 36480 7072 36544
rect 7088 36480 7152 36544
rect 7168 36480 7232 36544
rect 7248 36480 7312 36544
rect 7328 36480 7392 36544
rect 7408 36480 7472 36544
rect 7488 36480 7552 36544
rect 7568 36480 7632 36544
rect 7648 36480 7712 36544
rect 7728 36480 7792 36544
rect 7808 36480 7872 36544
rect 7888 36480 7952 36544
rect 7968 36480 8032 36544
rect 8048 36480 8112 36544
rect 8128 36480 8192 36544
rect 8208 36480 8272 36544
rect 8288 36480 8352 36544
rect 8368 36480 8432 36544
rect 8448 36480 8512 36544
rect 8528 36480 8592 36544
rect 8608 36480 8672 36544
rect 8688 36480 8752 36544
rect 8768 36480 8832 36544
rect 8848 36480 8912 36544
rect 8928 36480 8992 36544
rect 14112 36480 14176 36544
rect 14192 36480 14256 36544
rect 14272 36480 14336 36544
rect 14352 36480 14416 36544
rect 24112 36480 24176 36544
rect 24192 36480 24256 36544
rect 24272 36480 24336 36544
rect 24352 36480 24416 36544
rect 36376 36480 36440 36544
rect 36456 36480 36520 36544
rect 36536 36480 36600 36544
rect 36616 36480 36680 36544
rect 36696 36480 36760 36544
rect 36776 36480 36840 36544
rect 36856 36480 36920 36544
rect 36936 36480 37000 36544
rect 37016 36480 37080 36544
rect 37096 36480 37160 36544
rect 37176 36480 37240 36544
rect 37256 36480 37320 36544
rect 37336 36480 37400 36544
rect 37416 36480 37480 36544
rect 37496 36480 37560 36544
rect 37576 36480 37640 36544
rect 37656 36480 37720 36544
rect 37736 36480 37800 36544
rect 37816 36480 37880 36544
rect 37896 36480 37960 36544
rect 37976 36480 38040 36544
rect 38056 36480 38120 36544
rect 38136 36480 38200 36544
rect 38216 36480 38280 36544
rect 38296 36480 38360 36544
rect 38376 36480 38440 36544
rect 38456 36480 38520 36544
rect 38536 36480 38600 36544
rect 38616 36480 38680 36544
rect 38696 36480 38760 36544
rect 38776 36480 38840 36544
rect 38856 36480 38920 36544
rect 38936 36480 39000 36544
rect 39016 36480 39080 36544
rect 39096 36480 39160 36544
rect 39176 36480 39240 36544
rect 39256 36480 39320 36544
rect 39336 36480 39400 36544
rect 39416 36480 39480 36544
rect 39496 36480 39560 36544
rect 39576 36480 39640 36544
rect 39656 36480 39720 36544
rect 39736 36480 39800 36544
rect 39816 36480 39880 36544
rect 39896 36480 39960 36544
rect 39976 36480 40040 36544
rect 40056 36480 40120 36544
rect 40136 36480 40200 36544
rect 40216 36480 40280 36544
rect 40296 36480 40360 36544
rect 5008 36400 5072 36464
rect 5088 36400 5152 36464
rect 5168 36400 5232 36464
rect 5248 36400 5312 36464
rect 5328 36400 5392 36464
rect 5408 36400 5472 36464
rect 5488 36400 5552 36464
rect 5568 36400 5632 36464
rect 5648 36400 5712 36464
rect 5728 36400 5792 36464
rect 5808 36400 5872 36464
rect 5888 36400 5952 36464
rect 5968 36400 6032 36464
rect 6048 36400 6112 36464
rect 6128 36400 6192 36464
rect 6208 36400 6272 36464
rect 6288 36400 6352 36464
rect 6368 36400 6432 36464
rect 6448 36400 6512 36464
rect 6528 36400 6592 36464
rect 6608 36400 6672 36464
rect 6688 36400 6752 36464
rect 6768 36400 6832 36464
rect 6848 36400 6912 36464
rect 6928 36400 6992 36464
rect 7008 36400 7072 36464
rect 7088 36400 7152 36464
rect 7168 36400 7232 36464
rect 7248 36400 7312 36464
rect 7328 36400 7392 36464
rect 7408 36400 7472 36464
rect 7488 36400 7552 36464
rect 7568 36400 7632 36464
rect 7648 36400 7712 36464
rect 7728 36400 7792 36464
rect 7808 36400 7872 36464
rect 7888 36400 7952 36464
rect 7968 36400 8032 36464
rect 8048 36400 8112 36464
rect 8128 36400 8192 36464
rect 8208 36400 8272 36464
rect 8288 36400 8352 36464
rect 8368 36400 8432 36464
rect 8448 36400 8512 36464
rect 8528 36400 8592 36464
rect 8608 36400 8672 36464
rect 8688 36400 8752 36464
rect 8768 36400 8832 36464
rect 8848 36400 8912 36464
rect 8928 36400 8992 36464
rect 14112 36400 14176 36464
rect 14192 36400 14256 36464
rect 14272 36400 14336 36464
rect 14352 36400 14416 36464
rect 24112 36400 24176 36464
rect 24192 36400 24256 36464
rect 24272 36400 24336 36464
rect 24352 36400 24416 36464
rect 36376 36400 36440 36464
rect 36456 36400 36520 36464
rect 36536 36400 36600 36464
rect 36616 36400 36680 36464
rect 36696 36400 36760 36464
rect 36776 36400 36840 36464
rect 36856 36400 36920 36464
rect 36936 36400 37000 36464
rect 37016 36400 37080 36464
rect 37096 36400 37160 36464
rect 37176 36400 37240 36464
rect 37256 36400 37320 36464
rect 37336 36400 37400 36464
rect 37416 36400 37480 36464
rect 37496 36400 37560 36464
rect 37576 36400 37640 36464
rect 37656 36400 37720 36464
rect 37736 36400 37800 36464
rect 37816 36400 37880 36464
rect 37896 36400 37960 36464
rect 37976 36400 38040 36464
rect 38056 36400 38120 36464
rect 38136 36400 38200 36464
rect 38216 36400 38280 36464
rect 38296 36400 38360 36464
rect 38376 36400 38440 36464
rect 38456 36400 38520 36464
rect 38536 36400 38600 36464
rect 38616 36400 38680 36464
rect 38696 36400 38760 36464
rect 38776 36400 38840 36464
rect 38856 36400 38920 36464
rect 38936 36400 39000 36464
rect 39016 36400 39080 36464
rect 39096 36400 39160 36464
rect 39176 36400 39240 36464
rect 39256 36400 39320 36464
rect 39336 36400 39400 36464
rect 39416 36400 39480 36464
rect 39496 36400 39560 36464
rect 39576 36400 39640 36464
rect 39656 36400 39720 36464
rect 39736 36400 39800 36464
rect 39816 36400 39880 36464
rect 39896 36400 39960 36464
rect 39976 36400 40040 36464
rect 40056 36400 40120 36464
rect 40136 36400 40200 36464
rect 40216 36400 40280 36464
rect 40296 36400 40360 36464
rect 19112 34420 19176 34424
rect 19112 34364 19116 34420
rect 19116 34364 19172 34420
rect 19172 34364 19176 34420
rect 19112 34360 19176 34364
rect 19192 34420 19256 34424
rect 19192 34364 19196 34420
rect 19196 34364 19252 34420
rect 19252 34364 19256 34420
rect 19192 34360 19256 34364
rect 19272 34420 19336 34424
rect 19272 34364 19276 34420
rect 19276 34364 19332 34420
rect 19332 34364 19336 34420
rect 19272 34360 19336 34364
rect 19352 34420 19416 34424
rect 19352 34364 19356 34420
rect 19356 34364 19412 34420
rect 19412 34364 19416 34420
rect 19352 34360 19416 34364
rect 29112 34420 29176 34424
rect 29112 34364 29116 34420
rect 29116 34364 29172 34420
rect 29172 34364 29176 34420
rect 29112 34360 29176 34364
rect 29192 34420 29256 34424
rect 29192 34364 29196 34420
rect 29196 34364 29252 34420
rect 29252 34364 29256 34420
rect 29192 34360 29256 34364
rect 29272 34420 29336 34424
rect 29272 34364 29276 34420
rect 29276 34364 29332 34420
rect 29332 34364 29336 34420
rect 29272 34360 29336 34364
rect 29352 34420 29416 34424
rect 29352 34364 29356 34420
rect 29356 34364 29412 34420
rect 29412 34364 29416 34420
rect 29352 34360 29416 34364
rect 14112 33876 14176 33880
rect 14112 33820 14116 33876
rect 14116 33820 14172 33876
rect 14172 33820 14176 33876
rect 14112 33816 14176 33820
rect 14192 33876 14256 33880
rect 14192 33820 14196 33876
rect 14196 33820 14252 33876
rect 14252 33820 14256 33876
rect 14192 33816 14256 33820
rect 14272 33876 14336 33880
rect 14272 33820 14276 33876
rect 14276 33820 14332 33876
rect 14332 33820 14336 33876
rect 14272 33816 14336 33820
rect 14352 33876 14416 33880
rect 14352 33820 14356 33876
rect 14356 33820 14412 33876
rect 14412 33820 14416 33876
rect 14352 33816 14416 33820
rect 24112 33876 24176 33880
rect 24112 33820 24116 33876
rect 24116 33820 24172 33876
rect 24172 33820 24176 33876
rect 24112 33816 24176 33820
rect 24192 33876 24256 33880
rect 24192 33820 24196 33876
rect 24196 33820 24252 33876
rect 24252 33820 24256 33876
rect 24192 33816 24256 33820
rect 24272 33876 24336 33880
rect 24272 33820 24276 33876
rect 24276 33820 24332 33876
rect 24332 33820 24336 33876
rect 24272 33816 24336 33820
rect 24352 33876 24416 33880
rect 24352 33820 24356 33876
rect 24356 33820 24412 33876
rect 24412 33820 24416 33876
rect 24352 33816 24416 33820
rect 19112 33332 19176 33336
rect 19112 33276 19116 33332
rect 19116 33276 19172 33332
rect 19172 33276 19176 33332
rect 19112 33272 19176 33276
rect 19192 33332 19256 33336
rect 19192 33276 19196 33332
rect 19196 33276 19252 33332
rect 19252 33276 19256 33332
rect 19192 33272 19256 33276
rect 19272 33332 19336 33336
rect 19272 33276 19276 33332
rect 19276 33276 19332 33332
rect 19332 33276 19336 33332
rect 19272 33272 19336 33276
rect 19352 33332 19416 33336
rect 19352 33276 19356 33332
rect 19356 33276 19412 33332
rect 19412 33276 19416 33332
rect 19352 33272 19416 33276
rect 29112 33332 29176 33336
rect 29112 33276 29116 33332
rect 29116 33276 29172 33332
rect 29172 33276 29176 33332
rect 29112 33272 29176 33276
rect 29192 33332 29256 33336
rect 29192 33276 29196 33332
rect 29196 33276 29252 33332
rect 29252 33276 29256 33332
rect 29192 33272 29256 33276
rect 29272 33332 29336 33336
rect 29272 33276 29276 33332
rect 29276 33276 29332 33332
rect 29332 33276 29336 33332
rect 29272 33272 29336 33276
rect 29352 33332 29416 33336
rect 29352 33276 29356 33332
rect 29356 33276 29412 33332
rect 29412 33276 29416 33332
rect 29352 33272 29416 33276
rect 14112 32788 14176 32792
rect 14112 32732 14116 32788
rect 14116 32732 14172 32788
rect 14172 32732 14176 32788
rect 14112 32728 14176 32732
rect 14192 32788 14256 32792
rect 14192 32732 14196 32788
rect 14196 32732 14252 32788
rect 14252 32732 14256 32788
rect 14192 32728 14256 32732
rect 14272 32788 14336 32792
rect 14272 32732 14276 32788
rect 14276 32732 14332 32788
rect 14332 32732 14336 32788
rect 14272 32728 14336 32732
rect 14352 32788 14416 32792
rect 14352 32732 14356 32788
rect 14356 32732 14412 32788
rect 14412 32732 14416 32788
rect 14352 32728 14416 32732
rect 24112 32788 24176 32792
rect 24112 32732 24116 32788
rect 24116 32732 24172 32788
rect 24172 32732 24176 32788
rect 24112 32728 24176 32732
rect 24192 32788 24256 32792
rect 24192 32732 24196 32788
rect 24196 32732 24252 32788
rect 24252 32732 24256 32788
rect 24192 32728 24256 32732
rect 24272 32788 24336 32792
rect 24272 32732 24276 32788
rect 24276 32732 24332 32788
rect 24332 32732 24336 32788
rect 24272 32728 24336 32732
rect 24352 32788 24416 32792
rect 24352 32732 24356 32788
rect 24356 32732 24412 32788
rect 24412 32732 24416 32788
rect 24352 32728 24416 32732
rect 19112 32244 19176 32248
rect 19112 32188 19116 32244
rect 19116 32188 19172 32244
rect 19172 32188 19176 32244
rect 19112 32184 19176 32188
rect 19192 32244 19256 32248
rect 19192 32188 19196 32244
rect 19196 32188 19252 32244
rect 19252 32188 19256 32244
rect 19192 32184 19256 32188
rect 19272 32244 19336 32248
rect 19272 32188 19276 32244
rect 19276 32188 19332 32244
rect 19332 32188 19336 32244
rect 19272 32184 19336 32188
rect 19352 32244 19416 32248
rect 19352 32188 19356 32244
rect 19356 32188 19412 32244
rect 19412 32188 19416 32244
rect 19352 32184 19416 32188
rect 29112 32244 29176 32248
rect 29112 32188 29116 32244
rect 29116 32188 29172 32244
rect 29172 32188 29176 32244
rect 29112 32184 29176 32188
rect 29192 32244 29256 32248
rect 29192 32188 29196 32244
rect 29196 32188 29252 32244
rect 29252 32188 29256 32244
rect 29192 32184 29256 32188
rect 29272 32244 29336 32248
rect 29272 32188 29276 32244
rect 29276 32188 29332 32244
rect 29332 32188 29336 32244
rect 29272 32184 29336 32188
rect 29352 32244 29416 32248
rect 29352 32188 29356 32244
rect 29356 32188 29412 32244
rect 29412 32188 29416 32244
rect 29352 32184 29416 32188
rect 14112 31700 14176 31704
rect 14112 31644 14116 31700
rect 14116 31644 14172 31700
rect 14172 31644 14176 31700
rect 14112 31640 14176 31644
rect 14192 31700 14256 31704
rect 14192 31644 14196 31700
rect 14196 31644 14252 31700
rect 14252 31644 14256 31700
rect 14192 31640 14256 31644
rect 14272 31700 14336 31704
rect 14272 31644 14276 31700
rect 14276 31644 14332 31700
rect 14332 31644 14336 31700
rect 14272 31640 14336 31644
rect 14352 31700 14416 31704
rect 14352 31644 14356 31700
rect 14356 31644 14412 31700
rect 14412 31644 14416 31700
rect 14352 31640 14416 31644
rect 24112 31700 24176 31704
rect 24112 31644 24116 31700
rect 24116 31644 24172 31700
rect 24172 31644 24176 31700
rect 24112 31640 24176 31644
rect 24192 31700 24256 31704
rect 24192 31644 24196 31700
rect 24196 31644 24252 31700
rect 24252 31644 24256 31700
rect 24192 31640 24256 31644
rect 24272 31700 24336 31704
rect 24272 31644 24276 31700
rect 24276 31644 24332 31700
rect 24332 31644 24336 31700
rect 24272 31640 24336 31644
rect 24352 31700 24416 31704
rect 24352 31644 24356 31700
rect 24356 31644 24412 31700
rect 24412 31644 24416 31700
rect 24352 31640 24416 31644
rect 19112 31156 19176 31160
rect 19112 31100 19116 31156
rect 19116 31100 19172 31156
rect 19172 31100 19176 31156
rect 19112 31096 19176 31100
rect 19192 31156 19256 31160
rect 19192 31100 19196 31156
rect 19196 31100 19252 31156
rect 19252 31100 19256 31156
rect 19192 31096 19256 31100
rect 19272 31156 19336 31160
rect 19272 31100 19276 31156
rect 19276 31100 19332 31156
rect 19332 31100 19336 31156
rect 19272 31096 19336 31100
rect 19352 31156 19416 31160
rect 19352 31100 19356 31156
rect 19356 31100 19412 31156
rect 19412 31100 19416 31156
rect 19352 31096 19416 31100
rect 29112 31156 29176 31160
rect 29112 31100 29116 31156
rect 29116 31100 29172 31156
rect 29172 31100 29176 31156
rect 29112 31096 29176 31100
rect 29192 31156 29256 31160
rect 29192 31100 29196 31156
rect 29196 31100 29252 31156
rect 29252 31100 29256 31156
rect 29192 31096 29256 31100
rect 29272 31156 29336 31160
rect 29272 31100 29276 31156
rect 29276 31100 29332 31156
rect 29332 31100 29336 31156
rect 29272 31096 29336 31100
rect 29352 31156 29416 31160
rect 29352 31100 29356 31156
rect 29356 31100 29412 31156
rect 29412 31100 29416 31156
rect 29352 31096 29416 31100
rect 14112 30612 14176 30616
rect 14112 30556 14116 30612
rect 14116 30556 14172 30612
rect 14172 30556 14176 30612
rect 14112 30552 14176 30556
rect 14192 30612 14256 30616
rect 14192 30556 14196 30612
rect 14196 30556 14252 30612
rect 14252 30556 14256 30612
rect 14192 30552 14256 30556
rect 14272 30612 14336 30616
rect 14272 30556 14276 30612
rect 14276 30556 14332 30612
rect 14332 30556 14336 30612
rect 14272 30552 14336 30556
rect 14352 30612 14416 30616
rect 14352 30556 14356 30612
rect 14356 30556 14412 30612
rect 14412 30556 14416 30612
rect 14352 30552 14416 30556
rect 24112 30612 24176 30616
rect 24112 30556 24116 30612
rect 24116 30556 24172 30612
rect 24172 30556 24176 30612
rect 24112 30552 24176 30556
rect 24192 30612 24256 30616
rect 24192 30556 24196 30612
rect 24196 30556 24252 30612
rect 24252 30556 24256 30612
rect 24192 30552 24256 30556
rect 24272 30612 24336 30616
rect 24272 30556 24276 30612
rect 24276 30556 24332 30612
rect 24332 30556 24336 30612
rect 24272 30552 24336 30556
rect 24352 30612 24416 30616
rect 24352 30556 24356 30612
rect 24356 30556 24412 30612
rect 24412 30556 24416 30612
rect 24352 30552 24416 30556
rect 19112 30068 19176 30072
rect 19112 30012 19116 30068
rect 19116 30012 19172 30068
rect 19172 30012 19176 30068
rect 19112 30008 19176 30012
rect 19192 30068 19256 30072
rect 19192 30012 19196 30068
rect 19196 30012 19252 30068
rect 19252 30012 19256 30068
rect 19192 30008 19256 30012
rect 19272 30068 19336 30072
rect 19272 30012 19276 30068
rect 19276 30012 19332 30068
rect 19332 30012 19336 30068
rect 19272 30008 19336 30012
rect 19352 30068 19416 30072
rect 19352 30012 19356 30068
rect 19356 30012 19412 30068
rect 19412 30012 19416 30068
rect 19352 30008 19416 30012
rect 29112 30068 29176 30072
rect 29112 30012 29116 30068
rect 29116 30012 29172 30068
rect 29172 30012 29176 30068
rect 29112 30008 29176 30012
rect 29192 30068 29256 30072
rect 29192 30012 29196 30068
rect 29196 30012 29252 30068
rect 29252 30012 29256 30068
rect 29192 30008 29256 30012
rect 29272 30068 29336 30072
rect 29272 30012 29276 30068
rect 29276 30012 29332 30068
rect 29332 30012 29336 30068
rect 29272 30008 29336 30012
rect 29352 30068 29416 30072
rect 29352 30012 29356 30068
rect 29356 30012 29412 30068
rect 29412 30012 29416 30068
rect 29352 30008 29416 30012
rect 14112 29524 14176 29528
rect 14112 29468 14116 29524
rect 14116 29468 14172 29524
rect 14172 29468 14176 29524
rect 14112 29464 14176 29468
rect 14192 29524 14256 29528
rect 14192 29468 14196 29524
rect 14196 29468 14252 29524
rect 14252 29468 14256 29524
rect 14192 29464 14256 29468
rect 14272 29524 14336 29528
rect 14272 29468 14276 29524
rect 14276 29468 14332 29524
rect 14332 29468 14336 29524
rect 14272 29464 14336 29468
rect 14352 29524 14416 29528
rect 14352 29468 14356 29524
rect 14356 29468 14412 29524
rect 14412 29468 14416 29524
rect 14352 29464 14416 29468
rect 24112 29524 24176 29528
rect 24112 29468 24116 29524
rect 24116 29468 24172 29524
rect 24172 29468 24176 29524
rect 24112 29464 24176 29468
rect 24192 29524 24256 29528
rect 24192 29468 24196 29524
rect 24196 29468 24252 29524
rect 24252 29468 24256 29524
rect 24192 29464 24256 29468
rect 24272 29524 24336 29528
rect 24272 29468 24276 29524
rect 24276 29468 24332 29524
rect 24332 29468 24336 29524
rect 24272 29464 24336 29468
rect 24352 29524 24416 29528
rect 24352 29468 24356 29524
rect 24356 29468 24412 29524
rect 24412 29468 24416 29524
rect 24352 29464 24416 29468
rect 19112 28980 19176 28984
rect 19112 28924 19116 28980
rect 19116 28924 19172 28980
rect 19172 28924 19176 28980
rect 19112 28920 19176 28924
rect 19192 28980 19256 28984
rect 19192 28924 19196 28980
rect 19196 28924 19252 28980
rect 19252 28924 19256 28980
rect 19192 28920 19256 28924
rect 19272 28980 19336 28984
rect 19272 28924 19276 28980
rect 19276 28924 19332 28980
rect 19332 28924 19336 28980
rect 19272 28920 19336 28924
rect 19352 28980 19416 28984
rect 19352 28924 19356 28980
rect 19356 28924 19412 28980
rect 19412 28924 19416 28980
rect 19352 28920 19416 28924
rect 29112 28980 29176 28984
rect 29112 28924 29116 28980
rect 29116 28924 29172 28980
rect 29172 28924 29176 28980
rect 29112 28920 29176 28924
rect 29192 28980 29256 28984
rect 29192 28924 29196 28980
rect 29196 28924 29252 28980
rect 29252 28924 29256 28980
rect 29192 28920 29256 28924
rect 29272 28980 29336 28984
rect 29272 28924 29276 28980
rect 29276 28924 29332 28980
rect 29332 28924 29336 28980
rect 29272 28920 29336 28924
rect 29352 28980 29416 28984
rect 29352 28924 29356 28980
rect 29356 28924 29412 28980
rect 29412 28924 29416 28980
rect 29352 28920 29416 28924
rect 14112 28436 14176 28440
rect 14112 28380 14116 28436
rect 14116 28380 14172 28436
rect 14172 28380 14176 28436
rect 14112 28376 14176 28380
rect 14192 28436 14256 28440
rect 14192 28380 14196 28436
rect 14196 28380 14252 28436
rect 14252 28380 14256 28436
rect 14192 28376 14256 28380
rect 14272 28436 14336 28440
rect 14272 28380 14276 28436
rect 14276 28380 14332 28436
rect 14332 28380 14336 28436
rect 14272 28376 14336 28380
rect 14352 28436 14416 28440
rect 14352 28380 14356 28436
rect 14356 28380 14412 28436
rect 14412 28380 14416 28436
rect 14352 28376 14416 28380
rect 24112 28436 24176 28440
rect 24112 28380 24116 28436
rect 24116 28380 24172 28436
rect 24172 28380 24176 28436
rect 24112 28376 24176 28380
rect 24192 28436 24256 28440
rect 24192 28380 24196 28436
rect 24196 28380 24252 28436
rect 24252 28380 24256 28436
rect 24192 28376 24256 28380
rect 24272 28436 24336 28440
rect 24272 28380 24276 28436
rect 24276 28380 24332 28436
rect 24332 28380 24336 28436
rect 24272 28376 24336 28380
rect 24352 28436 24416 28440
rect 24352 28380 24356 28436
rect 24356 28380 24412 28436
rect 24412 28380 24416 28436
rect 24352 28376 24416 28380
rect 19112 27892 19176 27896
rect 19112 27836 19116 27892
rect 19116 27836 19172 27892
rect 19172 27836 19176 27892
rect 19112 27832 19176 27836
rect 19192 27892 19256 27896
rect 19192 27836 19196 27892
rect 19196 27836 19252 27892
rect 19252 27836 19256 27892
rect 19192 27832 19256 27836
rect 19272 27892 19336 27896
rect 19272 27836 19276 27892
rect 19276 27836 19332 27892
rect 19332 27836 19336 27892
rect 19272 27832 19336 27836
rect 19352 27892 19416 27896
rect 19352 27836 19356 27892
rect 19356 27836 19412 27892
rect 19412 27836 19416 27892
rect 19352 27832 19416 27836
rect 29112 27892 29176 27896
rect 29112 27836 29116 27892
rect 29116 27836 29172 27892
rect 29172 27836 29176 27892
rect 29112 27832 29176 27836
rect 29192 27892 29256 27896
rect 29192 27836 29196 27892
rect 29196 27836 29252 27892
rect 29252 27836 29256 27892
rect 29192 27832 29256 27836
rect 29272 27892 29336 27896
rect 29272 27836 29276 27892
rect 29276 27836 29332 27892
rect 29332 27836 29336 27892
rect 29272 27832 29336 27836
rect 29352 27892 29416 27896
rect 29352 27836 29356 27892
rect 29356 27836 29412 27892
rect 29412 27836 29416 27892
rect 29352 27832 29416 27836
rect 14112 27348 14176 27352
rect 14112 27292 14116 27348
rect 14116 27292 14172 27348
rect 14172 27292 14176 27348
rect 14112 27288 14176 27292
rect 14192 27348 14256 27352
rect 14192 27292 14196 27348
rect 14196 27292 14252 27348
rect 14252 27292 14256 27348
rect 14192 27288 14256 27292
rect 14272 27348 14336 27352
rect 14272 27292 14276 27348
rect 14276 27292 14332 27348
rect 14332 27292 14336 27348
rect 14272 27288 14336 27292
rect 14352 27348 14416 27352
rect 14352 27292 14356 27348
rect 14356 27292 14412 27348
rect 14412 27292 14416 27348
rect 14352 27288 14416 27292
rect 24112 27348 24176 27352
rect 24112 27292 24116 27348
rect 24116 27292 24172 27348
rect 24172 27292 24176 27348
rect 24112 27288 24176 27292
rect 24192 27348 24256 27352
rect 24192 27292 24196 27348
rect 24196 27292 24252 27348
rect 24252 27292 24256 27348
rect 24192 27288 24256 27292
rect 24272 27348 24336 27352
rect 24272 27292 24276 27348
rect 24276 27292 24332 27348
rect 24332 27292 24336 27348
rect 24272 27288 24336 27292
rect 24352 27348 24416 27352
rect 24352 27292 24356 27348
rect 24356 27292 24412 27348
rect 24412 27292 24416 27348
rect 24352 27288 24416 27292
rect 19112 26804 19176 26808
rect 19112 26748 19116 26804
rect 19116 26748 19172 26804
rect 19172 26748 19176 26804
rect 19112 26744 19176 26748
rect 19192 26804 19256 26808
rect 19192 26748 19196 26804
rect 19196 26748 19252 26804
rect 19252 26748 19256 26804
rect 19192 26744 19256 26748
rect 19272 26804 19336 26808
rect 19272 26748 19276 26804
rect 19276 26748 19332 26804
rect 19332 26748 19336 26804
rect 19272 26744 19336 26748
rect 19352 26804 19416 26808
rect 19352 26748 19356 26804
rect 19356 26748 19412 26804
rect 19412 26748 19416 26804
rect 19352 26744 19416 26748
rect 29112 26804 29176 26808
rect 29112 26748 29116 26804
rect 29116 26748 29172 26804
rect 29172 26748 29176 26804
rect 29112 26744 29176 26748
rect 29192 26804 29256 26808
rect 29192 26748 29196 26804
rect 29196 26748 29252 26804
rect 29252 26748 29256 26804
rect 29192 26744 29256 26748
rect 29272 26804 29336 26808
rect 29272 26748 29276 26804
rect 29276 26748 29332 26804
rect 29332 26748 29336 26804
rect 29272 26744 29336 26748
rect 29352 26804 29416 26808
rect 29352 26748 29356 26804
rect 29356 26748 29412 26804
rect 29412 26748 29416 26804
rect 29352 26744 29416 26748
rect 14112 26260 14176 26264
rect 14112 26204 14116 26260
rect 14116 26204 14172 26260
rect 14172 26204 14176 26260
rect 14112 26200 14176 26204
rect 14192 26260 14256 26264
rect 14192 26204 14196 26260
rect 14196 26204 14252 26260
rect 14252 26204 14256 26260
rect 14192 26200 14256 26204
rect 14272 26260 14336 26264
rect 14272 26204 14276 26260
rect 14276 26204 14332 26260
rect 14332 26204 14336 26260
rect 14272 26200 14336 26204
rect 14352 26260 14416 26264
rect 14352 26204 14356 26260
rect 14356 26204 14412 26260
rect 14412 26204 14416 26260
rect 14352 26200 14416 26204
rect 24112 26260 24176 26264
rect 24112 26204 24116 26260
rect 24116 26204 24172 26260
rect 24172 26204 24176 26260
rect 24112 26200 24176 26204
rect 24192 26260 24256 26264
rect 24192 26204 24196 26260
rect 24196 26204 24252 26260
rect 24252 26204 24256 26260
rect 24192 26200 24256 26204
rect 24272 26260 24336 26264
rect 24272 26204 24276 26260
rect 24276 26204 24332 26260
rect 24332 26204 24336 26260
rect 24272 26200 24336 26204
rect 24352 26260 24416 26264
rect 24352 26204 24356 26260
rect 24356 26204 24412 26260
rect 24412 26204 24416 26260
rect 24352 26200 24416 26204
rect 19112 25716 19176 25720
rect 19112 25660 19116 25716
rect 19116 25660 19172 25716
rect 19172 25660 19176 25716
rect 19112 25656 19176 25660
rect 19192 25716 19256 25720
rect 19192 25660 19196 25716
rect 19196 25660 19252 25716
rect 19252 25660 19256 25716
rect 19192 25656 19256 25660
rect 19272 25716 19336 25720
rect 19272 25660 19276 25716
rect 19276 25660 19332 25716
rect 19332 25660 19336 25716
rect 19272 25656 19336 25660
rect 19352 25716 19416 25720
rect 19352 25660 19356 25716
rect 19356 25660 19412 25716
rect 19412 25660 19416 25716
rect 19352 25656 19416 25660
rect 29112 25716 29176 25720
rect 29112 25660 29116 25716
rect 29116 25660 29172 25716
rect 29172 25660 29176 25716
rect 29112 25656 29176 25660
rect 29192 25716 29256 25720
rect 29192 25660 29196 25716
rect 29196 25660 29252 25716
rect 29252 25660 29256 25716
rect 29192 25656 29256 25660
rect 29272 25716 29336 25720
rect 29272 25660 29276 25716
rect 29276 25660 29332 25716
rect 29332 25660 29336 25716
rect 29272 25656 29336 25660
rect 29352 25716 29416 25720
rect 29352 25660 29356 25716
rect 29356 25660 29412 25716
rect 29412 25660 29416 25716
rect 29352 25656 29416 25660
rect 14112 25172 14176 25176
rect 14112 25116 14116 25172
rect 14116 25116 14172 25172
rect 14172 25116 14176 25172
rect 14112 25112 14176 25116
rect 14192 25172 14256 25176
rect 14192 25116 14196 25172
rect 14196 25116 14252 25172
rect 14252 25116 14256 25172
rect 14192 25112 14256 25116
rect 14272 25172 14336 25176
rect 14272 25116 14276 25172
rect 14276 25116 14332 25172
rect 14332 25116 14336 25172
rect 14272 25112 14336 25116
rect 14352 25172 14416 25176
rect 14352 25116 14356 25172
rect 14356 25116 14412 25172
rect 14412 25116 14416 25172
rect 14352 25112 14416 25116
rect 24112 25172 24176 25176
rect 24112 25116 24116 25172
rect 24116 25116 24172 25172
rect 24172 25116 24176 25172
rect 24112 25112 24176 25116
rect 24192 25172 24256 25176
rect 24192 25116 24196 25172
rect 24196 25116 24252 25172
rect 24252 25116 24256 25172
rect 24192 25112 24256 25116
rect 24272 25172 24336 25176
rect 24272 25116 24276 25172
rect 24276 25116 24332 25172
rect 24332 25116 24336 25172
rect 24272 25112 24336 25116
rect 24352 25172 24416 25176
rect 24352 25116 24356 25172
rect 24356 25116 24412 25172
rect 24412 25116 24416 25172
rect 24352 25112 24416 25116
rect 19112 24628 19176 24632
rect 19112 24572 19116 24628
rect 19116 24572 19172 24628
rect 19172 24572 19176 24628
rect 19112 24568 19176 24572
rect 19192 24628 19256 24632
rect 19192 24572 19196 24628
rect 19196 24572 19252 24628
rect 19252 24572 19256 24628
rect 19192 24568 19256 24572
rect 19272 24628 19336 24632
rect 19272 24572 19276 24628
rect 19276 24572 19332 24628
rect 19332 24572 19336 24628
rect 19272 24568 19336 24572
rect 19352 24628 19416 24632
rect 19352 24572 19356 24628
rect 19356 24572 19412 24628
rect 19412 24572 19416 24628
rect 19352 24568 19416 24572
rect 29112 24628 29176 24632
rect 29112 24572 29116 24628
rect 29116 24572 29172 24628
rect 29172 24572 29176 24628
rect 29112 24568 29176 24572
rect 29192 24628 29256 24632
rect 29192 24572 29196 24628
rect 29196 24572 29252 24628
rect 29252 24572 29256 24628
rect 29192 24568 29256 24572
rect 29272 24628 29336 24632
rect 29272 24572 29276 24628
rect 29276 24572 29332 24628
rect 29332 24572 29336 24628
rect 29272 24568 29336 24572
rect 29352 24628 29416 24632
rect 29352 24572 29356 24628
rect 29356 24572 29412 24628
rect 29412 24572 29416 24628
rect 29352 24568 29416 24572
rect 14112 24084 14176 24088
rect 14112 24028 14116 24084
rect 14116 24028 14172 24084
rect 14172 24028 14176 24084
rect 14112 24024 14176 24028
rect 14192 24084 14256 24088
rect 14192 24028 14196 24084
rect 14196 24028 14252 24084
rect 14252 24028 14256 24084
rect 14192 24024 14256 24028
rect 14272 24084 14336 24088
rect 14272 24028 14276 24084
rect 14276 24028 14332 24084
rect 14332 24028 14336 24084
rect 14272 24024 14336 24028
rect 14352 24084 14416 24088
rect 14352 24028 14356 24084
rect 14356 24028 14412 24084
rect 14412 24028 14416 24084
rect 14352 24024 14416 24028
rect 24112 24084 24176 24088
rect 24112 24028 24116 24084
rect 24116 24028 24172 24084
rect 24172 24028 24176 24084
rect 24112 24024 24176 24028
rect 24192 24084 24256 24088
rect 24192 24028 24196 24084
rect 24196 24028 24252 24084
rect 24252 24028 24256 24084
rect 24192 24024 24256 24028
rect 24272 24084 24336 24088
rect 24272 24028 24276 24084
rect 24276 24028 24332 24084
rect 24332 24028 24336 24084
rect 24272 24024 24336 24028
rect 24352 24084 24416 24088
rect 24352 24028 24356 24084
rect 24356 24028 24412 24084
rect 24412 24028 24416 24084
rect 24352 24024 24416 24028
rect 19112 23540 19176 23544
rect 19112 23484 19116 23540
rect 19116 23484 19172 23540
rect 19172 23484 19176 23540
rect 19112 23480 19176 23484
rect 19192 23540 19256 23544
rect 19192 23484 19196 23540
rect 19196 23484 19252 23540
rect 19252 23484 19256 23540
rect 19192 23480 19256 23484
rect 19272 23540 19336 23544
rect 19272 23484 19276 23540
rect 19276 23484 19332 23540
rect 19332 23484 19336 23540
rect 19272 23480 19336 23484
rect 19352 23540 19416 23544
rect 19352 23484 19356 23540
rect 19356 23484 19412 23540
rect 19412 23484 19416 23540
rect 19352 23480 19416 23484
rect 29112 23540 29176 23544
rect 29112 23484 29116 23540
rect 29116 23484 29172 23540
rect 29172 23484 29176 23540
rect 29112 23480 29176 23484
rect 29192 23540 29256 23544
rect 29192 23484 29196 23540
rect 29196 23484 29252 23540
rect 29252 23484 29256 23540
rect 29192 23480 29256 23484
rect 29272 23540 29336 23544
rect 29272 23484 29276 23540
rect 29276 23484 29332 23540
rect 29332 23484 29336 23540
rect 29272 23480 29336 23484
rect 29352 23540 29416 23544
rect 29352 23484 29356 23540
rect 29356 23484 29412 23540
rect 29412 23484 29416 23540
rect 29352 23480 29416 23484
rect 14112 22996 14176 23000
rect 14112 22940 14116 22996
rect 14116 22940 14172 22996
rect 14172 22940 14176 22996
rect 14112 22936 14176 22940
rect 14192 22996 14256 23000
rect 14192 22940 14196 22996
rect 14196 22940 14252 22996
rect 14252 22940 14256 22996
rect 14192 22936 14256 22940
rect 14272 22996 14336 23000
rect 14272 22940 14276 22996
rect 14276 22940 14332 22996
rect 14332 22940 14336 22996
rect 14272 22936 14336 22940
rect 14352 22996 14416 23000
rect 14352 22940 14356 22996
rect 14356 22940 14412 22996
rect 14412 22940 14416 22996
rect 14352 22936 14416 22940
rect 24112 22996 24176 23000
rect 24112 22940 24116 22996
rect 24116 22940 24172 22996
rect 24172 22940 24176 22996
rect 24112 22936 24176 22940
rect 24192 22996 24256 23000
rect 24192 22940 24196 22996
rect 24196 22940 24252 22996
rect 24252 22940 24256 22996
rect 24192 22936 24256 22940
rect 24272 22996 24336 23000
rect 24272 22940 24276 22996
rect 24276 22940 24332 22996
rect 24332 22940 24336 22996
rect 24272 22936 24336 22940
rect 24352 22996 24416 23000
rect 24352 22940 24356 22996
rect 24356 22940 24412 22996
rect 24412 22940 24416 22996
rect 24352 22936 24416 22940
rect 19112 22452 19176 22456
rect 19112 22396 19116 22452
rect 19116 22396 19172 22452
rect 19172 22396 19176 22452
rect 19112 22392 19176 22396
rect 19192 22452 19256 22456
rect 19192 22396 19196 22452
rect 19196 22396 19252 22452
rect 19252 22396 19256 22452
rect 19192 22392 19256 22396
rect 19272 22452 19336 22456
rect 19272 22396 19276 22452
rect 19276 22396 19332 22452
rect 19332 22396 19336 22452
rect 19272 22392 19336 22396
rect 19352 22452 19416 22456
rect 19352 22396 19356 22452
rect 19356 22396 19412 22452
rect 19412 22396 19416 22452
rect 19352 22392 19416 22396
rect 29112 22452 29176 22456
rect 29112 22396 29116 22452
rect 29116 22396 29172 22452
rect 29172 22396 29176 22452
rect 29112 22392 29176 22396
rect 29192 22452 29256 22456
rect 29192 22396 29196 22452
rect 29196 22396 29252 22452
rect 29252 22396 29256 22452
rect 29192 22392 29256 22396
rect 29272 22452 29336 22456
rect 29272 22396 29276 22452
rect 29276 22396 29332 22452
rect 29332 22396 29336 22452
rect 29272 22392 29336 22396
rect 29352 22452 29416 22456
rect 29352 22396 29356 22452
rect 29356 22396 29412 22452
rect 29412 22396 29416 22452
rect 29352 22392 29416 22396
rect 14112 21908 14176 21912
rect 14112 21852 14116 21908
rect 14116 21852 14172 21908
rect 14172 21852 14176 21908
rect 14112 21848 14176 21852
rect 14192 21908 14256 21912
rect 14192 21852 14196 21908
rect 14196 21852 14252 21908
rect 14252 21852 14256 21908
rect 14192 21848 14256 21852
rect 14272 21908 14336 21912
rect 14272 21852 14276 21908
rect 14276 21852 14332 21908
rect 14332 21852 14336 21908
rect 14272 21848 14336 21852
rect 14352 21908 14416 21912
rect 14352 21852 14356 21908
rect 14356 21852 14412 21908
rect 14412 21852 14416 21908
rect 14352 21848 14416 21852
rect 24112 21908 24176 21912
rect 24112 21852 24116 21908
rect 24116 21852 24172 21908
rect 24172 21852 24176 21908
rect 24112 21848 24176 21852
rect 24192 21908 24256 21912
rect 24192 21852 24196 21908
rect 24196 21852 24252 21908
rect 24252 21852 24256 21908
rect 24192 21848 24256 21852
rect 24272 21908 24336 21912
rect 24272 21852 24276 21908
rect 24276 21852 24332 21908
rect 24332 21852 24336 21908
rect 24272 21848 24336 21852
rect 24352 21908 24416 21912
rect 24352 21852 24356 21908
rect 24356 21852 24412 21908
rect 24412 21852 24416 21908
rect 24352 21848 24416 21852
rect 19112 21364 19176 21368
rect 19112 21308 19116 21364
rect 19116 21308 19172 21364
rect 19172 21308 19176 21364
rect 19112 21304 19176 21308
rect 19192 21364 19256 21368
rect 19192 21308 19196 21364
rect 19196 21308 19252 21364
rect 19252 21308 19256 21364
rect 19192 21304 19256 21308
rect 19272 21364 19336 21368
rect 19272 21308 19276 21364
rect 19276 21308 19332 21364
rect 19332 21308 19336 21364
rect 19272 21304 19336 21308
rect 19352 21364 19416 21368
rect 19352 21308 19356 21364
rect 19356 21308 19412 21364
rect 19412 21308 19416 21364
rect 19352 21304 19416 21308
rect 29112 21364 29176 21368
rect 29112 21308 29116 21364
rect 29116 21308 29172 21364
rect 29172 21308 29176 21364
rect 29112 21304 29176 21308
rect 29192 21364 29256 21368
rect 29192 21308 29196 21364
rect 29196 21308 29252 21364
rect 29252 21308 29256 21364
rect 29192 21304 29256 21308
rect 29272 21364 29336 21368
rect 29272 21308 29276 21364
rect 29276 21308 29332 21364
rect 29332 21308 29336 21364
rect 29272 21304 29336 21308
rect 29352 21364 29416 21368
rect 29352 21308 29356 21364
rect 29356 21308 29412 21364
rect 29412 21308 29416 21364
rect 29352 21304 29416 21308
rect 14112 20820 14176 20824
rect 14112 20764 14116 20820
rect 14116 20764 14172 20820
rect 14172 20764 14176 20820
rect 14112 20760 14176 20764
rect 14192 20820 14256 20824
rect 14192 20764 14196 20820
rect 14196 20764 14252 20820
rect 14252 20764 14256 20820
rect 14192 20760 14256 20764
rect 14272 20820 14336 20824
rect 14272 20764 14276 20820
rect 14276 20764 14332 20820
rect 14332 20764 14336 20820
rect 14272 20760 14336 20764
rect 14352 20820 14416 20824
rect 14352 20764 14356 20820
rect 14356 20764 14412 20820
rect 14412 20764 14416 20820
rect 14352 20760 14416 20764
rect 24112 20820 24176 20824
rect 24112 20764 24116 20820
rect 24116 20764 24172 20820
rect 24172 20764 24176 20820
rect 24112 20760 24176 20764
rect 24192 20820 24256 20824
rect 24192 20764 24196 20820
rect 24196 20764 24252 20820
rect 24252 20764 24256 20820
rect 24192 20760 24256 20764
rect 24272 20820 24336 20824
rect 24272 20764 24276 20820
rect 24276 20764 24332 20820
rect 24332 20764 24336 20820
rect 24272 20760 24336 20764
rect 24352 20820 24416 20824
rect 24352 20764 24356 20820
rect 24356 20764 24412 20820
rect 24412 20764 24416 20820
rect 24352 20760 24416 20764
rect 19112 20276 19176 20280
rect 19112 20220 19116 20276
rect 19116 20220 19172 20276
rect 19172 20220 19176 20276
rect 19112 20216 19176 20220
rect 19192 20276 19256 20280
rect 19192 20220 19196 20276
rect 19196 20220 19252 20276
rect 19252 20220 19256 20276
rect 19192 20216 19256 20220
rect 19272 20276 19336 20280
rect 19272 20220 19276 20276
rect 19276 20220 19332 20276
rect 19332 20220 19336 20276
rect 19272 20216 19336 20220
rect 19352 20276 19416 20280
rect 19352 20220 19356 20276
rect 19356 20220 19412 20276
rect 19412 20220 19416 20276
rect 19352 20216 19416 20220
rect 29112 20276 29176 20280
rect 29112 20220 29116 20276
rect 29116 20220 29172 20276
rect 29172 20220 29176 20276
rect 29112 20216 29176 20220
rect 29192 20276 29256 20280
rect 29192 20220 29196 20276
rect 29196 20220 29252 20276
rect 29252 20220 29256 20276
rect 29192 20216 29256 20220
rect 29272 20276 29336 20280
rect 29272 20220 29276 20276
rect 29276 20220 29332 20276
rect 29332 20220 29336 20276
rect 29272 20216 29336 20220
rect 29352 20276 29416 20280
rect 29352 20220 29356 20276
rect 29356 20220 29412 20276
rect 29412 20220 29416 20276
rect 29352 20216 29416 20220
rect 14112 19732 14176 19736
rect 14112 19676 14116 19732
rect 14116 19676 14172 19732
rect 14172 19676 14176 19732
rect 14112 19672 14176 19676
rect 14192 19732 14256 19736
rect 14192 19676 14196 19732
rect 14196 19676 14252 19732
rect 14252 19676 14256 19732
rect 14192 19672 14256 19676
rect 14272 19732 14336 19736
rect 14272 19676 14276 19732
rect 14276 19676 14332 19732
rect 14332 19676 14336 19732
rect 14272 19672 14336 19676
rect 14352 19732 14416 19736
rect 14352 19676 14356 19732
rect 14356 19676 14412 19732
rect 14412 19676 14416 19732
rect 14352 19672 14416 19676
rect 24112 19732 24176 19736
rect 24112 19676 24116 19732
rect 24116 19676 24172 19732
rect 24172 19676 24176 19732
rect 24112 19672 24176 19676
rect 24192 19732 24256 19736
rect 24192 19676 24196 19732
rect 24196 19676 24252 19732
rect 24252 19676 24256 19732
rect 24192 19672 24256 19676
rect 24272 19732 24336 19736
rect 24272 19676 24276 19732
rect 24276 19676 24332 19732
rect 24332 19676 24336 19732
rect 24272 19672 24336 19676
rect 24352 19732 24416 19736
rect 24352 19676 24356 19732
rect 24356 19676 24412 19732
rect 24412 19676 24416 19732
rect 24352 19672 24416 19676
rect 19112 19188 19176 19192
rect 19112 19132 19116 19188
rect 19116 19132 19172 19188
rect 19172 19132 19176 19188
rect 19112 19128 19176 19132
rect 19192 19188 19256 19192
rect 19192 19132 19196 19188
rect 19196 19132 19252 19188
rect 19252 19132 19256 19188
rect 19192 19128 19256 19132
rect 19272 19188 19336 19192
rect 19272 19132 19276 19188
rect 19276 19132 19332 19188
rect 19332 19132 19336 19188
rect 19272 19128 19336 19132
rect 19352 19188 19416 19192
rect 19352 19132 19356 19188
rect 19356 19132 19412 19188
rect 19412 19132 19416 19188
rect 19352 19128 19416 19132
rect 29112 19188 29176 19192
rect 29112 19132 29116 19188
rect 29116 19132 29172 19188
rect 29172 19132 29176 19188
rect 29112 19128 29176 19132
rect 29192 19188 29256 19192
rect 29192 19132 29196 19188
rect 29196 19132 29252 19188
rect 29252 19132 29256 19188
rect 29192 19128 29256 19132
rect 29272 19188 29336 19192
rect 29272 19132 29276 19188
rect 29276 19132 29332 19188
rect 29332 19132 29336 19188
rect 29272 19128 29336 19132
rect 29352 19188 29416 19192
rect 29352 19132 29356 19188
rect 29356 19132 29412 19188
rect 29412 19132 29416 19188
rect 29352 19128 29416 19132
rect 14112 18644 14176 18648
rect 14112 18588 14116 18644
rect 14116 18588 14172 18644
rect 14172 18588 14176 18644
rect 14112 18584 14176 18588
rect 14192 18644 14256 18648
rect 14192 18588 14196 18644
rect 14196 18588 14252 18644
rect 14252 18588 14256 18644
rect 14192 18584 14256 18588
rect 14272 18644 14336 18648
rect 14272 18588 14276 18644
rect 14276 18588 14332 18644
rect 14332 18588 14336 18644
rect 14272 18584 14336 18588
rect 14352 18644 14416 18648
rect 14352 18588 14356 18644
rect 14356 18588 14412 18644
rect 14412 18588 14416 18644
rect 14352 18584 14416 18588
rect 24112 18644 24176 18648
rect 24112 18588 24116 18644
rect 24116 18588 24172 18644
rect 24172 18588 24176 18644
rect 24112 18584 24176 18588
rect 24192 18644 24256 18648
rect 24192 18588 24196 18644
rect 24196 18588 24252 18644
rect 24252 18588 24256 18644
rect 24192 18584 24256 18588
rect 24272 18644 24336 18648
rect 24272 18588 24276 18644
rect 24276 18588 24332 18644
rect 24332 18588 24336 18644
rect 24272 18584 24336 18588
rect 24352 18644 24416 18648
rect 24352 18588 24356 18644
rect 24356 18588 24412 18644
rect 24412 18588 24416 18644
rect 24352 18584 24416 18588
rect 19112 18100 19176 18104
rect 19112 18044 19116 18100
rect 19116 18044 19172 18100
rect 19172 18044 19176 18100
rect 19112 18040 19176 18044
rect 19192 18100 19256 18104
rect 19192 18044 19196 18100
rect 19196 18044 19252 18100
rect 19252 18044 19256 18100
rect 19192 18040 19256 18044
rect 19272 18100 19336 18104
rect 19272 18044 19276 18100
rect 19276 18044 19332 18100
rect 19332 18044 19336 18100
rect 19272 18040 19336 18044
rect 19352 18100 19416 18104
rect 19352 18044 19356 18100
rect 19356 18044 19412 18100
rect 19412 18044 19416 18100
rect 19352 18040 19416 18044
rect 29112 18100 29176 18104
rect 29112 18044 29116 18100
rect 29116 18044 29172 18100
rect 29172 18044 29176 18100
rect 29112 18040 29176 18044
rect 29192 18100 29256 18104
rect 29192 18044 29196 18100
rect 29196 18044 29252 18100
rect 29252 18044 29256 18100
rect 29192 18040 29256 18044
rect 29272 18100 29336 18104
rect 29272 18044 29276 18100
rect 29276 18044 29332 18100
rect 29332 18044 29336 18100
rect 29272 18040 29336 18044
rect 29352 18100 29416 18104
rect 29352 18044 29356 18100
rect 29356 18044 29412 18100
rect 29412 18044 29416 18100
rect 29352 18040 29416 18044
rect 14112 17556 14176 17560
rect 14112 17500 14116 17556
rect 14116 17500 14172 17556
rect 14172 17500 14176 17556
rect 14112 17496 14176 17500
rect 14192 17556 14256 17560
rect 14192 17500 14196 17556
rect 14196 17500 14252 17556
rect 14252 17500 14256 17556
rect 14192 17496 14256 17500
rect 14272 17556 14336 17560
rect 14272 17500 14276 17556
rect 14276 17500 14332 17556
rect 14332 17500 14336 17556
rect 14272 17496 14336 17500
rect 14352 17556 14416 17560
rect 14352 17500 14356 17556
rect 14356 17500 14412 17556
rect 14412 17500 14416 17556
rect 14352 17496 14416 17500
rect 24112 17556 24176 17560
rect 24112 17500 24116 17556
rect 24116 17500 24172 17556
rect 24172 17500 24176 17556
rect 24112 17496 24176 17500
rect 24192 17556 24256 17560
rect 24192 17500 24196 17556
rect 24196 17500 24252 17556
rect 24252 17500 24256 17556
rect 24192 17496 24256 17500
rect 24272 17556 24336 17560
rect 24272 17500 24276 17556
rect 24276 17500 24332 17556
rect 24332 17500 24336 17556
rect 24272 17496 24336 17500
rect 24352 17556 24416 17560
rect 24352 17500 24356 17556
rect 24356 17500 24412 17556
rect 24412 17500 24416 17556
rect 24352 17496 24416 17500
rect 19112 17012 19176 17016
rect 19112 16956 19116 17012
rect 19116 16956 19172 17012
rect 19172 16956 19176 17012
rect 19112 16952 19176 16956
rect 19192 17012 19256 17016
rect 19192 16956 19196 17012
rect 19196 16956 19252 17012
rect 19252 16956 19256 17012
rect 19192 16952 19256 16956
rect 19272 17012 19336 17016
rect 19272 16956 19276 17012
rect 19276 16956 19332 17012
rect 19332 16956 19336 17012
rect 19272 16952 19336 16956
rect 19352 17012 19416 17016
rect 19352 16956 19356 17012
rect 19356 16956 19412 17012
rect 19412 16956 19416 17012
rect 19352 16952 19416 16956
rect 29112 17012 29176 17016
rect 29112 16956 29116 17012
rect 29116 16956 29172 17012
rect 29172 16956 29176 17012
rect 29112 16952 29176 16956
rect 29192 17012 29256 17016
rect 29192 16956 29196 17012
rect 29196 16956 29252 17012
rect 29252 16956 29256 17012
rect 29192 16952 29256 16956
rect 29272 17012 29336 17016
rect 29272 16956 29276 17012
rect 29276 16956 29332 17012
rect 29332 16956 29336 17012
rect 29272 16952 29336 16956
rect 29352 17012 29416 17016
rect 29352 16956 29356 17012
rect 29356 16956 29412 17012
rect 29412 16956 29416 17012
rect 29352 16952 29416 16956
rect 14112 16468 14176 16472
rect 14112 16412 14116 16468
rect 14116 16412 14172 16468
rect 14172 16412 14176 16468
rect 14112 16408 14176 16412
rect 14192 16468 14256 16472
rect 14192 16412 14196 16468
rect 14196 16412 14252 16468
rect 14252 16412 14256 16468
rect 14192 16408 14256 16412
rect 14272 16468 14336 16472
rect 14272 16412 14276 16468
rect 14276 16412 14332 16468
rect 14332 16412 14336 16468
rect 14272 16408 14336 16412
rect 14352 16468 14416 16472
rect 14352 16412 14356 16468
rect 14356 16412 14412 16468
rect 14412 16412 14416 16468
rect 14352 16408 14416 16412
rect 24112 16468 24176 16472
rect 24112 16412 24116 16468
rect 24116 16412 24172 16468
rect 24172 16412 24176 16468
rect 24112 16408 24176 16412
rect 24192 16468 24256 16472
rect 24192 16412 24196 16468
rect 24196 16412 24252 16468
rect 24252 16412 24256 16468
rect 24192 16408 24256 16412
rect 24272 16468 24336 16472
rect 24272 16412 24276 16468
rect 24276 16412 24332 16468
rect 24332 16412 24336 16468
rect 24272 16408 24336 16412
rect 24352 16468 24416 16472
rect 24352 16412 24356 16468
rect 24356 16412 24412 16468
rect 24412 16412 24416 16468
rect 24352 16408 24416 16412
rect 19112 15924 19176 15928
rect 19112 15868 19116 15924
rect 19116 15868 19172 15924
rect 19172 15868 19176 15924
rect 19112 15864 19176 15868
rect 19192 15924 19256 15928
rect 19192 15868 19196 15924
rect 19196 15868 19252 15924
rect 19252 15868 19256 15924
rect 19192 15864 19256 15868
rect 19272 15924 19336 15928
rect 19272 15868 19276 15924
rect 19276 15868 19332 15924
rect 19332 15868 19336 15924
rect 19272 15864 19336 15868
rect 19352 15924 19416 15928
rect 19352 15868 19356 15924
rect 19356 15868 19412 15924
rect 19412 15868 19416 15924
rect 19352 15864 19416 15868
rect 29112 15924 29176 15928
rect 29112 15868 29116 15924
rect 29116 15868 29172 15924
rect 29172 15868 29176 15924
rect 29112 15864 29176 15868
rect 29192 15924 29256 15928
rect 29192 15868 29196 15924
rect 29196 15868 29252 15924
rect 29252 15868 29256 15924
rect 29192 15864 29256 15868
rect 29272 15924 29336 15928
rect 29272 15868 29276 15924
rect 29276 15868 29332 15924
rect 29332 15868 29336 15924
rect 29272 15864 29336 15868
rect 29352 15924 29416 15928
rect 29352 15868 29356 15924
rect 29356 15868 29412 15924
rect 29412 15868 29416 15924
rect 29352 15864 29416 15868
rect 14112 15380 14176 15384
rect 14112 15324 14116 15380
rect 14116 15324 14172 15380
rect 14172 15324 14176 15380
rect 14112 15320 14176 15324
rect 14192 15380 14256 15384
rect 14192 15324 14196 15380
rect 14196 15324 14252 15380
rect 14252 15324 14256 15380
rect 14192 15320 14256 15324
rect 14272 15380 14336 15384
rect 14272 15324 14276 15380
rect 14276 15324 14332 15380
rect 14332 15324 14336 15380
rect 14272 15320 14336 15324
rect 14352 15380 14416 15384
rect 14352 15324 14356 15380
rect 14356 15324 14412 15380
rect 14412 15324 14416 15380
rect 14352 15320 14416 15324
rect 24112 15380 24176 15384
rect 24112 15324 24116 15380
rect 24116 15324 24172 15380
rect 24172 15324 24176 15380
rect 24112 15320 24176 15324
rect 24192 15380 24256 15384
rect 24192 15324 24196 15380
rect 24196 15324 24252 15380
rect 24252 15324 24256 15380
rect 24192 15320 24256 15324
rect 24272 15380 24336 15384
rect 24272 15324 24276 15380
rect 24276 15324 24332 15380
rect 24332 15324 24336 15380
rect 24272 15320 24336 15324
rect 24352 15380 24416 15384
rect 24352 15324 24356 15380
rect 24356 15324 24412 15380
rect 24412 15324 24416 15380
rect 24352 15320 24416 15324
rect 19112 14836 19176 14840
rect 19112 14780 19116 14836
rect 19116 14780 19172 14836
rect 19172 14780 19176 14836
rect 19112 14776 19176 14780
rect 19192 14836 19256 14840
rect 19192 14780 19196 14836
rect 19196 14780 19252 14836
rect 19252 14780 19256 14836
rect 19192 14776 19256 14780
rect 19272 14836 19336 14840
rect 19272 14780 19276 14836
rect 19276 14780 19332 14836
rect 19332 14780 19336 14836
rect 19272 14776 19336 14780
rect 19352 14836 19416 14840
rect 19352 14780 19356 14836
rect 19356 14780 19412 14836
rect 19412 14780 19416 14836
rect 19352 14776 19416 14780
rect 29112 14836 29176 14840
rect 29112 14780 29116 14836
rect 29116 14780 29172 14836
rect 29172 14780 29176 14836
rect 29112 14776 29176 14780
rect 29192 14836 29256 14840
rect 29192 14780 29196 14836
rect 29196 14780 29252 14836
rect 29252 14780 29256 14836
rect 29192 14776 29256 14780
rect 29272 14836 29336 14840
rect 29272 14780 29276 14836
rect 29276 14780 29332 14836
rect 29332 14780 29336 14836
rect 29272 14776 29336 14780
rect 29352 14836 29416 14840
rect 29352 14780 29356 14836
rect 29356 14780 29412 14836
rect 29412 14780 29416 14836
rect 29352 14776 29416 14780
rect 14112 14292 14176 14296
rect 14112 14236 14116 14292
rect 14116 14236 14172 14292
rect 14172 14236 14176 14292
rect 14112 14232 14176 14236
rect 14192 14292 14256 14296
rect 14192 14236 14196 14292
rect 14196 14236 14252 14292
rect 14252 14236 14256 14292
rect 14192 14232 14256 14236
rect 14272 14292 14336 14296
rect 14272 14236 14276 14292
rect 14276 14236 14332 14292
rect 14332 14236 14336 14292
rect 14272 14232 14336 14236
rect 14352 14292 14416 14296
rect 14352 14236 14356 14292
rect 14356 14236 14412 14292
rect 14412 14236 14416 14292
rect 14352 14232 14416 14236
rect 24112 14292 24176 14296
rect 24112 14236 24116 14292
rect 24116 14236 24172 14292
rect 24172 14236 24176 14292
rect 24112 14232 24176 14236
rect 24192 14292 24256 14296
rect 24192 14236 24196 14292
rect 24196 14236 24252 14292
rect 24252 14236 24256 14292
rect 24192 14232 24256 14236
rect 24272 14292 24336 14296
rect 24272 14236 24276 14292
rect 24276 14236 24332 14292
rect 24332 14236 24336 14292
rect 24272 14232 24336 14236
rect 24352 14292 24416 14296
rect 24352 14236 24356 14292
rect 24356 14236 24412 14292
rect 24412 14236 24416 14292
rect 24352 14232 24416 14236
rect 19112 13748 19176 13752
rect 19112 13692 19116 13748
rect 19116 13692 19172 13748
rect 19172 13692 19176 13748
rect 19112 13688 19176 13692
rect 19192 13748 19256 13752
rect 19192 13692 19196 13748
rect 19196 13692 19252 13748
rect 19252 13692 19256 13748
rect 19192 13688 19256 13692
rect 19272 13748 19336 13752
rect 19272 13692 19276 13748
rect 19276 13692 19332 13748
rect 19332 13692 19336 13748
rect 19272 13688 19336 13692
rect 19352 13748 19416 13752
rect 19352 13692 19356 13748
rect 19356 13692 19412 13748
rect 19412 13692 19416 13748
rect 19352 13688 19416 13692
rect 29112 13748 29176 13752
rect 29112 13692 29116 13748
rect 29116 13692 29172 13748
rect 29172 13692 29176 13748
rect 29112 13688 29176 13692
rect 29192 13748 29256 13752
rect 29192 13692 29196 13748
rect 29196 13692 29252 13748
rect 29252 13692 29256 13748
rect 29192 13688 29256 13692
rect 29272 13748 29336 13752
rect 29272 13692 29276 13748
rect 29276 13692 29332 13748
rect 29332 13692 29336 13748
rect 29272 13688 29336 13692
rect 29352 13748 29416 13752
rect 29352 13692 29356 13748
rect 29356 13692 29412 13748
rect 29412 13692 29416 13748
rect 29352 13688 29416 13692
rect 14112 13204 14176 13208
rect 14112 13148 14116 13204
rect 14116 13148 14172 13204
rect 14172 13148 14176 13204
rect 14112 13144 14176 13148
rect 14192 13204 14256 13208
rect 14192 13148 14196 13204
rect 14196 13148 14252 13204
rect 14252 13148 14256 13204
rect 14192 13144 14256 13148
rect 14272 13204 14336 13208
rect 14272 13148 14276 13204
rect 14276 13148 14332 13204
rect 14332 13148 14336 13204
rect 14272 13144 14336 13148
rect 14352 13204 14416 13208
rect 14352 13148 14356 13204
rect 14356 13148 14412 13204
rect 14412 13148 14416 13204
rect 14352 13144 14416 13148
rect 24112 13204 24176 13208
rect 24112 13148 24116 13204
rect 24116 13148 24172 13204
rect 24172 13148 24176 13204
rect 24112 13144 24176 13148
rect 24192 13204 24256 13208
rect 24192 13148 24196 13204
rect 24196 13148 24252 13204
rect 24252 13148 24256 13204
rect 24192 13144 24256 13148
rect 24272 13204 24336 13208
rect 24272 13148 24276 13204
rect 24276 13148 24332 13204
rect 24332 13148 24336 13204
rect 24272 13144 24336 13148
rect 24352 13204 24416 13208
rect 24352 13148 24356 13204
rect 24356 13148 24412 13204
rect 24412 13148 24416 13204
rect 24352 13144 24416 13148
rect 19112 12660 19176 12664
rect 19112 12604 19116 12660
rect 19116 12604 19172 12660
rect 19172 12604 19176 12660
rect 19112 12600 19176 12604
rect 19192 12660 19256 12664
rect 19192 12604 19196 12660
rect 19196 12604 19252 12660
rect 19252 12604 19256 12660
rect 19192 12600 19256 12604
rect 19272 12660 19336 12664
rect 19272 12604 19276 12660
rect 19276 12604 19332 12660
rect 19332 12604 19336 12660
rect 19272 12600 19336 12604
rect 19352 12660 19416 12664
rect 19352 12604 19356 12660
rect 19356 12604 19412 12660
rect 19412 12604 19416 12660
rect 19352 12600 19416 12604
rect 29112 12660 29176 12664
rect 29112 12604 29116 12660
rect 29116 12604 29172 12660
rect 29172 12604 29176 12660
rect 29112 12600 29176 12604
rect 29192 12660 29256 12664
rect 29192 12604 29196 12660
rect 29196 12604 29252 12660
rect 29252 12604 29256 12660
rect 29192 12600 29256 12604
rect 29272 12660 29336 12664
rect 29272 12604 29276 12660
rect 29276 12604 29332 12660
rect 29332 12604 29336 12660
rect 29272 12600 29336 12604
rect 29352 12660 29416 12664
rect 29352 12604 29356 12660
rect 29356 12604 29412 12660
rect 29412 12604 29416 12660
rect 29352 12600 29416 12604
rect 14112 12116 14176 12120
rect 14112 12060 14116 12116
rect 14116 12060 14172 12116
rect 14172 12060 14176 12116
rect 14112 12056 14176 12060
rect 14192 12116 14256 12120
rect 14192 12060 14196 12116
rect 14196 12060 14252 12116
rect 14252 12060 14256 12116
rect 14192 12056 14256 12060
rect 14272 12116 14336 12120
rect 14272 12060 14276 12116
rect 14276 12060 14332 12116
rect 14332 12060 14336 12116
rect 14272 12056 14336 12060
rect 14352 12116 14416 12120
rect 14352 12060 14356 12116
rect 14356 12060 14412 12116
rect 14412 12060 14416 12116
rect 14352 12056 14416 12060
rect 24112 12116 24176 12120
rect 24112 12060 24116 12116
rect 24116 12060 24172 12116
rect 24172 12060 24176 12116
rect 24112 12056 24176 12060
rect 24192 12116 24256 12120
rect 24192 12060 24196 12116
rect 24196 12060 24252 12116
rect 24252 12060 24256 12116
rect 24192 12056 24256 12060
rect 24272 12116 24336 12120
rect 24272 12060 24276 12116
rect 24276 12060 24332 12116
rect 24332 12060 24336 12116
rect 24272 12056 24336 12060
rect 24352 12116 24416 12120
rect 24352 12060 24356 12116
rect 24356 12060 24412 12116
rect 24412 12060 24416 12116
rect 24352 12056 24416 12060
rect 19112 11572 19176 11576
rect 19112 11516 19116 11572
rect 19116 11516 19172 11572
rect 19172 11516 19176 11572
rect 19112 11512 19176 11516
rect 19192 11572 19256 11576
rect 19192 11516 19196 11572
rect 19196 11516 19252 11572
rect 19252 11516 19256 11572
rect 19192 11512 19256 11516
rect 19272 11572 19336 11576
rect 19272 11516 19276 11572
rect 19276 11516 19332 11572
rect 19332 11516 19336 11572
rect 19272 11512 19336 11516
rect 19352 11572 19416 11576
rect 19352 11516 19356 11572
rect 19356 11516 19412 11572
rect 19412 11516 19416 11572
rect 19352 11512 19416 11516
rect 29112 11572 29176 11576
rect 29112 11516 29116 11572
rect 29116 11516 29172 11572
rect 29172 11516 29176 11572
rect 29112 11512 29176 11516
rect 29192 11572 29256 11576
rect 29192 11516 29196 11572
rect 29196 11516 29252 11572
rect 29252 11516 29256 11572
rect 29192 11512 29256 11516
rect 29272 11572 29336 11576
rect 29272 11516 29276 11572
rect 29276 11516 29332 11572
rect 29332 11516 29336 11572
rect 29272 11512 29336 11516
rect 29352 11572 29416 11576
rect 29352 11516 29356 11572
rect 29356 11516 29412 11572
rect 29412 11516 29416 11572
rect 29352 11512 29416 11516
rect 14112 11028 14176 11032
rect 14112 10972 14116 11028
rect 14116 10972 14172 11028
rect 14172 10972 14176 11028
rect 14112 10968 14176 10972
rect 14192 11028 14256 11032
rect 14192 10972 14196 11028
rect 14196 10972 14252 11028
rect 14252 10972 14256 11028
rect 14192 10968 14256 10972
rect 14272 11028 14336 11032
rect 14272 10972 14276 11028
rect 14276 10972 14332 11028
rect 14332 10972 14336 11028
rect 14272 10968 14336 10972
rect 14352 11028 14416 11032
rect 14352 10972 14356 11028
rect 14356 10972 14412 11028
rect 14412 10972 14416 11028
rect 14352 10968 14416 10972
rect 24112 11028 24176 11032
rect 24112 10972 24116 11028
rect 24116 10972 24172 11028
rect 24172 10972 24176 11028
rect 24112 10968 24176 10972
rect 24192 11028 24256 11032
rect 24192 10972 24196 11028
rect 24196 10972 24252 11028
rect 24252 10972 24256 11028
rect 24192 10968 24256 10972
rect 24272 11028 24336 11032
rect 24272 10972 24276 11028
rect 24276 10972 24332 11028
rect 24332 10972 24336 11028
rect 24272 10968 24336 10972
rect 24352 11028 24416 11032
rect 24352 10972 24356 11028
rect 24356 10972 24412 11028
rect 24412 10972 24416 11028
rect 24352 10968 24416 10972
rect 5008 8928 5072 8992
rect 5088 8928 5152 8992
rect 5168 8928 5232 8992
rect 5248 8928 5312 8992
rect 5328 8928 5392 8992
rect 5408 8928 5472 8992
rect 5488 8928 5552 8992
rect 5568 8928 5632 8992
rect 5648 8928 5712 8992
rect 5728 8928 5792 8992
rect 5808 8928 5872 8992
rect 5888 8928 5952 8992
rect 5968 8928 6032 8992
rect 6048 8928 6112 8992
rect 6128 8928 6192 8992
rect 6208 8928 6272 8992
rect 6288 8928 6352 8992
rect 6368 8928 6432 8992
rect 6448 8928 6512 8992
rect 6528 8928 6592 8992
rect 6608 8928 6672 8992
rect 6688 8928 6752 8992
rect 6768 8928 6832 8992
rect 6848 8928 6912 8992
rect 6928 8928 6992 8992
rect 7008 8928 7072 8992
rect 7088 8928 7152 8992
rect 7168 8928 7232 8992
rect 7248 8928 7312 8992
rect 7328 8928 7392 8992
rect 7408 8928 7472 8992
rect 7488 8928 7552 8992
rect 7568 8928 7632 8992
rect 7648 8928 7712 8992
rect 7728 8928 7792 8992
rect 7808 8928 7872 8992
rect 7888 8928 7952 8992
rect 7968 8928 8032 8992
rect 8048 8928 8112 8992
rect 8128 8928 8192 8992
rect 8208 8928 8272 8992
rect 8288 8928 8352 8992
rect 8368 8928 8432 8992
rect 8448 8928 8512 8992
rect 8528 8928 8592 8992
rect 8608 8928 8672 8992
rect 8688 8928 8752 8992
rect 8768 8928 8832 8992
rect 8848 8928 8912 8992
rect 8928 8928 8992 8992
rect 14112 8928 14176 8992
rect 14192 8928 14256 8992
rect 14272 8928 14336 8992
rect 14352 8928 14416 8992
rect 24112 8928 24176 8992
rect 24192 8928 24256 8992
rect 24272 8928 24336 8992
rect 24352 8928 24416 8992
rect 36376 8928 36440 8992
rect 36456 8928 36520 8992
rect 36536 8928 36600 8992
rect 36616 8928 36680 8992
rect 36696 8928 36760 8992
rect 36776 8928 36840 8992
rect 36856 8928 36920 8992
rect 36936 8928 37000 8992
rect 37016 8928 37080 8992
rect 37096 8928 37160 8992
rect 37176 8928 37240 8992
rect 37256 8928 37320 8992
rect 37336 8928 37400 8992
rect 37416 8928 37480 8992
rect 37496 8928 37560 8992
rect 37576 8928 37640 8992
rect 37656 8928 37720 8992
rect 37736 8928 37800 8992
rect 37816 8928 37880 8992
rect 37896 8928 37960 8992
rect 37976 8928 38040 8992
rect 38056 8928 38120 8992
rect 38136 8928 38200 8992
rect 38216 8928 38280 8992
rect 38296 8928 38360 8992
rect 38376 8928 38440 8992
rect 38456 8928 38520 8992
rect 38536 8928 38600 8992
rect 38616 8928 38680 8992
rect 38696 8928 38760 8992
rect 38776 8928 38840 8992
rect 38856 8928 38920 8992
rect 38936 8928 39000 8992
rect 39016 8928 39080 8992
rect 39096 8928 39160 8992
rect 39176 8928 39240 8992
rect 39256 8928 39320 8992
rect 39336 8928 39400 8992
rect 39416 8928 39480 8992
rect 39496 8928 39560 8992
rect 39576 8928 39640 8992
rect 39656 8928 39720 8992
rect 39736 8928 39800 8992
rect 39816 8928 39880 8992
rect 39896 8928 39960 8992
rect 39976 8928 40040 8992
rect 40056 8928 40120 8992
rect 40136 8928 40200 8992
rect 40216 8928 40280 8992
rect 40296 8928 40360 8992
rect 5008 8848 5072 8912
rect 5088 8848 5152 8912
rect 5168 8848 5232 8912
rect 5248 8848 5312 8912
rect 5328 8848 5392 8912
rect 5408 8848 5472 8912
rect 5488 8848 5552 8912
rect 5568 8848 5632 8912
rect 5648 8848 5712 8912
rect 5728 8848 5792 8912
rect 5808 8848 5872 8912
rect 5888 8848 5952 8912
rect 5968 8848 6032 8912
rect 6048 8848 6112 8912
rect 6128 8848 6192 8912
rect 6208 8848 6272 8912
rect 6288 8848 6352 8912
rect 6368 8848 6432 8912
rect 6448 8848 6512 8912
rect 6528 8848 6592 8912
rect 6608 8848 6672 8912
rect 6688 8848 6752 8912
rect 6768 8848 6832 8912
rect 6848 8848 6912 8912
rect 6928 8848 6992 8912
rect 7008 8848 7072 8912
rect 7088 8848 7152 8912
rect 7168 8848 7232 8912
rect 7248 8848 7312 8912
rect 7328 8848 7392 8912
rect 7408 8848 7472 8912
rect 7488 8848 7552 8912
rect 7568 8848 7632 8912
rect 7648 8848 7712 8912
rect 7728 8848 7792 8912
rect 7808 8848 7872 8912
rect 7888 8848 7952 8912
rect 7968 8848 8032 8912
rect 8048 8848 8112 8912
rect 8128 8848 8192 8912
rect 8208 8848 8272 8912
rect 8288 8848 8352 8912
rect 8368 8848 8432 8912
rect 8448 8848 8512 8912
rect 8528 8848 8592 8912
rect 8608 8848 8672 8912
rect 8688 8848 8752 8912
rect 8768 8848 8832 8912
rect 8848 8848 8912 8912
rect 8928 8848 8992 8912
rect 14112 8848 14176 8912
rect 14192 8848 14256 8912
rect 14272 8848 14336 8912
rect 14352 8848 14416 8912
rect 24112 8848 24176 8912
rect 24192 8848 24256 8912
rect 24272 8848 24336 8912
rect 24352 8848 24416 8912
rect 36376 8848 36440 8912
rect 36456 8848 36520 8912
rect 36536 8848 36600 8912
rect 36616 8848 36680 8912
rect 36696 8848 36760 8912
rect 36776 8848 36840 8912
rect 36856 8848 36920 8912
rect 36936 8848 37000 8912
rect 37016 8848 37080 8912
rect 37096 8848 37160 8912
rect 37176 8848 37240 8912
rect 37256 8848 37320 8912
rect 37336 8848 37400 8912
rect 37416 8848 37480 8912
rect 37496 8848 37560 8912
rect 37576 8848 37640 8912
rect 37656 8848 37720 8912
rect 37736 8848 37800 8912
rect 37816 8848 37880 8912
rect 37896 8848 37960 8912
rect 37976 8848 38040 8912
rect 38056 8848 38120 8912
rect 38136 8848 38200 8912
rect 38216 8848 38280 8912
rect 38296 8848 38360 8912
rect 38376 8848 38440 8912
rect 38456 8848 38520 8912
rect 38536 8848 38600 8912
rect 38616 8848 38680 8912
rect 38696 8848 38760 8912
rect 38776 8848 38840 8912
rect 38856 8848 38920 8912
rect 38936 8848 39000 8912
rect 39016 8848 39080 8912
rect 39096 8848 39160 8912
rect 39176 8848 39240 8912
rect 39256 8848 39320 8912
rect 39336 8848 39400 8912
rect 39416 8848 39480 8912
rect 39496 8848 39560 8912
rect 39576 8848 39640 8912
rect 39656 8848 39720 8912
rect 39736 8848 39800 8912
rect 39816 8848 39880 8912
rect 39896 8848 39960 8912
rect 39976 8848 40040 8912
rect 40056 8848 40120 8912
rect 40136 8848 40200 8912
rect 40216 8848 40280 8912
rect 40296 8848 40360 8912
rect 5008 8768 5072 8832
rect 5088 8768 5152 8832
rect 5168 8768 5232 8832
rect 5248 8768 5312 8832
rect 5328 8768 5392 8832
rect 5408 8768 5472 8832
rect 5488 8768 5552 8832
rect 5568 8768 5632 8832
rect 5648 8768 5712 8832
rect 5728 8768 5792 8832
rect 5808 8768 5872 8832
rect 5888 8768 5952 8832
rect 5968 8768 6032 8832
rect 6048 8768 6112 8832
rect 6128 8768 6192 8832
rect 6208 8768 6272 8832
rect 6288 8768 6352 8832
rect 6368 8768 6432 8832
rect 6448 8768 6512 8832
rect 6528 8768 6592 8832
rect 6608 8768 6672 8832
rect 6688 8768 6752 8832
rect 6768 8768 6832 8832
rect 6848 8768 6912 8832
rect 6928 8768 6992 8832
rect 7008 8768 7072 8832
rect 7088 8768 7152 8832
rect 7168 8768 7232 8832
rect 7248 8768 7312 8832
rect 7328 8768 7392 8832
rect 7408 8768 7472 8832
rect 7488 8768 7552 8832
rect 7568 8768 7632 8832
rect 7648 8768 7712 8832
rect 7728 8768 7792 8832
rect 7808 8768 7872 8832
rect 7888 8768 7952 8832
rect 7968 8768 8032 8832
rect 8048 8768 8112 8832
rect 8128 8768 8192 8832
rect 8208 8768 8272 8832
rect 8288 8768 8352 8832
rect 8368 8768 8432 8832
rect 8448 8768 8512 8832
rect 8528 8768 8592 8832
rect 8608 8768 8672 8832
rect 8688 8768 8752 8832
rect 8768 8768 8832 8832
rect 8848 8768 8912 8832
rect 8928 8768 8992 8832
rect 14112 8768 14176 8832
rect 14192 8768 14256 8832
rect 14272 8768 14336 8832
rect 14352 8768 14416 8832
rect 24112 8768 24176 8832
rect 24192 8768 24256 8832
rect 24272 8768 24336 8832
rect 24352 8768 24416 8832
rect 36376 8768 36440 8832
rect 36456 8768 36520 8832
rect 36536 8768 36600 8832
rect 36616 8768 36680 8832
rect 36696 8768 36760 8832
rect 36776 8768 36840 8832
rect 36856 8768 36920 8832
rect 36936 8768 37000 8832
rect 37016 8768 37080 8832
rect 37096 8768 37160 8832
rect 37176 8768 37240 8832
rect 37256 8768 37320 8832
rect 37336 8768 37400 8832
rect 37416 8768 37480 8832
rect 37496 8768 37560 8832
rect 37576 8768 37640 8832
rect 37656 8768 37720 8832
rect 37736 8768 37800 8832
rect 37816 8768 37880 8832
rect 37896 8768 37960 8832
rect 37976 8768 38040 8832
rect 38056 8768 38120 8832
rect 38136 8768 38200 8832
rect 38216 8768 38280 8832
rect 38296 8768 38360 8832
rect 38376 8768 38440 8832
rect 38456 8768 38520 8832
rect 38536 8768 38600 8832
rect 38616 8768 38680 8832
rect 38696 8768 38760 8832
rect 38776 8768 38840 8832
rect 38856 8768 38920 8832
rect 38936 8768 39000 8832
rect 39016 8768 39080 8832
rect 39096 8768 39160 8832
rect 39176 8768 39240 8832
rect 39256 8768 39320 8832
rect 39336 8768 39400 8832
rect 39416 8768 39480 8832
rect 39496 8768 39560 8832
rect 39576 8768 39640 8832
rect 39656 8768 39720 8832
rect 39736 8768 39800 8832
rect 39816 8768 39880 8832
rect 39896 8768 39960 8832
rect 39976 8768 40040 8832
rect 40056 8768 40120 8832
rect 40136 8768 40200 8832
rect 40216 8768 40280 8832
rect 40296 8768 40360 8832
rect 5008 8688 5072 8752
rect 5088 8688 5152 8752
rect 5168 8688 5232 8752
rect 5248 8688 5312 8752
rect 5328 8688 5392 8752
rect 5408 8688 5472 8752
rect 5488 8688 5552 8752
rect 5568 8688 5632 8752
rect 5648 8688 5712 8752
rect 5728 8688 5792 8752
rect 5808 8688 5872 8752
rect 5888 8688 5952 8752
rect 5968 8688 6032 8752
rect 6048 8688 6112 8752
rect 6128 8688 6192 8752
rect 6208 8688 6272 8752
rect 6288 8688 6352 8752
rect 6368 8688 6432 8752
rect 6448 8688 6512 8752
rect 6528 8688 6592 8752
rect 6608 8688 6672 8752
rect 6688 8688 6752 8752
rect 6768 8688 6832 8752
rect 6848 8688 6912 8752
rect 6928 8688 6992 8752
rect 7008 8688 7072 8752
rect 7088 8688 7152 8752
rect 7168 8688 7232 8752
rect 7248 8688 7312 8752
rect 7328 8688 7392 8752
rect 7408 8688 7472 8752
rect 7488 8688 7552 8752
rect 7568 8688 7632 8752
rect 7648 8688 7712 8752
rect 7728 8688 7792 8752
rect 7808 8688 7872 8752
rect 7888 8688 7952 8752
rect 7968 8688 8032 8752
rect 8048 8688 8112 8752
rect 8128 8688 8192 8752
rect 8208 8688 8272 8752
rect 8288 8688 8352 8752
rect 8368 8688 8432 8752
rect 8448 8688 8512 8752
rect 8528 8688 8592 8752
rect 8608 8688 8672 8752
rect 8688 8688 8752 8752
rect 8768 8688 8832 8752
rect 8848 8688 8912 8752
rect 8928 8688 8992 8752
rect 14112 8688 14176 8752
rect 14192 8688 14256 8752
rect 14272 8688 14336 8752
rect 14352 8688 14416 8752
rect 24112 8688 24176 8752
rect 24192 8688 24256 8752
rect 24272 8688 24336 8752
rect 24352 8688 24416 8752
rect 36376 8688 36440 8752
rect 36456 8688 36520 8752
rect 36536 8688 36600 8752
rect 36616 8688 36680 8752
rect 36696 8688 36760 8752
rect 36776 8688 36840 8752
rect 36856 8688 36920 8752
rect 36936 8688 37000 8752
rect 37016 8688 37080 8752
rect 37096 8688 37160 8752
rect 37176 8688 37240 8752
rect 37256 8688 37320 8752
rect 37336 8688 37400 8752
rect 37416 8688 37480 8752
rect 37496 8688 37560 8752
rect 37576 8688 37640 8752
rect 37656 8688 37720 8752
rect 37736 8688 37800 8752
rect 37816 8688 37880 8752
rect 37896 8688 37960 8752
rect 37976 8688 38040 8752
rect 38056 8688 38120 8752
rect 38136 8688 38200 8752
rect 38216 8688 38280 8752
rect 38296 8688 38360 8752
rect 38376 8688 38440 8752
rect 38456 8688 38520 8752
rect 38536 8688 38600 8752
rect 38616 8688 38680 8752
rect 38696 8688 38760 8752
rect 38776 8688 38840 8752
rect 38856 8688 38920 8752
rect 38936 8688 39000 8752
rect 39016 8688 39080 8752
rect 39096 8688 39160 8752
rect 39176 8688 39240 8752
rect 39256 8688 39320 8752
rect 39336 8688 39400 8752
rect 39416 8688 39480 8752
rect 39496 8688 39560 8752
rect 39576 8688 39640 8752
rect 39656 8688 39720 8752
rect 39736 8688 39800 8752
rect 39816 8688 39880 8752
rect 39896 8688 39960 8752
rect 39976 8688 40040 8752
rect 40056 8688 40120 8752
rect 40136 8688 40200 8752
rect 40216 8688 40280 8752
rect 40296 8688 40360 8752
rect 5008 8608 5072 8672
rect 5088 8608 5152 8672
rect 5168 8608 5232 8672
rect 5248 8608 5312 8672
rect 5328 8608 5392 8672
rect 5408 8608 5472 8672
rect 5488 8608 5552 8672
rect 5568 8608 5632 8672
rect 5648 8608 5712 8672
rect 5728 8608 5792 8672
rect 5808 8608 5872 8672
rect 5888 8608 5952 8672
rect 5968 8608 6032 8672
rect 6048 8608 6112 8672
rect 6128 8608 6192 8672
rect 6208 8608 6272 8672
rect 6288 8608 6352 8672
rect 6368 8608 6432 8672
rect 6448 8608 6512 8672
rect 6528 8608 6592 8672
rect 6608 8608 6672 8672
rect 6688 8608 6752 8672
rect 6768 8608 6832 8672
rect 6848 8608 6912 8672
rect 6928 8608 6992 8672
rect 7008 8608 7072 8672
rect 7088 8608 7152 8672
rect 7168 8608 7232 8672
rect 7248 8608 7312 8672
rect 7328 8608 7392 8672
rect 7408 8608 7472 8672
rect 7488 8608 7552 8672
rect 7568 8608 7632 8672
rect 7648 8608 7712 8672
rect 7728 8608 7792 8672
rect 7808 8608 7872 8672
rect 7888 8608 7952 8672
rect 7968 8608 8032 8672
rect 8048 8608 8112 8672
rect 8128 8608 8192 8672
rect 8208 8608 8272 8672
rect 8288 8608 8352 8672
rect 8368 8608 8432 8672
rect 8448 8608 8512 8672
rect 8528 8608 8592 8672
rect 8608 8608 8672 8672
rect 8688 8608 8752 8672
rect 8768 8608 8832 8672
rect 8848 8608 8912 8672
rect 8928 8608 8992 8672
rect 14112 8608 14176 8672
rect 14192 8608 14256 8672
rect 14272 8608 14336 8672
rect 14352 8608 14416 8672
rect 24112 8608 24176 8672
rect 24192 8608 24256 8672
rect 24272 8608 24336 8672
rect 24352 8608 24416 8672
rect 36376 8608 36440 8672
rect 36456 8608 36520 8672
rect 36536 8608 36600 8672
rect 36616 8608 36680 8672
rect 36696 8608 36760 8672
rect 36776 8608 36840 8672
rect 36856 8608 36920 8672
rect 36936 8608 37000 8672
rect 37016 8608 37080 8672
rect 37096 8608 37160 8672
rect 37176 8608 37240 8672
rect 37256 8608 37320 8672
rect 37336 8608 37400 8672
rect 37416 8608 37480 8672
rect 37496 8608 37560 8672
rect 37576 8608 37640 8672
rect 37656 8608 37720 8672
rect 37736 8608 37800 8672
rect 37816 8608 37880 8672
rect 37896 8608 37960 8672
rect 37976 8608 38040 8672
rect 38056 8608 38120 8672
rect 38136 8608 38200 8672
rect 38216 8608 38280 8672
rect 38296 8608 38360 8672
rect 38376 8608 38440 8672
rect 38456 8608 38520 8672
rect 38536 8608 38600 8672
rect 38616 8608 38680 8672
rect 38696 8608 38760 8672
rect 38776 8608 38840 8672
rect 38856 8608 38920 8672
rect 38936 8608 39000 8672
rect 39016 8608 39080 8672
rect 39096 8608 39160 8672
rect 39176 8608 39240 8672
rect 39256 8608 39320 8672
rect 39336 8608 39400 8672
rect 39416 8608 39480 8672
rect 39496 8608 39560 8672
rect 39576 8608 39640 8672
rect 39656 8608 39720 8672
rect 39736 8608 39800 8672
rect 39816 8608 39880 8672
rect 39896 8608 39960 8672
rect 39976 8608 40040 8672
rect 40056 8608 40120 8672
rect 40136 8608 40200 8672
rect 40216 8608 40280 8672
rect 40296 8608 40360 8672
rect 5008 8528 5072 8592
rect 5088 8528 5152 8592
rect 5168 8528 5232 8592
rect 5248 8528 5312 8592
rect 5328 8528 5392 8592
rect 5408 8528 5472 8592
rect 5488 8528 5552 8592
rect 5568 8528 5632 8592
rect 5648 8528 5712 8592
rect 5728 8528 5792 8592
rect 5808 8528 5872 8592
rect 5888 8528 5952 8592
rect 5968 8528 6032 8592
rect 6048 8528 6112 8592
rect 6128 8528 6192 8592
rect 6208 8528 6272 8592
rect 6288 8528 6352 8592
rect 6368 8528 6432 8592
rect 6448 8528 6512 8592
rect 6528 8528 6592 8592
rect 6608 8528 6672 8592
rect 6688 8528 6752 8592
rect 6768 8528 6832 8592
rect 6848 8528 6912 8592
rect 6928 8528 6992 8592
rect 7008 8528 7072 8592
rect 7088 8528 7152 8592
rect 7168 8528 7232 8592
rect 7248 8528 7312 8592
rect 7328 8528 7392 8592
rect 7408 8528 7472 8592
rect 7488 8528 7552 8592
rect 7568 8528 7632 8592
rect 7648 8528 7712 8592
rect 7728 8528 7792 8592
rect 7808 8528 7872 8592
rect 7888 8528 7952 8592
rect 7968 8528 8032 8592
rect 8048 8528 8112 8592
rect 8128 8528 8192 8592
rect 8208 8528 8272 8592
rect 8288 8528 8352 8592
rect 8368 8528 8432 8592
rect 8448 8528 8512 8592
rect 8528 8528 8592 8592
rect 8608 8528 8672 8592
rect 8688 8528 8752 8592
rect 8768 8528 8832 8592
rect 8848 8528 8912 8592
rect 8928 8528 8992 8592
rect 14112 8528 14176 8592
rect 14192 8528 14256 8592
rect 14272 8528 14336 8592
rect 14352 8528 14416 8592
rect 24112 8528 24176 8592
rect 24192 8528 24256 8592
rect 24272 8528 24336 8592
rect 24352 8528 24416 8592
rect 36376 8528 36440 8592
rect 36456 8528 36520 8592
rect 36536 8528 36600 8592
rect 36616 8528 36680 8592
rect 36696 8528 36760 8592
rect 36776 8528 36840 8592
rect 36856 8528 36920 8592
rect 36936 8528 37000 8592
rect 37016 8528 37080 8592
rect 37096 8528 37160 8592
rect 37176 8528 37240 8592
rect 37256 8528 37320 8592
rect 37336 8528 37400 8592
rect 37416 8528 37480 8592
rect 37496 8528 37560 8592
rect 37576 8528 37640 8592
rect 37656 8528 37720 8592
rect 37736 8528 37800 8592
rect 37816 8528 37880 8592
rect 37896 8528 37960 8592
rect 37976 8528 38040 8592
rect 38056 8528 38120 8592
rect 38136 8528 38200 8592
rect 38216 8528 38280 8592
rect 38296 8528 38360 8592
rect 38376 8528 38440 8592
rect 38456 8528 38520 8592
rect 38536 8528 38600 8592
rect 38616 8528 38680 8592
rect 38696 8528 38760 8592
rect 38776 8528 38840 8592
rect 38856 8528 38920 8592
rect 38936 8528 39000 8592
rect 39016 8528 39080 8592
rect 39096 8528 39160 8592
rect 39176 8528 39240 8592
rect 39256 8528 39320 8592
rect 39336 8528 39400 8592
rect 39416 8528 39480 8592
rect 39496 8528 39560 8592
rect 39576 8528 39640 8592
rect 39656 8528 39720 8592
rect 39736 8528 39800 8592
rect 39816 8528 39880 8592
rect 39896 8528 39960 8592
rect 39976 8528 40040 8592
rect 40056 8528 40120 8592
rect 40136 8528 40200 8592
rect 40216 8528 40280 8592
rect 40296 8528 40360 8592
rect 5008 8448 5072 8512
rect 5088 8448 5152 8512
rect 5168 8448 5232 8512
rect 5248 8448 5312 8512
rect 5328 8448 5392 8512
rect 5408 8448 5472 8512
rect 5488 8448 5552 8512
rect 5568 8448 5632 8512
rect 5648 8448 5712 8512
rect 5728 8448 5792 8512
rect 5808 8448 5872 8512
rect 5888 8448 5952 8512
rect 5968 8448 6032 8512
rect 6048 8448 6112 8512
rect 6128 8448 6192 8512
rect 6208 8448 6272 8512
rect 6288 8448 6352 8512
rect 6368 8448 6432 8512
rect 6448 8448 6512 8512
rect 6528 8448 6592 8512
rect 6608 8448 6672 8512
rect 6688 8448 6752 8512
rect 6768 8448 6832 8512
rect 6848 8448 6912 8512
rect 6928 8448 6992 8512
rect 7008 8448 7072 8512
rect 7088 8448 7152 8512
rect 7168 8448 7232 8512
rect 7248 8448 7312 8512
rect 7328 8448 7392 8512
rect 7408 8448 7472 8512
rect 7488 8448 7552 8512
rect 7568 8448 7632 8512
rect 7648 8448 7712 8512
rect 7728 8448 7792 8512
rect 7808 8448 7872 8512
rect 7888 8448 7952 8512
rect 7968 8448 8032 8512
rect 8048 8448 8112 8512
rect 8128 8448 8192 8512
rect 8208 8448 8272 8512
rect 8288 8448 8352 8512
rect 8368 8448 8432 8512
rect 8448 8448 8512 8512
rect 8528 8448 8592 8512
rect 8608 8448 8672 8512
rect 8688 8448 8752 8512
rect 8768 8448 8832 8512
rect 8848 8448 8912 8512
rect 8928 8448 8992 8512
rect 14112 8448 14176 8512
rect 14192 8448 14256 8512
rect 14272 8448 14336 8512
rect 14352 8448 14416 8512
rect 24112 8448 24176 8512
rect 24192 8448 24256 8512
rect 24272 8448 24336 8512
rect 24352 8448 24416 8512
rect 36376 8448 36440 8512
rect 36456 8448 36520 8512
rect 36536 8448 36600 8512
rect 36616 8448 36680 8512
rect 36696 8448 36760 8512
rect 36776 8448 36840 8512
rect 36856 8448 36920 8512
rect 36936 8448 37000 8512
rect 37016 8448 37080 8512
rect 37096 8448 37160 8512
rect 37176 8448 37240 8512
rect 37256 8448 37320 8512
rect 37336 8448 37400 8512
rect 37416 8448 37480 8512
rect 37496 8448 37560 8512
rect 37576 8448 37640 8512
rect 37656 8448 37720 8512
rect 37736 8448 37800 8512
rect 37816 8448 37880 8512
rect 37896 8448 37960 8512
rect 37976 8448 38040 8512
rect 38056 8448 38120 8512
rect 38136 8448 38200 8512
rect 38216 8448 38280 8512
rect 38296 8448 38360 8512
rect 38376 8448 38440 8512
rect 38456 8448 38520 8512
rect 38536 8448 38600 8512
rect 38616 8448 38680 8512
rect 38696 8448 38760 8512
rect 38776 8448 38840 8512
rect 38856 8448 38920 8512
rect 38936 8448 39000 8512
rect 39016 8448 39080 8512
rect 39096 8448 39160 8512
rect 39176 8448 39240 8512
rect 39256 8448 39320 8512
rect 39336 8448 39400 8512
rect 39416 8448 39480 8512
rect 39496 8448 39560 8512
rect 39576 8448 39640 8512
rect 39656 8448 39720 8512
rect 39736 8448 39800 8512
rect 39816 8448 39880 8512
rect 39896 8448 39960 8512
rect 39976 8448 40040 8512
rect 40056 8448 40120 8512
rect 40136 8448 40200 8512
rect 40216 8448 40280 8512
rect 40296 8448 40360 8512
rect 5008 8368 5072 8432
rect 5088 8368 5152 8432
rect 5168 8368 5232 8432
rect 5248 8368 5312 8432
rect 5328 8368 5392 8432
rect 5408 8368 5472 8432
rect 5488 8368 5552 8432
rect 5568 8368 5632 8432
rect 5648 8368 5712 8432
rect 5728 8368 5792 8432
rect 5808 8368 5872 8432
rect 5888 8368 5952 8432
rect 5968 8368 6032 8432
rect 6048 8368 6112 8432
rect 6128 8368 6192 8432
rect 6208 8368 6272 8432
rect 6288 8368 6352 8432
rect 6368 8368 6432 8432
rect 6448 8368 6512 8432
rect 6528 8368 6592 8432
rect 6608 8368 6672 8432
rect 6688 8368 6752 8432
rect 6768 8368 6832 8432
rect 6848 8368 6912 8432
rect 6928 8368 6992 8432
rect 7008 8368 7072 8432
rect 7088 8368 7152 8432
rect 7168 8368 7232 8432
rect 7248 8368 7312 8432
rect 7328 8368 7392 8432
rect 7408 8368 7472 8432
rect 7488 8368 7552 8432
rect 7568 8368 7632 8432
rect 7648 8368 7712 8432
rect 7728 8368 7792 8432
rect 7808 8368 7872 8432
rect 7888 8368 7952 8432
rect 7968 8368 8032 8432
rect 8048 8368 8112 8432
rect 8128 8368 8192 8432
rect 8208 8368 8272 8432
rect 8288 8368 8352 8432
rect 8368 8368 8432 8432
rect 8448 8368 8512 8432
rect 8528 8368 8592 8432
rect 8608 8368 8672 8432
rect 8688 8368 8752 8432
rect 8768 8368 8832 8432
rect 8848 8368 8912 8432
rect 8928 8368 8992 8432
rect 14112 8368 14176 8432
rect 14192 8368 14256 8432
rect 14272 8368 14336 8432
rect 14352 8368 14416 8432
rect 24112 8368 24176 8432
rect 24192 8368 24256 8432
rect 24272 8368 24336 8432
rect 24352 8368 24416 8432
rect 36376 8368 36440 8432
rect 36456 8368 36520 8432
rect 36536 8368 36600 8432
rect 36616 8368 36680 8432
rect 36696 8368 36760 8432
rect 36776 8368 36840 8432
rect 36856 8368 36920 8432
rect 36936 8368 37000 8432
rect 37016 8368 37080 8432
rect 37096 8368 37160 8432
rect 37176 8368 37240 8432
rect 37256 8368 37320 8432
rect 37336 8368 37400 8432
rect 37416 8368 37480 8432
rect 37496 8368 37560 8432
rect 37576 8368 37640 8432
rect 37656 8368 37720 8432
rect 37736 8368 37800 8432
rect 37816 8368 37880 8432
rect 37896 8368 37960 8432
rect 37976 8368 38040 8432
rect 38056 8368 38120 8432
rect 38136 8368 38200 8432
rect 38216 8368 38280 8432
rect 38296 8368 38360 8432
rect 38376 8368 38440 8432
rect 38456 8368 38520 8432
rect 38536 8368 38600 8432
rect 38616 8368 38680 8432
rect 38696 8368 38760 8432
rect 38776 8368 38840 8432
rect 38856 8368 38920 8432
rect 38936 8368 39000 8432
rect 39016 8368 39080 8432
rect 39096 8368 39160 8432
rect 39176 8368 39240 8432
rect 39256 8368 39320 8432
rect 39336 8368 39400 8432
rect 39416 8368 39480 8432
rect 39496 8368 39560 8432
rect 39576 8368 39640 8432
rect 39656 8368 39720 8432
rect 39736 8368 39800 8432
rect 39816 8368 39880 8432
rect 39896 8368 39960 8432
rect 39976 8368 40040 8432
rect 40056 8368 40120 8432
rect 40136 8368 40200 8432
rect 40216 8368 40280 8432
rect 40296 8368 40360 8432
rect 5008 8288 5072 8352
rect 5088 8288 5152 8352
rect 5168 8288 5232 8352
rect 5248 8288 5312 8352
rect 5328 8288 5392 8352
rect 5408 8288 5472 8352
rect 5488 8288 5552 8352
rect 5568 8288 5632 8352
rect 5648 8288 5712 8352
rect 5728 8288 5792 8352
rect 5808 8288 5872 8352
rect 5888 8288 5952 8352
rect 5968 8288 6032 8352
rect 6048 8288 6112 8352
rect 6128 8288 6192 8352
rect 6208 8288 6272 8352
rect 6288 8288 6352 8352
rect 6368 8288 6432 8352
rect 6448 8288 6512 8352
rect 6528 8288 6592 8352
rect 6608 8288 6672 8352
rect 6688 8288 6752 8352
rect 6768 8288 6832 8352
rect 6848 8288 6912 8352
rect 6928 8288 6992 8352
rect 7008 8288 7072 8352
rect 7088 8288 7152 8352
rect 7168 8288 7232 8352
rect 7248 8288 7312 8352
rect 7328 8288 7392 8352
rect 7408 8288 7472 8352
rect 7488 8288 7552 8352
rect 7568 8288 7632 8352
rect 7648 8288 7712 8352
rect 7728 8288 7792 8352
rect 7808 8288 7872 8352
rect 7888 8288 7952 8352
rect 7968 8288 8032 8352
rect 8048 8288 8112 8352
rect 8128 8288 8192 8352
rect 8208 8288 8272 8352
rect 8288 8288 8352 8352
rect 8368 8288 8432 8352
rect 8448 8288 8512 8352
rect 8528 8288 8592 8352
rect 8608 8288 8672 8352
rect 8688 8288 8752 8352
rect 8768 8288 8832 8352
rect 8848 8288 8912 8352
rect 8928 8288 8992 8352
rect 14112 8288 14176 8352
rect 14192 8288 14256 8352
rect 14272 8288 14336 8352
rect 14352 8288 14416 8352
rect 24112 8288 24176 8352
rect 24192 8288 24256 8352
rect 24272 8288 24336 8352
rect 24352 8288 24416 8352
rect 36376 8288 36440 8352
rect 36456 8288 36520 8352
rect 36536 8288 36600 8352
rect 36616 8288 36680 8352
rect 36696 8288 36760 8352
rect 36776 8288 36840 8352
rect 36856 8288 36920 8352
rect 36936 8288 37000 8352
rect 37016 8288 37080 8352
rect 37096 8288 37160 8352
rect 37176 8288 37240 8352
rect 37256 8288 37320 8352
rect 37336 8288 37400 8352
rect 37416 8288 37480 8352
rect 37496 8288 37560 8352
rect 37576 8288 37640 8352
rect 37656 8288 37720 8352
rect 37736 8288 37800 8352
rect 37816 8288 37880 8352
rect 37896 8288 37960 8352
rect 37976 8288 38040 8352
rect 38056 8288 38120 8352
rect 38136 8288 38200 8352
rect 38216 8288 38280 8352
rect 38296 8288 38360 8352
rect 38376 8288 38440 8352
rect 38456 8288 38520 8352
rect 38536 8288 38600 8352
rect 38616 8288 38680 8352
rect 38696 8288 38760 8352
rect 38776 8288 38840 8352
rect 38856 8288 38920 8352
rect 38936 8288 39000 8352
rect 39016 8288 39080 8352
rect 39096 8288 39160 8352
rect 39176 8288 39240 8352
rect 39256 8288 39320 8352
rect 39336 8288 39400 8352
rect 39416 8288 39480 8352
rect 39496 8288 39560 8352
rect 39576 8288 39640 8352
rect 39656 8288 39720 8352
rect 39736 8288 39800 8352
rect 39816 8288 39880 8352
rect 39896 8288 39960 8352
rect 39976 8288 40040 8352
rect 40056 8288 40120 8352
rect 40136 8288 40200 8352
rect 40216 8288 40280 8352
rect 40296 8288 40360 8352
rect 5008 8208 5072 8272
rect 5088 8208 5152 8272
rect 5168 8208 5232 8272
rect 5248 8208 5312 8272
rect 5328 8208 5392 8272
rect 5408 8208 5472 8272
rect 5488 8208 5552 8272
rect 5568 8208 5632 8272
rect 5648 8208 5712 8272
rect 5728 8208 5792 8272
rect 5808 8208 5872 8272
rect 5888 8208 5952 8272
rect 5968 8208 6032 8272
rect 6048 8208 6112 8272
rect 6128 8208 6192 8272
rect 6208 8208 6272 8272
rect 6288 8208 6352 8272
rect 6368 8208 6432 8272
rect 6448 8208 6512 8272
rect 6528 8208 6592 8272
rect 6608 8208 6672 8272
rect 6688 8208 6752 8272
rect 6768 8208 6832 8272
rect 6848 8208 6912 8272
rect 6928 8208 6992 8272
rect 7008 8208 7072 8272
rect 7088 8208 7152 8272
rect 7168 8208 7232 8272
rect 7248 8208 7312 8272
rect 7328 8208 7392 8272
rect 7408 8208 7472 8272
rect 7488 8208 7552 8272
rect 7568 8208 7632 8272
rect 7648 8208 7712 8272
rect 7728 8208 7792 8272
rect 7808 8208 7872 8272
rect 7888 8208 7952 8272
rect 7968 8208 8032 8272
rect 8048 8208 8112 8272
rect 8128 8208 8192 8272
rect 8208 8208 8272 8272
rect 8288 8208 8352 8272
rect 8368 8208 8432 8272
rect 8448 8208 8512 8272
rect 8528 8208 8592 8272
rect 8608 8208 8672 8272
rect 8688 8208 8752 8272
rect 8768 8208 8832 8272
rect 8848 8208 8912 8272
rect 8928 8208 8992 8272
rect 14112 8208 14176 8272
rect 14192 8208 14256 8272
rect 14272 8208 14336 8272
rect 14352 8208 14416 8272
rect 24112 8208 24176 8272
rect 24192 8208 24256 8272
rect 24272 8208 24336 8272
rect 24352 8208 24416 8272
rect 36376 8208 36440 8272
rect 36456 8208 36520 8272
rect 36536 8208 36600 8272
rect 36616 8208 36680 8272
rect 36696 8208 36760 8272
rect 36776 8208 36840 8272
rect 36856 8208 36920 8272
rect 36936 8208 37000 8272
rect 37016 8208 37080 8272
rect 37096 8208 37160 8272
rect 37176 8208 37240 8272
rect 37256 8208 37320 8272
rect 37336 8208 37400 8272
rect 37416 8208 37480 8272
rect 37496 8208 37560 8272
rect 37576 8208 37640 8272
rect 37656 8208 37720 8272
rect 37736 8208 37800 8272
rect 37816 8208 37880 8272
rect 37896 8208 37960 8272
rect 37976 8208 38040 8272
rect 38056 8208 38120 8272
rect 38136 8208 38200 8272
rect 38216 8208 38280 8272
rect 38296 8208 38360 8272
rect 38376 8208 38440 8272
rect 38456 8208 38520 8272
rect 38536 8208 38600 8272
rect 38616 8208 38680 8272
rect 38696 8208 38760 8272
rect 38776 8208 38840 8272
rect 38856 8208 38920 8272
rect 38936 8208 39000 8272
rect 39016 8208 39080 8272
rect 39096 8208 39160 8272
rect 39176 8208 39240 8272
rect 39256 8208 39320 8272
rect 39336 8208 39400 8272
rect 39416 8208 39480 8272
rect 39496 8208 39560 8272
rect 39576 8208 39640 8272
rect 39656 8208 39720 8272
rect 39736 8208 39800 8272
rect 39816 8208 39880 8272
rect 39896 8208 39960 8272
rect 39976 8208 40040 8272
rect 40056 8208 40120 8272
rect 40136 8208 40200 8272
rect 40216 8208 40280 8272
rect 40296 8208 40360 8272
rect 5008 8128 5072 8192
rect 5088 8128 5152 8192
rect 5168 8128 5232 8192
rect 5248 8128 5312 8192
rect 5328 8128 5392 8192
rect 5408 8128 5472 8192
rect 5488 8128 5552 8192
rect 5568 8128 5632 8192
rect 5648 8128 5712 8192
rect 5728 8128 5792 8192
rect 5808 8128 5872 8192
rect 5888 8128 5952 8192
rect 5968 8128 6032 8192
rect 6048 8128 6112 8192
rect 6128 8128 6192 8192
rect 6208 8128 6272 8192
rect 6288 8128 6352 8192
rect 6368 8128 6432 8192
rect 6448 8128 6512 8192
rect 6528 8128 6592 8192
rect 6608 8128 6672 8192
rect 6688 8128 6752 8192
rect 6768 8128 6832 8192
rect 6848 8128 6912 8192
rect 6928 8128 6992 8192
rect 7008 8128 7072 8192
rect 7088 8128 7152 8192
rect 7168 8128 7232 8192
rect 7248 8128 7312 8192
rect 7328 8128 7392 8192
rect 7408 8128 7472 8192
rect 7488 8128 7552 8192
rect 7568 8128 7632 8192
rect 7648 8128 7712 8192
rect 7728 8128 7792 8192
rect 7808 8128 7872 8192
rect 7888 8128 7952 8192
rect 7968 8128 8032 8192
rect 8048 8128 8112 8192
rect 8128 8128 8192 8192
rect 8208 8128 8272 8192
rect 8288 8128 8352 8192
rect 8368 8128 8432 8192
rect 8448 8128 8512 8192
rect 8528 8128 8592 8192
rect 8608 8128 8672 8192
rect 8688 8128 8752 8192
rect 8768 8128 8832 8192
rect 8848 8128 8912 8192
rect 8928 8128 8992 8192
rect 14112 8128 14176 8192
rect 14192 8128 14256 8192
rect 14272 8128 14336 8192
rect 14352 8128 14416 8192
rect 24112 8128 24176 8192
rect 24192 8128 24256 8192
rect 24272 8128 24336 8192
rect 24352 8128 24416 8192
rect 36376 8128 36440 8192
rect 36456 8128 36520 8192
rect 36536 8128 36600 8192
rect 36616 8128 36680 8192
rect 36696 8128 36760 8192
rect 36776 8128 36840 8192
rect 36856 8128 36920 8192
rect 36936 8128 37000 8192
rect 37016 8128 37080 8192
rect 37096 8128 37160 8192
rect 37176 8128 37240 8192
rect 37256 8128 37320 8192
rect 37336 8128 37400 8192
rect 37416 8128 37480 8192
rect 37496 8128 37560 8192
rect 37576 8128 37640 8192
rect 37656 8128 37720 8192
rect 37736 8128 37800 8192
rect 37816 8128 37880 8192
rect 37896 8128 37960 8192
rect 37976 8128 38040 8192
rect 38056 8128 38120 8192
rect 38136 8128 38200 8192
rect 38216 8128 38280 8192
rect 38296 8128 38360 8192
rect 38376 8128 38440 8192
rect 38456 8128 38520 8192
rect 38536 8128 38600 8192
rect 38616 8128 38680 8192
rect 38696 8128 38760 8192
rect 38776 8128 38840 8192
rect 38856 8128 38920 8192
rect 38936 8128 39000 8192
rect 39016 8128 39080 8192
rect 39096 8128 39160 8192
rect 39176 8128 39240 8192
rect 39256 8128 39320 8192
rect 39336 8128 39400 8192
rect 39416 8128 39480 8192
rect 39496 8128 39560 8192
rect 39576 8128 39640 8192
rect 39656 8128 39720 8192
rect 39736 8128 39800 8192
rect 39816 8128 39880 8192
rect 39896 8128 39960 8192
rect 39976 8128 40040 8192
rect 40056 8128 40120 8192
rect 40136 8128 40200 8192
rect 40216 8128 40280 8192
rect 40296 8128 40360 8192
rect 5008 8048 5072 8112
rect 5088 8048 5152 8112
rect 5168 8048 5232 8112
rect 5248 8048 5312 8112
rect 5328 8048 5392 8112
rect 5408 8048 5472 8112
rect 5488 8048 5552 8112
rect 5568 8048 5632 8112
rect 5648 8048 5712 8112
rect 5728 8048 5792 8112
rect 5808 8048 5872 8112
rect 5888 8048 5952 8112
rect 5968 8048 6032 8112
rect 6048 8048 6112 8112
rect 6128 8048 6192 8112
rect 6208 8048 6272 8112
rect 6288 8048 6352 8112
rect 6368 8048 6432 8112
rect 6448 8048 6512 8112
rect 6528 8048 6592 8112
rect 6608 8048 6672 8112
rect 6688 8048 6752 8112
rect 6768 8048 6832 8112
rect 6848 8048 6912 8112
rect 6928 8048 6992 8112
rect 7008 8048 7072 8112
rect 7088 8048 7152 8112
rect 7168 8048 7232 8112
rect 7248 8048 7312 8112
rect 7328 8048 7392 8112
rect 7408 8048 7472 8112
rect 7488 8048 7552 8112
rect 7568 8048 7632 8112
rect 7648 8048 7712 8112
rect 7728 8048 7792 8112
rect 7808 8048 7872 8112
rect 7888 8048 7952 8112
rect 7968 8048 8032 8112
rect 8048 8048 8112 8112
rect 8128 8048 8192 8112
rect 8208 8048 8272 8112
rect 8288 8048 8352 8112
rect 8368 8048 8432 8112
rect 8448 8048 8512 8112
rect 8528 8048 8592 8112
rect 8608 8048 8672 8112
rect 8688 8048 8752 8112
rect 8768 8048 8832 8112
rect 8848 8048 8912 8112
rect 8928 8048 8992 8112
rect 14112 8048 14176 8112
rect 14192 8048 14256 8112
rect 14272 8048 14336 8112
rect 14352 8048 14416 8112
rect 24112 8048 24176 8112
rect 24192 8048 24256 8112
rect 24272 8048 24336 8112
rect 24352 8048 24416 8112
rect 36376 8048 36440 8112
rect 36456 8048 36520 8112
rect 36536 8048 36600 8112
rect 36616 8048 36680 8112
rect 36696 8048 36760 8112
rect 36776 8048 36840 8112
rect 36856 8048 36920 8112
rect 36936 8048 37000 8112
rect 37016 8048 37080 8112
rect 37096 8048 37160 8112
rect 37176 8048 37240 8112
rect 37256 8048 37320 8112
rect 37336 8048 37400 8112
rect 37416 8048 37480 8112
rect 37496 8048 37560 8112
rect 37576 8048 37640 8112
rect 37656 8048 37720 8112
rect 37736 8048 37800 8112
rect 37816 8048 37880 8112
rect 37896 8048 37960 8112
rect 37976 8048 38040 8112
rect 38056 8048 38120 8112
rect 38136 8048 38200 8112
rect 38216 8048 38280 8112
rect 38296 8048 38360 8112
rect 38376 8048 38440 8112
rect 38456 8048 38520 8112
rect 38536 8048 38600 8112
rect 38616 8048 38680 8112
rect 38696 8048 38760 8112
rect 38776 8048 38840 8112
rect 38856 8048 38920 8112
rect 38936 8048 39000 8112
rect 39016 8048 39080 8112
rect 39096 8048 39160 8112
rect 39176 8048 39240 8112
rect 39256 8048 39320 8112
rect 39336 8048 39400 8112
rect 39416 8048 39480 8112
rect 39496 8048 39560 8112
rect 39576 8048 39640 8112
rect 39656 8048 39720 8112
rect 39736 8048 39800 8112
rect 39816 8048 39880 8112
rect 39896 8048 39960 8112
rect 39976 8048 40040 8112
rect 40056 8048 40120 8112
rect 40136 8048 40200 8112
rect 40216 8048 40280 8112
rect 40296 8048 40360 8112
rect 5008 7968 5072 8032
rect 5088 7968 5152 8032
rect 5168 7968 5232 8032
rect 5248 7968 5312 8032
rect 5328 7968 5392 8032
rect 5408 7968 5472 8032
rect 5488 7968 5552 8032
rect 5568 7968 5632 8032
rect 5648 7968 5712 8032
rect 5728 7968 5792 8032
rect 5808 7968 5872 8032
rect 5888 7968 5952 8032
rect 5968 7968 6032 8032
rect 6048 7968 6112 8032
rect 6128 7968 6192 8032
rect 6208 7968 6272 8032
rect 6288 7968 6352 8032
rect 6368 7968 6432 8032
rect 6448 7968 6512 8032
rect 6528 7968 6592 8032
rect 6608 7968 6672 8032
rect 6688 7968 6752 8032
rect 6768 7968 6832 8032
rect 6848 7968 6912 8032
rect 6928 7968 6992 8032
rect 7008 7968 7072 8032
rect 7088 7968 7152 8032
rect 7168 7968 7232 8032
rect 7248 7968 7312 8032
rect 7328 7968 7392 8032
rect 7408 7968 7472 8032
rect 7488 7968 7552 8032
rect 7568 7968 7632 8032
rect 7648 7968 7712 8032
rect 7728 7968 7792 8032
rect 7808 7968 7872 8032
rect 7888 7968 7952 8032
rect 7968 7968 8032 8032
rect 8048 7968 8112 8032
rect 8128 7968 8192 8032
rect 8208 7968 8272 8032
rect 8288 7968 8352 8032
rect 8368 7968 8432 8032
rect 8448 7968 8512 8032
rect 8528 7968 8592 8032
rect 8608 7968 8672 8032
rect 8688 7968 8752 8032
rect 8768 7968 8832 8032
rect 8848 7968 8912 8032
rect 8928 7968 8992 8032
rect 14112 7968 14176 8032
rect 14192 7968 14256 8032
rect 14272 7968 14336 8032
rect 14352 7968 14416 8032
rect 24112 7968 24176 8032
rect 24192 7968 24256 8032
rect 24272 7968 24336 8032
rect 24352 7968 24416 8032
rect 36376 7968 36440 8032
rect 36456 7968 36520 8032
rect 36536 7968 36600 8032
rect 36616 7968 36680 8032
rect 36696 7968 36760 8032
rect 36776 7968 36840 8032
rect 36856 7968 36920 8032
rect 36936 7968 37000 8032
rect 37016 7968 37080 8032
rect 37096 7968 37160 8032
rect 37176 7968 37240 8032
rect 37256 7968 37320 8032
rect 37336 7968 37400 8032
rect 37416 7968 37480 8032
rect 37496 7968 37560 8032
rect 37576 7968 37640 8032
rect 37656 7968 37720 8032
rect 37736 7968 37800 8032
rect 37816 7968 37880 8032
rect 37896 7968 37960 8032
rect 37976 7968 38040 8032
rect 38056 7968 38120 8032
rect 38136 7968 38200 8032
rect 38216 7968 38280 8032
rect 38296 7968 38360 8032
rect 38376 7968 38440 8032
rect 38456 7968 38520 8032
rect 38536 7968 38600 8032
rect 38616 7968 38680 8032
rect 38696 7968 38760 8032
rect 38776 7968 38840 8032
rect 38856 7968 38920 8032
rect 38936 7968 39000 8032
rect 39016 7968 39080 8032
rect 39096 7968 39160 8032
rect 39176 7968 39240 8032
rect 39256 7968 39320 8032
rect 39336 7968 39400 8032
rect 39416 7968 39480 8032
rect 39496 7968 39560 8032
rect 39576 7968 39640 8032
rect 39656 7968 39720 8032
rect 39736 7968 39800 8032
rect 39816 7968 39880 8032
rect 39896 7968 39960 8032
rect 39976 7968 40040 8032
rect 40056 7968 40120 8032
rect 40136 7968 40200 8032
rect 40216 7968 40280 8032
rect 40296 7968 40360 8032
rect 5008 7888 5072 7952
rect 5088 7888 5152 7952
rect 5168 7888 5232 7952
rect 5248 7888 5312 7952
rect 5328 7888 5392 7952
rect 5408 7888 5472 7952
rect 5488 7888 5552 7952
rect 5568 7888 5632 7952
rect 5648 7888 5712 7952
rect 5728 7888 5792 7952
rect 5808 7888 5872 7952
rect 5888 7888 5952 7952
rect 5968 7888 6032 7952
rect 6048 7888 6112 7952
rect 6128 7888 6192 7952
rect 6208 7888 6272 7952
rect 6288 7888 6352 7952
rect 6368 7888 6432 7952
rect 6448 7888 6512 7952
rect 6528 7888 6592 7952
rect 6608 7888 6672 7952
rect 6688 7888 6752 7952
rect 6768 7888 6832 7952
rect 6848 7888 6912 7952
rect 6928 7888 6992 7952
rect 7008 7888 7072 7952
rect 7088 7888 7152 7952
rect 7168 7888 7232 7952
rect 7248 7888 7312 7952
rect 7328 7888 7392 7952
rect 7408 7888 7472 7952
rect 7488 7888 7552 7952
rect 7568 7888 7632 7952
rect 7648 7888 7712 7952
rect 7728 7888 7792 7952
rect 7808 7888 7872 7952
rect 7888 7888 7952 7952
rect 7968 7888 8032 7952
rect 8048 7888 8112 7952
rect 8128 7888 8192 7952
rect 8208 7888 8272 7952
rect 8288 7888 8352 7952
rect 8368 7888 8432 7952
rect 8448 7888 8512 7952
rect 8528 7888 8592 7952
rect 8608 7888 8672 7952
rect 8688 7888 8752 7952
rect 8768 7888 8832 7952
rect 8848 7888 8912 7952
rect 8928 7888 8992 7952
rect 14112 7888 14176 7952
rect 14192 7888 14256 7952
rect 14272 7888 14336 7952
rect 14352 7888 14416 7952
rect 24112 7888 24176 7952
rect 24192 7888 24256 7952
rect 24272 7888 24336 7952
rect 24352 7888 24416 7952
rect 36376 7888 36440 7952
rect 36456 7888 36520 7952
rect 36536 7888 36600 7952
rect 36616 7888 36680 7952
rect 36696 7888 36760 7952
rect 36776 7888 36840 7952
rect 36856 7888 36920 7952
rect 36936 7888 37000 7952
rect 37016 7888 37080 7952
rect 37096 7888 37160 7952
rect 37176 7888 37240 7952
rect 37256 7888 37320 7952
rect 37336 7888 37400 7952
rect 37416 7888 37480 7952
rect 37496 7888 37560 7952
rect 37576 7888 37640 7952
rect 37656 7888 37720 7952
rect 37736 7888 37800 7952
rect 37816 7888 37880 7952
rect 37896 7888 37960 7952
rect 37976 7888 38040 7952
rect 38056 7888 38120 7952
rect 38136 7888 38200 7952
rect 38216 7888 38280 7952
rect 38296 7888 38360 7952
rect 38376 7888 38440 7952
rect 38456 7888 38520 7952
rect 38536 7888 38600 7952
rect 38616 7888 38680 7952
rect 38696 7888 38760 7952
rect 38776 7888 38840 7952
rect 38856 7888 38920 7952
rect 38936 7888 39000 7952
rect 39016 7888 39080 7952
rect 39096 7888 39160 7952
rect 39176 7888 39240 7952
rect 39256 7888 39320 7952
rect 39336 7888 39400 7952
rect 39416 7888 39480 7952
rect 39496 7888 39560 7952
rect 39576 7888 39640 7952
rect 39656 7888 39720 7952
rect 39736 7888 39800 7952
rect 39816 7888 39880 7952
rect 39896 7888 39960 7952
rect 39976 7888 40040 7952
rect 40056 7888 40120 7952
rect 40136 7888 40200 7952
rect 40216 7888 40280 7952
rect 40296 7888 40360 7952
rect 5008 7808 5072 7872
rect 5088 7808 5152 7872
rect 5168 7808 5232 7872
rect 5248 7808 5312 7872
rect 5328 7808 5392 7872
rect 5408 7808 5472 7872
rect 5488 7808 5552 7872
rect 5568 7808 5632 7872
rect 5648 7808 5712 7872
rect 5728 7808 5792 7872
rect 5808 7808 5872 7872
rect 5888 7808 5952 7872
rect 5968 7808 6032 7872
rect 6048 7808 6112 7872
rect 6128 7808 6192 7872
rect 6208 7808 6272 7872
rect 6288 7808 6352 7872
rect 6368 7808 6432 7872
rect 6448 7808 6512 7872
rect 6528 7808 6592 7872
rect 6608 7808 6672 7872
rect 6688 7808 6752 7872
rect 6768 7808 6832 7872
rect 6848 7808 6912 7872
rect 6928 7808 6992 7872
rect 7008 7808 7072 7872
rect 7088 7808 7152 7872
rect 7168 7808 7232 7872
rect 7248 7808 7312 7872
rect 7328 7808 7392 7872
rect 7408 7808 7472 7872
rect 7488 7808 7552 7872
rect 7568 7808 7632 7872
rect 7648 7808 7712 7872
rect 7728 7808 7792 7872
rect 7808 7808 7872 7872
rect 7888 7808 7952 7872
rect 7968 7808 8032 7872
rect 8048 7808 8112 7872
rect 8128 7808 8192 7872
rect 8208 7808 8272 7872
rect 8288 7808 8352 7872
rect 8368 7808 8432 7872
rect 8448 7808 8512 7872
rect 8528 7808 8592 7872
rect 8608 7808 8672 7872
rect 8688 7808 8752 7872
rect 8768 7808 8832 7872
rect 8848 7808 8912 7872
rect 8928 7808 8992 7872
rect 14112 7808 14176 7872
rect 14192 7808 14256 7872
rect 14272 7808 14336 7872
rect 14352 7808 14416 7872
rect 24112 7808 24176 7872
rect 24192 7808 24256 7872
rect 24272 7808 24336 7872
rect 24352 7808 24416 7872
rect 36376 7808 36440 7872
rect 36456 7808 36520 7872
rect 36536 7808 36600 7872
rect 36616 7808 36680 7872
rect 36696 7808 36760 7872
rect 36776 7808 36840 7872
rect 36856 7808 36920 7872
rect 36936 7808 37000 7872
rect 37016 7808 37080 7872
rect 37096 7808 37160 7872
rect 37176 7808 37240 7872
rect 37256 7808 37320 7872
rect 37336 7808 37400 7872
rect 37416 7808 37480 7872
rect 37496 7808 37560 7872
rect 37576 7808 37640 7872
rect 37656 7808 37720 7872
rect 37736 7808 37800 7872
rect 37816 7808 37880 7872
rect 37896 7808 37960 7872
rect 37976 7808 38040 7872
rect 38056 7808 38120 7872
rect 38136 7808 38200 7872
rect 38216 7808 38280 7872
rect 38296 7808 38360 7872
rect 38376 7808 38440 7872
rect 38456 7808 38520 7872
rect 38536 7808 38600 7872
rect 38616 7808 38680 7872
rect 38696 7808 38760 7872
rect 38776 7808 38840 7872
rect 38856 7808 38920 7872
rect 38936 7808 39000 7872
rect 39016 7808 39080 7872
rect 39096 7808 39160 7872
rect 39176 7808 39240 7872
rect 39256 7808 39320 7872
rect 39336 7808 39400 7872
rect 39416 7808 39480 7872
rect 39496 7808 39560 7872
rect 39576 7808 39640 7872
rect 39656 7808 39720 7872
rect 39736 7808 39800 7872
rect 39816 7808 39880 7872
rect 39896 7808 39960 7872
rect 39976 7808 40040 7872
rect 40056 7808 40120 7872
rect 40136 7808 40200 7872
rect 40216 7808 40280 7872
rect 40296 7808 40360 7872
rect 5008 7728 5072 7792
rect 5088 7728 5152 7792
rect 5168 7728 5232 7792
rect 5248 7728 5312 7792
rect 5328 7728 5392 7792
rect 5408 7728 5472 7792
rect 5488 7728 5552 7792
rect 5568 7728 5632 7792
rect 5648 7728 5712 7792
rect 5728 7728 5792 7792
rect 5808 7728 5872 7792
rect 5888 7728 5952 7792
rect 5968 7728 6032 7792
rect 6048 7728 6112 7792
rect 6128 7728 6192 7792
rect 6208 7728 6272 7792
rect 6288 7728 6352 7792
rect 6368 7728 6432 7792
rect 6448 7728 6512 7792
rect 6528 7728 6592 7792
rect 6608 7728 6672 7792
rect 6688 7728 6752 7792
rect 6768 7728 6832 7792
rect 6848 7728 6912 7792
rect 6928 7728 6992 7792
rect 7008 7728 7072 7792
rect 7088 7728 7152 7792
rect 7168 7728 7232 7792
rect 7248 7728 7312 7792
rect 7328 7728 7392 7792
rect 7408 7728 7472 7792
rect 7488 7728 7552 7792
rect 7568 7728 7632 7792
rect 7648 7728 7712 7792
rect 7728 7728 7792 7792
rect 7808 7728 7872 7792
rect 7888 7728 7952 7792
rect 7968 7728 8032 7792
rect 8048 7728 8112 7792
rect 8128 7728 8192 7792
rect 8208 7728 8272 7792
rect 8288 7728 8352 7792
rect 8368 7728 8432 7792
rect 8448 7728 8512 7792
rect 8528 7728 8592 7792
rect 8608 7728 8672 7792
rect 8688 7728 8752 7792
rect 8768 7728 8832 7792
rect 8848 7728 8912 7792
rect 8928 7728 8992 7792
rect 14112 7728 14176 7792
rect 14192 7728 14256 7792
rect 14272 7728 14336 7792
rect 14352 7728 14416 7792
rect 24112 7728 24176 7792
rect 24192 7728 24256 7792
rect 24272 7728 24336 7792
rect 24352 7728 24416 7792
rect 36376 7728 36440 7792
rect 36456 7728 36520 7792
rect 36536 7728 36600 7792
rect 36616 7728 36680 7792
rect 36696 7728 36760 7792
rect 36776 7728 36840 7792
rect 36856 7728 36920 7792
rect 36936 7728 37000 7792
rect 37016 7728 37080 7792
rect 37096 7728 37160 7792
rect 37176 7728 37240 7792
rect 37256 7728 37320 7792
rect 37336 7728 37400 7792
rect 37416 7728 37480 7792
rect 37496 7728 37560 7792
rect 37576 7728 37640 7792
rect 37656 7728 37720 7792
rect 37736 7728 37800 7792
rect 37816 7728 37880 7792
rect 37896 7728 37960 7792
rect 37976 7728 38040 7792
rect 38056 7728 38120 7792
rect 38136 7728 38200 7792
rect 38216 7728 38280 7792
rect 38296 7728 38360 7792
rect 38376 7728 38440 7792
rect 38456 7728 38520 7792
rect 38536 7728 38600 7792
rect 38616 7728 38680 7792
rect 38696 7728 38760 7792
rect 38776 7728 38840 7792
rect 38856 7728 38920 7792
rect 38936 7728 39000 7792
rect 39016 7728 39080 7792
rect 39096 7728 39160 7792
rect 39176 7728 39240 7792
rect 39256 7728 39320 7792
rect 39336 7728 39400 7792
rect 39416 7728 39480 7792
rect 39496 7728 39560 7792
rect 39576 7728 39640 7792
rect 39656 7728 39720 7792
rect 39736 7728 39800 7792
rect 39816 7728 39880 7792
rect 39896 7728 39960 7792
rect 39976 7728 40040 7792
rect 40056 7728 40120 7792
rect 40136 7728 40200 7792
rect 40216 7728 40280 7792
rect 40296 7728 40360 7792
rect 5008 7648 5072 7712
rect 5088 7648 5152 7712
rect 5168 7648 5232 7712
rect 5248 7648 5312 7712
rect 5328 7648 5392 7712
rect 5408 7648 5472 7712
rect 5488 7648 5552 7712
rect 5568 7648 5632 7712
rect 5648 7648 5712 7712
rect 5728 7648 5792 7712
rect 5808 7648 5872 7712
rect 5888 7648 5952 7712
rect 5968 7648 6032 7712
rect 6048 7648 6112 7712
rect 6128 7648 6192 7712
rect 6208 7648 6272 7712
rect 6288 7648 6352 7712
rect 6368 7648 6432 7712
rect 6448 7648 6512 7712
rect 6528 7648 6592 7712
rect 6608 7648 6672 7712
rect 6688 7648 6752 7712
rect 6768 7648 6832 7712
rect 6848 7648 6912 7712
rect 6928 7648 6992 7712
rect 7008 7648 7072 7712
rect 7088 7648 7152 7712
rect 7168 7648 7232 7712
rect 7248 7648 7312 7712
rect 7328 7648 7392 7712
rect 7408 7648 7472 7712
rect 7488 7648 7552 7712
rect 7568 7648 7632 7712
rect 7648 7648 7712 7712
rect 7728 7648 7792 7712
rect 7808 7648 7872 7712
rect 7888 7648 7952 7712
rect 7968 7648 8032 7712
rect 8048 7648 8112 7712
rect 8128 7648 8192 7712
rect 8208 7648 8272 7712
rect 8288 7648 8352 7712
rect 8368 7648 8432 7712
rect 8448 7648 8512 7712
rect 8528 7648 8592 7712
rect 8608 7648 8672 7712
rect 8688 7648 8752 7712
rect 8768 7648 8832 7712
rect 8848 7648 8912 7712
rect 8928 7648 8992 7712
rect 14112 7648 14176 7712
rect 14192 7648 14256 7712
rect 14272 7648 14336 7712
rect 14352 7648 14416 7712
rect 24112 7648 24176 7712
rect 24192 7648 24256 7712
rect 24272 7648 24336 7712
rect 24352 7648 24416 7712
rect 36376 7648 36440 7712
rect 36456 7648 36520 7712
rect 36536 7648 36600 7712
rect 36616 7648 36680 7712
rect 36696 7648 36760 7712
rect 36776 7648 36840 7712
rect 36856 7648 36920 7712
rect 36936 7648 37000 7712
rect 37016 7648 37080 7712
rect 37096 7648 37160 7712
rect 37176 7648 37240 7712
rect 37256 7648 37320 7712
rect 37336 7648 37400 7712
rect 37416 7648 37480 7712
rect 37496 7648 37560 7712
rect 37576 7648 37640 7712
rect 37656 7648 37720 7712
rect 37736 7648 37800 7712
rect 37816 7648 37880 7712
rect 37896 7648 37960 7712
rect 37976 7648 38040 7712
rect 38056 7648 38120 7712
rect 38136 7648 38200 7712
rect 38216 7648 38280 7712
rect 38296 7648 38360 7712
rect 38376 7648 38440 7712
rect 38456 7648 38520 7712
rect 38536 7648 38600 7712
rect 38616 7648 38680 7712
rect 38696 7648 38760 7712
rect 38776 7648 38840 7712
rect 38856 7648 38920 7712
rect 38936 7648 39000 7712
rect 39016 7648 39080 7712
rect 39096 7648 39160 7712
rect 39176 7648 39240 7712
rect 39256 7648 39320 7712
rect 39336 7648 39400 7712
rect 39416 7648 39480 7712
rect 39496 7648 39560 7712
rect 39576 7648 39640 7712
rect 39656 7648 39720 7712
rect 39736 7648 39800 7712
rect 39816 7648 39880 7712
rect 39896 7648 39960 7712
rect 39976 7648 40040 7712
rect 40056 7648 40120 7712
rect 40136 7648 40200 7712
rect 40216 7648 40280 7712
rect 40296 7648 40360 7712
rect 5008 7568 5072 7632
rect 5088 7568 5152 7632
rect 5168 7568 5232 7632
rect 5248 7568 5312 7632
rect 5328 7568 5392 7632
rect 5408 7568 5472 7632
rect 5488 7568 5552 7632
rect 5568 7568 5632 7632
rect 5648 7568 5712 7632
rect 5728 7568 5792 7632
rect 5808 7568 5872 7632
rect 5888 7568 5952 7632
rect 5968 7568 6032 7632
rect 6048 7568 6112 7632
rect 6128 7568 6192 7632
rect 6208 7568 6272 7632
rect 6288 7568 6352 7632
rect 6368 7568 6432 7632
rect 6448 7568 6512 7632
rect 6528 7568 6592 7632
rect 6608 7568 6672 7632
rect 6688 7568 6752 7632
rect 6768 7568 6832 7632
rect 6848 7568 6912 7632
rect 6928 7568 6992 7632
rect 7008 7568 7072 7632
rect 7088 7568 7152 7632
rect 7168 7568 7232 7632
rect 7248 7568 7312 7632
rect 7328 7568 7392 7632
rect 7408 7568 7472 7632
rect 7488 7568 7552 7632
rect 7568 7568 7632 7632
rect 7648 7568 7712 7632
rect 7728 7568 7792 7632
rect 7808 7568 7872 7632
rect 7888 7568 7952 7632
rect 7968 7568 8032 7632
rect 8048 7568 8112 7632
rect 8128 7568 8192 7632
rect 8208 7568 8272 7632
rect 8288 7568 8352 7632
rect 8368 7568 8432 7632
rect 8448 7568 8512 7632
rect 8528 7568 8592 7632
rect 8608 7568 8672 7632
rect 8688 7568 8752 7632
rect 8768 7568 8832 7632
rect 8848 7568 8912 7632
rect 8928 7568 8992 7632
rect 14112 7568 14176 7632
rect 14192 7568 14256 7632
rect 14272 7568 14336 7632
rect 14352 7568 14416 7632
rect 24112 7568 24176 7632
rect 24192 7568 24256 7632
rect 24272 7568 24336 7632
rect 24352 7568 24416 7632
rect 36376 7568 36440 7632
rect 36456 7568 36520 7632
rect 36536 7568 36600 7632
rect 36616 7568 36680 7632
rect 36696 7568 36760 7632
rect 36776 7568 36840 7632
rect 36856 7568 36920 7632
rect 36936 7568 37000 7632
rect 37016 7568 37080 7632
rect 37096 7568 37160 7632
rect 37176 7568 37240 7632
rect 37256 7568 37320 7632
rect 37336 7568 37400 7632
rect 37416 7568 37480 7632
rect 37496 7568 37560 7632
rect 37576 7568 37640 7632
rect 37656 7568 37720 7632
rect 37736 7568 37800 7632
rect 37816 7568 37880 7632
rect 37896 7568 37960 7632
rect 37976 7568 38040 7632
rect 38056 7568 38120 7632
rect 38136 7568 38200 7632
rect 38216 7568 38280 7632
rect 38296 7568 38360 7632
rect 38376 7568 38440 7632
rect 38456 7568 38520 7632
rect 38536 7568 38600 7632
rect 38616 7568 38680 7632
rect 38696 7568 38760 7632
rect 38776 7568 38840 7632
rect 38856 7568 38920 7632
rect 38936 7568 39000 7632
rect 39016 7568 39080 7632
rect 39096 7568 39160 7632
rect 39176 7568 39240 7632
rect 39256 7568 39320 7632
rect 39336 7568 39400 7632
rect 39416 7568 39480 7632
rect 39496 7568 39560 7632
rect 39576 7568 39640 7632
rect 39656 7568 39720 7632
rect 39736 7568 39800 7632
rect 39816 7568 39880 7632
rect 39896 7568 39960 7632
rect 39976 7568 40040 7632
rect 40056 7568 40120 7632
rect 40136 7568 40200 7632
rect 40216 7568 40280 7632
rect 40296 7568 40360 7632
rect 5008 7488 5072 7552
rect 5088 7488 5152 7552
rect 5168 7488 5232 7552
rect 5248 7488 5312 7552
rect 5328 7488 5392 7552
rect 5408 7488 5472 7552
rect 5488 7488 5552 7552
rect 5568 7488 5632 7552
rect 5648 7488 5712 7552
rect 5728 7488 5792 7552
rect 5808 7488 5872 7552
rect 5888 7488 5952 7552
rect 5968 7488 6032 7552
rect 6048 7488 6112 7552
rect 6128 7488 6192 7552
rect 6208 7488 6272 7552
rect 6288 7488 6352 7552
rect 6368 7488 6432 7552
rect 6448 7488 6512 7552
rect 6528 7488 6592 7552
rect 6608 7488 6672 7552
rect 6688 7488 6752 7552
rect 6768 7488 6832 7552
rect 6848 7488 6912 7552
rect 6928 7488 6992 7552
rect 7008 7488 7072 7552
rect 7088 7488 7152 7552
rect 7168 7488 7232 7552
rect 7248 7488 7312 7552
rect 7328 7488 7392 7552
rect 7408 7488 7472 7552
rect 7488 7488 7552 7552
rect 7568 7488 7632 7552
rect 7648 7488 7712 7552
rect 7728 7488 7792 7552
rect 7808 7488 7872 7552
rect 7888 7488 7952 7552
rect 7968 7488 8032 7552
rect 8048 7488 8112 7552
rect 8128 7488 8192 7552
rect 8208 7488 8272 7552
rect 8288 7488 8352 7552
rect 8368 7488 8432 7552
rect 8448 7488 8512 7552
rect 8528 7488 8592 7552
rect 8608 7488 8672 7552
rect 8688 7488 8752 7552
rect 8768 7488 8832 7552
rect 8848 7488 8912 7552
rect 8928 7488 8992 7552
rect 14112 7488 14176 7552
rect 14192 7488 14256 7552
rect 14272 7488 14336 7552
rect 14352 7488 14416 7552
rect 24112 7488 24176 7552
rect 24192 7488 24256 7552
rect 24272 7488 24336 7552
rect 24352 7488 24416 7552
rect 36376 7488 36440 7552
rect 36456 7488 36520 7552
rect 36536 7488 36600 7552
rect 36616 7488 36680 7552
rect 36696 7488 36760 7552
rect 36776 7488 36840 7552
rect 36856 7488 36920 7552
rect 36936 7488 37000 7552
rect 37016 7488 37080 7552
rect 37096 7488 37160 7552
rect 37176 7488 37240 7552
rect 37256 7488 37320 7552
rect 37336 7488 37400 7552
rect 37416 7488 37480 7552
rect 37496 7488 37560 7552
rect 37576 7488 37640 7552
rect 37656 7488 37720 7552
rect 37736 7488 37800 7552
rect 37816 7488 37880 7552
rect 37896 7488 37960 7552
rect 37976 7488 38040 7552
rect 38056 7488 38120 7552
rect 38136 7488 38200 7552
rect 38216 7488 38280 7552
rect 38296 7488 38360 7552
rect 38376 7488 38440 7552
rect 38456 7488 38520 7552
rect 38536 7488 38600 7552
rect 38616 7488 38680 7552
rect 38696 7488 38760 7552
rect 38776 7488 38840 7552
rect 38856 7488 38920 7552
rect 38936 7488 39000 7552
rect 39016 7488 39080 7552
rect 39096 7488 39160 7552
rect 39176 7488 39240 7552
rect 39256 7488 39320 7552
rect 39336 7488 39400 7552
rect 39416 7488 39480 7552
rect 39496 7488 39560 7552
rect 39576 7488 39640 7552
rect 39656 7488 39720 7552
rect 39736 7488 39800 7552
rect 39816 7488 39880 7552
rect 39896 7488 39960 7552
rect 39976 7488 40040 7552
rect 40056 7488 40120 7552
rect 40136 7488 40200 7552
rect 40216 7488 40280 7552
rect 40296 7488 40360 7552
rect 5008 7408 5072 7472
rect 5088 7408 5152 7472
rect 5168 7408 5232 7472
rect 5248 7408 5312 7472
rect 5328 7408 5392 7472
rect 5408 7408 5472 7472
rect 5488 7408 5552 7472
rect 5568 7408 5632 7472
rect 5648 7408 5712 7472
rect 5728 7408 5792 7472
rect 5808 7408 5872 7472
rect 5888 7408 5952 7472
rect 5968 7408 6032 7472
rect 6048 7408 6112 7472
rect 6128 7408 6192 7472
rect 6208 7408 6272 7472
rect 6288 7408 6352 7472
rect 6368 7408 6432 7472
rect 6448 7408 6512 7472
rect 6528 7408 6592 7472
rect 6608 7408 6672 7472
rect 6688 7408 6752 7472
rect 6768 7408 6832 7472
rect 6848 7408 6912 7472
rect 6928 7408 6992 7472
rect 7008 7408 7072 7472
rect 7088 7408 7152 7472
rect 7168 7408 7232 7472
rect 7248 7408 7312 7472
rect 7328 7408 7392 7472
rect 7408 7408 7472 7472
rect 7488 7408 7552 7472
rect 7568 7408 7632 7472
rect 7648 7408 7712 7472
rect 7728 7408 7792 7472
rect 7808 7408 7872 7472
rect 7888 7408 7952 7472
rect 7968 7408 8032 7472
rect 8048 7408 8112 7472
rect 8128 7408 8192 7472
rect 8208 7408 8272 7472
rect 8288 7408 8352 7472
rect 8368 7408 8432 7472
rect 8448 7408 8512 7472
rect 8528 7408 8592 7472
rect 8608 7408 8672 7472
rect 8688 7408 8752 7472
rect 8768 7408 8832 7472
rect 8848 7408 8912 7472
rect 8928 7408 8992 7472
rect 14112 7408 14176 7472
rect 14192 7408 14256 7472
rect 14272 7408 14336 7472
rect 14352 7408 14416 7472
rect 24112 7408 24176 7472
rect 24192 7408 24256 7472
rect 24272 7408 24336 7472
rect 24352 7408 24416 7472
rect 36376 7408 36440 7472
rect 36456 7408 36520 7472
rect 36536 7408 36600 7472
rect 36616 7408 36680 7472
rect 36696 7408 36760 7472
rect 36776 7408 36840 7472
rect 36856 7408 36920 7472
rect 36936 7408 37000 7472
rect 37016 7408 37080 7472
rect 37096 7408 37160 7472
rect 37176 7408 37240 7472
rect 37256 7408 37320 7472
rect 37336 7408 37400 7472
rect 37416 7408 37480 7472
rect 37496 7408 37560 7472
rect 37576 7408 37640 7472
rect 37656 7408 37720 7472
rect 37736 7408 37800 7472
rect 37816 7408 37880 7472
rect 37896 7408 37960 7472
rect 37976 7408 38040 7472
rect 38056 7408 38120 7472
rect 38136 7408 38200 7472
rect 38216 7408 38280 7472
rect 38296 7408 38360 7472
rect 38376 7408 38440 7472
rect 38456 7408 38520 7472
rect 38536 7408 38600 7472
rect 38616 7408 38680 7472
rect 38696 7408 38760 7472
rect 38776 7408 38840 7472
rect 38856 7408 38920 7472
rect 38936 7408 39000 7472
rect 39016 7408 39080 7472
rect 39096 7408 39160 7472
rect 39176 7408 39240 7472
rect 39256 7408 39320 7472
rect 39336 7408 39400 7472
rect 39416 7408 39480 7472
rect 39496 7408 39560 7472
rect 39576 7408 39640 7472
rect 39656 7408 39720 7472
rect 39736 7408 39800 7472
rect 39816 7408 39880 7472
rect 39896 7408 39960 7472
rect 39976 7408 40040 7472
rect 40056 7408 40120 7472
rect 40136 7408 40200 7472
rect 40216 7408 40280 7472
rect 40296 7408 40360 7472
rect 5008 7328 5072 7392
rect 5088 7328 5152 7392
rect 5168 7328 5232 7392
rect 5248 7328 5312 7392
rect 5328 7328 5392 7392
rect 5408 7328 5472 7392
rect 5488 7328 5552 7392
rect 5568 7328 5632 7392
rect 5648 7328 5712 7392
rect 5728 7328 5792 7392
rect 5808 7328 5872 7392
rect 5888 7328 5952 7392
rect 5968 7328 6032 7392
rect 6048 7328 6112 7392
rect 6128 7328 6192 7392
rect 6208 7328 6272 7392
rect 6288 7328 6352 7392
rect 6368 7328 6432 7392
rect 6448 7328 6512 7392
rect 6528 7328 6592 7392
rect 6608 7328 6672 7392
rect 6688 7328 6752 7392
rect 6768 7328 6832 7392
rect 6848 7328 6912 7392
rect 6928 7328 6992 7392
rect 7008 7328 7072 7392
rect 7088 7328 7152 7392
rect 7168 7328 7232 7392
rect 7248 7328 7312 7392
rect 7328 7328 7392 7392
rect 7408 7328 7472 7392
rect 7488 7328 7552 7392
rect 7568 7328 7632 7392
rect 7648 7328 7712 7392
rect 7728 7328 7792 7392
rect 7808 7328 7872 7392
rect 7888 7328 7952 7392
rect 7968 7328 8032 7392
rect 8048 7328 8112 7392
rect 8128 7328 8192 7392
rect 8208 7328 8272 7392
rect 8288 7328 8352 7392
rect 8368 7328 8432 7392
rect 8448 7328 8512 7392
rect 8528 7328 8592 7392
rect 8608 7328 8672 7392
rect 8688 7328 8752 7392
rect 8768 7328 8832 7392
rect 8848 7328 8912 7392
rect 8928 7328 8992 7392
rect 14112 7328 14176 7392
rect 14192 7328 14256 7392
rect 14272 7328 14336 7392
rect 14352 7328 14416 7392
rect 24112 7328 24176 7392
rect 24192 7328 24256 7392
rect 24272 7328 24336 7392
rect 24352 7328 24416 7392
rect 36376 7328 36440 7392
rect 36456 7328 36520 7392
rect 36536 7328 36600 7392
rect 36616 7328 36680 7392
rect 36696 7328 36760 7392
rect 36776 7328 36840 7392
rect 36856 7328 36920 7392
rect 36936 7328 37000 7392
rect 37016 7328 37080 7392
rect 37096 7328 37160 7392
rect 37176 7328 37240 7392
rect 37256 7328 37320 7392
rect 37336 7328 37400 7392
rect 37416 7328 37480 7392
rect 37496 7328 37560 7392
rect 37576 7328 37640 7392
rect 37656 7328 37720 7392
rect 37736 7328 37800 7392
rect 37816 7328 37880 7392
rect 37896 7328 37960 7392
rect 37976 7328 38040 7392
rect 38056 7328 38120 7392
rect 38136 7328 38200 7392
rect 38216 7328 38280 7392
rect 38296 7328 38360 7392
rect 38376 7328 38440 7392
rect 38456 7328 38520 7392
rect 38536 7328 38600 7392
rect 38616 7328 38680 7392
rect 38696 7328 38760 7392
rect 38776 7328 38840 7392
rect 38856 7328 38920 7392
rect 38936 7328 39000 7392
rect 39016 7328 39080 7392
rect 39096 7328 39160 7392
rect 39176 7328 39240 7392
rect 39256 7328 39320 7392
rect 39336 7328 39400 7392
rect 39416 7328 39480 7392
rect 39496 7328 39560 7392
rect 39576 7328 39640 7392
rect 39656 7328 39720 7392
rect 39736 7328 39800 7392
rect 39816 7328 39880 7392
rect 39896 7328 39960 7392
rect 39976 7328 40040 7392
rect 40056 7328 40120 7392
rect 40136 7328 40200 7392
rect 40216 7328 40280 7392
rect 40296 7328 40360 7392
rect 5008 7248 5072 7312
rect 5088 7248 5152 7312
rect 5168 7248 5232 7312
rect 5248 7248 5312 7312
rect 5328 7248 5392 7312
rect 5408 7248 5472 7312
rect 5488 7248 5552 7312
rect 5568 7248 5632 7312
rect 5648 7248 5712 7312
rect 5728 7248 5792 7312
rect 5808 7248 5872 7312
rect 5888 7248 5952 7312
rect 5968 7248 6032 7312
rect 6048 7248 6112 7312
rect 6128 7248 6192 7312
rect 6208 7248 6272 7312
rect 6288 7248 6352 7312
rect 6368 7248 6432 7312
rect 6448 7248 6512 7312
rect 6528 7248 6592 7312
rect 6608 7248 6672 7312
rect 6688 7248 6752 7312
rect 6768 7248 6832 7312
rect 6848 7248 6912 7312
rect 6928 7248 6992 7312
rect 7008 7248 7072 7312
rect 7088 7248 7152 7312
rect 7168 7248 7232 7312
rect 7248 7248 7312 7312
rect 7328 7248 7392 7312
rect 7408 7248 7472 7312
rect 7488 7248 7552 7312
rect 7568 7248 7632 7312
rect 7648 7248 7712 7312
rect 7728 7248 7792 7312
rect 7808 7248 7872 7312
rect 7888 7248 7952 7312
rect 7968 7248 8032 7312
rect 8048 7248 8112 7312
rect 8128 7248 8192 7312
rect 8208 7248 8272 7312
rect 8288 7248 8352 7312
rect 8368 7248 8432 7312
rect 8448 7248 8512 7312
rect 8528 7248 8592 7312
rect 8608 7248 8672 7312
rect 8688 7248 8752 7312
rect 8768 7248 8832 7312
rect 8848 7248 8912 7312
rect 8928 7248 8992 7312
rect 14112 7248 14176 7312
rect 14192 7248 14256 7312
rect 14272 7248 14336 7312
rect 14352 7248 14416 7312
rect 24112 7248 24176 7312
rect 24192 7248 24256 7312
rect 24272 7248 24336 7312
rect 24352 7248 24416 7312
rect 36376 7248 36440 7312
rect 36456 7248 36520 7312
rect 36536 7248 36600 7312
rect 36616 7248 36680 7312
rect 36696 7248 36760 7312
rect 36776 7248 36840 7312
rect 36856 7248 36920 7312
rect 36936 7248 37000 7312
rect 37016 7248 37080 7312
rect 37096 7248 37160 7312
rect 37176 7248 37240 7312
rect 37256 7248 37320 7312
rect 37336 7248 37400 7312
rect 37416 7248 37480 7312
rect 37496 7248 37560 7312
rect 37576 7248 37640 7312
rect 37656 7248 37720 7312
rect 37736 7248 37800 7312
rect 37816 7248 37880 7312
rect 37896 7248 37960 7312
rect 37976 7248 38040 7312
rect 38056 7248 38120 7312
rect 38136 7248 38200 7312
rect 38216 7248 38280 7312
rect 38296 7248 38360 7312
rect 38376 7248 38440 7312
rect 38456 7248 38520 7312
rect 38536 7248 38600 7312
rect 38616 7248 38680 7312
rect 38696 7248 38760 7312
rect 38776 7248 38840 7312
rect 38856 7248 38920 7312
rect 38936 7248 39000 7312
rect 39016 7248 39080 7312
rect 39096 7248 39160 7312
rect 39176 7248 39240 7312
rect 39256 7248 39320 7312
rect 39336 7248 39400 7312
rect 39416 7248 39480 7312
rect 39496 7248 39560 7312
rect 39576 7248 39640 7312
rect 39656 7248 39720 7312
rect 39736 7248 39800 7312
rect 39816 7248 39880 7312
rect 39896 7248 39960 7312
rect 39976 7248 40040 7312
rect 40056 7248 40120 7312
rect 40136 7248 40200 7312
rect 40216 7248 40280 7312
rect 40296 7248 40360 7312
rect 5008 7168 5072 7232
rect 5088 7168 5152 7232
rect 5168 7168 5232 7232
rect 5248 7168 5312 7232
rect 5328 7168 5392 7232
rect 5408 7168 5472 7232
rect 5488 7168 5552 7232
rect 5568 7168 5632 7232
rect 5648 7168 5712 7232
rect 5728 7168 5792 7232
rect 5808 7168 5872 7232
rect 5888 7168 5952 7232
rect 5968 7168 6032 7232
rect 6048 7168 6112 7232
rect 6128 7168 6192 7232
rect 6208 7168 6272 7232
rect 6288 7168 6352 7232
rect 6368 7168 6432 7232
rect 6448 7168 6512 7232
rect 6528 7168 6592 7232
rect 6608 7168 6672 7232
rect 6688 7168 6752 7232
rect 6768 7168 6832 7232
rect 6848 7168 6912 7232
rect 6928 7168 6992 7232
rect 7008 7168 7072 7232
rect 7088 7168 7152 7232
rect 7168 7168 7232 7232
rect 7248 7168 7312 7232
rect 7328 7168 7392 7232
rect 7408 7168 7472 7232
rect 7488 7168 7552 7232
rect 7568 7168 7632 7232
rect 7648 7168 7712 7232
rect 7728 7168 7792 7232
rect 7808 7168 7872 7232
rect 7888 7168 7952 7232
rect 7968 7168 8032 7232
rect 8048 7168 8112 7232
rect 8128 7168 8192 7232
rect 8208 7168 8272 7232
rect 8288 7168 8352 7232
rect 8368 7168 8432 7232
rect 8448 7168 8512 7232
rect 8528 7168 8592 7232
rect 8608 7168 8672 7232
rect 8688 7168 8752 7232
rect 8768 7168 8832 7232
rect 8848 7168 8912 7232
rect 8928 7168 8992 7232
rect 14112 7168 14176 7232
rect 14192 7168 14256 7232
rect 14272 7168 14336 7232
rect 14352 7168 14416 7232
rect 24112 7168 24176 7232
rect 24192 7168 24256 7232
rect 24272 7168 24336 7232
rect 24352 7168 24416 7232
rect 36376 7168 36440 7232
rect 36456 7168 36520 7232
rect 36536 7168 36600 7232
rect 36616 7168 36680 7232
rect 36696 7168 36760 7232
rect 36776 7168 36840 7232
rect 36856 7168 36920 7232
rect 36936 7168 37000 7232
rect 37016 7168 37080 7232
rect 37096 7168 37160 7232
rect 37176 7168 37240 7232
rect 37256 7168 37320 7232
rect 37336 7168 37400 7232
rect 37416 7168 37480 7232
rect 37496 7168 37560 7232
rect 37576 7168 37640 7232
rect 37656 7168 37720 7232
rect 37736 7168 37800 7232
rect 37816 7168 37880 7232
rect 37896 7168 37960 7232
rect 37976 7168 38040 7232
rect 38056 7168 38120 7232
rect 38136 7168 38200 7232
rect 38216 7168 38280 7232
rect 38296 7168 38360 7232
rect 38376 7168 38440 7232
rect 38456 7168 38520 7232
rect 38536 7168 38600 7232
rect 38616 7168 38680 7232
rect 38696 7168 38760 7232
rect 38776 7168 38840 7232
rect 38856 7168 38920 7232
rect 38936 7168 39000 7232
rect 39016 7168 39080 7232
rect 39096 7168 39160 7232
rect 39176 7168 39240 7232
rect 39256 7168 39320 7232
rect 39336 7168 39400 7232
rect 39416 7168 39480 7232
rect 39496 7168 39560 7232
rect 39576 7168 39640 7232
rect 39656 7168 39720 7232
rect 39736 7168 39800 7232
rect 39816 7168 39880 7232
rect 39896 7168 39960 7232
rect 39976 7168 40040 7232
rect 40056 7168 40120 7232
rect 40136 7168 40200 7232
rect 40216 7168 40280 7232
rect 40296 7168 40360 7232
rect 5008 7088 5072 7152
rect 5088 7088 5152 7152
rect 5168 7088 5232 7152
rect 5248 7088 5312 7152
rect 5328 7088 5392 7152
rect 5408 7088 5472 7152
rect 5488 7088 5552 7152
rect 5568 7088 5632 7152
rect 5648 7088 5712 7152
rect 5728 7088 5792 7152
rect 5808 7088 5872 7152
rect 5888 7088 5952 7152
rect 5968 7088 6032 7152
rect 6048 7088 6112 7152
rect 6128 7088 6192 7152
rect 6208 7088 6272 7152
rect 6288 7088 6352 7152
rect 6368 7088 6432 7152
rect 6448 7088 6512 7152
rect 6528 7088 6592 7152
rect 6608 7088 6672 7152
rect 6688 7088 6752 7152
rect 6768 7088 6832 7152
rect 6848 7088 6912 7152
rect 6928 7088 6992 7152
rect 7008 7088 7072 7152
rect 7088 7088 7152 7152
rect 7168 7088 7232 7152
rect 7248 7088 7312 7152
rect 7328 7088 7392 7152
rect 7408 7088 7472 7152
rect 7488 7088 7552 7152
rect 7568 7088 7632 7152
rect 7648 7088 7712 7152
rect 7728 7088 7792 7152
rect 7808 7088 7872 7152
rect 7888 7088 7952 7152
rect 7968 7088 8032 7152
rect 8048 7088 8112 7152
rect 8128 7088 8192 7152
rect 8208 7088 8272 7152
rect 8288 7088 8352 7152
rect 8368 7088 8432 7152
rect 8448 7088 8512 7152
rect 8528 7088 8592 7152
rect 8608 7088 8672 7152
rect 8688 7088 8752 7152
rect 8768 7088 8832 7152
rect 8848 7088 8912 7152
rect 8928 7088 8992 7152
rect 14112 7088 14176 7152
rect 14192 7088 14256 7152
rect 14272 7088 14336 7152
rect 14352 7088 14416 7152
rect 24112 7088 24176 7152
rect 24192 7088 24256 7152
rect 24272 7088 24336 7152
rect 24352 7088 24416 7152
rect 36376 7088 36440 7152
rect 36456 7088 36520 7152
rect 36536 7088 36600 7152
rect 36616 7088 36680 7152
rect 36696 7088 36760 7152
rect 36776 7088 36840 7152
rect 36856 7088 36920 7152
rect 36936 7088 37000 7152
rect 37016 7088 37080 7152
rect 37096 7088 37160 7152
rect 37176 7088 37240 7152
rect 37256 7088 37320 7152
rect 37336 7088 37400 7152
rect 37416 7088 37480 7152
rect 37496 7088 37560 7152
rect 37576 7088 37640 7152
rect 37656 7088 37720 7152
rect 37736 7088 37800 7152
rect 37816 7088 37880 7152
rect 37896 7088 37960 7152
rect 37976 7088 38040 7152
rect 38056 7088 38120 7152
rect 38136 7088 38200 7152
rect 38216 7088 38280 7152
rect 38296 7088 38360 7152
rect 38376 7088 38440 7152
rect 38456 7088 38520 7152
rect 38536 7088 38600 7152
rect 38616 7088 38680 7152
rect 38696 7088 38760 7152
rect 38776 7088 38840 7152
rect 38856 7088 38920 7152
rect 38936 7088 39000 7152
rect 39016 7088 39080 7152
rect 39096 7088 39160 7152
rect 39176 7088 39240 7152
rect 39256 7088 39320 7152
rect 39336 7088 39400 7152
rect 39416 7088 39480 7152
rect 39496 7088 39560 7152
rect 39576 7088 39640 7152
rect 39656 7088 39720 7152
rect 39736 7088 39800 7152
rect 39816 7088 39880 7152
rect 39896 7088 39960 7152
rect 39976 7088 40040 7152
rect 40056 7088 40120 7152
rect 40136 7088 40200 7152
rect 40216 7088 40280 7152
rect 40296 7088 40360 7152
rect 5008 7008 5072 7072
rect 5088 7008 5152 7072
rect 5168 7008 5232 7072
rect 5248 7008 5312 7072
rect 5328 7008 5392 7072
rect 5408 7008 5472 7072
rect 5488 7008 5552 7072
rect 5568 7008 5632 7072
rect 5648 7008 5712 7072
rect 5728 7008 5792 7072
rect 5808 7008 5872 7072
rect 5888 7008 5952 7072
rect 5968 7008 6032 7072
rect 6048 7008 6112 7072
rect 6128 7008 6192 7072
rect 6208 7008 6272 7072
rect 6288 7008 6352 7072
rect 6368 7008 6432 7072
rect 6448 7008 6512 7072
rect 6528 7008 6592 7072
rect 6608 7008 6672 7072
rect 6688 7008 6752 7072
rect 6768 7008 6832 7072
rect 6848 7008 6912 7072
rect 6928 7008 6992 7072
rect 7008 7008 7072 7072
rect 7088 7008 7152 7072
rect 7168 7008 7232 7072
rect 7248 7008 7312 7072
rect 7328 7008 7392 7072
rect 7408 7008 7472 7072
rect 7488 7008 7552 7072
rect 7568 7008 7632 7072
rect 7648 7008 7712 7072
rect 7728 7008 7792 7072
rect 7808 7008 7872 7072
rect 7888 7008 7952 7072
rect 7968 7008 8032 7072
rect 8048 7008 8112 7072
rect 8128 7008 8192 7072
rect 8208 7008 8272 7072
rect 8288 7008 8352 7072
rect 8368 7008 8432 7072
rect 8448 7008 8512 7072
rect 8528 7008 8592 7072
rect 8608 7008 8672 7072
rect 8688 7008 8752 7072
rect 8768 7008 8832 7072
rect 8848 7008 8912 7072
rect 8928 7008 8992 7072
rect 14112 7008 14176 7072
rect 14192 7008 14256 7072
rect 14272 7008 14336 7072
rect 14352 7008 14416 7072
rect 24112 7008 24176 7072
rect 24192 7008 24256 7072
rect 24272 7008 24336 7072
rect 24352 7008 24416 7072
rect 36376 7008 36440 7072
rect 36456 7008 36520 7072
rect 36536 7008 36600 7072
rect 36616 7008 36680 7072
rect 36696 7008 36760 7072
rect 36776 7008 36840 7072
rect 36856 7008 36920 7072
rect 36936 7008 37000 7072
rect 37016 7008 37080 7072
rect 37096 7008 37160 7072
rect 37176 7008 37240 7072
rect 37256 7008 37320 7072
rect 37336 7008 37400 7072
rect 37416 7008 37480 7072
rect 37496 7008 37560 7072
rect 37576 7008 37640 7072
rect 37656 7008 37720 7072
rect 37736 7008 37800 7072
rect 37816 7008 37880 7072
rect 37896 7008 37960 7072
rect 37976 7008 38040 7072
rect 38056 7008 38120 7072
rect 38136 7008 38200 7072
rect 38216 7008 38280 7072
rect 38296 7008 38360 7072
rect 38376 7008 38440 7072
rect 38456 7008 38520 7072
rect 38536 7008 38600 7072
rect 38616 7008 38680 7072
rect 38696 7008 38760 7072
rect 38776 7008 38840 7072
rect 38856 7008 38920 7072
rect 38936 7008 39000 7072
rect 39016 7008 39080 7072
rect 39096 7008 39160 7072
rect 39176 7008 39240 7072
rect 39256 7008 39320 7072
rect 39336 7008 39400 7072
rect 39416 7008 39480 7072
rect 39496 7008 39560 7072
rect 39576 7008 39640 7072
rect 39656 7008 39720 7072
rect 39736 7008 39800 7072
rect 39816 7008 39880 7072
rect 39896 7008 39960 7072
rect 39976 7008 40040 7072
rect 40056 7008 40120 7072
rect 40136 7008 40200 7072
rect 40216 7008 40280 7072
rect 40296 7008 40360 7072
rect 5008 6928 5072 6992
rect 5088 6928 5152 6992
rect 5168 6928 5232 6992
rect 5248 6928 5312 6992
rect 5328 6928 5392 6992
rect 5408 6928 5472 6992
rect 5488 6928 5552 6992
rect 5568 6928 5632 6992
rect 5648 6928 5712 6992
rect 5728 6928 5792 6992
rect 5808 6928 5872 6992
rect 5888 6928 5952 6992
rect 5968 6928 6032 6992
rect 6048 6928 6112 6992
rect 6128 6928 6192 6992
rect 6208 6928 6272 6992
rect 6288 6928 6352 6992
rect 6368 6928 6432 6992
rect 6448 6928 6512 6992
rect 6528 6928 6592 6992
rect 6608 6928 6672 6992
rect 6688 6928 6752 6992
rect 6768 6928 6832 6992
rect 6848 6928 6912 6992
rect 6928 6928 6992 6992
rect 7008 6928 7072 6992
rect 7088 6928 7152 6992
rect 7168 6928 7232 6992
rect 7248 6928 7312 6992
rect 7328 6928 7392 6992
rect 7408 6928 7472 6992
rect 7488 6928 7552 6992
rect 7568 6928 7632 6992
rect 7648 6928 7712 6992
rect 7728 6928 7792 6992
rect 7808 6928 7872 6992
rect 7888 6928 7952 6992
rect 7968 6928 8032 6992
rect 8048 6928 8112 6992
rect 8128 6928 8192 6992
rect 8208 6928 8272 6992
rect 8288 6928 8352 6992
rect 8368 6928 8432 6992
rect 8448 6928 8512 6992
rect 8528 6928 8592 6992
rect 8608 6928 8672 6992
rect 8688 6928 8752 6992
rect 8768 6928 8832 6992
rect 8848 6928 8912 6992
rect 8928 6928 8992 6992
rect 14112 6928 14176 6992
rect 14192 6928 14256 6992
rect 14272 6928 14336 6992
rect 14352 6928 14416 6992
rect 24112 6928 24176 6992
rect 24192 6928 24256 6992
rect 24272 6928 24336 6992
rect 24352 6928 24416 6992
rect 36376 6928 36440 6992
rect 36456 6928 36520 6992
rect 36536 6928 36600 6992
rect 36616 6928 36680 6992
rect 36696 6928 36760 6992
rect 36776 6928 36840 6992
rect 36856 6928 36920 6992
rect 36936 6928 37000 6992
rect 37016 6928 37080 6992
rect 37096 6928 37160 6992
rect 37176 6928 37240 6992
rect 37256 6928 37320 6992
rect 37336 6928 37400 6992
rect 37416 6928 37480 6992
rect 37496 6928 37560 6992
rect 37576 6928 37640 6992
rect 37656 6928 37720 6992
rect 37736 6928 37800 6992
rect 37816 6928 37880 6992
rect 37896 6928 37960 6992
rect 37976 6928 38040 6992
rect 38056 6928 38120 6992
rect 38136 6928 38200 6992
rect 38216 6928 38280 6992
rect 38296 6928 38360 6992
rect 38376 6928 38440 6992
rect 38456 6928 38520 6992
rect 38536 6928 38600 6992
rect 38616 6928 38680 6992
rect 38696 6928 38760 6992
rect 38776 6928 38840 6992
rect 38856 6928 38920 6992
rect 38936 6928 39000 6992
rect 39016 6928 39080 6992
rect 39096 6928 39160 6992
rect 39176 6928 39240 6992
rect 39256 6928 39320 6992
rect 39336 6928 39400 6992
rect 39416 6928 39480 6992
rect 39496 6928 39560 6992
rect 39576 6928 39640 6992
rect 39656 6928 39720 6992
rect 39736 6928 39800 6992
rect 39816 6928 39880 6992
rect 39896 6928 39960 6992
rect 39976 6928 40040 6992
rect 40056 6928 40120 6992
rect 40136 6928 40200 6992
rect 40216 6928 40280 6992
rect 40296 6928 40360 6992
rect 5008 6848 5072 6912
rect 5088 6848 5152 6912
rect 5168 6848 5232 6912
rect 5248 6848 5312 6912
rect 5328 6848 5392 6912
rect 5408 6848 5472 6912
rect 5488 6848 5552 6912
rect 5568 6848 5632 6912
rect 5648 6848 5712 6912
rect 5728 6848 5792 6912
rect 5808 6848 5872 6912
rect 5888 6848 5952 6912
rect 5968 6848 6032 6912
rect 6048 6848 6112 6912
rect 6128 6848 6192 6912
rect 6208 6848 6272 6912
rect 6288 6848 6352 6912
rect 6368 6848 6432 6912
rect 6448 6848 6512 6912
rect 6528 6848 6592 6912
rect 6608 6848 6672 6912
rect 6688 6848 6752 6912
rect 6768 6848 6832 6912
rect 6848 6848 6912 6912
rect 6928 6848 6992 6912
rect 7008 6848 7072 6912
rect 7088 6848 7152 6912
rect 7168 6848 7232 6912
rect 7248 6848 7312 6912
rect 7328 6848 7392 6912
rect 7408 6848 7472 6912
rect 7488 6848 7552 6912
rect 7568 6848 7632 6912
rect 7648 6848 7712 6912
rect 7728 6848 7792 6912
rect 7808 6848 7872 6912
rect 7888 6848 7952 6912
rect 7968 6848 8032 6912
rect 8048 6848 8112 6912
rect 8128 6848 8192 6912
rect 8208 6848 8272 6912
rect 8288 6848 8352 6912
rect 8368 6848 8432 6912
rect 8448 6848 8512 6912
rect 8528 6848 8592 6912
rect 8608 6848 8672 6912
rect 8688 6848 8752 6912
rect 8768 6848 8832 6912
rect 8848 6848 8912 6912
rect 8928 6848 8992 6912
rect 14112 6848 14176 6912
rect 14192 6848 14256 6912
rect 14272 6848 14336 6912
rect 14352 6848 14416 6912
rect 24112 6848 24176 6912
rect 24192 6848 24256 6912
rect 24272 6848 24336 6912
rect 24352 6848 24416 6912
rect 36376 6848 36440 6912
rect 36456 6848 36520 6912
rect 36536 6848 36600 6912
rect 36616 6848 36680 6912
rect 36696 6848 36760 6912
rect 36776 6848 36840 6912
rect 36856 6848 36920 6912
rect 36936 6848 37000 6912
rect 37016 6848 37080 6912
rect 37096 6848 37160 6912
rect 37176 6848 37240 6912
rect 37256 6848 37320 6912
rect 37336 6848 37400 6912
rect 37416 6848 37480 6912
rect 37496 6848 37560 6912
rect 37576 6848 37640 6912
rect 37656 6848 37720 6912
rect 37736 6848 37800 6912
rect 37816 6848 37880 6912
rect 37896 6848 37960 6912
rect 37976 6848 38040 6912
rect 38056 6848 38120 6912
rect 38136 6848 38200 6912
rect 38216 6848 38280 6912
rect 38296 6848 38360 6912
rect 38376 6848 38440 6912
rect 38456 6848 38520 6912
rect 38536 6848 38600 6912
rect 38616 6848 38680 6912
rect 38696 6848 38760 6912
rect 38776 6848 38840 6912
rect 38856 6848 38920 6912
rect 38936 6848 39000 6912
rect 39016 6848 39080 6912
rect 39096 6848 39160 6912
rect 39176 6848 39240 6912
rect 39256 6848 39320 6912
rect 39336 6848 39400 6912
rect 39416 6848 39480 6912
rect 39496 6848 39560 6912
rect 39576 6848 39640 6912
rect 39656 6848 39720 6912
rect 39736 6848 39800 6912
rect 39816 6848 39880 6912
rect 39896 6848 39960 6912
rect 39976 6848 40040 6912
rect 40056 6848 40120 6912
rect 40136 6848 40200 6912
rect 40216 6848 40280 6912
rect 40296 6848 40360 6912
rect 5008 6768 5072 6832
rect 5088 6768 5152 6832
rect 5168 6768 5232 6832
rect 5248 6768 5312 6832
rect 5328 6768 5392 6832
rect 5408 6768 5472 6832
rect 5488 6768 5552 6832
rect 5568 6768 5632 6832
rect 5648 6768 5712 6832
rect 5728 6768 5792 6832
rect 5808 6768 5872 6832
rect 5888 6768 5952 6832
rect 5968 6768 6032 6832
rect 6048 6768 6112 6832
rect 6128 6768 6192 6832
rect 6208 6768 6272 6832
rect 6288 6768 6352 6832
rect 6368 6768 6432 6832
rect 6448 6768 6512 6832
rect 6528 6768 6592 6832
rect 6608 6768 6672 6832
rect 6688 6768 6752 6832
rect 6768 6768 6832 6832
rect 6848 6768 6912 6832
rect 6928 6768 6992 6832
rect 7008 6768 7072 6832
rect 7088 6768 7152 6832
rect 7168 6768 7232 6832
rect 7248 6768 7312 6832
rect 7328 6768 7392 6832
rect 7408 6768 7472 6832
rect 7488 6768 7552 6832
rect 7568 6768 7632 6832
rect 7648 6768 7712 6832
rect 7728 6768 7792 6832
rect 7808 6768 7872 6832
rect 7888 6768 7952 6832
rect 7968 6768 8032 6832
rect 8048 6768 8112 6832
rect 8128 6768 8192 6832
rect 8208 6768 8272 6832
rect 8288 6768 8352 6832
rect 8368 6768 8432 6832
rect 8448 6768 8512 6832
rect 8528 6768 8592 6832
rect 8608 6768 8672 6832
rect 8688 6768 8752 6832
rect 8768 6768 8832 6832
rect 8848 6768 8912 6832
rect 8928 6768 8992 6832
rect 14112 6768 14176 6832
rect 14192 6768 14256 6832
rect 14272 6768 14336 6832
rect 14352 6768 14416 6832
rect 24112 6768 24176 6832
rect 24192 6768 24256 6832
rect 24272 6768 24336 6832
rect 24352 6768 24416 6832
rect 36376 6768 36440 6832
rect 36456 6768 36520 6832
rect 36536 6768 36600 6832
rect 36616 6768 36680 6832
rect 36696 6768 36760 6832
rect 36776 6768 36840 6832
rect 36856 6768 36920 6832
rect 36936 6768 37000 6832
rect 37016 6768 37080 6832
rect 37096 6768 37160 6832
rect 37176 6768 37240 6832
rect 37256 6768 37320 6832
rect 37336 6768 37400 6832
rect 37416 6768 37480 6832
rect 37496 6768 37560 6832
rect 37576 6768 37640 6832
rect 37656 6768 37720 6832
rect 37736 6768 37800 6832
rect 37816 6768 37880 6832
rect 37896 6768 37960 6832
rect 37976 6768 38040 6832
rect 38056 6768 38120 6832
rect 38136 6768 38200 6832
rect 38216 6768 38280 6832
rect 38296 6768 38360 6832
rect 38376 6768 38440 6832
rect 38456 6768 38520 6832
rect 38536 6768 38600 6832
rect 38616 6768 38680 6832
rect 38696 6768 38760 6832
rect 38776 6768 38840 6832
rect 38856 6768 38920 6832
rect 38936 6768 39000 6832
rect 39016 6768 39080 6832
rect 39096 6768 39160 6832
rect 39176 6768 39240 6832
rect 39256 6768 39320 6832
rect 39336 6768 39400 6832
rect 39416 6768 39480 6832
rect 39496 6768 39560 6832
rect 39576 6768 39640 6832
rect 39656 6768 39720 6832
rect 39736 6768 39800 6832
rect 39816 6768 39880 6832
rect 39896 6768 39960 6832
rect 39976 6768 40040 6832
rect 40056 6768 40120 6832
rect 40136 6768 40200 6832
rect 40216 6768 40280 6832
rect 40296 6768 40360 6832
rect 5008 6688 5072 6752
rect 5088 6688 5152 6752
rect 5168 6688 5232 6752
rect 5248 6688 5312 6752
rect 5328 6688 5392 6752
rect 5408 6688 5472 6752
rect 5488 6688 5552 6752
rect 5568 6688 5632 6752
rect 5648 6688 5712 6752
rect 5728 6688 5792 6752
rect 5808 6688 5872 6752
rect 5888 6688 5952 6752
rect 5968 6688 6032 6752
rect 6048 6688 6112 6752
rect 6128 6688 6192 6752
rect 6208 6688 6272 6752
rect 6288 6688 6352 6752
rect 6368 6688 6432 6752
rect 6448 6688 6512 6752
rect 6528 6688 6592 6752
rect 6608 6688 6672 6752
rect 6688 6688 6752 6752
rect 6768 6688 6832 6752
rect 6848 6688 6912 6752
rect 6928 6688 6992 6752
rect 7008 6688 7072 6752
rect 7088 6688 7152 6752
rect 7168 6688 7232 6752
rect 7248 6688 7312 6752
rect 7328 6688 7392 6752
rect 7408 6688 7472 6752
rect 7488 6688 7552 6752
rect 7568 6688 7632 6752
rect 7648 6688 7712 6752
rect 7728 6688 7792 6752
rect 7808 6688 7872 6752
rect 7888 6688 7952 6752
rect 7968 6688 8032 6752
rect 8048 6688 8112 6752
rect 8128 6688 8192 6752
rect 8208 6688 8272 6752
rect 8288 6688 8352 6752
rect 8368 6688 8432 6752
rect 8448 6688 8512 6752
rect 8528 6688 8592 6752
rect 8608 6688 8672 6752
rect 8688 6688 8752 6752
rect 8768 6688 8832 6752
rect 8848 6688 8912 6752
rect 8928 6688 8992 6752
rect 14112 6688 14176 6752
rect 14192 6688 14256 6752
rect 14272 6688 14336 6752
rect 14352 6688 14416 6752
rect 24112 6688 24176 6752
rect 24192 6688 24256 6752
rect 24272 6688 24336 6752
rect 24352 6688 24416 6752
rect 36376 6688 36440 6752
rect 36456 6688 36520 6752
rect 36536 6688 36600 6752
rect 36616 6688 36680 6752
rect 36696 6688 36760 6752
rect 36776 6688 36840 6752
rect 36856 6688 36920 6752
rect 36936 6688 37000 6752
rect 37016 6688 37080 6752
rect 37096 6688 37160 6752
rect 37176 6688 37240 6752
rect 37256 6688 37320 6752
rect 37336 6688 37400 6752
rect 37416 6688 37480 6752
rect 37496 6688 37560 6752
rect 37576 6688 37640 6752
rect 37656 6688 37720 6752
rect 37736 6688 37800 6752
rect 37816 6688 37880 6752
rect 37896 6688 37960 6752
rect 37976 6688 38040 6752
rect 38056 6688 38120 6752
rect 38136 6688 38200 6752
rect 38216 6688 38280 6752
rect 38296 6688 38360 6752
rect 38376 6688 38440 6752
rect 38456 6688 38520 6752
rect 38536 6688 38600 6752
rect 38616 6688 38680 6752
rect 38696 6688 38760 6752
rect 38776 6688 38840 6752
rect 38856 6688 38920 6752
rect 38936 6688 39000 6752
rect 39016 6688 39080 6752
rect 39096 6688 39160 6752
rect 39176 6688 39240 6752
rect 39256 6688 39320 6752
rect 39336 6688 39400 6752
rect 39416 6688 39480 6752
rect 39496 6688 39560 6752
rect 39576 6688 39640 6752
rect 39656 6688 39720 6752
rect 39736 6688 39800 6752
rect 39816 6688 39880 6752
rect 39896 6688 39960 6752
rect 39976 6688 40040 6752
rect 40056 6688 40120 6752
rect 40136 6688 40200 6752
rect 40216 6688 40280 6752
rect 40296 6688 40360 6752
rect 5008 6608 5072 6672
rect 5088 6608 5152 6672
rect 5168 6608 5232 6672
rect 5248 6608 5312 6672
rect 5328 6608 5392 6672
rect 5408 6608 5472 6672
rect 5488 6608 5552 6672
rect 5568 6608 5632 6672
rect 5648 6608 5712 6672
rect 5728 6608 5792 6672
rect 5808 6608 5872 6672
rect 5888 6608 5952 6672
rect 5968 6608 6032 6672
rect 6048 6608 6112 6672
rect 6128 6608 6192 6672
rect 6208 6608 6272 6672
rect 6288 6608 6352 6672
rect 6368 6608 6432 6672
rect 6448 6608 6512 6672
rect 6528 6608 6592 6672
rect 6608 6608 6672 6672
rect 6688 6608 6752 6672
rect 6768 6608 6832 6672
rect 6848 6608 6912 6672
rect 6928 6608 6992 6672
rect 7008 6608 7072 6672
rect 7088 6608 7152 6672
rect 7168 6608 7232 6672
rect 7248 6608 7312 6672
rect 7328 6608 7392 6672
rect 7408 6608 7472 6672
rect 7488 6608 7552 6672
rect 7568 6608 7632 6672
rect 7648 6608 7712 6672
rect 7728 6608 7792 6672
rect 7808 6608 7872 6672
rect 7888 6608 7952 6672
rect 7968 6608 8032 6672
rect 8048 6608 8112 6672
rect 8128 6608 8192 6672
rect 8208 6608 8272 6672
rect 8288 6608 8352 6672
rect 8368 6608 8432 6672
rect 8448 6608 8512 6672
rect 8528 6608 8592 6672
rect 8608 6608 8672 6672
rect 8688 6608 8752 6672
rect 8768 6608 8832 6672
rect 8848 6608 8912 6672
rect 8928 6608 8992 6672
rect 14112 6608 14176 6672
rect 14192 6608 14256 6672
rect 14272 6608 14336 6672
rect 14352 6608 14416 6672
rect 24112 6608 24176 6672
rect 24192 6608 24256 6672
rect 24272 6608 24336 6672
rect 24352 6608 24416 6672
rect 36376 6608 36440 6672
rect 36456 6608 36520 6672
rect 36536 6608 36600 6672
rect 36616 6608 36680 6672
rect 36696 6608 36760 6672
rect 36776 6608 36840 6672
rect 36856 6608 36920 6672
rect 36936 6608 37000 6672
rect 37016 6608 37080 6672
rect 37096 6608 37160 6672
rect 37176 6608 37240 6672
rect 37256 6608 37320 6672
rect 37336 6608 37400 6672
rect 37416 6608 37480 6672
rect 37496 6608 37560 6672
rect 37576 6608 37640 6672
rect 37656 6608 37720 6672
rect 37736 6608 37800 6672
rect 37816 6608 37880 6672
rect 37896 6608 37960 6672
rect 37976 6608 38040 6672
rect 38056 6608 38120 6672
rect 38136 6608 38200 6672
rect 38216 6608 38280 6672
rect 38296 6608 38360 6672
rect 38376 6608 38440 6672
rect 38456 6608 38520 6672
rect 38536 6608 38600 6672
rect 38616 6608 38680 6672
rect 38696 6608 38760 6672
rect 38776 6608 38840 6672
rect 38856 6608 38920 6672
rect 38936 6608 39000 6672
rect 39016 6608 39080 6672
rect 39096 6608 39160 6672
rect 39176 6608 39240 6672
rect 39256 6608 39320 6672
rect 39336 6608 39400 6672
rect 39416 6608 39480 6672
rect 39496 6608 39560 6672
rect 39576 6608 39640 6672
rect 39656 6608 39720 6672
rect 39736 6608 39800 6672
rect 39816 6608 39880 6672
rect 39896 6608 39960 6672
rect 39976 6608 40040 6672
rect 40056 6608 40120 6672
rect 40136 6608 40200 6672
rect 40216 6608 40280 6672
rect 40296 6608 40360 6672
rect 5008 6528 5072 6592
rect 5088 6528 5152 6592
rect 5168 6528 5232 6592
rect 5248 6528 5312 6592
rect 5328 6528 5392 6592
rect 5408 6528 5472 6592
rect 5488 6528 5552 6592
rect 5568 6528 5632 6592
rect 5648 6528 5712 6592
rect 5728 6528 5792 6592
rect 5808 6528 5872 6592
rect 5888 6528 5952 6592
rect 5968 6528 6032 6592
rect 6048 6528 6112 6592
rect 6128 6528 6192 6592
rect 6208 6528 6272 6592
rect 6288 6528 6352 6592
rect 6368 6528 6432 6592
rect 6448 6528 6512 6592
rect 6528 6528 6592 6592
rect 6608 6528 6672 6592
rect 6688 6528 6752 6592
rect 6768 6528 6832 6592
rect 6848 6528 6912 6592
rect 6928 6528 6992 6592
rect 7008 6528 7072 6592
rect 7088 6528 7152 6592
rect 7168 6528 7232 6592
rect 7248 6528 7312 6592
rect 7328 6528 7392 6592
rect 7408 6528 7472 6592
rect 7488 6528 7552 6592
rect 7568 6528 7632 6592
rect 7648 6528 7712 6592
rect 7728 6528 7792 6592
rect 7808 6528 7872 6592
rect 7888 6528 7952 6592
rect 7968 6528 8032 6592
rect 8048 6528 8112 6592
rect 8128 6528 8192 6592
rect 8208 6528 8272 6592
rect 8288 6528 8352 6592
rect 8368 6528 8432 6592
rect 8448 6528 8512 6592
rect 8528 6528 8592 6592
rect 8608 6528 8672 6592
rect 8688 6528 8752 6592
rect 8768 6528 8832 6592
rect 8848 6528 8912 6592
rect 8928 6528 8992 6592
rect 14112 6528 14176 6592
rect 14192 6528 14256 6592
rect 14272 6528 14336 6592
rect 14352 6528 14416 6592
rect 24112 6528 24176 6592
rect 24192 6528 24256 6592
rect 24272 6528 24336 6592
rect 24352 6528 24416 6592
rect 36376 6528 36440 6592
rect 36456 6528 36520 6592
rect 36536 6528 36600 6592
rect 36616 6528 36680 6592
rect 36696 6528 36760 6592
rect 36776 6528 36840 6592
rect 36856 6528 36920 6592
rect 36936 6528 37000 6592
rect 37016 6528 37080 6592
rect 37096 6528 37160 6592
rect 37176 6528 37240 6592
rect 37256 6528 37320 6592
rect 37336 6528 37400 6592
rect 37416 6528 37480 6592
rect 37496 6528 37560 6592
rect 37576 6528 37640 6592
rect 37656 6528 37720 6592
rect 37736 6528 37800 6592
rect 37816 6528 37880 6592
rect 37896 6528 37960 6592
rect 37976 6528 38040 6592
rect 38056 6528 38120 6592
rect 38136 6528 38200 6592
rect 38216 6528 38280 6592
rect 38296 6528 38360 6592
rect 38376 6528 38440 6592
rect 38456 6528 38520 6592
rect 38536 6528 38600 6592
rect 38616 6528 38680 6592
rect 38696 6528 38760 6592
rect 38776 6528 38840 6592
rect 38856 6528 38920 6592
rect 38936 6528 39000 6592
rect 39016 6528 39080 6592
rect 39096 6528 39160 6592
rect 39176 6528 39240 6592
rect 39256 6528 39320 6592
rect 39336 6528 39400 6592
rect 39416 6528 39480 6592
rect 39496 6528 39560 6592
rect 39576 6528 39640 6592
rect 39656 6528 39720 6592
rect 39736 6528 39800 6592
rect 39816 6528 39880 6592
rect 39896 6528 39960 6592
rect 39976 6528 40040 6592
rect 40056 6528 40120 6592
rect 40136 6528 40200 6592
rect 40216 6528 40280 6592
rect 40296 6528 40360 6592
rect 5008 6448 5072 6512
rect 5088 6448 5152 6512
rect 5168 6448 5232 6512
rect 5248 6448 5312 6512
rect 5328 6448 5392 6512
rect 5408 6448 5472 6512
rect 5488 6448 5552 6512
rect 5568 6448 5632 6512
rect 5648 6448 5712 6512
rect 5728 6448 5792 6512
rect 5808 6448 5872 6512
rect 5888 6448 5952 6512
rect 5968 6448 6032 6512
rect 6048 6448 6112 6512
rect 6128 6448 6192 6512
rect 6208 6448 6272 6512
rect 6288 6448 6352 6512
rect 6368 6448 6432 6512
rect 6448 6448 6512 6512
rect 6528 6448 6592 6512
rect 6608 6448 6672 6512
rect 6688 6448 6752 6512
rect 6768 6448 6832 6512
rect 6848 6448 6912 6512
rect 6928 6448 6992 6512
rect 7008 6448 7072 6512
rect 7088 6448 7152 6512
rect 7168 6448 7232 6512
rect 7248 6448 7312 6512
rect 7328 6448 7392 6512
rect 7408 6448 7472 6512
rect 7488 6448 7552 6512
rect 7568 6448 7632 6512
rect 7648 6448 7712 6512
rect 7728 6448 7792 6512
rect 7808 6448 7872 6512
rect 7888 6448 7952 6512
rect 7968 6448 8032 6512
rect 8048 6448 8112 6512
rect 8128 6448 8192 6512
rect 8208 6448 8272 6512
rect 8288 6448 8352 6512
rect 8368 6448 8432 6512
rect 8448 6448 8512 6512
rect 8528 6448 8592 6512
rect 8608 6448 8672 6512
rect 8688 6448 8752 6512
rect 8768 6448 8832 6512
rect 8848 6448 8912 6512
rect 8928 6448 8992 6512
rect 14112 6448 14176 6512
rect 14192 6448 14256 6512
rect 14272 6448 14336 6512
rect 14352 6448 14416 6512
rect 24112 6448 24176 6512
rect 24192 6448 24256 6512
rect 24272 6448 24336 6512
rect 24352 6448 24416 6512
rect 36376 6448 36440 6512
rect 36456 6448 36520 6512
rect 36536 6448 36600 6512
rect 36616 6448 36680 6512
rect 36696 6448 36760 6512
rect 36776 6448 36840 6512
rect 36856 6448 36920 6512
rect 36936 6448 37000 6512
rect 37016 6448 37080 6512
rect 37096 6448 37160 6512
rect 37176 6448 37240 6512
rect 37256 6448 37320 6512
rect 37336 6448 37400 6512
rect 37416 6448 37480 6512
rect 37496 6448 37560 6512
rect 37576 6448 37640 6512
rect 37656 6448 37720 6512
rect 37736 6448 37800 6512
rect 37816 6448 37880 6512
rect 37896 6448 37960 6512
rect 37976 6448 38040 6512
rect 38056 6448 38120 6512
rect 38136 6448 38200 6512
rect 38216 6448 38280 6512
rect 38296 6448 38360 6512
rect 38376 6448 38440 6512
rect 38456 6448 38520 6512
rect 38536 6448 38600 6512
rect 38616 6448 38680 6512
rect 38696 6448 38760 6512
rect 38776 6448 38840 6512
rect 38856 6448 38920 6512
rect 38936 6448 39000 6512
rect 39016 6448 39080 6512
rect 39096 6448 39160 6512
rect 39176 6448 39240 6512
rect 39256 6448 39320 6512
rect 39336 6448 39400 6512
rect 39416 6448 39480 6512
rect 39496 6448 39560 6512
rect 39576 6448 39640 6512
rect 39656 6448 39720 6512
rect 39736 6448 39800 6512
rect 39816 6448 39880 6512
rect 39896 6448 39960 6512
rect 39976 6448 40040 6512
rect 40056 6448 40120 6512
rect 40136 6448 40200 6512
rect 40216 6448 40280 6512
rect 40296 6448 40360 6512
rect 5008 6368 5072 6432
rect 5088 6368 5152 6432
rect 5168 6368 5232 6432
rect 5248 6368 5312 6432
rect 5328 6368 5392 6432
rect 5408 6368 5472 6432
rect 5488 6368 5552 6432
rect 5568 6368 5632 6432
rect 5648 6368 5712 6432
rect 5728 6368 5792 6432
rect 5808 6368 5872 6432
rect 5888 6368 5952 6432
rect 5968 6368 6032 6432
rect 6048 6368 6112 6432
rect 6128 6368 6192 6432
rect 6208 6368 6272 6432
rect 6288 6368 6352 6432
rect 6368 6368 6432 6432
rect 6448 6368 6512 6432
rect 6528 6368 6592 6432
rect 6608 6368 6672 6432
rect 6688 6368 6752 6432
rect 6768 6368 6832 6432
rect 6848 6368 6912 6432
rect 6928 6368 6992 6432
rect 7008 6368 7072 6432
rect 7088 6368 7152 6432
rect 7168 6368 7232 6432
rect 7248 6368 7312 6432
rect 7328 6368 7392 6432
rect 7408 6368 7472 6432
rect 7488 6368 7552 6432
rect 7568 6368 7632 6432
rect 7648 6368 7712 6432
rect 7728 6368 7792 6432
rect 7808 6368 7872 6432
rect 7888 6368 7952 6432
rect 7968 6368 8032 6432
rect 8048 6368 8112 6432
rect 8128 6368 8192 6432
rect 8208 6368 8272 6432
rect 8288 6368 8352 6432
rect 8368 6368 8432 6432
rect 8448 6368 8512 6432
rect 8528 6368 8592 6432
rect 8608 6368 8672 6432
rect 8688 6368 8752 6432
rect 8768 6368 8832 6432
rect 8848 6368 8912 6432
rect 8928 6368 8992 6432
rect 14112 6368 14176 6432
rect 14192 6368 14256 6432
rect 14272 6368 14336 6432
rect 14352 6368 14416 6432
rect 24112 6368 24176 6432
rect 24192 6368 24256 6432
rect 24272 6368 24336 6432
rect 24352 6368 24416 6432
rect 36376 6368 36440 6432
rect 36456 6368 36520 6432
rect 36536 6368 36600 6432
rect 36616 6368 36680 6432
rect 36696 6368 36760 6432
rect 36776 6368 36840 6432
rect 36856 6368 36920 6432
rect 36936 6368 37000 6432
rect 37016 6368 37080 6432
rect 37096 6368 37160 6432
rect 37176 6368 37240 6432
rect 37256 6368 37320 6432
rect 37336 6368 37400 6432
rect 37416 6368 37480 6432
rect 37496 6368 37560 6432
rect 37576 6368 37640 6432
rect 37656 6368 37720 6432
rect 37736 6368 37800 6432
rect 37816 6368 37880 6432
rect 37896 6368 37960 6432
rect 37976 6368 38040 6432
rect 38056 6368 38120 6432
rect 38136 6368 38200 6432
rect 38216 6368 38280 6432
rect 38296 6368 38360 6432
rect 38376 6368 38440 6432
rect 38456 6368 38520 6432
rect 38536 6368 38600 6432
rect 38616 6368 38680 6432
rect 38696 6368 38760 6432
rect 38776 6368 38840 6432
rect 38856 6368 38920 6432
rect 38936 6368 39000 6432
rect 39016 6368 39080 6432
rect 39096 6368 39160 6432
rect 39176 6368 39240 6432
rect 39256 6368 39320 6432
rect 39336 6368 39400 6432
rect 39416 6368 39480 6432
rect 39496 6368 39560 6432
rect 39576 6368 39640 6432
rect 39656 6368 39720 6432
rect 39736 6368 39800 6432
rect 39816 6368 39880 6432
rect 39896 6368 39960 6432
rect 39976 6368 40040 6432
rect 40056 6368 40120 6432
rect 40136 6368 40200 6432
rect 40216 6368 40280 6432
rect 40296 6368 40360 6432
rect 5008 6288 5072 6352
rect 5088 6288 5152 6352
rect 5168 6288 5232 6352
rect 5248 6288 5312 6352
rect 5328 6288 5392 6352
rect 5408 6288 5472 6352
rect 5488 6288 5552 6352
rect 5568 6288 5632 6352
rect 5648 6288 5712 6352
rect 5728 6288 5792 6352
rect 5808 6288 5872 6352
rect 5888 6288 5952 6352
rect 5968 6288 6032 6352
rect 6048 6288 6112 6352
rect 6128 6288 6192 6352
rect 6208 6288 6272 6352
rect 6288 6288 6352 6352
rect 6368 6288 6432 6352
rect 6448 6288 6512 6352
rect 6528 6288 6592 6352
rect 6608 6288 6672 6352
rect 6688 6288 6752 6352
rect 6768 6288 6832 6352
rect 6848 6288 6912 6352
rect 6928 6288 6992 6352
rect 7008 6288 7072 6352
rect 7088 6288 7152 6352
rect 7168 6288 7232 6352
rect 7248 6288 7312 6352
rect 7328 6288 7392 6352
rect 7408 6288 7472 6352
rect 7488 6288 7552 6352
rect 7568 6288 7632 6352
rect 7648 6288 7712 6352
rect 7728 6288 7792 6352
rect 7808 6288 7872 6352
rect 7888 6288 7952 6352
rect 7968 6288 8032 6352
rect 8048 6288 8112 6352
rect 8128 6288 8192 6352
rect 8208 6288 8272 6352
rect 8288 6288 8352 6352
rect 8368 6288 8432 6352
rect 8448 6288 8512 6352
rect 8528 6288 8592 6352
rect 8608 6288 8672 6352
rect 8688 6288 8752 6352
rect 8768 6288 8832 6352
rect 8848 6288 8912 6352
rect 8928 6288 8992 6352
rect 14112 6288 14176 6352
rect 14192 6288 14256 6352
rect 14272 6288 14336 6352
rect 14352 6288 14416 6352
rect 24112 6288 24176 6352
rect 24192 6288 24256 6352
rect 24272 6288 24336 6352
rect 24352 6288 24416 6352
rect 36376 6288 36440 6352
rect 36456 6288 36520 6352
rect 36536 6288 36600 6352
rect 36616 6288 36680 6352
rect 36696 6288 36760 6352
rect 36776 6288 36840 6352
rect 36856 6288 36920 6352
rect 36936 6288 37000 6352
rect 37016 6288 37080 6352
rect 37096 6288 37160 6352
rect 37176 6288 37240 6352
rect 37256 6288 37320 6352
rect 37336 6288 37400 6352
rect 37416 6288 37480 6352
rect 37496 6288 37560 6352
rect 37576 6288 37640 6352
rect 37656 6288 37720 6352
rect 37736 6288 37800 6352
rect 37816 6288 37880 6352
rect 37896 6288 37960 6352
rect 37976 6288 38040 6352
rect 38056 6288 38120 6352
rect 38136 6288 38200 6352
rect 38216 6288 38280 6352
rect 38296 6288 38360 6352
rect 38376 6288 38440 6352
rect 38456 6288 38520 6352
rect 38536 6288 38600 6352
rect 38616 6288 38680 6352
rect 38696 6288 38760 6352
rect 38776 6288 38840 6352
rect 38856 6288 38920 6352
rect 38936 6288 39000 6352
rect 39016 6288 39080 6352
rect 39096 6288 39160 6352
rect 39176 6288 39240 6352
rect 39256 6288 39320 6352
rect 39336 6288 39400 6352
rect 39416 6288 39480 6352
rect 39496 6288 39560 6352
rect 39576 6288 39640 6352
rect 39656 6288 39720 6352
rect 39736 6288 39800 6352
rect 39816 6288 39880 6352
rect 39896 6288 39960 6352
rect 39976 6288 40040 6352
rect 40056 6288 40120 6352
rect 40136 6288 40200 6352
rect 40216 6288 40280 6352
rect 40296 6288 40360 6352
rect 5008 6208 5072 6272
rect 5088 6208 5152 6272
rect 5168 6208 5232 6272
rect 5248 6208 5312 6272
rect 5328 6208 5392 6272
rect 5408 6208 5472 6272
rect 5488 6208 5552 6272
rect 5568 6208 5632 6272
rect 5648 6208 5712 6272
rect 5728 6208 5792 6272
rect 5808 6208 5872 6272
rect 5888 6208 5952 6272
rect 5968 6208 6032 6272
rect 6048 6208 6112 6272
rect 6128 6208 6192 6272
rect 6208 6208 6272 6272
rect 6288 6208 6352 6272
rect 6368 6208 6432 6272
rect 6448 6208 6512 6272
rect 6528 6208 6592 6272
rect 6608 6208 6672 6272
rect 6688 6208 6752 6272
rect 6768 6208 6832 6272
rect 6848 6208 6912 6272
rect 6928 6208 6992 6272
rect 7008 6208 7072 6272
rect 7088 6208 7152 6272
rect 7168 6208 7232 6272
rect 7248 6208 7312 6272
rect 7328 6208 7392 6272
rect 7408 6208 7472 6272
rect 7488 6208 7552 6272
rect 7568 6208 7632 6272
rect 7648 6208 7712 6272
rect 7728 6208 7792 6272
rect 7808 6208 7872 6272
rect 7888 6208 7952 6272
rect 7968 6208 8032 6272
rect 8048 6208 8112 6272
rect 8128 6208 8192 6272
rect 8208 6208 8272 6272
rect 8288 6208 8352 6272
rect 8368 6208 8432 6272
rect 8448 6208 8512 6272
rect 8528 6208 8592 6272
rect 8608 6208 8672 6272
rect 8688 6208 8752 6272
rect 8768 6208 8832 6272
rect 8848 6208 8912 6272
rect 8928 6208 8992 6272
rect 14112 6208 14176 6272
rect 14192 6208 14256 6272
rect 14272 6208 14336 6272
rect 14352 6208 14416 6272
rect 24112 6208 24176 6272
rect 24192 6208 24256 6272
rect 24272 6208 24336 6272
rect 24352 6208 24416 6272
rect 36376 6208 36440 6272
rect 36456 6208 36520 6272
rect 36536 6208 36600 6272
rect 36616 6208 36680 6272
rect 36696 6208 36760 6272
rect 36776 6208 36840 6272
rect 36856 6208 36920 6272
rect 36936 6208 37000 6272
rect 37016 6208 37080 6272
rect 37096 6208 37160 6272
rect 37176 6208 37240 6272
rect 37256 6208 37320 6272
rect 37336 6208 37400 6272
rect 37416 6208 37480 6272
rect 37496 6208 37560 6272
rect 37576 6208 37640 6272
rect 37656 6208 37720 6272
rect 37736 6208 37800 6272
rect 37816 6208 37880 6272
rect 37896 6208 37960 6272
rect 37976 6208 38040 6272
rect 38056 6208 38120 6272
rect 38136 6208 38200 6272
rect 38216 6208 38280 6272
rect 38296 6208 38360 6272
rect 38376 6208 38440 6272
rect 38456 6208 38520 6272
rect 38536 6208 38600 6272
rect 38616 6208 38680 6272
rect 38696 6208 38760 6272
rect 38776 6208 38840 6272
rect 38856 6208 38920 6272
rect 38936 6208 39000 6272
rect 39016 6208 39080 6272
rect 39096 6208 39160 6272
rect 39176 6208 39240 6272
rect 39256 6208 39320 6272
rect 39336 6208 39400 6272
rect 39416 6208 39480 6272
rect 39496 6208 39560 6272
rect 39576 6208 39640 6272
rect 39656 6208 39720 6272
rect 39736 6208 39800 6272
rect 39816 6208 39880 6272
rect 39896 6208 39960 6272
rect 39976 6208 40040 6272
rect 40056 6208 40120 6272
rect 40136 6208 40200 6272
rect 40216 6208 40280 6272
rect 40296 6208 40360 6272
rect 5008 6128 5072 6192
rect 5088 6128 5152 6192
rect 5168 6128 5232 6192
rect 5248 6128 5312 6192
rect 5328 6128 5392 6192
rect 5408 6128 5472 6192
rect 5488 6128 5552 6192
rect 5568 6128 5632 6192
rect 5648 6128 5712 6192
rect 5728 6128 5792 6192
rect 5808 6128 5872 6192
rect 5888 6128 5952 6192
rect 5968 6128 6032 6192
rect 6048 6128 6112 6192
rect 6128 6128 6192 6192
rect 6208 6128 6272 6192
rect 6288 6128 6352 6192
rect 6368 6128 6432 6192
rect 6448 6128 6512 6192
rect 6528 6128 6592 6192
rect 6608 6128 6672 6192
rect 6688 6128 6752 6192
rect 6768 6128 6832 6192
rect 6848 6128 6912 6192
rect 6928 6128 6992 6192
rect 7008 6128 7072 6192
rect 7088 6128 7152 6192
rect 7168 6128 7232 6192
rect 7248 6128 7312 6192
rect 7328 6128 7392 6192
rect 7408 6128 7472 6192
rect 7488 6128 7552 6192
rect 7568 6128 7632 6192
rect 7648 6128 7712 6192
rect 7728 6128 7792 6192
rect 7808 6128 7872 6192
rect 7888 6128 7952 6192
rect 7968 6128 8032 6192
rect 8048 6128 8112 6192
rect 8128 6128 8192 6192
rect 8208 6128 8272 6192
rect 8288 6128 8352 6192
rect 8368 6128 8432 6192
rect 8448 6128 8512 6192
rect 8528 6128 8592 6192
rect 8608 6128 8672 6192
rect 8688 6128 8752 6192
rect 8768 6128 8832 6192
rect 8848 6128 8912 6192
rect 8928 6128 8992 6192
rect 14112 6128 14176 6192
rect 14192 6128 14256 6192
rect 14272 6128 14336 6192
rect 14352 6128 14416 6192
rect 24112 6128 24176 6192
rect 24192 6128 24256 6192
rect 24272 6128 24336 6192
rect 24352 6128 24416 6192
rect 36376 6128 36440 6192
rect 36456 6128 36520 6192
rect 36536 6128 36600 6192
rect 36616 6128 36680 6192
rect 36696 6128 36760 6192
rect 36776 6128 36840 6192
rect 36856 6128 36920 6192
rect 36936 6128 37000 6192
rect 37016 6128 37080 6192
rect 37096 6128 37160 6192
rect 37176 6128 37240 6192
rect 37256 6128 37320 6192
rect 37336 6128 37400 6192
rect 37416 6128 37480 6192
rect 37496 6128 37560 6192
rect 37576 6128 37640 6192
rect 37656 6128 37720 6192
rect 37736 6128 37800 6192
rect 37816 6128 37880 6192
rect 37896 6128 37960 6192
rect 37976 6128 38040 6192
rect 38056 6128 38120 6192
rect 38136 6128 38200 6192
rect 38216 6128 38280 6192
rect 38296 6128 38360 6192
rect 38376 6128 38440 6192
rect 38456 6128 38520 6192
rect 38536 6128 38600 6192
rect 38616 6128 38680 6192
rect 38696 6128 38760 6192
rect 38776 6128 38840 6192
rect 38856 6128 38920 6192
rect 38936 6128 39000 6192
rect 39016 6128 39080 6192
rect 39096 6128 39160 6192
rect 39176 6128 39240 6192
rect 39256 6128 39320 6192
rect 39336 6128 39400 6192
rect 39416 6128 39480 6192
rect 39496 6128 39560 6192
rect 39576 6128 39640 6192
rect 39656 6128 39720 6192
rect 39736 6128 39800 6192
rect 39816 6128 39880 6192
rect 39896 6128 39960 6192
rect 39976 6128 40040 6192
rect 40056 6128 40120 6192
rect 40136 6128 40200 6192
rect 40216 6128 40280 6192
rect 40296 6128 40360 6192
rect 5008 6048 5072 6112
rect 5088 6048 5152 6112
rect 5168 6048 5232 6112
rect 5248 6048 5312 6112
rect 5328 6048 5392 6112
rect 5408 6048 5472 6112
rect 5488 6048 5552 6112
rect 5568 6048 5632 6112
rect 5648 6048 5712 6112
rect 5728 6048 5792 6112
rect 5808 6048 5872 6112
rect 5888 6048 5952 6112
rect 5968 6048 6032 6112
rect 6048 6048 6112 6112
rect 6128 6048 6192 6112
rect 6208 6048 6272 6112
rect 6288 6048 6352 6112
rect 6368 6048 6432 6112
rect 6448 6048 6512 6112
rect 6528 6048 6592 6112
rect 6608 6048 6672 6112
rect 6688 6048 6752 6112
rect 6768 6048 6832 6112
rect 6848 6048 6912 6112
rect 6928 6048 6992 6112
rect 7008 6048 7072 6112
rect 7088 6048 7152 6112
rect 7168 6048 7232 6112
rect 7248 6048 7312 6112
rect 7328 6048 7392 6112
rect 7408 6048 7472 6112
rect 7488 6048 7552 6112
rect 7568 6048 7632 6112
rect 7648 6048 7712 6112
rect 7728 6048 7792 6112
rect 7808 6048 7872 6112
rect 7888 6048 7952 6112
rect 7968 6048 8032 6112
rect 8048 6048 8112 6112
rect 8128 6048 8192 6112
rect 8208 6048 8272 6112
rect 8288 6048 8352 6112
rect 8368 6048 8432 6112
rect 8448 6048 8512 6112
rect 8528 6048 8592 6112
rect 8608 6048 8672 6112
rect 8688 6048 8752 6112
rect 8768 6048 8832 6112
rect 8848 6048 8912 6112
rect 8928 6048 8992 6112
rect 14112 6048 14176 6112
rect 14192 6048 14256 6112
rect 14272 6048 14336 6112
rect 14352 6048 14416 6112
rect 24112 6048 24176 6112
rect 24192 6048 24256 6112
rect 24272 6048 24336 6112
rect 24352 6048 24416 6112
rect 36376 6048 36440 6112
rect 36456 6048 36520 6112
rect 36536 6048 36600 6112
rect 36616 6048 36680 6112
rect 36696 6048 36760 6112
rect 36776 6048 36840 6112
rect 36856 6048 36920 6112
rect 36936 6048 37000 6112
rect 37016 6048 37080 6112
rect 37096 6048 37160 6112
rect 37176 6048 37240 6112
rect 37256 6048 37320 6112
rect 37336 6048 37400 6112
rect 37416 6048 37480 6112
rect 37496 6048 37560 6112
rect 37576 6048 37640 6112
rect 37656 6048 37720 6112
rect 37736 6048 37800 6112
rect 37816 6048 37880 6112
rect 37896 6048 37960 6112
rect 37976 6048 38040 6112
rect 38056 6048 38120 6112
rect 38136 6048 38200 6112
rect 38216 6048 38280 6112
rect 38296 6048 38360 6112
rect 38376 6048 38440 6112
rect 38456 6048 38520 6112
rect 38536 6048 38600 6112
rect 38616 6048 38680 6112
rect 38696 6048 38760 6112
rect 38776 6048 38840 6112
rect 38856 6048 38920 6112
rect 38936 6048 39000 6112
rect 39016 6048 39080 6112
rect 39096 6048 39160 6112
rect 39176 6048 39240 6112
rect 39256 6048 39320 6112
rect 39336 6048 39400 6112
rect 39416 6048 39480 6112
rect 39496 6048 39560 6112
rect 39576 6048 39640 6112
rect 39656 6048 39720 6112
rect 39736 6048 39800 6112
rect 39816 6048 39880 6112
rect 39896 6048 39960 6112
rect 39976 6048 40040 6112
rect 40056 6048 40120 6112
rect 40136 6048 40200 6112
rect 40216 6048 40280 6112
rect 40296 6048 40360 6112
rect 5008 5968 5072 6032
rect 5088 5968 5152 6032
rect 5168 5968 5232 6032
rect 5248 5968 5312 6032
rect 5328 5968 5392 6032
rect 5408 5968 5472 6032
rect 5488 5968 5552 6032
rect 5568 5968 5632 6032
rect 5648 5968 5712 6032
rect 5728 5968 5792 6032
rect 5808 5968 5872 6032
rect 5888 5968 5952 6032
rect 5968 5968 6032 6032
rect 6048 5968 6112 6032
rect 6128 5968 6192 6032
rect 6208 5968 6272 6032
rect 6288 5968 6352 6032
rect 6368 5968 6432 6032
rect 6448 5968 6512 6032
rect 6528 5968 6592 6032
rect 6608 5968 6672 6032
rect 6688 5968 6752 6032
rect 6768 5968 6832 6032
rect 6848 5968 6912 6032
rect 6928 5968 6992 6032
rect 7008 5968 7072 6032
rect 7088 5968 7152 6032
rect 7168 5968 7232 6032
rect 7248 5968 7312 6032
rect 7328 5968 7392 6032
rect 7408 5968 7472 6032
rect 7488 5968 7552 6032
rect 7568 5968 7632 6032
rect 7648 5968 7712 6032
rect 7728 5968 7792 6032
rect 7808 5968 7872 6032
rect 7888 5968 7952 6032
rect 7968 5968 8032 6032
rect 8048 5968 8112 6032
rect 8128 5968 8192 6032
rect 8208 5968 8272 6032
rect 8288 5968 8352 6032
rect 8368 5968 8432 6032
rect 8448 5968 8512 6032
rect 8528 5968 8592 6032
rect 8608 5968 8672 6032
rect 8688 5968 8752 6032
rect 8768 5968 8832 6032
rect 8848 5968 8912 6032
rect 8928 5968 8992 6032
rect 14112 5968 14176 6032
rect 14192 5968 14256 6032
rect 14272 5968 14336 6032
rect 14352 5968 14416 6032
rect 24112 5968 24176 6032
rect 24192 5968 24256 6032
rect 24272 5968 24336 6032
rect 24352 5968 24416 6032
rect 36376 5968 36440 6032
rect 36456 5968 36520 6032
rect 36536 5968 36600 6032
rect 36616 5968 36680 6032
rect 36696 5968 36760 6032
rect 36776 5968 36840 6032
rect 36856 5968 36920 6032
rect 36936 5968 37000 6032
rect 37016 5968 37080 6032
rect 37096 5968 37160 6032
rect 37176 5968 37240 6032
rect 37256 5968 37320 6032
rect 37336 5968 37400 6032
rect 37416 5968 37480 6032
rect 37496 5968 37560 6032
rect 37576 5968 37640 6032
rect 37656 5968 37720 6032
rect 37736 5968 37800 6032
rect 37816 5968 37880 6032
rect 37896 5968 37960 6032
rect 37976 5968 38040 6032
rect 38056 5968 38120 6032
rect 38136 5968 38200 6032
rect 38216 5968 38280 6032
rect 38296 5968 38360 6032
rect 38376 5968 38440 6032
rect 38456 5968 38520 6032
rect 38536 5968 38600 6032
rect 38616 5968 38680 6032
rect 38696 5968 38760 6032
rect 38776 5968 38840 6032
rect 38856 5968 38920 6032
rect 38936 5968 39000 6032
rect 39016 5968 39080 6032
rect 39096 5968 39160 6032
rect 39176 5968 39240 6032
rect 39256 5968 39320 6032
rect 39336 5968 39400 6032
rect 39416 5968 39480 6032
rect 39496 5968 39560 6032
rect 39576 5968 39640 6032
rect 39656 5968 39720 6032
rect 39736 5968 39800 6032
rect 39816 5968 39880 6032
rect 39896 5968 39960 6032
rect 39976 5968 40040 6032
rect 40056 5968 40120 6032
rect 40136 5968 40200 6032
rect 40216 5968 40280 6032
rect 40296 5968 40360 6032
rect 5008 5888 5072 5952
rect 5088 5888 5152 5952
rect 5168 5888 5232 5952
rect 5248 5888 5312 5952
rect 5328 5888 5392 5952
rect 5408 5888 5472 5952
rect 5488 5888 5552 5952
rect 5568 5888 5632 5952
rect 5648 5888 5712 5952
rect 5728 5888 5792 5952
rect 5808 5888 5872 5952
rect 5888 5888 5952 5952
rect 5968 5888 6032 5952
rect 6048 5888 6112 5952
rect 6128 5888 6192 5952
rect 6208 5888 6272 5952
rect 6288 5888 6352 5952
rect 6368 5888 6432 5952
rect 6448 5888 6512 5952
rect 6528 5888 6592 5952
rect 6608 5888 6672 5952
rect 6688 5888 6752 5952
rect 6768 5888 6832 5952
rect 6848 5888 6912 5952
rect 6928 5888 6992 5952
rect 7008 5888 7072 5952
rect 7088 5888 7152 5952
rect 7168 5888 7232 5952
rect 7248 5888 7312 5952
rect 7328 5888 7392 5952
rect 7408 5888 7472 5952
rect 7488 5888 7552 5952
rect 7568 5888 7632 5952
rect 7648 5888 7712 5952
rect 7728 5888 7792 5952
rect 7808 5888 7872 5952
rect 7888 5888 7952 5952
rect 7968 5888 8032 5952
rect 8048 5888 8112 5952
rect 8128 5888 8192 5952
rect 8208 5888 8272 5952
rect 8288 5888 8352 5952
rect 8368 5888 8432 5952
rect 8448 5888 8512 5952
rect 8528 5888 8592 5952
rect 8608 5888 8672 5952
rect 8688 5888 8752 5952
rect 8768 5888 8832 5952
rect 8848 5888 8912 5952
rect 8928 5888 8992 5952
rect 14112 5888 14176 5952
rect 14192 5888 14256 5952
rect 14272 5888 14336 5952
rect 14352 5888 14416 5952
rect 24112 5888 24176 5952
rect 24192 5888 24256 5952
rect 24272 5888 24336 5952
rect 24352 5888 24416 5952
rect 36376 5888 36440 5952
rect 36456 5888 36520 5952
rect 36536 5888 36600 5952
rect 36616 5888 36680 5952
rect 36696 5888 36760 5952
rect 36776 5888 36840 5952
rect 36856 5888 36920 5952
rect 36936 5888 37000 5952
rect 37016 5888 37080 5952
rect 37096 5888 37160 5952
rect 37176 5888 37240 5952
rect 37256 5888 37320 5952
rect 37336 5888 37400 5952
rect 37416 5888 37480 5952
rect 37496 5888 37560 5952
rect 37576 5888 37640 5952
rect 37656 5888 37720 5952
rect 37736 5888 37800 5952
rect 37816 5888 37880 5952
rect 37896 5888 37960 5952
rect 37976 5888 38040 5952
rect 38056 5888 38120 5952
rect 38136 5888 38200 5952
rect 38216 5888 38280 5952
rect 38296 5888 38360 5952
rect 38376 5888 38440 5952
rect 38456 5888 38520 5952
rect 38536 5888 38600 5952
rect 38616 5888 38680 5952
rect 38696 5888 38760 5952
rect 38776 5888 38840 5952
rect 38856 5888 38920 5952
rect 38936 5888 39000 5952
rect 39016 5888 39080 5952
rect 39096 5888 39160 5952
rect 39176 5888 39240 5952
rect 39256 5888 39320 5952
rect 39336 5888 39400 5952
rect 39416 5888 39480 5952
rect 39496 5888 39560 5952
rect 39576 5888 39640 5952
rect 39656 5888 39720 5952
rect 39736 5888 39800 5952
rect 39816 5888 39880 5952
rect 39896 5888 39960 5952
rect 39976 5888 40040 5952
rect 40056 5888 40120 5952
rect 40136 5888 40200 5952
rect 40216 5888 40280 5952
rect 40296 5888 40360 5952
rect 5008 5808 5072 5872
rect 5088 5808 5152 5872
rect 5168 5808 5232 5872
rect 5248 5808 5312 5872
rect 5328 5808 5392 5872
rect 5408 5808 5472 5872
rect 5488 5808 5552 5872
rect 5568 5808 5632 5872
rect 5648 5808 5712 5872
rect 5728 5808 5792 5872
rect 5808 5808 5872 5872
rect 5888 5808 5952 5872
rect 5968 5808 6032 5872
rect 6048 5808 6112 5872
rect 6128 5808 6192 5872
rect 6208 5808 6272 5872
rect 6288 5808 6352 5872
rect 6368 5808 6432 5872
rect 6448 5808 6512 5872
rect 6528 5808 6592 5872
rect 6608 5808 6672 5872
rect 6688 5808 6752 5872
rect 6768 5808 6832 5872
rect 6848 5808 6912 5872
rect 6928 5808 6992 5872
rect 7008 5808 7072 5872
rect 7088 5808 7152 5872
rect 7168 5808 7232 5872
rect 7248 5808 7312 5872
rect 7328 5808 7392 5872
rect 7408 5808 7472 5872
rect 7488 5808 7552 5872
rect 7568 5808 7632 5872
rect 7648 5808 7712 5872
rect 7728 5808 7792 5872
rect 7808 5808 7872 5872
rect 7888 5808 7952 5872
rect 7968 5808 8032 5872
rect 8048 5808 8112 5872
rect 8128 5808 8192 5872
rect 8208 5808 8272 5872
rect 8288 5808 8352 5872
rect 8368 5808 8432 5872
rect 8448 5808 8512 5872
rect 8528 5808 8592 5872
rect 8608 5808 8672 5872
rect 8688 5808 8752 5872
rect 8768 5808 8832 5872
rect 8848 5808 8912 5872
rect 8928 5808 8992 5872
rect 14112 5808 14176 5872
rect 14192 5808 14256 5872
rect 14272 5808 14336 5872
rect 14352 5808 14416 5872
rect 24112 5808 24176 5872
rect 24192 5808 24256 5872
rect 24272 5808 24336 5872
rect 24352 5808 24416 5872
rect 36376 5808 36440 5872
rect 36456 5808 36520 5872
rect 36536 5808 36600 5872
rect 36616 5808 36680 5872
rect 36696 5808 36760 5872
rect 36776 5808 36840 5872
rect 36856 5808 36920 5872
rect 36936 5808 37000 5872
rect 37016 5808 37080 5872
rect 37096 5808 37160 5872
rect 37176 5808 37240 5872
rect 37256 5808 37320 5872
rect 37336 5808 37400 5872
rect 37416 5808 37480 5872
rect 37496 5808 37560 5872
rect 37576 5808 37640 5872
rect 37656 5808 37720 5872
rect 37736 5808 37800 5872
rect 37816 5808 37880 5872
rect 37896 5808 37960 5872
rect 37976 5808 38040 5872
rect 38056 5808 38120 5872
rect 38136 5808 38200 5872
rect 38216 5808 38280 5872
rect 38296 5808 38360 5872
rect 38376 5808 38440 5872
rect 38456 5808 38520 5872
rect 38536 5808 38600 5872
rect 38616 5808 38680 5872
rect 38696 5808 38760 5872
rect 38776 5808 38840 5872
rect 38856 5808 38920 5872
rect 38936 5808 39000 5872
rect 39016 5808 39080 5872
rect 39096 5808 39160 5872
rect 39176 5808 39240 5872
rect 39256 5808 39320 5872
rect 39336 5808 39400 5872
rect 39416 5808 39480 5872
rect 39496 5808 39560 5872
rect 39576 5808 39640 5872
rect 39656 5808 39720 5872
rect 39736 5808 39800 5872
rect 39816 5808 39880 5872
rect 39896 5808 39960 5872
rect 39976 5808 40040 5872
rect 40056 5808 40120 5872
rect 40136 5808 40200 5872
rect 40216 5808 40280 5872
rect 40296 5808 40360 5872
rect 5008 5728 5072 5792
rect 5088 5728 5152 5792
rect 5168 5728 5232 5792
rect 5248 5728 5312 5792
rect 5328 5728 5392 5792
rect 5408 5728 5472 5792
rect 5488 5728 5552 5792
rect 5568 5728 5632 5792
rect 5648 5728 5712 5792
rect 5728 5728 5792 5792
rect 5808 5728 5872 5792
rect 5888 5728 5952 5792
rect 5968 5728 6032 5792
rect 6048 5728 6112 5792
rect 6128 5728 6192 5792
rect 6208 5728 6272 5792
rect 6288 5728 6352 5792
rect 6368 5728 6432 5792
rect 6448 5728 6512 5792
rect 6528 5728 6592 5792
rect 6608 5728 6672 5792
rect 6688 5728 6752 5792
rect 6768 5728 6832 5792
rect 6848 5728 6912 5792
rect 6928 5728 6992 5792
rect 7008 5728 7072 5792
rect 7088 5728 7152 5792
rect 7168 5728 7232 5792
rect 7248 5728 7312 5792
rect 7328 5728 7392 5792
rect 7408 5728 7472 5792
rect 7488 5728 7552 5792
rect 7568 5728 7632 5792
rect 7648 5728 7712 5792
rect 7728 5728 7792 5792
rect 7808 5728 7872 5792
rect 7888 5728 7952 5792
rect 7968 5728 8032 5792
rect 8048 5728 8112 5792
rect 8128 5728 8192 5792
rect 8208 5728 8272 5792
rect 8288 5728 8352 5792
rect 8368 5728 8432 5792
rect 8448 5728 8512 5792
rect 8528 5728 8592 5792
rect 8608 5728 8672 5792
rect 8688 5728 8752 5792
rect 8768 5728 8832 5792
rect 8848 5728 8912 5792
rect 8928 5728 8992 5792
rect 14112 5728 14176 5792
rect 14192 5728 14256 5792
rect 14272 5728 14336 5792
rect 14352 5728 14416 5792
rect 24112 5728 24176 5792
rect 24192 5728 24256 5792
rect 24272 5728 24336 5792
rect 24352 5728 24416 5792
rect 36376 5728 36440 5792
rect 36456 5728 36520 5792
rect 36536 5728 36600 5792
rect 36616 5728 36680 5792
rect 36696 5728 36760 5792
rect 36776 5728 36840 5792
rect 36856 5728 36920 5792
rect 36936 5728 37000 5792
rect 37016 5728 37080 5792
rect 37096 5728 37160 5792
rect 37176 5728 37240 5792
rect 37256 5728 37320 5792
rect 37336 5728 37400 5792
rect 37416 5728 37480 5792
rect 37496 5728 37560 5792
rect 37576 5728 37640 5792
rect 37656 5728 37720 5792
rect 37736 5728 37800 5792
rect 37816 5728 37880 5792
rect 37896 5728 37960 5792
rect 37976 5728 38040 5792
rect 38056 5728 38120 5792
rect 38136 5728 38200 5792
rect 38216 5728 38280 5792
rect 38296 5728 38360 5792
rect 38376 5728 38440 5792
rect 38456 5728 38520 5792
rect 38536 5728 38600 5792
rect 38616 5728 38680 5792
rect 38696 5728 38760 5792
rect 38776 5728 38840 5792
rect 38856 5728 38920 5792
rect 38936 5728 39000 5792
rect 39016 5728 39080 5792
rect 39096 5728 39160 5792
rect 39176 5728 39240 5792
rect 39256 5728 39320 5792
rect 39336 5728 39400 5792
rect 39416 5728 39480 5792
rect 39496 5728 39560 5792
rect 39576 5728 39640 5792
rect 39656 5728 39720 5792
rect 39736 5728 39800 5792
rect 39816 5728 39880 5792
rect 39896 5728 39960 5792
rect 39976 5728 40040 5792
rect 40056 5728 40120 5792
rect 40136 5728 40200 5792
rect 40216 5728 40280 5792
rect 40296 5728 40360 5792
rect 5008 5648 5072 5712
rect 5088 5648 5152 5712
rect 5168 5648 5232 5712
rect 5248 5648 5312 5712
rect 5328 5648 5392 5712
rect 5408 5648 5472 5712
rect 5488 5648 5552 5712
rect 5568 5648 5632 5712
rect 5648 5648 5712 5712
rect 5728 5648 5792 5712
rect 5808 5648 5872 5712
rect 5888 5648 5952 5712
rect 5968 5648 6032 5712
rect 6048 5648 6112 5712
rect 6128 5648 6192 5712
rect 6208 5648 6272 5712
rect 6288 5648 6352 5712
rect 6368 5648 6432 5712
rect 6448 5648 6512 5712
rect 6528 5648 6592 5712
rect 6608 5648 6672 5712
rect 6688 5648 6752 5712
rect 6768 5648 6832 5712
rect 6848 5648 6912 5712
rect 6928 5648 6992 5712
rect 7008 5648 7072 5712
rect 7088 5648 7152 5712
rect 7168 5648 7232 5712
rect 7248 5648 7312 5712
rect 7328 5648 7392 5712
rect 7408 5648 7472 5712
rect 7488 5648 7552 5712
rect 7568 5648 7632 5712
rect 7648 5648 7712 5712
rect 7728 5648 7792 5712
rect 7808 5648 7872 5712
rect 7888 5648 7952 5712
rect 7968 5648 8032 5712
rect 8048 5648 8112 5712
rect 8128 5648 8192 5712
rect 8208 5648 8272 5712
rect 8288 5648 8352 5712
rect 8368 5648 8432 5712
rect 8448 5648 8512 5712
rect 8528 5648 8592 5712
rect 8608 5648 8672 5712
rect 8688 5648 8752 5712
rect 8768 5648 8832 5712
rect 8848 5648 8912 5712
rect 8928 5648 8992 5712
rect 14112 5648 14176 5712
rect 14192 5648 14256 5712
rect 14272 5648 14336 5712
rect 14352 5648 14416 5712
rect 24112 5648 24176 5712
rect 24192 5648 24256 5712
rect 24272 5648 24336 5712
rect 24352 5648 24416 5712
rect 36376 5648 36440 5712
rect 36456 5648 36520 5712
rect 36536 5648 36600 5712
rect 36616 5648 36680 5712
rect 36696 5648 36760 5712
rect 36776 5648 36840 5712
rect 36856 5648 36920 5712
rect 36936 5648 37000 5712
rect 37016 5648 37080 5712
rect 37096 5648 37160 5712
rect 37176 5648 37240 5712
rect 37256 5648 37320 5712
rect 37336 5648 37400 5712
rect 37416 5648 37480 5712
rect 37496 5648 37560 5712
rect 37576 5648 37640 5712
rect 37656 5648 37720 5712
rect 37736 5648 37800 5712
rect 37816 5648 37880 5712
rect 37896 5648 37960 5712
rect 37976 5648 38040 5712
rect 38056 5648 38120 5712
rect 38136 5648 38200 5712
rect 38216 5648 38280 5712
rect 38296 5648 38360 5712
rect 38376 5648 38440 5712
rect 38456 5648 38520 5712
rect 38536 5648 38600 5712
rect 38616 5648 38680 5712
rect 38696 5648 38760 5712
rect 38776 5648 38840 5712
rect 38856 5648 38920 5712
rect 38936 5648 39000 5712
rect 39016 5648 39080 5712
rect 39096 5648 39160 5712
rect 39176 5648 39240 5712
rect 39256 5648 39320 5712
rect 39336 5648 39400 5712
rect 39416 5648 39480 5712
rect 39496 5648 39560 5712
rect 39576 5648 39640 5712
rect 39656 5648 39720 5712
rect 39736 5648 39800 5712
rect 39816 5648 39880 5712
rect 39896 5648 39960 5712
rect 39976 5648 40040 5712
rect 40056 5648 40120 5712
rect 40136 5648 40200 5712
rect 40216 5648 40280 5712
rect 40296 5648 40360 5712
rect 5008 5568 5072 5632
rect 5088 5568 5152 5632
rect 5168 5568 5232 5632
rect 5248 5568 5312 5632
rect 5328 5568 5392 5632
rect 5408 5568 5472 5632
rect 5488 5568 5552 5632
rect 5568 5568 5632 5632
rect 5648 5568 5712 5632
rect 5728 5568 5792 5632
rect 5808 5568 5872 5632
rect 5888 5568 5952 5632
rect 5968 5568 6032 5632
rect 6048 5568 6112 5632
rect 6128 5568 6192 5632
rect 6208 5568 6272 5632
rect 6288 5568 6352 5632
rect 6368 5568 6432 5632
rect 6448 5568 6512 5632
rect 6528 5568 6592 5632
rect 6608 5568 6672 5632
rect 6688 5568 6752 5632
rect 6768 5568 6832 5632
rect 6848 5568 6912 5632
rect 6928 5568 6992 5632
rect 7008 5568 7072 5632
rect 7088 5568 7152 5632
rect 7168 5568 7232 5632
rect 7248 5568 7312 5632
rect 7328 5568 7392 5632
rect 7408 5568 7472 5632
rect 7488 5568 7552 5632
rect 7568 5568 7632 5632
rect 7648 5568 7712 5632
rect 7728 5568 7792 5632
rect 7808 5568 7872 5632
rect 7888 5568 7952 5632
rect 7968 5568 8032 5632
rect 8048 5568 8112 5632
rect 8128 5568 8192 5632
rect 8208 5568 8272 5632
rect 8288 5568 8352 5632
rect 8368 5568 8432 5632
rect 8448 5568 8512 5632
rect 8528 5568 8592 5632
rect 8608 5568 8672 5632
rect 8688 5568 8752 5632
rect 8768 5568 8832 5632
rect 8848 5568 8912 5632
rect 8928 5568 8992 5632
rect 14112 5568 14176 5632
rect 14192 5568 14256 5632
rect 14272 5568 14336 5632
rect 14352 5568 14416 5632
rect 24112 5568 24176 5632
rect 24192 5568 24256 5632
rect 24272 5568 24336 5632
rect 24352 5568 24416 5632
rect 36376 5568 36440 5632
rect 36456 5568 36520 5632
rect 36536 5568 36600 5632
rect 36616 5568 36680 5632
rect 36696 5568 36760 5632
rect 36776 5568 36840 5632
rect 36856 5568 36920 5632
rect 36936 5568 37000 5632
rect 37016 5568 37080 5632
rect 37096 5568 37160 5632
rect 37176 5568 37240 5632
rect 37256 5568 37320 5632
rect 37336 5568 37400 5632
rect 37416 5568 37480 5632
rect 37496 5568 37560 5632
rect 37576 5568 37640 5632
rect 37656 5568 37720 5632
rect 37736 5568 37800 5632
rect 37816 5568 37880 5632
rect 37896 5568 37960 5632
rect 37976 5568 38040 5632
rect 38056 5568 38120 5632
rect 38136 5568 38200 5632
rect 38216 5568 38280 5632
rect 38296 5568 38360 5632
rect 38376 5568 38440 5632
rect 38456 5568 38520 5632
rect 38536 5568 38600 5632
rect 38616 5568 38680 5632
rect 38696 5568 38760 5632
rect 38776 5568 38840 5632
rect 38856 5568 38920 5632
rect 38936 5568 39000 5632
rect 39016 5568 39080 5632
rect 39096 5568 39160 5632
rect 39176 5568 39240 5632
rect 39256 5568 39320 5632
rect 39336 5568 39400 5632
rect 39416 5568 39480 5632
rect 39496 5568 39560 5632
rect 39576 5568 39640 5632
rect 39656 5568 39720 5632
rect 39736 5568 39800 5632
rect 39816 5568 39880 5632
rect 39896 5568 39960 5632
rect 39976 5568 40040 5632
rect 40056 5568 40120 5632
rect 40136 5568 40200 5632
rect 40216 5568 40280 5632
rect 40296 5568 40360 5632
rect 5008 5488 5072 5552
rect 5088 5488 5152 5552
rect 5168 5488 5232 5552
rect 5248 5488 5312 5552
rect 5328 5488 5392 5552
rect 5408 5488 5472 5552
rect 5488 5488 5552 5552
rect 5568 5488 5632 5552
rect 5648 5488 5712 5552
rect 5728 5488 5792 5552
rect 5808 5488 5872 5552
rect 5888 5488 5952 5552
rect 5968 5488 6032 5552
rect 6048 5488 6112 5552
rect 6128 5488 6192 5552
rect 6208 5488 6272 5552
rect 6288 5488 6352 5552
rect 6368 5488 6432 5552
rect 6448 5488 6512 5552
rect 6528 5488 6592 5552
rect 6608 5488 6672 5552
rect 6688 5488 6752 5552
rect 6768 5488 6832 5552
rect 6848 5488 6912 5552
rect 6928 5488 6992 5552
rect 7008 5488 7072 5552
rect 7088 5488 7152 5552
rect 7168 5488 7232 5552
rect 7248 5488 7312 5552
rect 7328 5488 7392 5552
rect 7408 5488 7472 5552
rect 7488 5488 7552 5552
rect 7568 5488 7632 5552
rect 7648 5488 7712 5552
rect 7728 5488 7792 5552
rect 7808 5488 7872 5552
rect 7888 5488 7952 5552
rect 7968 5488 8032 5552
rect 8048 5488 8112 5552
rect 8128 5488 8192 5552
rect 8208 5488 8272 5552
rect 8288 5488 8352 5552
rect 8368 5488 8432 5552
rect 8448 5488 8512 5552
rect 8528 5488 8592 5552
rect 8608 5488 8672 5552
rect 8688 5488 8752 5552
rect 8768 5488 8832 5552
rect 8848 5488 8912 5552
rect 8928 5488 8992 5552
rect 14112 5488 14176 5552
rect 14192 5488 14256 5552
rect 14272 5488 14336 5552
rect 14352 5488 14416 5552
rect 24112 5488 24176 5552
rect 24192 5488 24256 5552
rect 24272 5488 24336 5552
rect 24352 5488 24416 5552
rect 36376 5488 36440 5552
rect 36456 5488 36520 5552
rect 36536 5488 36600 5552
rect 36616 5488 36680 5552
rect 36696 5488 36760 5552
rect 36776 5488 36840 5552
rect 36856 5488 36920 5552
rect 36936 5488 37000 5552
rect 37016 5488 37080 5552
rect 37096 5488 37160 5552
rect 37176 5488 37240 5552
rect 37256 5488 37320 5552
rect 37336 5488 37400 5552
rect 37416 5488 37480 5552
rect 37496 5488 37560 5552
rect 37576 5488 37640 5552
rect 37656 5488 37720 5552
rect 37736 5488 37800 5552
rect 37816 5488 37880 5552
rect 37896 5488 37960 5552
rect 37976 5488 38040 5552
rect 38056 5488 38120 5552
rect 38136 5488 38200 5552
rect 38216 5488 38280 5552
rect 38296 5488 38360 5552
rect 38376 5488 38440 5552
rect 38456 5488 38520 5552
rect 38536 5488 38600 5552
rect 38616 5488 38680 5552
rect 38696 5488 38760 5552
rect 38776 5488 38840 5552
rect 38856 5488 38920 5552
rect 38936 5488 39000 5552
rect 39016 5488 39080 5552
rect 39096 5488 39160 5552
rect 39176 5488 39240 5552
rect 39256 5488 39320 5552
rect 39336 5488 39400 5552
rect 39416 5488 39480 5552
rect 39496 5488 39560 5552
rect 39576 5488 39640 5552
rect 39656 5488 39720 5552
rect 39736 5488 39800 5552
rect 39816 5488 39880 5552
rect 39896 5488 39960 5552
rect 39976 5488 40040 5552
rect 40056 5488 40120 5552
rect 40136 5488 40200 5552
rect 40216 5488 40280 5552
rect 40296 5488 40360 5552
rect 5008 5408 5072 5472
rect 5088 5408 5152 5472
rect 5168 5408 5232 5472
rect 5248 5408 5312 5472
rect 5328 5408 5392 5472
rect 5408 5408 5472 5472
rect 5488 5408 5552 5472
rect 5568 5408 5632 5472
rect 5648 5408 5712 5472
rect 5728 5408 5792 5472
rect 5808 5408 5872 5472
rect 5888 5408 5952 5472
rect 5968 5408 6032 5472
rect 6048 5408 6112 5472
rect 6128 5408 6192 5472
rect 6208 5408 6272 5472
rect 6288 5408 6352 5472
rect 6368 5408 6432 5472
rect 6448 5408 6512 5472
rect 6528 5408 6592 5472
rect 6608 5408 6672 5472
rect 6688 5408 6752 5472
rect 6768 5408 6832 5472
rect 6848 5408 6912 5472
rect 6928 5408 6992 5472
rect 7008 5408 7072 5472
rect 7088 5408 7152 5472
rect 7168 5408 7232 5472
rect 7248 5408 7312 5472
rect 7328 5408 7392 5472
rect 7408 5408 7472 5472
rect 7488 5408 7552 5472
rect 7568 5408 7632 5472
rect 7648 5408 7712 5472
rect 7728 5408 7792 5472
rect 7808 5408 7872 5472
rect 7888 5408 7952 5472
rect 7968 5408 8032 5472
rect 8048 5408 8112 5472
rect 8128 5408 8192 5472
rect 8208 5408 8272 5472
rect 8288 5408 8352 5472
rect 8368 5408 8432 5472
rect 8448 5408 8512 5472
rect 8528 5408 8592 5472
rect 8608 5408 8672 5472
rect 8688 5408 8752 5472
rect 8768 5408 8832 5472
rect 8848 5408 8912 5472
rect 8928 5408 8992 5472
rect 14112 5408 14176 5472
rect 14192 5408 14256 5472
rect 14272 5408 14336 5472
rect 14352 5408 14416 5472
rect 24112 5408 24176 5472
rect 24192 5408 24256 5472
rect 24272 5408 24336 5472
rect 24352 5408 24416 5472
rect 36376 5408 36440 5472
rect 36456 5408 36520 5472
rect 36536 5408 36600 5472
rect 36616 5408 36680 5472
rect 36696 5408 36760 5472
rect 36776 5408 36840 5472
rect 36856 5408 36920 5472
rect 36936 5408 37000 5472
rect 37016 5408 37080 5472
rect 37096 5408 37160 5472
rect 37176 5408 37240 5472
rect 37256 5408 37320 5472
rect 37336 5408 37400 5472
rect 37416 5408 37480 5472
rect 37496 5408 37560 5472
rect 37576 5408 37640 5472
rect 37656 5408 37720 5472
rect 37736 5408 37800 5472
rect 37816 5408 37880 5472
rect 37896 5408 37960 5472
rect 37976 5408 38040 5472
rect 38056 5408 38120 5472
rect 38136 5408 38200 5472
rect 38216 5408 38280 5472
rect 38296 5408 38360 5472
rect 38376 5408 38440 5472
rect 38456 5408 38520 5472
rect 38536 5408 38600 5472
rect 38616 5408 38680 5472
rect 38696 5408 38760 5472
rect 38776 5408 38840 5472
rect 38856 5408 38920 5472
rect 38936 5408 39000 5472
rect 39016 5408 39080 5472
rect 39096 5408 39160 5472
rect 39176 5408 39240 5472
rect 39256 5408 39320 5472
rect 39336 5408 39400 5472
rect 39416 5408 39480 5472
rect 39496 5408 39560 5472
rect 39576 5408 39640 5472
rect 39656 5408 39720 5472
rect 39736 5408 39800 5472
rect 39816 5408 39880 5472
rect 39896 5408 39960 5472
rect 39976 5408 40040 5472
rect 40056 5408 40120 5472
rect 40136 5408 40200 5472
rect 40216 5408 40280 5472
rect 40296 5408 40360 5472
rect 5008 5328 5072 5392
rect 5088 5328 5152 5392
rect 5168 5328 5232 5392
rect 5248 5328 5312 5392
rect 5328 5328 5392 5392
rect 5408 5328 5472 5392
rect 5488 5328 5552 5392
rect 5568 5328 5632 5392
rect 5648 5328 5712 5392
rect 5728 5328 5792 5392
rect 5808 5328 5872 5392
rect 5888 5328 5952 5392
rect 5968 5328 6032 5392
rect 6048 5328 6112 5392
rect 6128 5328 6192 5392
rect 6208 5328 6272 5392
rect 6288 5328 6352 5392
rect 6368 5328 6432 5392
rect 6448 5328 6512 5392
rect 6528 5328 6592 5392
rect 6608 5328 6672 5392
rect 6688 5328 6752 5392
rect 6768 5328 6832 5392
rect 6848 5328 6912 5392
rect 6928 5328 6992 5392
rect 7008 5328 7072 5392
rect 7088 5328 7152 5392
rect 7168 5328 7232 5392
rect 7248 5328 7312 5392
rect 7328 5328 7392 5392
rect 7408 5328 7472 5392
rect 7488 5328 7552 5392
rect 7568 5328 7632 5392
rect 7648 5328 7712 5392
rect 7728 5328 7792 5392
rect 7808 5328 7872 5392
rect 7888 5328 7952 5392
rect 7968 5328 8032 5392
rect 8048 5328 8112 5392
rect 8128 5328 8192 5392
rect 8208 5328 8272 5392
rect 8288 5328 8352 5392
rect 8368 5328 8432 5392
rect 8448 5328 8512 5392
rect 8528 5328 8592 5392
rect 8608 5328 8672 5392
rect 8688 5328 8752 5392
rect 8768 5328 8832 5392
rect 8848 5328 8912 5392
rect 8928 5328 8992 5392
rect 14112 5328 14176 5392
rect 14192 5328 14256 5392
rect 14272 5328 14336 5392
rect 14352 5328 14416 5392
rect 24112 5328 24176 5392
rect 24192 5328 24256 5392
rect 24272 5328 24336 5392
rect 24352 5328 24416 5392
rect 36376 5328 36440 5392
rect 36456 5328 36520 5392
rect 36536 5328 36600 5392
rect 36616 5328 36680 5392
rect 36696 5328 36760 5392
rect 36776 5328 36840 5392
rect 36856 5328 36920 5392
rect 36936 5328 37000 5392
rect 37016 5328 37080 5392
rect 37096 5328 37160 5392
rect 37176 5328 37240 5392
rect 37256 5328 37320 5392
rect 37336 5328 37400 5392
rect 37416 5328 37480 5392
rect 37496 5328 37560 5392
rect 37576 5328 37640 5392
rect 37656 5328 37720 5392
rect 37736 5328 37800 5392
rect 37816 5328 37880 5392
rect 37896 5328 37960 5392
rect 37976 5328 38040 5392
rect 38056 5328 38120 5392
rect 38136 5328 38200 5392
rect 38216 5328 38280 5392
rect 38296 5328 38360 5392
rect 38376 5328 38440 5392
rect 38456 5328 38520 5392
rect 38536 5328 38600 5392
rect 38616 5328 38680 5392
rect 38696 5328 38760 5392
rect 38776 5328 38840 5392
rect 38856 5328 38920 5392
rect 38936 5328 39000 5392
rect 39016 5328 39080 5392
rect 39096 5328 39160 5392
rect 39176 5328 39240 5392
rect 39256 5328 39320 5392
rect 39336 5328 39400 5392
rect 39416 5328 39480 5392
rect 39496 5328 39560 5392
rect 39576 5328 39640 5392
rect 39656 5328 39720 5392
rect 39736 5328 39800 5392
rect 39816 5328 39880 5392
rect 39896 5328 39960 5392
rect 39976 5328 40040 5392
rect 40056 5328 40120 5392
rect 40136 5328 40200 5392
rect 40216 5328 40280 5392
rect 40296 5328 40360 5392
rect 5008 5248 5072 5312
rect 5088 5248 5152 5312
rect 5168 5248 5232 5312
rect 5248 5248 5312 5312
rect 5328 5248 5392 5312
rect 5408 5248 5472 5312
rect 5488 5248 5552 5312
rect 5568 5248 5632 5312
rect 5648 5248 5712 5312
rect 5728 5248 5792 5312
rect 5808 5248 5872 5312
rect 5888 5248 5952 5312
rect 5968 5248 6032 5312
rect 6048 5248 6112 5312
rect 6128 5248 6192 5312
rect 6208 5248 6272 5312
rect 6288 5248 6352 5312
rect 6368 5248 6432 5312
rect 6448 5248 6512 5312
rect 6528 5248 6592 5312
rect 6608 5248 6672 5312
rect 6688 5248 6752 5312
rect 6768 5248 6832 5312
rect 6848 5248 6912 5312
rect 6928 5248 6992 5312
rect 7008 5248 7072 5312
rect 7088 5248 7152 5312
rect 7168 5248 7232 5312
rect 7248 5248 7312 5312
rect 7328 5248 7392 5312
rect 7408 5248 7472 5312
rect 7488 5248 7552 5312
rect 7568 5248 7632 5312
rect 7648 5248 7712 5312
rect 7728 5248 7792 5312
rect 7808 5248 7872 5312
rect 7888 5248 7952 5312
rect 7968 5248 8032 5312
rect 8048 5248 8112 5312
rect 8128 5248 8192 5312
rect 8208 5248 8272 5312
rect 8288 5248 8352 5312
rect 8368 5248 8432 5312
rect 8448 5248 8512 5312
rect 8528 5248 8592 5312
rect 8608 5248 8672 5312
rect 8688 5248 8752 5312
rect 8768 5248 8832 5312
rect 8848 5248 8912 5312
rect 8928 5248 8992 5312
rect 14112 5248 14176 5312
rect 14192 5248 14256 5312
rect 14272 5248 14336 5312
rect 14352 5248 14416 5312
rect 24112 5248 24176 5312
rect 24192 5248 24256 5312
rect 24272 5248 24336 5312
rect 24352 5248 24416 5312
rect 36376 5248 36440 5312
rect 36456 5248 36520 5312
rect 36536 5248 36600 5312
rect 36616 5248 36680 5312
rect 36696 5248 36760 5312
rect 36776 5248 36840 5312
rect 36856 5248 36920 5312
rect 36936 5248 37000 5312
rect 37016 5248 37080 5312
rect 37096 5248 37160 5312
rect 37176 5248 37240 5312
rect 37256 5248 37320 5312
rect 37336 5248 37400 5312
rect 37416 5248 37480 5312
rect 37496 5248 37560 5312
rect 37576 5248 37640 5312
rect 37656 5248 37720 5312
rect 37736 5248 37800 5312
rect 37816 5248 37880 5312
rect 37896 5248 37960 5312
rect 37976 5248 38040 5312
rect 38056 5248 38120 5312
rect 38136 5248 38200 5312
rect 38216 5248 38280 5312
rect 38296 5248 38360 5312
rect 38376 5248 38440 5312
rect 38456 5248 38520 5312
rect 38536 5248 38600 5312
rect 38616 5248 38680 5312
rect 38696 5248 38760 5312
rect 38776 5248 38840 5312
rect 38856 5248 38920 5312
rect 38936 5248 39000 5312
rect 39016 5248 39080 5312
rect 39096 5248 39160 5312
rect 39176 5248 39240 5312
rect 39256 5248 39320 5312
rect 39336 5248 39400 5312
rect 39416 5248 39480 5312
rect 39496 5248 39560 5312
rect 39576 5248 39640 5312
rect 39656 5248 39720 5312
rect 39736 5248 39800 5312
rect 39816 5248 39880 5312
rect 39896 5248 39960 5312
rect 39976 5248 40040 5312
rect 40056 5248 40120 5312
rect 40136 5248 40200 5312
rect 40216 5248 40280 5312
rect 40296 5248 40360 5312
rect 5008 5168 5072 5232
rect 5088 5168 5152 5232
rect 5168 5168 5232 5232
rect 5248 5168 5312 5232
rect 5328 5168 5392 5232
rect 5408 5168 5472 5232
rect 5488 5168 5552 5232
rect 5568 5168 5632 5232
rect 5648 5168 5712 5232
rect 5728 5168 5792 5232
rect 5808 5168 5872 5232
rect 5888 5168 5952 5232
rect 5968 5168 6032 5232
rect 6048 5168 6112 5232
rect 6128 5168 6192 5232
rect 6208 5168 6272 5232
rect 6288 5168 6352 5232
rect 6368 5168 6432 5232
rect 6448 5168 6512 5232
rect 6528 5168 6592 5232
rect 6608 5168 6672 5232
rect 6688 5168 6752 5232
rect 6768 5168 6832 5232
rect 6848 5168 6912 5232
rect 6928 5168 6992 5232
rect 7008 5168 7072 5232
rect 7088 5168 7152 5232
rect 7168 5168 7232 5232
rect 7248 5168 7312 5232
rect 7328 5168 7392 5232
rect 7408 5168 7472 5232
rect 7488 5168 7552 5232
rect 7568 5168 7632 5232
rect 7648 5168 7712 5232
rect 7728 5168 7792 5232
rect 7808 5168 7872 5232
rect 7888 5168 7952 5232
rect 7968 5168 8032 5232
rect 8048 5168 8112 5232
rect 8128 5168 8192 5232
rect 8208 5168 8272 5232
rect 8288 5168 8352 5232
rect 8368 5168 8432 5232
rect 8448 5168 8512 5232
rect 8528 5168 8592 5232
rect 8608 5168 8672 5232
rect 8688 5168 8752 5232
rect 8768 5168 8832 5232
rect 8848 5168 8912 5232
rect 8928 5168 8992 5232
rect 14112 5168 14176 5232
rect 14192 5168 14256 5232
rect 14272 5168 14336 5232
rect 14352 5168 14416 5232
rect 24112 5168 24176 5232
rect 24192 5168 24256 5232
rect 24272 5168 24336 5232
rect 24352 5168 24416 5232
rect 36376 5168 36440 5232
rect 36456 5168 36520 5232
rect 36536 5168 36600 5232
rect 36616 5168 36680 5232
rect 36696 5168 36760 5232
rect 36776 5168 36840 5232
rect 36856 5168 36920 5232
rect 36936 5168 37000 5232
rect 37016 5168 37080 5232
rect 37096 5168 37160 5232
rect 37176 5168 37240 5232
rect 37256 5168 37320 5232
rect 37336 5168 37400 5232
rect 37416 5168 37480 5232
rect 37496 5168 37560 5232
rect 37576 5168 37640 5232
rect 37656 5168 37720 5232
rect 37736 5168 37800 5232
rect 37816 5168 37880 5232
rect 37896 5168 37960 5232
rect 37976 5168 38040 5232
rect 38056 5168 38120 5232
rect 38136 5168 38200 5232
rect 38216 5168 38280 5232
rect 38296 5168 38360 5232
rect 38376 5168 38440 5232
rect 38456 5168 38520 5232
rect 38536 5168 38600 5232
rect 38616 5168 38680 5232
rect 38696 5168 38760 5232
rect 38776 5168 38840 5232
rect 38856 5168 38920 5232
rect 38936 5168 39000 5232
rect 39016 5168 39080 5232
rect 39096 5168 39160 5232
rect 39176 5168 39240 5232
rect 39256 5168 39320 5232
rect 39336 5168 39400 5232
rect 39416 5168 39480 5232
rect 39496 5168 39560 5232
rect 39576 5168 39640 5232
rect 39656 5168 39720 5232
rect 39736 5168 39800 5232
rect 39816 5168 39880 5232
rect 39896 5168 39960 5232
rect 39976 5168 40040 5232
rect 40056 5168 40120 5232
rect 40136 5168 40200 5232
rect 40216 5168 40280 5232
rect 40296 5168 40360 5232
rect 5008 5088 5072 5152
rect 5088 5088 5152 5152
rect 5168 5088 5232 5152
rect 5248 5088 5312 5152
rect 5328 5088 5392 5152
rect 5408 5088 5472 5152
rect 5488 5088 5552 5152
rect 5568 5088 5632 5152
rect 5648 5088 5712 5152
rect 5728 5088 5792 5152
rect 5808 5088 5872 5152
rect 5888 5088 5952 5152
rect 5968 5088 6032 5152
rect 6048 5088 6112 5152
rect 6128 5088 6192 5152
rect 6208 5088 6272 5152
rect 6288 5088 6352 5152
rect 6368 5088 6432 5152
rect 6448 5088 6512 5152
rect 6528 5088 6592 5152
rect 6608 5088 6672 5152
rect 6688 5088 6752 5152
rect 6768 5088 6832 5152
rect 6848 5088 6912 5152
rect 6928 5088 6992 5152
rect 7008 5088 7072 5152
rect 7088 5088 7152 5152
rect 7168 5088 7232 5152
rect 7248 5088 7312 5152
rect 7328 5088 7392 5152
rect 7408 5088 7472 5152
rect 7488 5088 7552 5152
rect 7568 5088 7632 5152
rect 7648 5088 7712 5152
rect 7728 5088 7792 5152
rect 7808 5088 7872 5152
rect 7888 5088 7952 5152
rect 7968 5088 8032 5152
rect 8048 5088 8112 5152
rect 8128 5088 8192 5152
rect 8208 5088 8272 5152
rect 8288 5088 8352 5152
rect 8368 5088 8432 5152
rect 8448 5088 8512 5152
rect 8528 5088 8592 5152
rect 8608 5088 8672 5152
rect 8688 5088 8752 5152
rect 8768 5088 8832 5152
rect 8848 5088 8912 5152
rect 8928 5088 8992 5152
rect 14112 5088 14176 5152
rect 14192 5088 14256 5152
rect 14272 5088 14336 5152
rect 14352 5088 14416 5152
rect 24112 5088 24176 5152
rect 24192 5088 24256 5152
rect 24272 5088 24336 5152
rect 24352 5088 24416 5152
rect 36376 5088 36440 5152
rect 36456 5088 36520 5152
rect 36536 5088 36600 5152
rect 36616 5088 36680 5152
rect 36696 5088 36760 5152
rect 36776 5088 36840 5152
rect 36856 5088 36920 5152
rect 36936 5088 37000 5152
rect 37016 5088 37080 5152
rect 37096 5088 37160 5152
rect 37176 5088 37240 5152
rect 37256 5088 37320 5152
rect 37336 5088 37400 5152
rect 37416 5088 37480 5152
rect 37496 5088 37560 5152
rect 37576 5088 37640 5152
rect 37656 5088 37720 5152
rect 37736 5088 37800 5152
rect 37816 5088 37880 5152
rect 37896 5088 37960 5152
rect 37976 5088 38040 5152
rect 38056 5088 38120 5152
rect 38136 5088 38200 5152
rect 38216 5088 38280 5152
rect 38296 5088 38360 5152
rect 38376 5088 38440 5152
rect 38456 5088 38520 5152
rect 38536 5088 38600 5152
rect 38616 5088 38680 5152
rect 38696 5088 38760 5152
rect 38776 5088 38840 5152
rect 38856 5088 38920 5152
rect 38936 5088 39000 5152
rect 39016 5088 39080 5152
rect 39096 5088 39160 5152
rect 39176 5088 39240 5152
rect 39256 5088 39320 5152
rect 39336 5088 39400 5152
rect 39416 5088 39480 5152
rect 39496 5088 39560 5152
rect 39576 5088 39640 5152
rect 39656 5088 39720 5152
rect 39736 5088 39800 5152
rect 39816 5088 39880 5152
rect 39896 5088 39960 5152
rect 39976 5088 40040 5152
rect 40056 5088 40120 5152
rect 40136 5088 40200 5152
rect 40216 5088 40280 5152
rect 40296 5088 40360 5152
rect 5008 5008 5072 5072
rect 5088 5008 5152 5072
rect 5168 5008 5232 5072
rect 5248 5008 5312 5072
rect 5328 5008 5392 5072
rect 5408 5008 5472 5072
rect 5488 5008 5552 5072
rect 5568 5008 5632 5072
rect 5648 5008 5712 5072
rect 5728 5008 5792 5072
rect 5808 5008 5872 5072
rect 5888 5008 5952 5072
rect 5968 5008 6032 5072
rect 6048 5008 6112 5072
rect 6128 5008 6192 5072
rect 6208 5008 6272 5072
rect 6288 5008 6352 5072
rect 6368 5008 6432 5072
rect 6448 5008 6512 5072
rect 6528 5008 6592 5072
rect 6608 5008 6672 5072
rect 6688 5008 6752 5072
rect 6768 5008 6832 5072
rect 6848 5008 6912 5072
rect 6928 5008 6992 5072
rect 7008 5008 7072 5072
rect 7088 5008 7152 5072
rect 7168 5008 7232 5072
rect 7248 5008 7312 5072
rect 7328 5008 7392 5072
rect 7408 5008 7472 5072
rect 7488 5008 7552 5072
rect 7568 5008 7632 5072
rect 7648 5008 7712 5072
rect 7728 5008 7792 5072
rect 7808 5008 7872 5072
rect 7888 5008 7952 5072
rect 7968 5008 8032 5072
rect 8048 5008 8112 5072
rect 8128 5008 8192 5072
rect 8208 5008 8272 5072
rect 8288 5008 8352 5072
rect 8368 5008 8432 5072
rect 8448 5008 8512 5072
rect 8528 5008 8592 5072
rect 8608 5008 8672 5072
rect 8688 5008 8752 5072
rect 8768 5008 8832 5072
rect 8848 5008 8912 5072
rect 8928 5008 8992 5072
rect 14112 5008 14176 5072
rect 14192 5008 14256 5072
rect 14272 5008 14336 5072
rect 14352 5008 14416 5072
rect 24112 5008 24176 5072
rect 24192 5008 24256 5072
rect 24272 5008 24336 5072
rect 24352 5008 24416 5072
rect 36376 5008 36440 5072
rect 36456 5008 36520 5072
rect 36536 5008 36600 5072
rect 36616 5008 36680 5072
rect 36696 5008 36760 5072
rect 36776 5008 36840 5072
rect 36856 5008 36920 5072
rect 36936 5008 37000 5072
rect 37016 5008 37080 5072
rect 37096 5008 37160 5072
rect 37176 5008 37240 5072
rect 37256 5008 37320 5072
rect 37336 5008 37400 5072
rect 37416 5008 37480 5072
rect 37496 5008 37560 5072
rect 37576 5008 37640 5072
rect 37656 5008 37720 5072
rect 37736 5008 37800 5072
rect 37816 5008 37880 5072
rect 37896 5008 37960 5072
rect 37976 5008 38040 5072
rect 38056 5008 38120 5072
rect 38136 5008 38200 5072
rect 38216 5008 38280 5072
rect 38296 5008 38360 5072
rect 38376 5008 38440 5072
rect 38456 5008 38520 5072
rect 38536 5008 38600 5072
rect 38616 5008 38680 5072
rect 38696 5008 38760 5072
rect 38776 5008 38840 5072
rect 38856 5008 38920 5072
rect 38936 5008 39000 5072
rect 39016 5008 39080 5072
rect 39096 5008 39160 5072
rect 39176 5008 39240 5072
rect 39256 5008 39320 5072
rect 39336 5008 39400 5072
rect 39416 5008 39480 5072
rect 39496 5008 39560 5072
rect 39576 5008 39640 5072
rect 39656 5008 39720 5072
rect 39736 5008 39800 5072
rect 39816 5008 39880 5072
rect 39896 5008 39960 5072
rect 39976 5008 40040 5072
rect 40056 5008 40120 5072
rect 40136 5008 40200 5072
rect 40216 5008 40280 5072
rect 40296 5008 40360 5072
rect 8 3928 72 3992
rect 88 3928 152 3992
rect 168 3928 232 3992
rect 248 3928 312 3992
rect 328 3928 392 3992
rect 408 3928 472 3992
rect 488 3928 552 3992
rect 568 3928 632 3992
rect 648 3928 712 3992
rect 728 3928 792 3992
rect 808 3928 872 3992
rect 888 3928 952 3992
rect 968 3928 1032 3992
rect 1048 3928 1112 3992
rect 1128 3928 1192 3992
rect 1208 3928 1272 3992
rect 1288 3928 1352 3992
rect 1368 3928 1432 3992
rect 1448 3928 1512 3992
rect 1528 3928 1592 3992
rect 1608 3928 1672 3992
rect 1688 3928 1752 3992
rect 1768 3928 1832 3992
rect 1848 3928 1912 3992
rect 1928 3928 1992 3992
rect 2008 3928 2072 3992
rect 2088 3928 2152 3992
rect 2168 3928 2232 3992
rect 2248 3928 2312 3992
rect 2328 3928 2392 3992
rect 2408 3928 2472 3992
rect 2488 3928 2552 3992
rect 2568 3928 2632 3992
rect 2648 3928 2712 3992
rect 2728 3928 2792 3992
rect 2808 3928 2872 3992
rect 2888 3928 2952 3992
rect 2968 3928 3032 3992
rect 3048 3928 3112 3992
rect 3128 3928 3192 3992
rect 3208 3928 3272 3992
rect 3288 3928 3352 3992
rect 3368 3928 3432 3992
rect 3448 3928 3512 3992
rect 3528 3928 3592 3992
rect 3608 3928 3672 3992
rect 3688 3928 3752 3992
rect 3768 3928 3832 3992
rect 3848 3928 3912 3992
rect 3928 3928 3992 3992
rect 19112 3928 19176 3992
rect 19192 3928 19256 3992
rect 19272 3928 19336 3992
rect 19352 3928 19416 3992
rect 29112 3928 29176 3992
rect 29192 3928 29256 3992
rect 29272 3928 29336 3992
rect 29352 3928 29416 3992
rect 41376 3928 41440 3992
rect 41456 3928 41520 3992
rect 41536 3928 41600 3992
rect 41616 3928 41680 3992
rect 41696 3928 41760 3992
rect 41776 3928 41840 3992
rect 41856 3928 41920 3992
rect 41936 3928 42000 3992
rect 42016 3928 42080 3992
rect 42096 3928 42160 3992
rect 42176 3928 42240 3992
rect 42256 3928 42320 3992
rect 42336 3928 42400 3992
rect 42416 3928 42480 3992
rect 42496 3928 42560 3992
rect 42576 3928 42640 3992
rect 42656 3928 42720 3992
rect 42736 3928 42800 3992
rect 42816 3928 42880 3992
rect 42896 3928 42960 3992
rect 42976 3928 43040 3992
rect 43056 3928 43120 3992
rect 43136 3928 43200 3992
rect 43216 3928 43280 3992
rect 43296 3928 43360 3992
rect 43376 3928 43440 3992
rect 43456 3928 43520 3992
rect 43536 3928 43600 3992
rect 43616 3928 43680 3992
rect 43696 3928 43760 3992
rect 43776 3928 43840 3992
rect 43856 3928 43920 3992
rect 43936 3928 44000 3992
rect 44016 3928 44080 3992
rect 44096 3928 44160 3992
rect 44176 3928 44240 3992
rect 44256 3928 44320 3992
rect 44336 3928 44400 3992
rect 44416 3928 44480 3992
rect 44496 3928 44560 3992
rect 44576 3928 44640 3992
rect 44656 3928 44720 3992
rect 44736 3928 44800 3992
rect 44816 3928 44880 3992
rect 44896 3928 44960 3992
rect 44976 3928 45040 3992
rect 45056 3928 45120 3992
rect 45136 3928 45200 3992
rect 45216 3928 45280 3992
rect 45296 3928 45360 3992
rect 8 3848 72 3912
rect 88 3848 152 3912
rect 168 3848 232 3912
rect 248 3848 312 3912
rect 328 3848 392 3912
rect 408 3848 472 3912
rect 488 3848 552 3912
rect 568 3848 632 3912
rect 648 3848 712 3912
rect 728 3848 792 3912
rect 808 3848 872 3912
rect 888 3848 952 3912
rect 968 3848 1032 3912
rect 1048 3848 1112 3912
rect 1128 3848 1192 3912
rect 1208 3848 1272 3912
rect 1288 3848 1352 3912
rect 1368 3848 1432 3912
rect 1448 3848 1512 3912
rect 1528 3848 1592 3912
rect 1608 3848 1672 3912
rect 1688 3848 1752 3912
rect 1768 3848 1832 3912
rect 1848 3848 1912 3912
rect 1928 3848 1992 3912
rect 2008 3848 2072 3912
rect 2088 3848 2152 3912
rect 2168 3848 2232 3912
rect 2248 3848 2312 3912
rect 2328 3848 2392 3912
rect 2408 3848 2472 3912
rect 2488 3848 2552 3912
rect 2568 3848 2632 3912
rect 2648 3848 2712 3912
rect 2728 3848 2792 3912
rect 2808 3848 2872 3912
rect 2888 3848 2952 3912
rect 2968 3848 3032 3912
rect 3048 3848 3112 3912
rect 3128 3848 3192 3912
rect 3208 3848 3272 3912
rect 3288 3848 3352 3912
rect 3368 3848 3432 3912
rect 3448 3848 3512 3912
rect 3528 3848 3592 3912
rect 3608 3848 3672 3912
rect 3688 3848 3752 3912
rect 3768 3848 3832 3912
rect 3848 3848 3912 3912
rect 3928 3848 3992 3912
rect 19112 3848 19176 3912
rect 19192 3848 19256 3912
rect 19272 3848 19336 3912
rect 19352 3848 19416 3912
rect 29112 3848 29176 3912
rect 29192 3848 29256 3912
rect 29272 3848 29336 3912
rect 29352 3848 29416 3912
rect 41376 3848 41440 3912
rect 41456 3848 41520 3912
rect 41536 3848 41600 3912
rect 41616 3848 41680 3912
rect 41696 3848 41760 3912
rect 41776 3848 41840 3912
rect 41856 3848 41920 3912
rect 41936 3848 42000 3912
rect 42016 3848 42080 3912
rect 42096 3848 42160 3912
rect 42176 3848 42240 3912
rect 42256 3848 42320 3912
rect 42336 3848 42400 3912
rect 42416 3848 42480 3912
rect 42496 3848 42560 3912
rect 42576 3848 42640 3912
rect 42656 3848 42720 3912
rect 42736 3848 42800 3912
rect 42816 3848 42880 3912
rect 42896 3848 42960 3912
rect 42976 3848 43040 3912
rect 43056 3848 43120 3912
rect 43136 3848 43200 3912
rect 43216 3848 43280 3912
rect 43296 3848 43360 3912
rect 43376 3848 43440 3912
rect 43456 3848 43520 3912
rect 43536 3848 43600 3912
rect 43616 3848 43680 3912
rect 43696 3848 43760 3912
rect 43776 3848 43840 3912
rect 43856 3848 43920 3912
rect 43936 3848 44000 3912
rect 44016 3848 44080 3912
rect 44096 3848 44160 3912
rect 44176 3848 44240 3912
rect 44256 3848 44320 3912
rect 44336 3848 44400 3912
rect 44416 3848 44480 3912
rect 44496 3848 44560 3912
rect 44576 3848 44640 3912
rect 44656 3848 44720 3912
rect 44736 3848 44800 3912
rect 44816 3848 44880 3912
rect 44896 3848 44960 3912
rect 44976 3848 45040 3912
rect 45056 3848 45120 3912
rect 45136 3848 45200 3912
rect 45216 3848 45280 3912
rect 45296 3848 45360 3912
rect 8 3768 72 3832
rect 88 3768 152 3832
rect 168 3768 232 3832
rect 248 3768 312 3832
rect 328 3768 392 3832
rect 408 3768 472 3832
rect 488 3768 552 3832
rect 568 3768 632 3832
rect 648 3768 712 3832
rect 728 3768 792 3832
rect 808 3768 872 3832
rect 888 3768 952 3832
rect 968 3768 1032 3832
rect 1048 3768 1112 3832
rect 1128 3768 1192 3832
rect 1208 3768 1272 3832
rect 1288 3768 1352 3832
rect 1368 3768 1432 3832
rect 1448 3768 1512 3832
rect 1528 3768 1592 3832
rect 1608 3768 1672 3832
rect 1688 3768 1752 3832
rect 1768 3768 1832 3832
rect 1848 3768 1912 3832
rect 1928 3768 1992 3832
rect 2008 3768 2072 3832
rect 2088 3768 2152 3832
rect 2168 3768 2232 3832
rect 2248 3768 2312 3832
rect 2328 3768 2392 3832
rect 2408 3768 2472 3832
rect 2488 3768 2552 3832
rect 2568 3768 2632 3832
rect 2648 3768 2712 3832
rect 2728 3768 2792 3832
rect 2808 3768 2872 3832
rect 2888 3768 2952 3832
rect 2968 3768 3032 3832
rect 3048 3768 3112 3832
rect 3128 3768 3192 3832
rect 3208 3768 3272 3832
rect 3288 3768 3352 3832
rect 3368 3768 3432 3832
rect 3448 3768 3512 3832
rect 3528 3768 3592 3832
rect 3608 3768 3672 3832
rect 3688 3768 3752 3832
rect 3768 3768 3832 3832
rect 3848 3768 3912 3832
rect 3928 3768 3992 3832
rect 19112 3768 19176 3832
rect 19192 3768 19256 3832
rect 19272 3768 19336 3832
rect 19352 3768 19416 3832
rect 29112 3768 29176 3832
rect 29192 3768 29256 3832
rect 29272 3768 29336 3832
rect 29352 3768 29416 3832
rect 41376 3768 41440 3832
rect 41456 3768 41520 3832
rect 41536 3768 41600 3832
rect 41616 3768 41680 3832
rect 41696 3768 41760 3832
rect 41776 3768 41840 3832
rect 41856 3768 41920 3832
rect 41936 3768 42000 3832
rect 42016 3768 42080 3832
rect 42096 3768 42160 3832
rect 42176 3768 42240 3832
rect 42256 3768 42320 3832
rect 42336 3768 42400 3832
rect 42416 3768 42480 3832
rect 42496 3768 42560 3832
rect 42576 3768 42640 3832
rect 42656 3768 42720 3832
rect 42736 3768 42800 3832
rect 42816 3768 42880 3832
rect 42896 3768 42960 3832
rect 42976 3768 43040 3832
rect 43056 3768 43120 3832
rect 43136 3768 43200 3832
rect 43216 3768 43280 3832
rect 43296 3768 43360 3832
rect 43376 3768 43440 3832
rect 43456 3768 43520 3832
rect 43536 3768 43600 3832
rect 43616 3768 43680 3832
rect 43696 3768 43760 3832
rect 43776 3768 43840 3832
rect 43856 3768 43920 3832
rect 43936 3768 44000 3832
rect 44016 3768 44080 3832
rect 44096 3768 44160 3832
rect 44176 3768 44240 3832
rect 44256 3768 44320 3832
rect 44336 3768 44400 3832
rect 44416 3768 44480 3832
rect 44496 3768 44560 3832
rect 44576 3768 44640 3832
rect 44656 3768 44720 3832
rect 44736 3768 44800 3832
rect 44816 3768 44880 3832
rect 44896 3768 44960 3832
rect 44976 3768 45040 3832
rect 45056 3768 45120 3832
rect 45136 3768 45200 3832
rect 45216 3768 45280 3832
rect 45296 3768 45360 3832
rect 8 3688 72 3752
rect 88 3688 152 3752
rect 168 3688 232 3752
rect 248 3688 312 3752
rect 328 3688 392 3752
rect 408 3688 472 3752
rect 488 3688 552 3752
rect 568 3688 632 3752
rect 648 3688 712 3752
rect 728 3688 792 3752
rect 808 3688 872 3752
rect 888 3688 952 3752
rect 968 3688 1032 3752
rect 1048 3688 1112 3752
rect 1128 3688 1192 3752
rect 1208 3688 1272 3752
rect 1288 3688 1352 3752
rect 1368 3688 1432 3752
rect 1448 3688 1512 3752
rect 1528 3688 1592 3752
rect 1608 3688 1672 3752
rect 1688 3688 1752 3752
rect 1768 3688 1832 3752
rect 1848 3688 1912 3752
rect 1928 3688 1992 3752
rect 2008 3688 2072 3752
rect 2088 3688 2152 3752
rect 2168 3688 2232 3752
rect 2248 3688 2312 3752
rect 2328 3688 2392 3752
rect 2408 3688 2472 3752
rect 2488 3688 2552 3752
rect 2568 3688 2632 3752
rect 2648 3688 2712 3752
rect 2728 3688 2792 3752
rect 2808 3688 2872 3752
rect 2888 3688 2952 3752
rect 2968 3688 3032 3752
rect 3048 3688 3112 3752
rect 3128 3688 3192 3752
rect 3208 3688 3272 3752
rect 3288 3688 3352 3752
rect 3368 3688 3432 3752
rect 3448 3688 3512 3752
rect 3528 3688 3592 3752
rect 3608 3688 3672 3752
rect 3688 3688 3752 3752
rect 3768 3688 3832 3752
rect 3848 3688 3912 3752
rect 3928 3688 3992 3752
rect 19112 3688 19176 3752
rect 19192 3688 19256 3752
rect 19272 3688 19336 3752
rect 19352 3688 19416 3752
rect 29112 3688 29176 3752
rect 29192 3688 29256 3752
rect 29272 3688 29336 3752
rect 29352 3688 29416 3752
rect 41376 3688 41440 3752
rect 41456 3688 41520 3752
rect 41536 3688 41600 3752
rect 41616 3688 41680 3752
rect 41696 3688 41760 3752
rect 41776 3688 41840 3752
rect 41856 3688 41920 3752
rect 41936 3688 42000 3752
rect 42016 3688 42080 3752
rect 42096 3688 42160 3752
rect 42176 3688 42240 3752
rect 42256 3688 42320 3752
rect 42336 3688 42400 3752
rect 42416 3688 42480 3752
rect 42496 3688 42560 3752
rect 42576 3688 42640 3752
rect 42656 3688 42720 3752
rect 42736 3688 42800 3752
rect 42816 3688 42880 3752
rect 42896 3688 42960 3752
rect 42976 3688 43040 3752
rect 43056 3688 43120 3752
rect 43136 3688 43200 3752
rect 43216 3688 43280 3752
rect 43296 3688 43360 3752
rect 43376 3688 43440 3752
rect 43456 3688 43520 3752
rect 43536 3688 43600 3752
rect 43616 3688 43680 3752
rect 43696 3688 43760 3752
rect 43776 3688 43840 3752
rect 43856 3688 43920 3752
rect 43936 3688 44000 3752
rect 44016 3688 44080 3752
rect 44096 3688 44160 3752
rect 44176 3688 44240 3752
rect 44256 3688 44320 3752
rect 44336 3688 44400 3752
rect 44416 3688 44480 3752
rect 44496 3688 44560 3752
rect 44576 3688 44640 3752
rect 44656 3688 44720 3752
rect 44736 3688 44800 3752
rect 44816 3688 44880 3752
rect 44896 3688 44960 3752
rect 44976 3688 45040 3752
rect 45056 3688 45120 3752
rect 45136 3688 45200 3752
rect 45216 3688 45280 3752
rect 45296 3688 45360 3752
rect 8 3608 72 3672
rect 88 3608 152 3672
rect 168 3608 232 3672
rect 248 3608 312 3672
rect 328 3608 392 3672
rect 408 3608 472 3672
rect 488 3608 552 3672
rect 568 3608 632 3672
rect 648 3608 712 3672
rect 728 3608 792 3672
rect 808 3608 872 3672
rect 888 3608 952 3672
rect 968 3608 1032 3672
rect 1048 3608 1112 3672
rect 1128 3608 1192 3672
rect 1208 3608 1272 3672
rect 1288 3608 1352 3672
rect 1368 3608 1432 3672
rect 1448 3608 1512 3672
rect 1528 3608 1592 3672
rect 1608 3608 1672 3672
rect 1688 3608 1752 3672
rect 1768 3608 1832 3672
rect 1848 3608 1912 3672
rect 1928 3608 1992 3672
rect 2008 3608 2072 3672
rect 2088 3608 2152 3672
rect 2168 3608 2232 3672
rect 2248 3608 2312 3672
rect 2328 3608 2392 3672
rect 2408 3608 2472 3672
rect 2488 3608 2552 3672
rect 2568 3608 2632 3672
rect 2648 3608 2712 3672
rect 2728 3608 2792 3672
rect 2808 3608 2872 3672
rect 2888 3608 2952 3672
rect 2968 3608 3032 3672
rect 3048 3608 3112 3672
rect 3128 3608 3192 3672
rect 3208 3608 3272 3672
rect 3288 3608 3352 3672
rect 3368 3608 3432 3672
rect 3448 3608 3512 3672
rect 3528 3608 3592 3672
rect 3608 3608 3672 3672
rect 3688 3608 3752 3672
rect 3768 3608 3832 3672
rect 3848 3608 3912 3672
rect 3928 3608 3992 3672
rect 19112 3608 19176 3672
rect 19192 3608 19256 3672
rect 19272 3608 19336 3672
rect 19352 3608 19416 3672
rect 29112 3608 29176 3672
rect 29192 3608 29256 3672
rect 29272 3608 29336 3672
rect 29352 3608 29416 3672
rect 41376 3608 41440 3672
rect 41456 3608 41520 3672
rect 41536 3608 41600 3672
rect 41616 3608 41680 3672
rect 41696 3608 41760 3672
rect 41776 3608 41840 3672
rect 41856 3608 41920 3672
rect 41936 3608 42000 3672
rect 42016 3608 42080 3672
rect 42096 3608 42160 3672
rect 42176 3608 42240 3672
rect 42256 3608 42320 3672
rect 42336 3608 42400 3672
rect 42416 3608 42480 3672
rect 42496 3608 42560 3672
rect 42576 3608 42640 3672
rect 42656 3608 42720 3672
rect 42736 3608 42800 3672
rect 42816 3608 42880 3672
rect 42896 3608 42960 3672
rect 42976 3608 43040 3672
rect 43056 3608 43120 3672
rect 43136 3608 43200 3672
rect 43216 3608 43280 3672
rect 43296 3608 43360 3672
rect 43376 3608 43440 3672
rect 43456 3608 43520 3672
rect 43536 3608 43600 3672
rect 43616 3608 43680 3672
rect 43696 3608 43760 3672
rect 43776 3608 43840 3672
rect 43856 3608 43920 3672
rect 43936 3608 44000 3672
rect 44016 3608 44080 3672
rect 44096 3608 44160 3672
rect 44176 3608 44240 3672
rect 44256 3608 44320 3672
rect 44336 3608 44400 3672
rect 44416 3608 44480 3672
rect 44496 3608 44560 3672
rect 44576 3608 44640 3672
rect 44656 3608 44720 3672
rect 44736 3608 44800 3672
rect 44816 3608 44880 3672
rect 44896 3608 44960 3672
rect 44976 3608 45040 3672
rect 45056 3608 45120 3672
rect 45136 3608 45200 3672
rect 45216 3608 45280 3672
rect 45296 3608 45360 3672
rect 8 3528 72 3592
rect 88 3528 152 3592
rect 168 3528 232 3592
rect 248 3528 312 3592
rect 328 3528 392 3592
rect 408 3528 472 3592
rect 488 3528 552 3592
rect 568 3528 632 3592
rect 648 3528 712 3592
rect 728 3528 792 3592
rect 808 3528 872 3592
rect 888 3528 952 3592
rect 968 3528 1032 3592
rect 1048 3528 1112 3592
rect 1128 3528 1192 3592
rect 1208 3528 1272 3592
rect 1288 3528 1352 3592
rect 1368 3528 1432 3592
rect 1448 3528 1512 3592
rect 1528 3528 1592 3592
rect 1608 3528 1672 3592
rect 1688 3528 1752 3592
rect 1768 3528 1832 3592
rect 1848 3528 1912 3592
rect 1928 3528 1992 3592
rect 2008 3528 2072 3592
rect 2088 3528 2152 3592
rect 2168 3528 2232 3592
rect 2248 3528 2312 3592
rect 2328 3528 2392 3592
rect 2408 3528 2472 3592
rect 2488 3528 2552 3592
rect 2568 3528 2632 3592
rect 2648 3528 2712 3592
rect 2728 3528 2792 3592
rect 2808 3528 2872 3592
rect 2888 3528 2952 3592
rect 2968 3528 3032 3592
rect 3048 3528 3112 3592
rect 3128 3528 3192 3592
rect 3208 3528 3272 3592
rect 3288 3528 3352 3592
rect 3368 3528 3432 3592
rect 3448 3528 3512 3592
rect 3528 3528 3592 3592
rect 3608 3528 3672 3592
rect 3688 3528 3752 3592
rect 3768 3528 3832 3592
rect 3848 3528 3912 3592
rect 3928 3528 3992 3592
rect 19112 3528 19176 3592
rect 19192 3528 19256 3592
rect 19272 3528 19336 3592
rect 19352 3528 19416 3592
rect 29112 3528 29176 3592
rect 29192 3528 29256 3592
rect 29272 3528 29336 3592
rect 29352 3528 29416 3592
rect 41376 3528 41440 3592
rect 41456 3528 41520 3592
rect 41536 3528 41600 3592
rect 41616 3528 41680 3592
rect 41696 3528 41760 3592
rect 41776 3528 41840 3592
rect 41856 3528 41920 3592
rect 41936 3528 42000 3592
rect 42016 3528 42080 3592
rect 42096 3528 42160 3592
rect 42176 3528 42240 3592
rect 42256 3528 42320 3592
rect 42336 3528 42400 3592
rect 42416 3528 42480 3592
rect 42496 3528 42560 3592
rect 42576 3528 42640 3592
rect 42656 3528 42720 3592
rect 42736 3528 42800 3592
rect 42816 3528 42880 3592
rect 42896 3528 42960 3592
rect 42976 3528 43040 3592
rect 43056 3528 43120 3592
rect 43136 3528 43200 3592
rect 43216 3528 43280 3592
rect 43296 3528 43360 3592
rect 43376 3528 43440 3592
rect 43456 3528 43520 3592
rect 43536 3528 43600 3592
rect 43616 3528 43680 3592
rect 43696 3528 43760 3592
rect 43776 3528 43840 3592
rect 43856 3528 43920 3592
rect 43936 3528 44000 3592
rect 44016 3528 44080 3592
rect 44096 3528 44160 3592
rect 44176 3528 44240 3592
rect 44256 3528 44320 3592
rect 44336 3528 44400 3592
rect 44416 3528 44480 3592
rect 44496 3528 44560 3592
rect 44576 3528 44640 3592
rect 44656 3528 44720 3592
rect 44736 3528 44800 3592
rect 44816 3528 44880 3592
rect 44896 3528 44960 3592
rect 44976 3528 45040 3592
rect 45056 3528 45120 3592
rect 45136 3528 45200 3592
rect 45216 3528 45280 3592
rect 45296 3528 45360 3592
rect 8 3448 72 3512
rect 88 3448 152 3512
rect 168 3448 232 3512
rect 248 3448 312 3512
rect 328 3448 392 3512
rect 408 3448 472 3512
rect 488 3448 552 3512
rect 568 3448 632 3512
rect 648 3448 712 3512
rect 728 3448 792 3512
rect 808 3448 872 3512
rect 888 3448 952 3512
rect 968 3448 1032 3512
rect 1048 3448 1112 3512
rect 1128 3448 1192 3512
rect 1208 3448 1272 3512
rect 1288 3448 1352 3512
rect 1368 3448 1432 3512
rect 1448 3448 1512 3512
rect 1528 3448 1592 3512
rect 1608 3448 1672 3512
rect 1688 3448 1752 3512
rect 1768 3448 1832 3512
rect 1848 3448 1912 3512
rect 1928 3448 1992 3512
rect 2008 3448 2072 3512
rect 2088 3448 2152 3512
rect 2168 3448 2232 3512
rect 2248 3448 2312 3512
rect 2328 3448 2392 3512
rect 2408 3448 2472 3512
rect 2488 3448 2552 3512
rect 2568 3448 2632 3512
rect 2648 3448 2712 3512
rect 2728 3448 2792 3512
rect 2808 3448 2872 3512
rect 2888 3448 2952 3512
rect 2968 3448 3032 3512
rect 3048 3448 3112 3512
rect 3128 3448 3192 3512
rect 3208 3448 3272 3512
rect 3288 3448 3352 3512
rect 3368 3448 3432 3512
rect 3448 3448 3512 3512
rect 3528 3448 3592 3512
rect 3608 3448 3672 3512
rect 3688 3448 3752 3512
rect 3768 3448 3832 3512
rect 3848 3448 3912 3512
rect 3928 3448 3992 3512
rect 19112 3448 19176 3512
rect 19192 3448 19256 3512
rect 19272 3448 19336 3512
rect 19352 3448 19416 3512
rect 29112 3448 29176 3512
rect 29192 3448 29256 3512
rect 29272 3448 29336 3512
rect 29352 3448 29416 3512
rect 41376 3448 41440 3512
rect 41456 3448 41520 3512
rect 41536 3448 41600 3512
rect 41616 3448 41680 3512
rect 41696 3448 41760 3512
rect 41776 3448 41840 3512
rect 41856 3448 41920 3512
rect 41936 3448 42000 3512
rect 42016 3448 42080 3512
rect 42096 3448 42160 3512
rect 42176 3448 42240 3512
rect 42256 3448 42320 3512
rect 42336 3448 42400 3512
rect 42416 3448 42480 3512
rect 42496 3448 42560 3512
rect 42576 3448 42640 3512
rect 42656 3448 42720 3512
rect 42736 3448 42800 3512
rect 42816 3448 42880 3512
rect 42896 3448 42960 3512
rect 42976 3448 43040 3512
rect 43056 3448 43120 3512
rect 43136 3448 43200 3512
rect 43216 3448 43280 3512
rect 43296 3448 43360 3512
rect 43376 3448 43440 3512
rect 43456 3448 43520 3512
rect 43536 3448 43600 3512
rect 43616 3448 43680 3512
rect 43696 3448 43760 3512
rect 43776 3448 43840 3512
rect 43856 3448 43920 3512
rect 43936 3448 44000 3512
rect 44016 3448 44080 3512
rect 44096 3448 44160 3512
rect 44176 3448 44240 3512
rect 44256 3448 44320 3512
rect 44336 3448 44400 3512
rect 44416 3448 44480 3512
rect 44496 3448 44560 3512
rect 44576 3448 44640 3512
rect 44656 3448 44720 3512
rect 44736 3448 44800 3512
rect 44816 3448 44880 3512
rect 44896 3448 44960 3512
rect 44976 3448 45040 3512
rect 45056 3448 45120 3512
rect 45136 3448 45200 3512
rect 45216 3448 45280 3512
rect 45296 3448 45360 3512
rect 8 3368 72 3432
rect 88 3368 152 3432
rect 168 3368 232 3432
rect 248 3368 312 3432
rect 328 3368 392 3432
rect 408 3368 472 3432
rect 488 3368 552 3432
rect 568 3368 632 3432
rect 648 3368 712 3432
rect 728 3368 792 3432
rect 808 3368 872 3432
rect 888 3368 952 3432
rect 968 3368 1032 3432
rect 1048 3368 1112 3432
rect 1128 3368 1192 3432
rect 1208 3368 1272 3432
rect 1288 3368 1352 3432
rect 1368 3368 1432 3432
rect 1448 3368 1512 3432
rect 1528 3368 1592 3432
rect 1608 3368 1672 3432
rect 1688 3368 1752 3432
rect 1768 3368 1832 3432
rect 1848 3368 1912 3432
rect 1928 3368 1992 3432
rect 2008 3368 2072 3432
rect 2088 3368 2152 3432
rect 2168 3368 2232 3432
rect 2248 3368 2312 3432
rect 2328 3368 2392 3432
rect 2408 3368 2472 3432
rect 2488 3368 2552 3432
rect 2568 3368 2632 3432
rect 2648 3368 2712 3432
rect 2728 3368 2792 3432
rect 2808 3368 2872 3432
rect 2888 3368 2952 3432
rect 2968 3368 3032 3432
rect 3048 3368 3112 3432
rect 3128 3368 3192 3432
rect 3208 3368 3272 3432
rect 3288 3368 3352 3432
rect 3368 3368 3432 3432
rect 3448 3368 3512 3432
rect 3528 3368 3592 3432
rect 3608 3368 3672 3432
rect 3688 3368 3752 3432
rect 3768 3368 3832 3432
rect 3848 3368 3912 3432
rect 3928 3368 3992 3432
rect 19112 3368 19176 3432
rect 19192 3368 19256 3432
rect 19272 3368 19336 3432
rect 19352 3368 19416 3432
rect 29112 3368 29176 3432
rect 29192 3368 29256 3432
rect 29272 3368 29336 3432
rect 29352 3368 29416 3432
rect 41376 3368 41440 3432
rect 41456 3368 41520 3432
rect 41536 3368 41600 3432
rect 41616 3368 41680 3432
rect 41696 3368 41760 3432
rect 41776 3368 41840 3432
rect 41856 3368 41920 3432
rect 41936 3368 42000 3432
rect 42016 3368 42080 3432
rect 42096 3368 42160 3432
rect 42176 3368 42240 3432
rect 42256 3368 42320 3432
rect 42336 3368 42400 3432
rect 42416 3368 42480 3432
rect 42496 3368 42560 3432
rect 42576 3368 42640 3432
rect 42656 3368 42720 3432
rect 42736 3368 42800 3432
rect 42816 3368 42880 3432
rect 42896 3368 42960 3432
rect 42976 3368 43040 3432
rect 43056 3368 43120 3432
rect 43136 3368 43200 3432
rect 43216 3368 43280 3432
rect 43296 3368 43360 3432
rect 43376 3368 43440 3432
rect 43456 3368 43520 3432
rect 43536 3368 43600 3432
rect 43616 3368 43680 3432
rect 43696 3368 43760 3432
rect 43776 3368 43840 3432
rect 43856 3368 43920 3432
rect 43936 3368 44000 3432
rect 44016 3368 44080 3432
rect 44096 3368 44160 3432
rect 44176 3368 44240 3432
rect 44256 3368 44320 3432
rect 44336 3368 44400 3432
rect 44416 3368 44480 3432
rect 44496 3368 44560 3432
rect 44576 3368 44640 3432
rect 44656 3368 44720 3432
rect 44736 3368 44800 3432
rect 44816 3368 44880 3432
rect 44896 3368 44960 3432
rect 44976 3368 45040 3432
rect 45056 3368 45120 3432
rect 45136 3368 45200 3432
rect 45216 3368 45280 3432
rect 45296 3368 45360 3432
rect 8 3288 72 3352
rect 88 3288 152 3352
rect 168 3288 232 3352
rect 248 3288 312 3352
rect 328 3288 392 3352
rect 408 3288 472 3352
rect 488 3288 552 3352
rect 568 3288 632 3352
rect 648 3288 712 3352
rect 728 3288 792 3352
rect 808 3288 872 3352
rect 888 3288 952 3352
rect 968 3288 1032 3352
rect 1048 3288 1112 3352
rect 1128 3288 1192 3352
rect 1208 3288 1272 3352
rect 1288 3288 1352 3352
rect 1368 3288 1432 3352
rect 1448 3288 1512 3352
rect 1528 3288 1592 3352
rect 1608 3288 1672 3352
rect 1688 3288 1752 3352
rect 1768 3288 1832 3352
rect 1848 3288 1912 3352
rect 1928 3288 1992 3352
rect 2008 3288 2072 3352
rect 2088 3288 2152 3352
rect 2168 3288 2232 3352
rect 2248 3288 2312 3352
rect 2328 3288 2392 3352
rect 2408 3288 2472 3352
rect 2488 3288 2552 3352
rect 2568 3288 2632 3352
rect 2648 3288 2712 3352
rect 2728 3288 2792 3352
rect 2808 3288 2872 3352
rect 2888 3288 2952 3352
rect 2968 3288 3032 3352
rect 3048 3288 3112 3352
rect 3128 3288 3192 3352
rect 3208 3288 3272 3352
rect 3288 3288 3352 3352
rect 3368 3288 3432 3352
rect 3448 3288 3512 3352
rect 3528 3288 3592 3352
rect 3608 3288 3672 3352
rect 3688 3288 3752 3352
rect 3768 3288 3832 3352
rect 3848 3288 3912 3352
rect 3928 3288 3992 3352
rect 19112 3288 19176 3352
rect 19192 3288 19256 3352
rect 19272 3288 19336 3352
rect 19352 3288 19416 3352
rect 29112 3288 29176 3352
rect 29192 3288 29256 3352
rect 29272 3288 29336 3352
rect 29352 3288 29416 3352
rect 41376 3288 41440 3352
rect 41456 3288 41520 3352
rect 41536 3288 41600 3352
rect 41616 3288 41680 3352
rect 41696 3288 41760 3352
rect 41776 3288 41840 3352
rect 41856 3288 41920 3352
rect 41936 3288 42000 3352
rect 42016 3288 42080 3352
rect 42096 3288 42160 3352
rect 42176 3288 42240 3352
rect 42256 3288 42320 3352
rect 42336 3288 42400 3352
rect 42416 3288 42480 3352
rect 42496 3288 42560 3352
rect 42576 3288 42640 3352
rect 42656 3288 42720 3352
rect 42736 3288 42800 3352
rect 42816 3288 42880 3352
rect 42896 3288 42960 3352
rect 42976 3288 43040 3352
rect 43056 3288 43120 3352
rect 43136 3288 43200 3352
rect 43216 3288 43280 3352
rect 43296 3288 43360 3352
rect 43376 3288 43440 3352
rect 43456 3288 43520 3352
rect 43536 3288 43600 3352
rect 43616 3288 43680 3352
rect 43696 3288 43760 3352
rect 43776 3288 43840 3352
rect 43856 3288 43920 3352
rect 43936 3288 44000 3352
rect 44016 3288 44080 3352
rect 44096 3288 44160 3352
rect 44176 3288 44240 3352
rect 44256 3288 44320 3352
rect 44336 3288 44400 3352
rect 44416 3288 44480 3352
rect 44496 3288 44560 3352
rect 44576 3288 44640 3352
rect 44656 3288 44720 3352
rect 44736 3288 44800 3352
rect 44816 3288 44880 3352
rect 44896 3288 44960 3352
rect 44976 3288 45040 3352
rect 45056 3288 45120 3352
rect 45136 3288 45200 3352
rect 45216 3288 45280 3352
rect 45296 3288 45360 3352
rect 8 3208 72 3272
rect 88 3208 152 3272
rect 168 3208 232 3272
rect 248 3208 312 3272
rect 328 3208 392 3272
rect 408 3208 472 3272
rect 488 3208 552 3272
rect 568 3208 632 3272
rect 648 3208 712 3272
rect 728 3208 792 3272
rect 808 3208 872 3272
rect 888 3208 952 3272
rect 968 3208 1032 3272
rect 1048 3208 1112 3272
rect 1128 3208 1192 3272
rect 1208 3208 1272 3272
rect 1288 3208 1352 3272
rect 1368 3208 1432 3272
rect 1448 3208 1512 3272
rect 1528 3208 1592 3272
rect 1608 3208 1672 3272
rect 1688 3208 1752 3272
rect 1768 3208 1832 3272
rect 1848 3208 1912 3272
rect 1928 3208 1992 3272
rect 2008 3208 2072 3272
rect 2088 3208 2152 3272
rect 2168 3208 2232 3272
rect 2248 3208 2312 3272
rect 2328 3208 2392 3272
rect 2408 3208 2472 3272
rect 2488 3208 2552 3272
rect 2568 3208 2632 3272
rect 2648 3208 2712 3272
rect 2728 3208 2792 3272
rect 2808 3208 2872 3272
rect 2888 3208 2952 3272
rect 2968 3208 3032 3272
rect 3048 3208 3112 3272
rect 3128 3208 3192 3272
rect 3208 3208 3272 3272
rect 3288 3208 3352 3272
rect 3368 3208 3432 3272
rect 3448 3208 3512 3272
rect 3528 3208 3592 3272
rect 3608 3208 3672 3272
rect 3688 3208 3752 3272
rect 3768 3208 3832 3272
rect 3848 3208 3912 3272
rect 3928 3208 3992 3272
rect 19112 3208 19176 3272
rect 19192 3208 19256 3272
rect 19272 3208 19336 3272
rect 19352 3208 19416 3272
rect 29112 3208 29176 3272
rect 29192 3208 29256 3272
rect 29272 3208 29336 3272
rect 29352 3208 29416 3272
rect 41376 3208 41440 3272
rect 41456 3208 41520 3272
rect 41536 3208 41600 3272
rect 41616 3208 41680 3272
rect 41696 3208 41760 3272
rect 41776 3208 41840 3272
rect 41856 3208 41920 3272
rect 41936 3208 42000 3272
rect 42016 3208 42080 3272
rect 42096 3208 42160 3272
rect 42176 3208 42240 3272
rect 42256 3208 42320 3272
rect 42336 3208 42400 3272
rect 42416 3208 42480 3272
rect 42496 3208 42560 3272
rect 42576 3208 42640 3272
rect 42656 3208 42720 3272
rect 42736 3208 42800 3272
rect 42816 3208 42880 3272
rect 42896 3208 42960 3272
rect 42976 3208 43040 3272
rect 43056 3208 43120 3272
rect 43136 3208 43200 3272
rect 43216 3208 43280 3272
rect 43296 3208 43360 3272
rect 43376 3208 43440 3272
rect 43456 3208 43520 3272
rect 43536 3208 43600 3272
rect 43616 3208 43680 3272
rect 43696 3208 43760 3272
rect 43776 3208 43840 3272
rect 43856 3208 43920 3272
rect 43936 3208 44000 3272
rect 44016 3208 44080 3272
rect 44096 3208 44160 3272
rect 44176 3208 44240 3272
rect 44256 3208 44320 3272
rect 44336 3208 44400 3272
rect 44416 3208 44480 3272
rect 44496 3208 44560 3272
rect 44576 3208 44640 3272
rect 44656 3208 44720 3272
rect 44736 3208 44800 3272
rect 44816 3208 44880 3272
rect 44896 3208 44960 3272
rect 44976 3208 45040 3272
rect 45056 3208 45120 3272
rect 45136 3208 45200 3272
rect 45216 3208 45280 3272
rect 45296 3208 45360 3272
rect 8 3128 72 3192
rect 88 3128 152 3192
rect 168 3128 232 3192
rect 248 3128 312 3192
rect 328 3128 392 3192
rect 408 3128 472 3192
rect 488 3128 552 3192
rect 568 3128 632 3192
rect 648 3128 712 3192
rect 728 3128 792 3192
rect 808 3128 872 3192
rect 888 3128 952 3192
rect 968 3128 1032 3192
rect 1048 3128 1112 3192
rect 1128 3128 1192 3192
rect 1208 3128 1272 3192
rect 1288 3128 1352 3192
rect 1368 3128 1432 3192
rect 1448 3128 1512 3192
rect 1528 3128 1592 3192
rect 1608 3128 1672 3192
rect 1688 3128 1752 3192
rect 1768 3128 1832 3192
rect 1848 3128 1912 3192
rect 1928 3128 1992 3192
rect 2008 3128 2072 3192
rect 2088 3128 2152 3192
rect 2168 3128 2232 3192
rect 2248 3128 2312 3192
rect 2328 3128 2392 3192
rect 2408 3128 2472 3192
rect 2488 3128 2552 3192
rect 2568 3128 2632 3192
rect 2648 3128 2712 3192
rect 2728 3128 2792 3192
rect 2808 3128 2872 3192
rect 2888 3128 2952 3192
rect 2968 3128 3032 3192
rect 3048 3128 3112 3192
rect 3128 3128 3192 3192
rect 3208 3128 3272 3192
rect 3288 3128 3352 3192
rect 3368 3128 3432 3192
rect 3448 3128 3512 3192
rect 3528 3128 3592 3192
rect 3608 3128 3672 3192
rect 3688 3128 3752 3192
rect 3768 3128 3832 3192
rect 3848 3128 3912 3192
rect 3928 3128 3992 3192
rect 19112 3128 19176 3192
rect 19192 3128 19256 3192
rect 19272 3128 19336 3192
rect 19352 3128 19416 3192
rect 29112 3128 29176 3192
rect 29192 3128 29256 3192
rect 29272 3128 29336 3192
rect 29352 3128 29416 3192
rect 41376 3128 41440 3192
rect 41456 3128 41520 3192
rect 41536 3128 41600 3192
rect 41616 3128 41680 3192
rect 41696 3128 41760 3192
rect 41776 3128 41840 3192
rect 41856 3128 41920 3192
rect 41936 3128 42000 3192
rect 42016 3128 42080 3192
rect 42096 3128 42160 3192
rect 42176 3128 42240 3192
rect 42256 3128 42320 3192
rect 42336 3128 42400 3192
rect 42416 3128 42480 3192
rect 42496 3128 42560 3192
rect 42576 3128 42640 3192
rect 42656 3128 42720 3192
rect 42736 3128 42800 3192
rect 42816 3128 42880 3192
rect 42896 3128 42960 3192
rect 42976 3128 43040 3192
rect 43056 3128 43120 3192
rect 43136 3128 43200 3192
rect 43216 3128 43280 3192
rect 43296 3128 43360 3192
rect 43376 3128 43440 3192
rect 43456 3128 43520 3192
rect 43536 3128 43600 3192
rect 43616 3128 43680 3192
rect 43696 3128 43760 3192
rect 43776 3128 43840 3192
rect 43856 3128 43920 3192
rect 43936 3128 44000 3192
rect 44016 3128 44080 3192
rect 44096 3128 44160 3192
rect 44176 3128 44240 3192
rect 44256 3128 44320 3192
rect 44336 3128 44400 3192
rect 44416 3128 44480 3192
rect 44496 3128 44560 3192
rect 44576 3128 44640 3192
rect 44656 3128 44720 3192
rect 44736 3128 44800 3192
rect 44816 3128 44880 3192
rect 44896 3128 44960 3192
rect 44976 3128 45040 3192
rect 45056 3128 45120 3192
rect 45136 3128 45200 3192
rect 45216 3128 45280 3192
rect 45296 3128 45360 3192
rect 8 3048 72 3112
rect 88 3048 152 3112
rect 168 3048 232 3112
rect 248 3048 312 3112
rect 328 3048 392 3112
rect 408 3048 472 3112
rect 488 3048 552 3112
rect 568 3048 632 3112
rect 648 3048 712 3112
rect 728 3048 792 3112
rect 808 3048 872 3112
rect 888 3048 952 3112
rect 968 3048 1032 3112
rect 1048 3048 1112 3112
rect 1128 3048 1192 3112
rect 1208 3048 1272 3112
rect 1288 3048 1352 3112
rect 1368 3048 1432 3112
rect 1448 3048 1512 3112
rect 1528 3048 1592 3112
rect 1608 3048 1672 3112
rect 1688 3048 1752 3112
rect 1768 3048 1832 3112
rect 1848 3048 1912 3112
rect 1928 3048 1992 3112
rect 2008 3048 2072 3112
rect 2088 3048 2152 3112
rect 2168 3048 2232 3112
rect 2248 3048 2312 3112
rect 2328 3048 2392 3112
rect 2408 3048 2472 3112
rect 2488 3048 2552 3112
rect 2568 3048 2632 3112
rect 2648 3048 2712 3112
rect 2728 3048 2792 3112
rect 2808 3048 2872 3112
rect 2888 3048 2952 3112
rect 2968 3048 3032 3112
rect 3048 3048 3112 3112
rect 3128 3048 3192 3112
rect 3208 3048 3272 3112
rect 3288 3048 3352 3112
rect 3368 3048 3432 3112
rect 3448 3048 3512 3112
rect 3528 3048 3592 3112
rect 3608 3048 3672 3112
rect 3688 3048 3752 3112
rect 3768 3048 3832 3112
rect 3848 3048 3912 3112
rect 3928 3048 3992 3112
rect 19112 3048 19176 3112
rect 19192 3048 19256 3112
rect 19272 3048 19336 3112
rect 19352 3048 19416 3112
rect 29112 3048 29176 3112
rect 29192 3048 29256 3112
rect 29272 3048 29336 3112
rect 29352 3048 29416 3112
rect 41376 3048 41440 3112
rect 41456 3048 41520 3112
rect 41536 3048 41600 3112
rect 41616 3048 41680 3112
rect 41696 3048 41760 3112
rect 41776 3048 41840 3112
rect 41856 3048 41920 3112
rect 41936 3048 42000 3112
rect 42016 3048 42080 3112
rect 42096 3048 42160 3112
rect 42176 3048 42240 3112
rect 42256 3048 42320 3112
rect 42336 3048 42400 3112
rect 42416 3048 42480 3112
rect 42496 3048 42560 3112
rect 42576 3048 42640 3112
rect 42656 3048 42720 3112
rect 42736 3048 42800 3112
rect 42816 3048 42880 3112
rect 42896 3048 42960 3112
rect 42976 3048 43040 3112
rect 43056 3048 43120 3112
rect 43136 3048 43200 3112
rect 43216 3048 43280 3112
rect 43296 3048 43360 3112
rect 43376 3048 43440 3112
rect 43456 3048 43520 3112
rect 43536 3048 43600 3112
rect 43616 3048 43680 3112
rect 43696 3048 43760 3112
rect 43776 3048 43840 3112
rect 43856 3048 43920 3112
rect 43936 3048 44000 3112
rect 44016 3048 44080 3112
rect 44096 3048 44160 3112
rect 44176 3048 44240 3112
rect 44256 3048 44320 3112
rect 44336 3048 44400 3112
rect 44416 3048 44480 3112
rect 44496 3048 44560 3112
rect 44576 3048 44640 3112
rect 44656 3048 44720 3112
rect 44736 3048 44800 3112
rect 44816 3048 44880 3112
rect 44896 3048 44960 3112
rect 44976 3048 45040 3112
rect 45056 3048 45120 3112
rect 45136 3048 45200 3112
rect 45216 3048 45280 3112
rect 45296 3048 45360 3112
rect 8 2968 72 3032
rect 88 2968 152 3032
rect 168 2968 232 3032
rect 248 2968 312 3032
rect 328 2968 392 3032
rect 408 2968 472 3032
rect 488 2968 552 3032
rect 568 2968 632 3032
rect 648 2968 712 3032
rect 728 2968 792 3032
rect 808 2968 872 3032
rect 888 2968 952 3032
rect 968 2968 1032 3032
rect 1048 2968 1112 3032
rect 1128 2968 1192 3032
rect 1208 2968 1272 3032
rect 1288 2968 1352 3032
rect 1368 2968 1432 3032
rect 1448 2968 1512 3032
rect 1528 2968 1592 3032
rect 1608 2968 1672 3032
rect 1688 2968 1752 3032
rect 1768 2968 1832 3032
rect 1848 2968 1912 3032
rect 1928 2968 1992 3032
rect 2008 2968 2072 3032
rect 2088 2968 2152 3032
rect 2168 2968 2232 3032
rect 2248 2968 2312 3032
rect 2328 2968 2392 3032
rect 2408 2968 2472 3032
rect 2488 2968 2552 3032
rect 2568 2968 2632 3032
rect 2648 2968 2712 3032
rect 2728 2968 2792 3032
rect 2808 2968 2872 3032
rect 2888 2968 2952 3032
rect 2968 2968 3032 3032
rect 3048 2968 3112 3032
rect 3128 2968 3192 3032
rect 3208 2968 3272 3032
rect 3288 2968 3352 3032
rect 3368 2968 3432 3032
rect 3448 2968 3512 3032
rect 3528 2968 3592 3032
rect 3608 2968 3672 3032
rect 3688 2968 3752 3032
rect 3768 2968 3832 3032
rect 3848 2968 3912 3032
rect 3928 2968 3992 3032
rect 19112 2968 19176 3032
rect 19192 2968 19256 3032
rect 19272 2968 19336 3032
rect 19352 2968 19416 3032
rect 29112 2968 29176 3032
rect 29192 2968 29256 3032
rect 29272 2968 29336 3032
rect 29352 2968 29416 3032
rect 41376 2968 41440 3032
rect 41456 2968 41520 3032
rect 41536 2968 41600 3032
rect 41616 2968 41680 3032
rect 41696 2968 41760 3032
rect 41776 2968 41840 3032
rect 41856 2968 41920 3032
rect 41936 2968 42000 3032
rect 42016 2968 42080 3032
rect 42096 2968 42160 3032
rect 42176 2968 42240 3032
rect 42256 2968 42320 3032
rect 42336 2968 42400 3032
rect 42416 2968 42480 3032
rect 42496 2968 42560 3032
rect 42576 2968 42640 3032
rect 42656 2968 42720 3032
rect 42736 2968 42800 3032
rect 42816 2968 42880 3032
rect 42896 2968 42960 3032
rect 42976 2968 43040 3032
rect 43056 2968 43120 3032
rect 43136 2968 43200 3032
rect 43216 2968 43280 3032
rect 43296 2968 43360 3032
rect 43376 2968 43440 3032
rect 43456 2968 43520 3032
rect 43536 2968 43600 3032
rect 43616 2968 43680 3032
rect 43696 2968 43760 3032
rect 43776 2968 43840 3032
rect 43856 2968 43920 3032
rect 43936 2968 44000 3032
rect 44016 2968 44080 3032
rect 44096 2968 44160 3032
rect 44176 2968 44240 3032
rect 44256 2968 44320 3032
rect 44336 2968 44400 3032
rect 44416 2968 44480 3032
rect 44496 2968 44560 3032
rect 44576 2968 44640 3032
rect 44656 2968 44720 3032
rect 44736 2968 44800 3032
rect 44816 2968 44880 3032
rect 44896 2968 44960 3032
rect 44976 2968 45040 3032
rect 45056 2968 45120 3032
rect 45136 2968 45200 3032
rect 45216 2968 45280 3032
rect 45296 2968 45360 3032
rect 8 2888 72 2952
rect 88 2888 152 2952
rect 168 2888 232 2952
rect 248 2888 312 2952
rect 328 2888 392 2952
rect 408 2888 472 2952
rect 488 2888 552 2952
rect 568 2888 632 2952
rect 648 2888 712 2952
rect 728 2888 792 2952
rect 808 2888 872 2952
rect 888 2888 952 2952
rect 968 2888 1032 2952
rect 1048 2888 1112 2952
rect 1128 2888 1192 2952
rect 1208 2888 1272 2952
rect 1288 2888 1352 2952
rect 1368 2888 1432 2952
rect 1448 2888 1512 2952
rect 1528 2888 1592 2952
rect 1608 2888 1672 2952
rect 1688 2888 1752 2952
rect 1768 2888 1832 2952
rect 1848 2888 1912 2952
rect 1928 2888 1992 2952
rect 2008 2888 2072 2952
rect 2088 2888 2152 2952
rect 2168 2888 2232 2952
rect 2248 2888 2312 2952
rect 2328 2888 2392 2952
rect 2408 2888 2472 2952
rect 2488 2888 2552 2952
rect 2568 2888 2632 2952
rect 2648 2888 2712 2952
rect 2728 2888 2792 2952
rect 2808 2888 2872 2952
rect 2888 2888 2952 2952
rect 2968 2888 3032 2952
rect 3048 2888 3112 2952
rect 3128 2888 3192 2952
rect 3208 2888 3272 2952
rect 3288 2888 3352 2952
rect 3368 2888 3432 2952
rect 3448 2888 3512 2952
rect 3528 2888 3592 2952
rect 3608 2888 3672 2952
rect 3688 2888 3752 2952
rect 3768 2888 3832 2952
rect 3848 2888 3912 2952
rect 3928 2888 3992 2952
rect 19112 2888 19176 2952
rect 19192 2888 19256 2952
rect 19272 2888 19336 2952
rect 19352 2888 19416 2952
rect 29112 2888 29176 2952
rect 29192 2888 29256 2952
rect 29272 2888 29336 2952
rect 29352 2888 29416 2952
rect 41376 2888 41440 2952
rect 41456 2888 41520 2952
rect 41536 2888 41600 2952
rect 41616 2888 41680 2952
rect 41696 2888 41760 2952
rect 41776 2888 41840 2952
rect 41856 2888 41920 2952
rect 41936 2888 42000 2952
rect 42016 2888 42080 2952
rect 42096 2888 42160 2952
rect 42176 2888 42240 2952
rect 42256 2888 42320 2952
rect 42336 2888 42400 2952
rect 42416 2888 42480 2952
rect 42496 2888 42560 2952
rect 42576 2888 42640 2952
rect 42656 2888 42720 2952
rect 42736 2888 42800 2952
rect 42816 2888 42880 2952
rect 42896 2888 42960 2952
rect 42976 2888 43040 2952
rect 43056 2888 43120 2952
rect 43136 2888 43200 2952
rect 43216 2888 43280 2952
rect 43296 2888 43360 2952
rect 43376 2888 43440 2952
rect 43456 2888 43520 2952
rect 43536 2888 43600 2952
rect 43616 2888 43680 2952
rect 43696 2888 43760 2952
rect 43776 2888 43840 2952
rect 43856 2888 43920 2952
rect 43936 2888 44000 2952
rect 44016 2888 44080 2952
rect 44096 2888 44160 2952
rect 44176 2888 44240 2952
rect 44256 2888 44320 2952
rect 44336 2888 44400 2952
rect 44416 2888 44480 2952
rect 44496 2888 44560 2952
rect 44576 2888 44640 2952
rect 44656 2888 44720 2952
rect 44736 2888 44800 2952
rect 44816 2888 44880 2952
rect 44896 2888 44960 2952
rect 44976 2888 45040 2952
rect 45056 2888 45120 2952
rect 45136 2888 45200 2952
rect 45216 2888 45280 2952
rect 45296 2888 45360 2952
rect 8 2808 72 2872
rect 88 2808 152 2872
rect 168 2808 232 2872
rect 248 2808 312 2872
rect 328 2808 392 2872
rect 408 2808 472 2872
rect 488 2808 552 2872
rect 568 2808 632 2872
rect 648 2808 712 2872
rect 728 2808 792 2872
rect 808 2808 872 2872
rect 888 2808 952 2872
rect 968 2808 1032 2872
rect 1048 2808 1112 2872
rect 1128 2808 1192 2872
rect 1208 2808 1272 2872
rect 1288 2808 1352 2872
rect 1368 2808 1432 2872
rect 1448 2808 1512 2872
rect 1528 2808 1592 2872
rect 1608 2808 1672 2872
rect 1688 2808 1752 2872
rect 1768 2808 1832 2872
rect 1848 2808 1912 2872
rect 1928 2808 1992 2872
rect 2008 2808 2072 2872
rect 2088 2808 2152 2872
rect 2168 2808 2232 2872
rect 2248 2808 2312 2872
rect 2328 2808 2392 2872
rect 2408 2808 2472 2872
rect 2488 2808 2552 2872
rect 2568 2808 2632 2872
rect 2648 2808 2712 2872
rect 2728 2808 2792 2872
rect 2808 2808 2872 2872
rect 2888 2808 2952 2872
rect 2968 2808 3032 2872
rect 3048 2808 3112 2872
rect 3128 2808 3192 2872
rect 3208 2808 3272 2872
rect 3288 2808 3352 2872
rect 3368 2808 3432 2872
rect 3448 2808 3512 2872
rect 3528 2808 3592 2872
rect 3608 2808 3672 2872
rect 3688 2808 3752 2872
rect 3768 2808 3832 2872
rect 3848 2808 3912 2872
rect 3928 2808 3992 2872
rect 19112 2808 19176 2872
rect 19192 2808 19256 2872
rect 19272 2808 19336 2872
rect 19352 2808 19416 2872
rect 29112 2808 29176 2872
rect 29192 2808 29256 2872
rect 29272 2808 29336 2872
rect 29352 2808 29416 2872
rect 41376 2808 41440 2872
rect 41456 2808 41520 2872
rect 41536 2808 41600 2872
rect 41616 2808 41680 2872
rect 41696 2808 41760 2872
rect 41776 2808 41840 2872
rect 41856 2808 41920 2872
rect 41936 2808 42000 2872
rect 42016 2808 42080 2872
rect 42096 2808 42160 2872
rect 42176 2808 42240 2872
rect 42256 2808 42320 2872
rect 42336 2808 42400 2872
rect 42416 2808 42480 2872
rect 42496 2808 42560 2872
rect 42576 2808 42640 2872
rect 42656 2808 42720 2872
rect 42736 2808 42800 2872
rect 42816 2808 42880 2872
rect 42896 2808 42960 2872
rect 42976 2808 43040 2872
rect 43056 2808 43120 2872
rect 43136 2808 43200 2872
rect 43216 2808 43280 2872
rect 43296 2808 43360 2872
rect 43376 2808 43440 2872
rect 43456 2808 43520 2872
rect 43536 2808 43600 2872
rect 43616 2808 43680 2872
rect 43696 2808 43760 2872
rect 43776 2808 43840 2872
rect 43856 2808 43920 2872
rect 43936 2808 44000 2872
rect 44016 2808 44080 2872
rect 44096 2808 44160 2872
rect 44176 2808 44240 2872
rect 44256 2808 44320 2872
rect 44336 2808 44400 2872
rect 44416 2808 44480 2872
rect 44496 2808 44560 2872
rect 44576 2808 44640 2872
rect 44656 2808 44720 2872
rect 44736 2808 44800 2872
rect 44816 2808 44880 2872
rect 44896 2808 44960 2872
rect 44976 2808 45040 2872
rect 45056 2808 45120 2872
rect 45136 2808 45200 2872
rect 45216 2808 45280 2872
rect 45296 2808 45360 2872
rect 8 2728 72 2792
rect 88 2728 152 2792
rect 168 2728 232 2792
rect 248 2728 312 2792
rect 328 2728 392 2792
rect 408 2728 472 2792
rect 488 2728 552 2792
rect 568 2728 632 2792
rect 648 2728 712 2792
rect 728 2728 792 2792
rect 808 2728 872 2792
rect 888 2728 952 2792
rect 968 2728 1032 2792
rect 1048 2728 1112 2792
rect 1128 2728 1192 2792
rect 1208 2728 1272 2792
rect 1288 2728 1352 2792
rect 1368 2728 1432 2792
rect 1448 2728 1512 2792
rect 1528 2728 1592 2792
rect 1608 2728 1672 2792
rect 1688 2728 1752 2792
rect 1768 2728 1832 2792
rect 1848 2728 1912 2792
rect 1928 2728 1992 2792
rect 2008 2728 2072 2792
rect 2088 2728 2152 2792
rect 2168 2728 2232 2792
rect 2248 2728 2312 2792
rect 2328 2728 2392 2792
rect 2408 2728 2472 2792
rect 2488 2728 2552 2792
rect 2568 2728 2632 2792
rect 2648 2728 2712 2792
rect 2728 2728 2792 2792
rect 2808 2728 2872 2792
rect 2888 2728 2952 2792
rect 2968 2728 3032 2792
rect 3048 2728 3112 2792
rect 3128 2728 3192 2792
rect 3208 2728 3272 2792
rect 3288 2728 3352 2792
rect 3368 2728 3432 2792
rect 3448 2728 3512 2792
rect 3528 2728 3592 2792
rect 3608 2728 3672 2792
rect 3688 2728 3752 2792
rect 3768 2728 3832 2792
rect 3848 2728 3912 2792
rect 3928 2728 3992 2792
rect 19112 2728 19176 2792
rect 19192 2728 19256 2792
rect 19272 2728 19336 2792
rect 19352 2728 19416 2792
rect 29112 2728 29176 2792
rect 29192 2728 29256 2792
rect 29272 2728 29336 2792
rect 29352 2728 29416 2792
rect 41376 2728 41440 2792
rect 41456 2728 41520 2792
rect 41536 2728 41600 2792
rect 41616 2728 41680 2792
rect 41696 2728 41760 2792
rect 41776 2728 41840 2792
rect 41856 2728 41920 2792
rect 41936 2728 42000 2792
rect 42016 2728 42080 2792
rect 42096 2728 42160 2792
rect 42176 2728 42240 2792
rect 42256 2728 42320 2792
rect 42336 2728 42400 2792
rect 42416 2728 42480 2792
rect 42496 2728 42560 2792
rect 42576 2728 42640 2792
rect 42656 2728 42720 2792
rect 42736 2728 42800 2792
rect 42816 2728 42880 2792
rect 42896 2728 42960 2792
rect 42976 2728 43040 2792
rect 43056 2728 43120 2792
rect 43136 2728 43200 2792
rect 43216 2728 43280 2792
rect 43296 2728 43360 2792
rect 43376 2728 43440 2792
rect 43456 2728 43520 2792
rect 43536 2728 43600 2792
rect 43616 2728 43680 2792
rect 43696 2728 43760 2792
rect 43776 2728 43840 2792
rect 43856 2728 43920 2792
rect 43936 2728 44000 2792
rect 44016 2728 44080 2792
rect 44096 2728 44160 2792
rect 44176 2728 44240 2792
rect 44256 2728 44320 2792
rect 44336 2728 44400 2792
rect 44416 2728 44480 2792
rect 44496 2728 44560 2792
rect 44576 2728 44640 2792
rect 44656 2728 44720 2792
rect 44736 2728 44800 2792
rect 44816 2728 44880 2792
rect 44896 2728 44960 2792
rect 44976 2728 45040 2792
rect 45056 2728 45120 2792
rect 45136 2728 45200 2792
rect 45216 2728 45280 2792
rect 45296 2728 45360 2792
rect 8 2648 72 2712
rect 88 2648 152 2712
rect 168 2648 232 2712
rect 248 2648 312 2712
rect 328 2648 392 2712
rect 408 2648 472 2712
rect 488 2648 552 2712
rect 568 2648 632 2712
rect 648 2648 712 2712
rect 728 2648 792 2712
rect 808 2648 872 2712
rect 888 2648 952 2712
rect 968 2648 1032 2712
rect 1048 2648 1112 2712
rect 1128 2648 1192 2712
rect 1208 2648 1272 2712
rect 1288 2648 1352 2712
rect 1368 2648 1432 2712
rect 1448 2648 1512 2712
rect 1528 2648 1592 2712
rect 1608 2648 1672 2712
rect 1688 2648 1752 2712
rect 1768 2648 1832 2712
rect 1848 2648 1912 2712
rect 1928 2648 1992 2712
rect 2008 2648 2072 2712
rect 2088 2648 2152 2712
rect 2168 2648 2232 2712
rect 2248 2648 2312 2712
rect 2328 2648 2392 2712
rect 2408 2648 2472 2712
rect 2488 2648 2552 2712
rect 2568 2648 2632 2712
rect 2648 2648 2712 2712
rect 2728 2648 2792 2712
rect 2808 2648 2872 2712
rect 2888 2648 2952 2712
rect 2968 2648 3032 2712
rect 3048 2648 3112 2712
rect 3128 2648 3192 2712
rect 3208 2648 3272 2712
rect 3288 2648 3352 2712
rect 3368 2648 3432 2712
rect 3448 2648 3512 2712
rect 3528 2648 3592 2712
rect 3608 2648 3672 2712
rect 3688 2648 3752 2712
rect 3768 2648 3832 2712
rect 3848 2648 3912 2712
rect 3928 2648 3992 2712
rect 19112 2648 19176 2712
rect 19192 2648 19256 2712
rect 19272 2648 19336 2712
rect 19352 2648 19416 2712
rect 29112 2648 29176 2712
rect 29192 2648 29256 2712
rect 29272 2648 29336 2712
rect 29352 2648 29416 2712
rect 41376 2648 41440 2712
rect 41456 2648 41520 2712
rect 41536 2648 41600 2712
rect 41616 2648 41680 2712
rect 41696 2648 41760 2712
rect 41776 2648 41840 2712
rect 41856 2648 41920 2712
rect 41936 2648 42000 2712
rect 42016 2648 42080 2712
rect 42096 2648 42160 2712
rect 42176 2648 42240 2712
rect 42256 2648 42320 2712
rect 42336 2648 42400 2712
rect 42416 2648 42480 2712
rect 42496 2648 42560 2712
rect 42576 2648 42640 2712
rect 42656 2648 42720 2712
rect 42736 2648 42800 2712
rect 42816 2648 42880 2712
rect 42896 2648 42960 2712
rect 42976 2648 43040 2712
rect 43056 2648 43120 2712
rect 43136 2648 43200 2712
rect 43216 2648 43280 2712
rect 43296 2648 43360 2712
rect 43376 2648 43440 2712
rect 43456 2648 43520 2712
rect 43536 2648 43600 2712
rect 43616 2648 43680 2712
rect 43696 2648 43760 2712
rect 43776 2648 43840 2712
rect 43856 2648 43920 2712
rect 43936 2648 44000 2712
rect 44016 2648 44080 2712
rect 44096 2648 44160 2712
rect 44176 2648 44240 2712
rect 44256 2648 44320 2712
rect 44336 2648 44400 2712
rect 44416 2648 44480 2712
rect 44496 2648 44560 2712
rect 44576 2648 44640 2712
rect 44656 2648 44720 2712
rect 44736 2648 44800 2712
rect 44816 2648 44880 2712
rect 44896 2648 44960 2712
rect 44976 2648 45040 2712
rect 45056 2648 45120 2712
rect 45136 2648 45200 2712
rect 45216 2648 45280 2712
rect 45296 2648 45360 2712
rect 8 2568 72 2632
rect 88 2568 152 2632
rect 168 2568 232 2632
rect 248 2568 312 2632
rect 328 2568 392 2632
rect 408 2568 472 2632
rect 488 2568 552 2632
rect 568 2568 632 2632
rect 648 2568 712 2632
rect 728 2568 792 2632
rect 808 2568 872 2632
rect 888 2568 952 2632
rect 968 2568 1032 2632
rect 1048 2568 1112 2632
rect 1128 2568 1192 2632
rect 1208 2568 1272 2632
rect 1288 2568 1352 2632
rect 1368 2568 1432 2632
rect 1448 2568 1512 2632
rect 1528 2568 1592 2632
rect 1608 2568 1672 2632
rect 1688 2568 1752 2632
rect 1768 2568 1832 2632
rect 1848 2568 1912 2632
rect 1928 2568 1992 2632
rect 2008 2568 2072 2632
rect 2088 2568 2152 2632
rect 2168 2568 2232 2632
rect 2248 2568 2312 2632
rect 2328 2568 2392 2632
rect 2408 2568 2472 2632
rect 2488 2568 2552 2632
rect 2568 2568 2632 2632
rect 2648 2568 2712 2632
rect 2728 2568 2792 2632
rect 2808 2568 2872 2632
rect 2888 2568 2952 2632
rect 2968 2568 3032 2632
rect 3048 2568 3112 2632
rect 3128 2568 3192 2632
rect 3208 2568 3272 2632
rect 3288 2568 3352 2632
rect 3368 2568 3432 2632
rect 3448 2568 3512 2632
rect 3528 2568 3592 2632
rect 3608 2568 3672 2632
rect 3688 2568 3752 2632
rect 3768 2568 3832 2632
rect 3848 2568 3912 2632
rect 3928 2568 3992 2632
rect 19112 2568 19176 2632
rect 19192 2568 19256 2632
rect 19272 2568 19336 2632
rect 19352 2568 19416 2632
rect 29112 2568 29176 2632
rect 29192 2568 29256 2632
rect 29272 2568 29336 2632
rect 29352 2568 29416 2632
rect 41376 2568 41440 2632
rect 41456 2568 41520 2632
rect 41536 2568 41600 2632
rect 41616 2568 41680 2632
rect 41696 2568 41760 2632
rect 41776 2568 41840 2632
rect 41856 2568 41920 2632
rect 41936 2568 42000 2632
rect 42016 2568 42080 2632
rect 42096 2568 42160 2632
rect 42176 2568 42240 2632
rect 42256 2568 42320 2632
rect 42336 2568 42400 2632
rect 42416 2568 42480 2632
rect 42496 2568 42560 2632
rect 42576 2568 42640 2632
rect 42656 2568 42720 2632
rect 42736 2568 42800 2632
rect 42816 2568 42880 2632
rect 42896 2568 42960 2632
rect 42976 2568 43040 2632
rect 43056 2568 43120 2632
rect 43136 2568 43200 2632
rect 43216 2568 43280 2632
rect 43296 2568 43360 2632
rect 43376 2568 43440 2632
rect 43456 2568 43520 2632
rect 43536 2568 43600 2632
rect 43616 2568 43680 2632
rect 43696 2568 43760 2632
rect 43776 2568 43840 2632
rect 43856 2568 43920 2632
rect 43936 2568 44000 2632
rect 44016 2568 44080 2632
rect 44096 2568 44160 2632
rect 44176 2568 44240 2632
rect 44256 2568 44320 2632
rect 44336 2568 44400 2632
rect 44416 2568 44480 2632
rect 44496 2568 44560 2632
rect 44576 2568 44640 2632
rect 44656 2568 44720 2632
rect 44736 2568 44800 2632
rect 44816 2568 44880 2632
rect 44896 2568 44960 2632
rect 44976 2568 45040 2632
rect 45056 2568 45120 2632
rect 45136 2568 45200 2632
rect 45216 2568 45280 2632
rect 45296 2568 45360 2632
rect 8 2488 72 2552
rect 88 2488 152 2552
rect 168 2488 232 2552
rect 248 2488 312 2552
rect 328 2488 392 2552
rect 408 2488 472 2552
rect 488 2488 552 2552
rect 568 2488 632 2552
rect 648 2488 712 2552
rect 728 2488 792 2552
rect 808 2488 872 2552
rect 888 2488 952 2552
rect 968 2488 1032 2552
rect 1048 2488 1112 2552
rect 1128 2488 1192 2552
rect 1208 2488 1272 2552
rect 1288 2488 1352 2552
rect 1368 2488 1432 2552
rect 1448 2488 1512 2552
rect 1528 2488 1592 2552
rect 1608 2488 1672 2552
rect 1688 2488 1752 2552
rect 1768 2488 1832 2552
rect 1848 2488 1912 2552
rect 1928 2488 1992 2552
rect 2008 2488 2072 2552
rect 2088 2488 2152 2552
rect 2168 2488 2232 2552
rect 2248 2488 2312 2552
rect 2328 2488 2392 2552
rect 2408 2488 2472 2552
rect 2488 2488 2552 2552
rect 2568 2488 2632 2552
rect 2648 2488 2712 2552
rect 2728 2488 2792 2552
rect 2808 2488 2872 2552
rect 2888 2488 2952 2552
rect 2968 2488 3032 2552
rect 3048 2488 3112 2552
rect 3128 2488 3192 2552
rect 3208 2488 3272 2552
rect 3288 2488 3352 2552
rect 3368 2488 3432 2552
rect 3448 2488 3512 2552
rect 3528 2488 3592 2552
rect 3608 2488 3672 2552
rect 3688 2488 3752 2552
rect 3768 2488 3832 2552
rect 3848 2488 3912 2552
rect 3928 2488 3992 2552
rect 19112 2488 19176 2552
rect 19192 2488 19256 2552
rect 19272 2488 19336 2552
rect 19352 2488 19416 2552
rect 29112 2488 29176 2552
rect 29192 2488 29256 2552
rect 29272 2488 29336 2552
rect 29352 2488 29416 2552
rect 41376 2488 41440 2552
rect 41456 2488 41520 2552
rect 41536 2488 41600 2552
rect 41616 2488 41680 2552
rect 41696 2488 41760 2552
rect 41776 2488 41840 2552
rect 41856 2488 41920 2552
rect 41936 2488 42000 2552
rect 42016 2488 42080 2552
rect 42096 2488 42160 2552
rect 42176 2488 42240 2552
rect 42256 2488 42320 2552
rect 42336 2488 42400 2552
rect 42416 2488 42480 2552
rect 42496 2488 42560 2552
rect 42576 2488 42640 2552
rect 42656 2488 42720 2552
rect 42736 2488 42800 2552
rect 42816 2488 42880 2552
rect 42896 2488 42960 2552
rect 42976 2488 43040 2552
rect 43056 2488 43120 2552
rect 43136 2488 43200 2552
rect 43216 2488 43280 2552
rect 43296 2488 43360 2552
rect 43376 2488 43440 2552
rect 43456 2488 43520 2552
rect 43536 2488 43600 2552
rect 43616 2488 43680 2552
rect 43696 2488 43760 2552
rect 43776 2488 43840 2552
rect 43856 2488 43920 2552
rect 43936 2488 44000 2552
rect 44016 2488 44080 2552
rect 44096 2488 44160 2552
rect 44176 2488 44240 2552
rect 44256 2488 44320 2552
rect 44336 2488 44400 2552
rect 44416 2488 44480 2552
rect 44496 2488 44560 2552
rect 44576 2488 44640 2552
rect 44656 2488 44720 2552
rect 44736 2488 44800 2552
rect 44816 2488 44880 2552
rect 44896 2488 44960 2552
rect 44976 2488 45040 2552
rect 45056 2488 45120 2552
rect 45136 2488 45200 2552
rect 45216 2488 45280 2552
rect 45296 2488 45360 2552
rect 8 2408 72 2472
rect 88 2408 152 2472
rect 168 2408 232 2472
rect 248 2408 312 2472
rect 328 2408 392 2472
rect 408 2408 472 2472
rect 488 2408 552 2472
rect 568 2408 632 2472
rect 648 2408 712 2472
rect 728 2408 792 2472
rect 808 2408 872 2472
rect 888 2408 952 2472
rect 968 2408 1032 2472
rect 1048 2408 1112 2472
rect 1128 2408 1192 2472
rect 1208 2408 1272 2472
rect 1288 2408 1352 2472
rect 1368 2408 1432 2472
rect 1448 2408 1512 2472
rect 1528 2408 1592 2472
rect 1608 2408 1672 2472
rect 1688 2408 1752 2472
rect 1768 2408 1832 2472
rect 1848 2408 1912 2472
rect 1928 2408 1992 2472
rect 2008 2408 2072 2472
rect 2088 2408 2152 2472
rect 2168 2408 2232 2472
rect 2248 2408 2312 2472
rect 2328 2408 2392 2472
rect 2408 2408 2472 2472
rect 2488 2408 2552 2472
rect 2568 2408 2632 2472
rect 2648 2408 2712 2472
rect 2728 2408 2792 2472
rect 2808 2408 2872 2472
rect 2888 2408 2952 2472
rect 2968 2408 3032 2472
rect 3048 2408 3112 2472
rect 3128 2408 3192 2472
rect 3208 2408 3272 2472
rect 3288 2408 3352 2472
rect 3368 2408 3432 2472
rect 3448 2408 3512 2472
rect 3528 2408 3592 2472
rect 3608 2408 3672 2472
rect 3688 2408 3752 2472
rect 3768 2408 3832 2472
rect 3848 2408 3912 2472
rect 3928 2408 3992 2472
rect 19112 2408 19176 2472
rect 19192 2408 19256 2472
rect 19272 2408 19336 2472
rect 19352 2408 19416 2472
rect 29112 2408 29176 2472
rect 29192 2408 29256 2472
rect 29272 2408 29336 2472
rect 29352 2408 29416 2472
rect 41376 2408 41440 2472
rect 41456 2408 41520 2472
rect 41536 2408 41600 2472
rect 41616 2408 41680 2472
rect 41696 2408 41760 2472
rect 41776 2408 41840 2472
rect 41856 2408 41920 2472
rect 41936 2408 42000 2472
rect 42016 2408 42080 2472
rect 42096 2408 42160 2472
rect 42176 2408 42240 2472
rect 42256 2408 42320 2472
rect 42336 2408 42400 2472
rect 42416 2408 42480 2472
rect 42496 2408 42560 2472
rect 42576 2408 42640 2472
rect 42656 2408 42720 2472
rect 42736 2408 42800 2472
rect 42816 2408 42880 2472
rect 42896 2408 42960 2472
rect 42976 2408 43040 2472
rect 43056 2408 43120 2472
rect 43136 2408 43200 2472
rect 43216 2408 43280 2472
rect 43296 2408 43360 2472
rect 43376 2408 43440 2472
rect 43456 2408 43520 2472
rect 43536 2408 43600 2472
rect 43616 2408 43680 2472
rect 43696 2408 43760 2472
rect 43776 2408 43840 2472
rect 43856 2408 43920 2472
rect 43936 2408 44000 2472
rect 44016 2408 44080 2472
rect 44096 2408 44160 2472
rect 44176 2408 44240 2472
rect 44256 2408 44320 2472
rect 44336 2408 44400 2472
rect 44416 2408 44480 2472
rect 44496 2408 44560 2472
rect 44576 2408 44640 2472
rect 44656 2408 44720 2472
rect 44736 2408 44800 2472
rect 44816 2408 44880 2472
rect 44896 2408 44960 2472
rect 44976 2408 45040 2472
rect 45056 2408 45120 2472
rect 45136 2408 45200 2472
rect 45216 2408 45280 2472
rect 45296 2408 45360 2472
rect 8 2328 72 2392
rect 88 2328 152 2392
rect 168 2328 232 2392
rect 248 2328 312 2392
rect 328 2328 392 2392
rect 408 2328 472 2392
rect 488 2328 552 2392
rect 568 2328 632 2392
rect 648 2328 712 2392
rect 728 2328 792 2392
rect 808 2328 872 2392
rect 888 2328 952 2392
rect 968 2328 1032 2392
rect 1048 2328 1112 2392
rect 1128 2328 1192 2392
rect 1208 2328 1272 2392
rect 1288 2328 1352 2392
rect 1368 2328 1432 2392
rect 1448 2328 1512 2392
rect 1528 2328 1592 2392
rect 1608 2328 1672 2392
rect 1688 2328 1752 2392
rect 1768 2328 1832 2392
rect 1848 2328 1912 2392
rect 1928 2328 1992 2392
rect 2008 2328 2072 2392
rect 2088 2328 2152 2392
rect 2168 2328 2232 2392
rect 2248 2328 2312 2392
rect 2328 2328 2392 2392
rect 2408 2328 2472 2392
rect 2488 2328 2552 2392
rect 2568 2328 2632 2392
rect 2648 2328 2712 2392
rect 2728 2328 2792 2392
rect 2808 2328 2872 2392
rect 2888 2328 2952 2392
rect 2968 2328 3032 2392
rect 3048 2328 3112 2392
rect 3128 2328 3192 2392
rect 3208 2328 3272 2392
rect 3288 2328 3352 2392
rect 3368 2328 3432 2392
rect 3448 2328 3512 2392
rect 3528 2328 3592 2392
rect 3608 2328 3672 2392
rect 3688 2328 3752 2392
rect 3768 2328 3832 2392
rect 3848 2328 3912 2392
rect 3928 2328 3992 2392
rect 19112 2328 19176 2392
rect 19192 2328 19256 2392
rect 19272 2328 19336 2392
rect 19352 2328 19416 2392
rect 29112 2328 29176 2392
rect 29192 2328 29256 2392
rect 29272 2328 29336 2392
rect 29352 2328 29416 2392
rect 41376 2328 41440 2392
rect 41456 2328 41520 2392
rect 41536 2328 41600 2392
rect 41616 2328 41680 2392
rect 41696 2328 41760 2392
rect 41776 2328 41840 2392
rect 41856 2328 41920 2392
rect 41936 2328 42000 2392
rect 42016 2328 42080 2392
rect 42096 2328 42160 2392
rect 42176 2328 42240 2392
rect 42256 2328 42320 2392
rect 42336 2328 42400 2392
rect 42416 2328 42480 2392
rect 42496 2328 42560 2392
rect 42576 2328 42640 2392
rect 42656 2328 42720 2392
rect 42736 2328 42800 2392
rect 42816 2328 42880 2392
rect 42896 2328 42960 2392
rect 42976 2328 43040 2392
rect 43056 2328 43120 2392
rect 43136 2328 43200 2392
rect 43216 2328 43280 2392
rect 43296 2328 43360 2392
rect 43376 2328 43440 2392
rect 43456 2328 43520 2392
rect 43536 2328 43600 2392
rect 43616 2328 43680 2392
rect 43696 2328 43760 2392
rect 43776 2328 43840 2392
rect 43856 2328 43920 2392
rect 43936 2328 44000 2392
rect 44016 2328 44080 2392
rect 44096 2328 44160 2392
rect 44176 2328 44240 2392
rect 44256 2328 44320 2392
rect 44336 2328 44400 2392
rect 44416 2328 44480 2392
rect 44496 2328 44560 2392
rect 44576 2328 44640 2392
rect 44656 2328 44720 2392
rect 44736 2328 44800 2392
rect 44816 2328 44880 2392
rect 44896 2328 44960 2392
rect 44976 2328 45040 2392
rect 45056 2328 45120 2392
rect 45136 2328 45200 2392
rect 45216 2328 45280 2392
rect 45296 2328 45360 2392
rect 8 2248 72 2312
rect 88 2248 152 2312
rect 168 2248 232 2312
rect 248 2248 312 2312
rect 328 2248 392 2312
rect 408 2248 472 2312
rect 488 2248 552 2312
rect 568 2248 632 2312
rect 648 2248 712 2312
rect 728 2248 792 2312
rect 808 2248 872 2312
rect 888 2248 952 2312
rect 968 2248 1032 2312
rect 1048 2248 1112 2312
rect 1128 2248 1192 2312
rect 1208 2248 1272 2312
rect 1288 2248 1352 2312
rect 1368 2248 1432 2312
rect 1448 2248 1512 2312
rect 1528 2248 1592 2312
rect 1608 2248 1672 2312
rect 1688 2248 1752 2312
rect 1768 2248 1832 2312
rect 1848 2248 1912 2312
rect 1928 2248 1992 2312
rect 2008 2248 2072 2312
rect 2088 2248 2152 2312
rect 2168 2248 2232 2312
rect 2248 2248 2312 2312
rect 2328 2248 2392 2312
rect 2408 2248 2472 2312
rect 2488 2248 2552 2312
rect 2568 2248 2632 2312
rect 2648 2248 2712 2312
rect 2728 2248 2792 2312
rect 2808 2248 2872 2312
rect 2888 2248 2952 2312
rect 2968 2248 3032 2312
rect 3048 2248 3112 2312
rect 3128 2248 3192 2312
rect 3208 2248 3272 2312
rect 3288 2248 3352 2312
rect 3368 2248 3432 2312
rect 3448 2248 3512 2312
rect 3528 2248 3592 2312
rect 3608 2248 3672 2312
rect 3688 2248 3752 2312
rect 3768 2248 3832 2312
rect 3848 2248 3912 2312
rect 3928 2248 3992 2312
rect 19112 2248 19176 2312
rect 19192 2248 19256 2312
rect 19272 2248 19336 2312
rect 19352 2248 19416 2312
rect 29112 2248 29176 2312
rect 29192 2248 29256 2312
rect 29272 2248 29336 2312
rect 29352 2248 29416 2312
rect 41376 2248 41440 2312
rect 41456 2248 41520 2312
rect 41536 2248 41600 2312
rect 41616 2248 41680 2312
rect 41696 2248 41760 2312
rect 41776 2248 41840 2312
rect 41856 2248 41920 2312
rect 41936 2248 42000 2312
rect 42016 2248 42080 2312
rect 42096 2248 42160 2312
rect 42176 2248 42240 2312
rect 42256 2248 42320 2312
rect 42336 2248 42400 2312
rect 42416 2248 42480 2312
rect 42496 2248 42560 2312
rect 42576 2248 42640 2312
rect 42656 2248 42720 2312
rect 42736 2248 42800 2312
rect 42816 2248 42880 2312
rect 42896 2248 42960 2312
rect 42976 2248 43040 2312
rect 43056 2248 43120 2312
rect 43136 2248 43200 2312
rect 43216 2248 43280 2312
rect 43296 2248 43360 2312
rect 43376 2248 43440 2312
rect 43456 2248 43520 2312
rect 43536 2248 43600 2312
rect 43616 2248 43680 2312
rect 43696 2248 43760 2312
rect 43776 2248 43840 2312
rect 43856 2248 43920 2312
rect 43936 2248 44000 2312
rect 44016 2248 44080 2312
rect 44096 2248 44160 2312
rect 44176 2248 44240 2312
rect 44256 2248 44320 2312
rect 44336 2248 44400 2312
rect 44416 2248 44480 2312
rect 44496 2248 44560 2312
rect 44576 2248 44640 2312
rect 44656 2248 44720 2312
rect 44736 2248 44800 2312
rect 44816 2248 44880 2312
rect 44896 2248 44960 2312
rect 44976 2248 45040 2312
rect 45056 2248 45120 2312
rect 45136 2248 45200 2312
rect 45216 2248 45280 2312
rect 45296 2248 45360 2312
rect 8 2168 72 2232
rect 88 2168 152 2232
rect 168 2168 232 2232
rect 248 2168 312 2232
rect 328 2168 392 2232
rect 408 2168 472 2232
rect 488 2168 552 2232
rect 568 2168 632 2232
rect 648 2168 712 2232
rect 728 2168 792 2232
rect 808 2168 872 2232
rect 888 2168 952 2232
rect 968 2168 1032 2232
rect 1048 2168 1112 2232
rect 1128 2168 1192 2232
rect 1208 2168 1272 2232
rect 1288 2168 1352 2232
rect 1368 2168 1432 2232
rect 1448 2168 1512 2232
rect 1528 2168 1592 2232
rect 1608 2168 1672 2232
rect 1688 2168 1752 2232
rect 1768 2168 1832 2232
rect 1848 2168 1912 2232
rect 1928 2168 1992 2232
rect 2008 2168 2072 2232
rect 2088 2168 2152 2232
rect 2168 2168 2232 2232
rect 2248 2168 2312 2232
rect 2328 2168 2392 2232
rect 2408 2168 2472 2232
rect 2488 2168 2552 2232
rect 2568 2168 2632 2232
rect 2648 2168 2712 2232
rect 2728 2168 2792 2232
rect 2808 2168 2872 2232
rect 2888 2168 2952 2232
rect 2968 2168 3032 2232
rect 3048 2168 3112 2232
rect 3128 2168 3192 2232
rect 3208 2168 3272 2232
rect 3288 2168 3352 2232
rect 3368 2168 3432 2232
rect 3448 2168 3512 2232
rect 3528 2168 3592 2232
rect 3608 2168 3672 2232
rect 3688 2168 3752 2232
rect 3768 2168 3832 2232
rect 3848 2168 3912 2232
rect 3928 2168 3992 2232
rect 19112 2168 19176 2232
rect 19192 2168 19256 2232
rect 19272 2168 19336 2232
rect 19352 2168 19416 2232
rect 29112 2168 29176 2232
rect 29192 2168 29256 2232
rect 29272 2168 29336 2232
rect 29352 2168 29416 2232
rect 41376 2168 41440 2232
rect 41456 2168 41520 2232
rect 41536 2168 41600 2232
rect 41616 2168 41680 2232
rect 41696 2168 41760 2232
rect 41776 2168 41840 2232
rect 41856 2168 41920 2232
rect 41936 2168 42000 2232
rect 42016 2168 42080 2232
rect 42096 2168 42160 2232
rect 42176 2168 42240 2232
rect 42256 2168 42320 2232
rect 42336 2168 42400 2232
rect 42416 2168 42480 2232
rect 42496 2168 42560 2232
rect 42576 2168 42640 2232
rect 42656 2168 42720 2232
rect 42736 2168 42800 2232
rect 42816 2168 42880 2232
rect 42896 2168 42960 2232
rect 42976 2168 43040 2232
rect 43056 2168 43120 2232
rect 43136 2168 43200 2232
rect 43216 2168 43280 2232
rect 43296 2168 43360 2232
rect 43376 2168 43440 2232
rect 43456 2168 43520 2232
rect 43536 2168 43600 2232
rect 43616 2168 43680 2232
rect 43696 2168 43760 2232
rect 43776 2168 43840 2232
rect 43856 2168 43920 2232
rect 43936 2168 44000 2232
rect 44016 2168 44080 2232
rect 44096 2168 44160 2232
rect 44176 2168 44240 2232
rect 44256 2168 44320 2232
rect 44336 2168 44400 2232
rect 44416 2168 44480 2232
rect 44496 2168 44560 2232
rect 44576 2168 44640 2232
rect 44656 2168 44720 2232
rect 44736 2168 44800 2232
rect 44816 2168 44880 2232
rect 44896 2168 44960 2232
rect 44976 2168 45040 2232
rect 45056 2168 45120 2232
rect 45136 2168 45200 2232
rect 45216 2168 45280 2232
rect 45296 2168 45360 2232
rect 8 2088 72 2152
rect 88 2088 152 2152
rect 168 2088 232 2152
rect 248 2088 312 2152
rect 328 2088 392 2152
rect 408 2088 472 2152
rect 488 2088 552 2152
rect 568 2088 632 2152
rect 648 2088 712 2152
rect 728 2088 792 2152
rect 808 2088 872 2152
rect 888 2088 952 2152
rect 968 2088 1032 2152
rect 1048 2088 1112 2152
rect 1128 2088 1192 2152
rect 1208 2088 1272 2152
rect 1288 2088 1352 2152
rect 1368 2088 1432 2152
rect 1448 2088 1512 2152
rect 1528 2088 1592 2152
rect 1608 2088 1672 2152
rect 1688 2088 1752 2152
rect 1768 2088 1832 2152
rect 1848 2088 1912 2152
rect 1928 2088 1992 2152
rect 2008 2088 2072 2152
rect 2088 2088 2152 2152
rect 2168 2088 2232 2152
rect 2248 2088 2312 2152
rect 2328 2088 2392 2152
rect 2408 2088 2472 2152
rect 2488 2088 2552 2152
rect 2568 2088 2632 2152
rect 2648 2088 2712 2152
rect 2728 2088 2792 2152
rect 2808 2088 2872 2152
rect 2888 2088 2952 2152
rect 2968 2088 3032 2152
rect 3048 2088 3112 2152
rect 3128 2088 3192 2152
rect 3208 2088 3272 2152
rect 3288 2088 3352 2152
rect 3368 2088 3432 2152
rect 3448 2088 3512 2152
rect 3528 2088 3592 2152
rect 3608 2088 3672 2152
rect 3688 2088 3752 2152
rect 3768 2088 3832 2152
rect 3848 2088 3912 2152
rect 3928 2088 3992 2152
rect 19112 2088 19176 2152
rect 19192 2088 19256 2152
rect 19272 2088 19336 2152
rect 19352 2088 19416 2152
rect 29112 2088 29176 2152
rect 29192 2088 29256 2152
rect 29272 2088 29336 2152
rect 29352 2088 29416 2152
rect 41376 2088 41440 2152
rect 41456 2088 41520 2152
rect 41536 2088 41600 2152
rect 41616 2088 41680 2152
rect 41696 2088 41760 2152
rect 41776 2088 41840 2152
rect 41856 2088 41920 2152
rect 41936 2088 42000 2152
rect 42016 2088 42080 2152
rect 42096 2088 42160 2152
rect 42176 2088 42240 2152
rect 42256 2088 42320 2152
rect 42336 2088 42400 2152
rect 42416 2088 42480 2152
rect 42496 2088 42560 2152
rect 42576 2088 42640 2152
rect 42656 2088 42720 2152
rect 42736 2088 42800 2152
rect 42816 2088 42880 2152
rect 42896 2088 42960 2152
rect 42976 2088 43040 2152
rect 43056 2088 43120 2152
rect 43136 2088 43200 2152
rect 43216 2088 43280 2152
rect 43296 2088 43360 2152
rect 43376 2088 43440 2152
rect 43456 2088 43520 2152
rect 43536 2088 43600 2152
rect 43616 2088 43680 2152
rect 43696 2088 43760 2152
rect 43776 2088 43840 2152
rect 43856 2088 43920 2152
rect 43936 2088 44000 2152
rect 44016 2088 44080 2152
rect 44096 2088 44160 2152
rect 44176 2088 44240 2152
rect 44256 2088 44320 2152
rect 44336 2088 44400 2152
rect 44416 2088 44480 2152
rect 44496 2088 44560 2152
rect 44576 2088 44640 2152
rect 44656 2088 44720 2152
rect 44736 2088 44800 2152
rect 44816 2088 44880 2152
rect 44896 2088 44960 2152
rect 44976 2088 45040 2152
rect 45056 2088 45120 2152
rect 45136 2088 45200 2152
rect 45216 2088 45280 2152
rect 45296 2088 45360 2152
rect 8 2008 72 2072
rect 88 2008 152 2072
rect 168 2008 232 2072
rect 248 2008 312 2072
rect 328 2008 392 2072
rect 408 2008 472 2072
rect 488 2008 552 2072
rect 568 2008 632 2072
rect 648 2008 712 2072
rect 728 2008 792 2072
rect 808 2008 872 2072
rect 888 2008 952 2072
rect 968 2008 1032 2072
rect 1048 2008 1112 2072
rect 1128 2008 1192 2072
rect 1208 2008 1272 2072
rect 1288 2008 1352 2072
rect 1368 2008 1432 2072
rect 1448 2008 1512 2072
rect 1528 2008 1592 2072
rect 1608 2008 1672 2072
rect 1688 2008 1752 2072
rect 1768 2008 1832 2072
rect 1848 2008 1912 2072
rect 1928 2008 1992 2072
rect 2008 2008 2072 2072
rect 2088 2008 2152 2072
rect 2168 2008 2232 2072
rect 2248 2008 2312 2072
rect 2328 2008 2392 2072
rect 2408 2008 2472 2072
rect 2488 2008 2552 2072
rect 2568 2008 2632 2072
rect 2648 2008 2712 2072
rect 2728 2008 2792 2072
rect 2808 2008 2872 2072
rect 2888 2008 2952 2072
rect 2968 2008 3032 2072
rect 3048 2008 3112 2072
rect 3128 2008 3192 2072
rect 3208 2008 3272 2072
rect 3288 2008 3352 2072
rect 3368 2008 3432 2072
rect 3448 2008 3512 2072
rect 3528 2008 3592 2072
rect 3608 2008 3672 2072
rect 3688 2008 3752 2072
rect 3768 2008 3832 2072
rect 3848 2008 3912 2072
rect 3928 2008 3992 2072
rect 19112 2008 19176 2072
rect 19192 2008 19256 2072
rect 19272 2008 19336 2072
rect 19352 2008 19416 2072
rect 29112 2008 29176 2072
rect 29192 2008 29256 2072
rect 29272 2008 29336 2072
rect 29352 2008 29416 2072
rect 41376 2008 41440 2072
rect 41456 2008 41520 2072
rect 41536 2008 41600 2072
rect 41616 2008 41680 2072
rect 41696 2008 41760 2072
rect 41776 2008 41840 2072
rect 41856 2008 41920 2072
rect 41936 2008 42000 2072
rect 42016 2008 42080 2072
rect 42096 2008 42160 2072
rect 42176 2008 42240 2072
rect 42256 2008 42320 2072
rect 42336 2008 42400 2072
rect 42416 2008 42480 2072
rect 42496 2008 42560 2072
rect 42576 2008 42640 2072
rect 42656 2008 42720 2072
rect 42736 2008 42800 2072
rect 42816 2008 42880 2072
rect 42896 2008 42960 2072
rect 42976 2008 43040 2072
rect 43056 2008 43120 2072
rect 43136 2008 43200 2072
rect 43216 2008 43280 2072
rect 43296 2008 43360 2072
rect 43376 2008 43440 2072
rect 43456 2008 43520 2072
rect 43536 2008 43600 2072
rect 43616 2008 43680 2072
rect 43696 2008 43760 2072
rect 43776 2008 43840 2072
rect 43856 2008 43920 2072
rect 43936 2008 44000 2072
rect 44016 2008 44080 2072
rect 44096 2008 44160 2072
rect 44176 2008 44240 2072
rect 44256 2008 44320 2072
rect 44336 2008 44400 2072
rect 44416 2008 44480 2072
rect 44496 2008 44560 2072
rect 44576 2008 44640 2072
rect 44656 2008 44720 2072
rect 44736 2008 44800 2072
rect 44816 2008 44880 2072
rect 44896 2008 44960 2072
rect 44976 2008 45040 2072
rect 45056 2008 45120 2072
rect 45136 2008 45200 2072
rect 45216 2008 45280 2072
rect 45296 2008 45360 2072
rect 8 1928 72 1992
rect 88 1928 152 1992
rect 168 1928 232 1992
rect 248 1928 312 1992
rect 328 1928 392 1992
rect 408 1928 472 1992
rect 488 1928 552 1992
rect 568 1928 632 1992
rect 648 1928 712 1992
rect 728 1928 792 1992
rect 808 1928 872 1992
rect 888 1928 952 1992
rect 968 1928 1032 1992
rect 1048 1928 1112 1992
rect 1128 1928 1192 1992
rect 1208 1928 1272 1992
rect 1288 1928 1352 1992
rect 1368 1928 1432 1992
rect 1448 1928 1512 1992
rect 1528 1928 1592 1992
rect 1608 1928 1672 1992
rect 1688 1928 1752 1992
rect 1768 1928 1832 1992
rect 1848 1928 1912 1992
rect 1928 1928 1992 1992
rect 2008 1928 2072 1992
rect 2088 1928 2152 1992
rect 2168 1928 2232 1992
rect 2248 1928 2312 1992
rect 2328 1928 2392 1992
rect 2408 1928 2472 1992
rect 2488 1928 2552 1992
rect 2568 1928 2632 1992
rect 2648 1928 2712 1992
rect 2728 1928 2792 1992
rect 2808 1928 2872 1992
rect 2888 1928 2952 1992
rect 2968 1928 3032 1992
rect 3048 1928 3112 1992
rect 3128 1928 3192 1992
rect 3208 1928 3272 1992
rect 3288 1928 3352 1992
rect 3368 1928 3432 1992
rect 3448 1928 3512 1992
rect 3528 1928 3592 1992
rect 3608 1928 3672 1992
rect 3688 1928 3752 1992
rect 3768 1928 3832 1992
rect 3848 1928 3912 1992
rect 3928 1928 3992 1992
rect 19112 1928 19176 1992
rect 19192 1928 19256 1992
rect 19272 1928 19336 1992
rect 19352 1928 19416 1992
rect 29112 1928 29176 1992
rect 29192 1928 29256 1992
rect 29272 1928 29336 1992
rect 29352 1928 29416 1992
rect 41376 1928 41440 1992
rect 41456 1928 41520 1992
rect 41536 1928 41600 1992
rect 41616 1928 41680 1992
rect 41696 1928 41760 1992
rect 41776 1928 41840 1992
rect 41856 1928 41920 1992
rect 41936 1928 42000 1992
rect 42016 1928 42080 1992
rect 42096 1928 42160 1992
rect 42176 1928 42240 1992
rect 42256 1928 42320 1992
rect 42336 1928 42400 1992
rect 42416 1928 42480 1992
rect 42496 1928 42560 1992
rect 42576 1928 42640 1992
rect 42656 1928 42720 1992
rect 42736 1928 42800 1992
rect 42816 1928 42880 1992
rect 42896 1928 42960 1992
rect 42976 1928 43040 1992
rect 43056 1928 43120 1992
rect 43136 1928 43200 1992
rect 43216 1928 43280 1992
rect 43296 1928 43360 1992
rect 43376 1928 43440 1992
rect 43456 1928 43520 1992
rect 43536 1928 43600 1992
rect 43616 1928 43680 1992
rect 43696 1928 43760 1992
rect 43776 1928 43840 1992
rect 43856 1928 43920 1992
rect 43936 1928 44000 1992
rect 44016 1928 44080 1992
rect 44096 1928 44160 1992
rect 44176 1928 44240 1992
rect 44256 1928 44320 1992
rect 44336 1928 44400 1992
rect 44416 1928 44480 1992
rect 44496 1928 44560 1992
rect 44576 1928 44640 1992
rect 44656 1928 44720 1992
rect 44736 1928 44800 1992
rect 44816 1928 44880 1992
rect 44896 1928 44960 1992
rect 44976 1928 45040 1992
rect 45056 1928 45120 1992
rect 45136 1928 45200 1992
rect 45216 1928 45280 1992
rect 45296 1928 45360 1992
rect 8 1848 72 1912
rect 88 1848 152 1912
rect 168 1848 232 1912
rect 248 1848 312 1912
rect 328 1848 392 1912
rect 408 1848 472 1912
rect 488 1848 552 1912
rect 568 1848 632 1912
rect 648 1848 712 1912
rect 728 1848 792 1912
rect 808 1848 872 1912
rect 888 1848 952 1912
rect 968 1848 1032 1912
rect 1048 1848 1112 1912
rect 1128 1848 1192 1912
rect 1208 1848 1272 1912
rect 1288 1848 1352 1912
rect 1368 1848 1432 1912
rect 1448 1848 1512 1912
rect 1528 1848 1592 1912
rect 1608 1848 1672 1912
rect 1688 1848 1752 1912
rect 1768 1848 1832 1912
rect 1848 1848 1912 1912
rect 1928 1848 1992 1912
rect 2008 1848 2072 1912
rect 2088 1848 2152 1912
rect 2168 1848 2232 1912
rect 2248 1848 2312 1912
rect 2328 1848 2392 1912
rect 2408 1848 2472 1912
rect 2488 1848 2552 1912
rect 2568 1848 2632 1912
rect 2648 1848 2712 1912
rect 2728 1848 2792 1912
rect 2808 1848 2872 1912
rect 2888 1848 2952 1912
rect 2968 1848 3032 1912
rect 3048 1848 3112 1912
rect 3128 1848 3192 1912
rect 3208 1848 3272 1912
rect 3288 1848 3352 1912
rect 3368 1848 3432 1912
rect 3448 1848 3512 1912
rect 3528 1848 3592 1912
rect 3608 1848 3672 1912
rect 3688 1848 3752 1912
rect 3768 1848 3832 1912
rect 3848 1848 3912 1912
rect 3928 1848 3992 1912
rect 19112 1848 19176 1912
rect 19192 1848 19256 1912
rect 19272 1848 19336 1912
rect 19352 1848 19416 1912
rect 29112 1848 29176 1912
rect 29192 1848 29256 1912
rect 29272 1848 29336 1912
rect 29352 1848 29416 1912
rect 41376 1848 41440 1912
rect 41456 1848 41520 1912
rect 41536 1848 41600 1912
rect 41616 1848 41680 1912
rect 41696 1848 41760 1912
rect 41776 1848 41840 1912
rect 41856 1848 41920 1912
rect 41936 1848 42000 1912
rect 42016 1848 42080 1912
rect 42096 1848 42160 1912
rect 42176 1848 42240 1912
rect 42256 1848 42320 1912
rect 42336 1848 42400 1912
rect 42416 1848 42480 1912
rect 42496 1848 42560 1912
rect 42576 1848 42640 1912
rect 42656 1848 42720 1912
rect 42736 1848 42800 1912
rect 42816 1848 42880 1912
rect 42896 1848 42960 1912
rect 42976 1848 43040 1912
rect 43056 1848 43120 1912
rect 43136 1848 43200 1912
rect 43216 1848 43280 1912
rect 43296 1848 43360 1912
rect 43376 1848 43440 1912
rect 43456 1848 43520 1912
rect 43536 1848 43600 1912
rect 43616 1848 43680 1912
rect 43696 1848 43760 1912
rect 43776 1848 43840 1912
rect 43856 1848 43920 1912
rect 43936 1848 44000 1912
rect 44016 1848 44080 1912
rect 44096 1848 44160 1912
rect 44176 1848 44240 1912
rect 44256 1848 44320 1912
rect 44336 1848 44400 1912
rect 44416 1848 44480 1912
rect 44496 1848 44560 1912
rect 44576 1848 44640 1912
rect 44656 1848 44720 1912
rect 44736 1848 44800 1912
rect 44816 1848 44880 1912
rect 44896 1848 44960 1912
rect 44976 1848 45040 1912
rect 45056 1848 45120 1912
rect 45136 1848 45200 1912
rect 45216 1848 45280 1912
rect 45296 1848 45360 1912
rect 8 1768 72 1832
rect 88 1768 152 1832
rect 168 1768 232 1832
rect 248 1768 312 1832
rect 328 1768 392 1832
rect 408 1768 472 1832
rect 488 1768 552 1832
rect 568 1768 632 1832
rect 648 1768 712 1832
rect 728 1768 792 1832
rect 808 1768 872 1832
rect 888 1768 952 1832
rect 968 1768 1032 1832
rect 1048 1768 1112 1832
rect 1128 1768 1192 1832
rect 1208 1768 1272 1832
rect 1288 1768 1352 1832
rect 1368 1768 1432 1832
rect 1448 1768 1512 1832
rect 1528 1768 1592 1832
rect 1608 1768 1672 1832
rect 1688 1768 1752 1832
rect 1768 1768 1832 1832
rect 1848 1768 1912 1832
rect 1928 1768 1992 1832
rect 2008 1768 2072 1832
rect 2088 1768 2152 1832
rect 2168 1768 2232 1832
rect 2248 1768 2312 1832
rect 2328 1768 2392 1832
rect 2408 1768 2472 1832
rect 2488 1768 2552 1832
rect 2568 1768 2632 1832
rect 2648 1768 2712 1832
rect 2728 1768 2792 1832
rect 2808 1768 2872 1832
rect 2888 1768 2952 1832
rect 2968 1768 3032 1832
rect 3048 1768 3112 1832
rect 3128 1768 3192 1832
rect 3208 1768 3272 1832
rect 3288 1768 3352 1832
rect 3368 1768 3432 1832
rect 3448 1768 3512 1832
rect 3528 1768 3592 1832
rect 3608 1768 3672 1832
rect 3688 1768 3752 1832
rect 3768 1768 3832 1832
rect 3848 1768 3912 1832
rect 3928 1768 3992 1832
rect 19112 1768 19176 1832
rect 19192 1768 19256 1832
rect 19272 1768 19336 1832
rect 19352 1768 19416 1832
rect 29112 1768 29176 1832
rect 29192 1768 29256 1832
rect 29272 1768 29336 1832
rect 29352 1768 29416 1832
rect 41376 1768 41440 1832
rect 41456 1768 41520 1832
rect 41536 1768 41600 1832
rect 41616 1768 41680 1832
rect 41696 1768 41760 1832
rect 41776 1768 41840 1832
rect 41856 1768 41920 1832
rect 41936 1768 42000 1832
rect 42016 1768 42080 1832
rect 42096 1768 42160 1832
rect 42176 1768 42240 1832
rect 42256 1768 42320 1832
rect 42336 1768 42400 1832
rect 42416 1768 42480 1832
rect 42496 1768 42560 1832
rect 42576 1768 42640 1832
rect 42656 1768 42720 1832
rect 42736 1768 42800 1832
rect 42816 1768 42880 1832
rect 42896 1768 42960 1832
rect 42976 1768 43040 1832
rect 43056 1768 43120 1832
rect 43136 1768 43200 1832
rect 43216 1768 43280 1832
rect 43296 1768 43360 1832
rect 43376 1768 43440 1832
rect 43456 1768 43520 1832
rect 43536 1768 43600 1832
rect 43616 1768 43680 1832
rect 43696 1768 43760 1832
rect 43776 1768 43840 1832
rect 43856 1768 43920 1832
rect 43936 1768 44000 1832
rect 44016 1768 44080 1832
rect 44096 1768 44160 1832
rect 44176 1768 44240 1832
rect 44256 1768 44320 1832
rect 44336 1768 44400 1832
rect 44416 1768 44480 1832
rect 44496 1768 44560 1832
rect 44576 1768 44640 1832
rect 44656 1768 44720 1832
rect 44736 1768 44800 1832
rect 44816 1768 44880 1832
rect 44896 1768 44960 1832
rect 44976 1768 45040 1832
rect 45056 1768 45120 1832
rect 45136 1768 45200 1832
rect 45216 1768 45280 1832
rect 45296 1768 45360 1832
rect 8 1688 72 1752
rect 88 1688 152 1752
rect 168 1688 232 1752
rect 248 1688 312 1752
rect 328 1688 392 1752
rect 408 1688 472 1752
rect 488 1688 552 1752
rect 568 1688 632 1752
rect 648 1688 712 1752
rect 728 1688 792 1752
rect 808 1688 872 1752
rect 888 1688 952 1752
rect 968 1688 1032 1752
rect 1048 1688 1112 1752
rect 1128 1688 1192 1752
rect 1208 1688 1272 1752
rect 1288 1688 1352 1752
rect 1368 1688 1432 1752
rect 1448 1688 1512 1752
rect 1528 1688 1592 1752
rect 1608 1688 1672 1752
rect 1688 1688 1752 1752
rect 1768 1688 1832 1752
rect 1848 1688 1912 1752
rect 1928 1688 1992 1752
rect 2008 1688 2072 1752
rect 2088 1688 2152 1752
rect 2168 1688 2232 1752
rect 2248 1688 2312 1752
rect 2328 1688 2392 1752
rect 2408 1688 2472 1752
rect 2488 1688 2552 1752
rect 2568 1688 2632 1752
rect 2648 1688 2712 1752
rect 2728 1688 2792 1752
rect 2808 1688 2872 1752
rect 2888 1688 2952 1752
rect 2968 1688 3032 1752
rect 3048 1688 3112 1752
rect 3128 1688 3192 1752
rect 3208 1688 3272 1752
rect 3288 1688 3352 1752
rect 3368 1688 3432 1752
rect 3448 1688 3512 1752
rect 3528 1688 3592 1752
rect 3608 1688 3672 1752
rect 3688 1688 3752 1752
rect 3768 1688 3832 1752
rect 3848 1688 3912 1752
rect 3928 1688 3992 1752
rect 19112 1688 19176 1752
rect 19192 1688 19256 1752
rect 19272 1688 19336 1752
rect 19352 1688 19416 1752
rect 29112 1688 29176 1752
rect 29192 1688 29256 1752
rect 29272 1688 29336 1752
rect 29352 1688 29416 1752
rect 41376 1688 41440 1752
rect 41456 1688 41520 1752
rect 41536 1688 41600 1752
rect 41616 1688 41680 1752
rect 41696 1688 41760 1752
rect 41776 1688 41840 1752
rect 41856 1688 41920 1752
rect 41936 1688 42000 1752
rect 42016 1688 42080 1752
rect 42096 1688 42160 1752
rect 42176 1688 42240 1752
rect 42256 1688 42320 1752
rect 42336 1688 42400 1752
rect 42416 1688 42480 1752
rect 42496 1688 42560 1752
rect 42576 1688 42640 1752
rect 42656 1688 42720 1752
rect 42736 1688 42800 1752
rect 42816 1688 42880 1752
rect 42896 1688 42960 1752
rect 42976 1688 43040 1752
rect 43056 1688 43120 1752
rect 43136 1688 43200 1752
rect 43216 1688 43280 1752
rect 43296 1688 43360 1752
rect 43376 1688 43440 1752
rect 43456 1688 43520 1752
rect 43536 1688 43600 1752
rect 43616 1688 43680 1752
rect 43696 1688 43760 1752
rect 43776 1688 43840 1752
rect 43856 1688 43920 1752
rect 43936 1688 44000 1752
rect 44016 1688 44080 1752
rect 44096 1688 44160 1752
rect 44176 1688 44240 1752
rect 44256 1688 44320 1752
rect 44336 1688 44400 1752
rect 44416 1688 44480 1752
rect 44496 1688 44560 1752
rect 44576 1688 44640 1752
rect 44656 1688 44720 1752
rect 44736 1688 44800 1752
rect 44816 1688 44880 1752
rect 44896 1688 44960 1752
rect 44976 1688 45040 1752
rect 45056 1688 45120 1752
rect 45136 1688 45200 1752
rect 45216 1688 45280 1752
rect 45296 1688 45360 1752
rect 8 1608 72 1672
rect 88 1608 152 1672
rect 168 1608 232 1672
rect 248 1608 312 1672
rect 328 1608 392 1672
rect 408 1608 472 1672
rect 488 1608 552 1672
rect 568 1608 632 1672
rect 648 1608 712 1672
rect 728 1608 792 1672
rect 808 1608 872 1672
rect 888 1608 952 1672
rect 968 1608 1032 1672
rect 1048 1608 1112 1672
rect 1128 1608 1192 1672
rect 1208 1608 1272 1672
rect 1288 1608 1352 1672
rect 1368 1608 1432 1672
rect 1448 1608 1512 1672
rect 1528 1608 1592 1672
rect 1608 1608 1672 1672
rect 1688 1608 1752 1672
rect 1768 1608 1832 1672
rect 1848 1608 1912 1672
rect 1928 1608 1992 1672
rect 2008 1608 2072 1672
rect 2088 1608 2152 1672
rect 2168 1608 2232 1672
rect 2248 1608 2312 1672
rect 2328 1608 2392 1672
rect 2408 1608 2472 1672
rect 2488 1608 2552 1672
rect 2568 1608 2632 1672
rect 2648 1608 2712 1672
rect 2728 1608 2792 1672
rect 2808 1608 2872 1672
rect 2888 1608 2952 1672
rect 2968 1608 3032 1672
rect 3048 1608 3112 1672
rect 3128 1608 3192 1672
rect 3208 1608 3272 1672
rect 3288 1608 3352 1672
rect 3368 1608 3432 1672
rect 3448 1608 3512 1672
rect 3528 1608 3592 1672
rect 3608 1608 3672 1672
rect 3688 1608 3752 1672
rect 3768 1608 3832 1672
rect 3848 1608 3912 1672
rect 3928 1608 3992 1672
rect 19112 1608 19176 1672
rect 19192 1608 19256 1672
rect 19272 1608 19336 1672
rect 19352 1608 19416 1672
rect 29112 1608 29176 1672
rect 29192 1608 29256 1672
rect 29272 1608 29336 1672
rect 29352 1608 29416 1672
rect 41376 1608 41440 1672
rect 41456 1608 41520 1672
rect 41536 1608 41600 1672
rect 41616 1608 41680 1672
rect 41696 1608 41760 1672
rect 41776 1608 41840 1672
rect 41856 1608 41920 1672
rect 41936 1608 42000 1672
rect 42016 1608 42080 1672
rect 42096 1608 42160 1672
rect 42176 1608 42240 1672
rect 42256 1608 42320 1672
rect 42336 1608 42400 1672
rect 42416 1608 42480 1672
rect 42496 1608 42560 1672
rect 42576 1608 42640 1672
rect 42656 1608 42720 1672
rect 42736 1608 42800 1672
rect 42816 1608 42880 1672
rect 42896 1608 42960 1672
rect 42976 1608 43040 1672
rect 43056 1608 43120 1672
rect 43136 1608 43200 1672
rect 43216 1608 43280 1672
rect 43296 1608 43360 1672
rect 43376 1608 43440 1672
rect 43456 1608 43520 1672
rect 43536 1608 43600 1672
rect 43616 1608 43680 1672
rect 43696 1608 43760 1672
rect 43776 1608 43840 1672
rect 43856 1608 43920 1672
rect 43936 1608 44000 1672
rect 44016 1608 44080 1672
rect 44096 1608 44160 1672
rect 44176 1608 44240 1672
rect 44256 1608 44320 1672
rect 44336 1608 44400 1672
rect 44416 1608 44480 1672
rect 44496 1608 44560 1672
rect 44576 1608 44640 1672
rect 44656 1608 44720 1672
rect 44736 1608 44800 1672
rect 44816 1608 44880 1672
rect 44896 1608 44960 1672
rect 44976 1608 45040 1672
rect 45056 1608 45120 1672
rect 45136 1608 45200 1672
rect 45216 1608 45280 1672
rect 45296 1608 45360 1672
rect 8 1528 72 1592
rect 88 1528 152 1592
rect 168 1528 232 1592
rect 248 1528 312 1592
rect 328 1528 392 1592
rect 408 1528 472 1592
rect 488 1528 552 1592
rect 568 1528 632 1592
rect 648 1528 712 1592
rect 728 1528 792 1592
rect 808 1528 872 1592
rect 888 1528 952 1592
rect 968 1528 1032 1592
rect 1048 1528 1112 1592
rect 1128 1528 1192 1592
rect 1208 1528 1272 1592
rect 1288 1528 1352 1592
rect 1368 1528 1432 1592
rect 1448 1528 1512 1592
rect 1528 1528 1592 1592
rect 1608 1528 1672 1592
rect 1688 1528 1752 1592
rect 1768 1528 1832 1592
rect 1848 1528 1912 1592
rect 1928 1528 1992 1592
rect 2008 1528 2072 1592
rect 2088 1528 2152 1592
rect 2168 1528 2232 1592
rect 2248 1528 2312 1592
rect 2328 1528 2392 1592
rect 2408 1528 2472 1592
rect 2488 1528 2552 1592
rect 2568 1528 2632 1592
rect 2648 1528 2712 1592
rect 2728 1528 2792 1592
rect 2808 1528 2872 1592
rect 2888 1528 2952 1592
rect 2968 1528 3032 1592
rect 3048 1528 3112 1592
rect 3128 1528 3192 1592
rect 3208 1528 3272 1592
rect 3288 1528 3352 1592
rect 3368 1528 3432 1592
rect 3448 1528 3512 1592
rect 3528 1528 3592 1592
rect 3608 1528 3672 1592
rect 3688 1528 3752 1592
rect 3768 1528 3832 1592
rect 3848 1528 3912 1592
rect 3928 1528 3992 1592
rect 19112 1528 19176 1592
rect 19192 1528 19256 1592
rect 19272 1528 19336 1592
rect 19352 1528 19416 1592
rect 29112 1528 29176 1592
rect 29192 1528 29256 1592
rect 29272 1528 29336 1592
rect 29352 1528 29416 1592
rect 41376 1528 41440 1592
rect 41456 1528 41520 1592
rect 41536 1528 41600 1592
rect 41616 1528 41680 1592
rect 41696 1528 41760 1592
rect 41776 1528 41840 1592
rect 41856 1528 41920 1592
rect 41936 1528 42000 1592
rect 42016 1528 42080 1592
rect 42096 1528 42160 1592
rect 42176 1528 42240 1592
rect 42256 1528 42320 1592
rect 42336 1528 42400 1592
rect 42416 1528 42480 1592
rect 42496 1528 42560 1592
rect 42576 1528 42640 1592
rect 42656 1528 42720 1592
rect 42736 1528 42800 1592
rect 42816 1528 42880 1592
rect 42896 1528 42960 1592
rect 42976 1528 43040 1592
rect 43056 1528 43120 1592
rect 43136 1528 43200 1592
rect 43216 1528 43280 1592
rect 43296 1528 43360 1592
rect 43376 1528 43440 1592
rect 43456 1528 43520 1592
rect 43536 1528 43600 1592
rect 43616 1528 43680 1592
rect 43696 1528 43760 1592
rect 43776 1528 43840 1592
rect 43856 1528 43920 1592
rect 43936 1528 44000 1592
rect 44016 1528 44080 1592
rect 44096 1528 44160 1592
rect 44176 1528 44240 1592
rect 44256 1528 44320 1592
rect 44336 1528 44400 1592
rect 44416 1528 44480 1592
rect 44496 1528 44560 1592
rect 44576 1528 44640 1592
rect 44656 1528 44720 1592
rect 44736 1528 44800 1592
rect 44816 1528 44880 1592
rect 44896 1528 44960 1592
rect 44976 1528 45040 1592
rect 45056 1528 45120 1592
rect 45136 1528 45200 1592
rect 45216 1528 45280 1592
rect 45296 1528 45360 1592
rect 8 1448 72 1512
rect 88 1448 152 1512
rect 168 1448 232 1512
rect 248 1448 312 1512
rect 328 1448 392 1512
rect 408 1448 472 1512
rect 488 1448 552 1512
rect 568 1448 632 1512
rect 648 1448 712 1512
rect 728 1448 792 1512
rect 808 1448 872 1512
rect 888 1448 952 1512
rect 968 1448 1032 1512
rect 1048 1448 1112 1512
rect 1128 1448 1192 1512
rect 1208 1448 1272 1512
rect 1288 1448 1352 1512
rect 1368 1448 1432 1512
rect 1448 1448 1512 1512
rect 1528 1448 1592 1512
rect 1608 1448 1672 1512
rect 1688 1448 1752 1512
rect 1768 1448 1832 1512
rect 1848 1448 1912 1512
rect 1928 1448 1992 1512
rect 2008 1448 2072 1512
rect 2088 1448 2152 1512
rect 2168 1448 2232 1512
rect 2248 1448 2312 1512
rect 2328 1448 2392 1512
rect 2408 1448 2472 1512
rect 2488 1448 2552 1512
rect 2568 1448 2632 1512
rect 2648 1448 2712 1512
rect 2728 1448 2792 1512
rect 2808 1448 2872 1512
rect 2888 1448 2952 1512
rect 2968 1448 3032 1512
rect 3048 1448 3112 1512
rect 3128 1448 3192 1512
rect 3208 1448 3272 1512
rect 3288 1448 3352 1512
rect 3368 1448 3432 1512
rect 3448 1448 3512 1512
rect 3528 1448 3592 1512
rect 3608 1448 3672 1512
rect 3688 1448 3752 1512
rect 3768 1448 3832 1512
rect 3848 1448 3912 1512
rect 3928 1448 3992 1512
rect 19112 1448 19176 1512
rect 19192 1448 19256 1512
rect 19272 1448 19336 1512
rect 19352 1448 19416 1512
rect 29112 1448 29176 1512
rect 29192 1448 29256 1512
rect 29272 1448 29336 1512
rect 29352 1448 29416 1512
rect 41376 1448 41440 1512
rect 41456 1448 41520 1512
rect 41536 1448 41600 1512
rect 41616 1448 41680 1512
rect 41696 1448 41760 1512
rect 41776 1448 41840 1512
rect 41856 1448 41920 1512
rect 41936 1448 42000 1512
rect 42016 1448 42080 1512
rect 42096 1448 42160 1512
rect 42176 1448 42240 1512
rect 42256 1448 42320 1512
rect 42336 1448 42400 1512
rect 42416 1448 42480 1512
rect 42496 1448 42560 1512
rect 42576 1448 42640 1512
rect 42656 1448 42720 1512
rect 42736 1448 42800 1512
rect 42816 1448 42880 1512
rect 42896 1448 42960 1512
rect 42976 1448 43040 1512
rect 43056 1448 43120 1512
rect 43136 1448 43200 1512
rect 43216 1448 43280 1512
rect 43296 1448 43360 1512
rect 43376 1448 43440 1512
rect 43456 1448 43520 1512
rect 43536 1448 43600 1512
rect 43616 1448 43680 1512
rect 43696 1448 43760 1512
rect 43776 1448 43840 1512
rect 43856 1448 43920 1512
rect 43936 1448 44000 1512
rect 44016 1448 44080 1512
rect 44096 1448 44160 1512
rect 44176 1448 44240 1512
rect 44256 1448 44320 1512
rect 44336 1448 44400 1512
rect 44416 1448 44480 1512
rect 44496 1448 44560 1512
rect 44576 1448 44640 1512
rect 44656 1448 44720 1512
rect 44736 1448 44800 1512
rect 44816 1448 44880 1512
rect 44896 1448 44960 1512
rect 44976 1448 45040 1512
rect 45056 1448 45120 1512
rect 45136 1448 45200 1512
rect 45216 1448 45280 1512
rect 45296 1448 45360 1512
rect 8 1368 72 1432
rect 88 1368 152 1432
rect 168 1368 232 1432
rect 248 1368 312 1432
rect 328 1368 392 1432
rect 408 1368 472 1432
rect 488 1368 552 1432
rect 568 1368 632 1432
rect 648 1368 712 1432
rect 728 1368 792 1432
rect 808 1368 872 1432
rect 888 1368 952 1432
rect 968 1368 1032 1432
rect 1048 1368 1112 1432
rect 1128 1368 1192 1432
rect 1208 1368 1272 1432
rect 1288 1368 1352 1432
rect 1368 1368 1432 1432
rect 1448 1368 1512 1432
rect 1528 1368 1592 1432
rect 1608 1368 1672 1432
rect 1688 1368 1752 1432
rect 1768 1368 1832 1432
rect 1848 1368 1912 1432
rect 1928 1368 1992 1432
rect 2008 1368 2072 1432
rect 2088 1368 2152 1432
rect 2168 1368 2232 1432
rect 2248 1368 2312 1432
rect 2328 1368 2392 1432
rect 2408 1368 2472 1432
rect 2488 1368 2552 1432
rect 2568 1368 2632 1432
rect 2648 1368 2712 1432
rect 2728 1368 2792 1432
rect 2808 1368 2872 1432
rect 2888 1368 2952 1432
rect 2968 1368 3032 1432
rect 3048 1368 3112 1432
rect 3128 1368 3192 1432
rect 3208 1368 3272 1432
rect 3288 1368 3352 1432
rect 3368 1368 3432 1432
rect 3448 1368 3512 1432
rect 3528 1368 3592 1432
rect 3608 1368 3672 1432
rect 3688 1368 3752 1432
rect 3768 1368 3832 1432
rect 3848 1368 3912 1432
rect 3928 1368 3992 1432
rect 19112 1368 19176 1432
rect 19192 1368 19256 1432
rect 19272 1368 19336 1432
rect 19352 1368 19416 1432
rect 29112 1368 29176 1432
rect 29192 1368 29256 1432
rect 29272 1368 29336 1432
rect 29352 1368 29416 1432
rect 41376 1368 41440 1432
rect 41456 1368 41520 1432
rect 41536 1368 41600 1432
rect 41616 1368 41680 1432
rect 41696 1368 41760 1432
rect 41776 1368 41840 1432
rect 41856 1368 41920 1432
rect 41936 1368 42000 1432
rect 42016 1368 42080 1432
rect 42096 1368 42160 1432
rect 42176 1368 42240 1432
rect 42256 1368 42320 1432
rect 42336 1368 42400 1432
rect 42416 1368 42480 1432
rect 42496 1368 42560 1432
rect 42576 1368 42640 1432
rect 42656 1368 42720 1432
rect 42736 1368 42800 1432
rect 42816 1368 42880 1432
rect 42896 1368 42960 1432
rect 42976 1368 43040 1432
rect 43056 1368 43120 1432
rect 43136 1368 43200 1432
rect 43216 1368 43280 1432
rect 43296 1368 43360 1432
rect 43376 1368 43440 1432
rect 43456 1368 43520 1432
rect 43536 1368 43600 1432
rect 43616 1368 43680 1432
rect 43696 1368 43760 1432
rect 43776 1368 43840 1432
rect 43856 1368 43920 1432
rect 43936 1368 44000 1432
rect 44016 1368 44080 1432
rect 44096 1368 44160 1432
rect 44176 1368 44240 1432
rect 44256 1368 44320 1432
rect 44336 1368 44400 1432
rect 44416 1368 44480 1432
rect 44496 1368 44560 1432
rect 44576 1368 44640 1432
rect 44656 1368 44720 1432
rect 44736 1368 44800 1432
rect 44816 1368 44880 1432
rect 44896 1368 44960 1432
rect 44976 1368 45040 1432
rect 45056 1368 45120 1432
rect 45136 1368 45200 1432
rect 45216 1368 45280 1432
rect 45296 1368 45360 1432
rect 8 1288 72 1352
rect 88 1288 152 1352
rect 168 1288 232 1352
rect 248 1288 312 1352
rect 328 1288 392 1352
rect 408 1288 472 1352
rect 488 1288 552 1352
rect 568 1288 632 1352
rect 648 1288 712 1352
rect 728 1288 792 1352
rect 808 1288 872 1352
rect 888 1288 952 1352
rect 968 1288 1032 1352
rect 1048 1288 1112 1352
rect 1128 1288 1192 1352
rect 1208 1288 1272 1352
rect 1288 1288 1352 1352
rect 1368 1288 1432 1352
rect 1448 1288 1512 1352
rect 1528 1288 1592 1352
rect 1608 1288 1672 1352
rect 1688 1288 1752 1352
rect 1768 1288 1832 1352
rect 1848 1288 1912 1352
rect 1928 1288 1992 1352
rect 2008 1288 2072 1352
rect 2088 1288 2152 1352
rect 2168 1288 2232 1352
rect 2248 1288 2312 1352
rect 2328 1288 2392 1352
rect 2408 1288 2472 1352
rect 2488 1288 2552 1352
rect 2568 1288 2632 1352
rect 2648 1288 2712 1352
rect 2728 1288 2792 1352
rect 2808 1288 2872 1352
rect 2888 1288 2952 1352
rect 2968 1288 3032 1352
rect 3048 1288 3112 1352
rect 3128 1288 3192 1352
rect 3208 1288 3272 1352
rect 3288 1288 3352 1352
rect 3368 1288 3432 1352
rect 3448 1288 3512 1352
rect 3528 1288 3592 1352
rect 3608 1288 3672 1352
rect 3688 1288 3752 1352
rect 3768 1288 3832 1352
rect 3848 1288 3912 1352
rect 3928 1288 3992 1352
rect 19112 1288 19176 1352
rect 19192 1288 19256 1352
rect 19272 1288 19336 1352
rect 19352 1288 19416 1352
rect 29112 1288 29176 1352
rect 29192 1288 29256 1352
rect 29272 1288 29336 1352
rect 29352 1288 29416 1352
rect 41376 1288 41440 1352
rect 41456 1288 41520 1352
rect 41536 1288 41600 1352
rect 41616 1288 41680 1352
rect 41696 1288 41760 1352
rect 41776 1288 41840 1352
rect 41856 1288 41920 1352
rect 41936 1288 42000 1352
rect 42016 1288 42080 1352
rect 42096 1288 42160 1352
rect 42176 1288 42240 1352
rect 42256 1288 42320 1352
rect 42336 1288 42400 1352
rect 42416 1288 42480 1352
rect 42496 1288 42560 1352
rect 42576 1288 42640 1352
rect 42656 1288 42720 1352
rect 42736 1288 42800 1352
rect 42816 1288 42880 1352
rect 42896 1288 42960 1352
rect 42976 1288 43040 1352
rect 43056 1288 43120 1352
rect 43136 1288 43200 1352
rect 43216 1288 43280 1352
rect 43296 1288 43360 1352
rect 43376 1288 43440 1352
rect 43456 1288 43520 1352
rect 43536 1288 43600 1352
rect 43616 1288 43680 1352
rect 43696 1288 43760 1352
rect 43776 1288 43840 1352
rect 43856 1288 43920 1352
rect 43936 1288 44000 1352
rect 44016 1288 44080 1352
rect 44096 1288 44160 1352
rect 44176 1288 44240 1352
rect 44256 1288 44320 1352
rect 44336 1288 44400 1352
rect 44416 1288 44480 1352
rect 44496 1288 44560 1352
rect 44576 1288 44640 1352
rect 44656 1288 44720 1352
rect 44736 1288 44800 1352
rect 44816 1288 44880 1352
rect 44896 1288 44960 1352
rect 44976 1288 45040 1352
rect 45056 1288 45120 1352
rect 45136 1288 45200 1352
rect 45216 1288 45280 1352
rect 45296 1288 45360 1352
rect 8 1208 72 1272
rect 88 1208 152 1272
rect 168 1208 232 1272
rect 248 1208 312 1272
rect 328 1208 392 1272
rect 408 1208 472 1272
rect 488 1208 552 1272
rect 568 1208 632 1272
rect 648 1208 712 1272
rect 728 1208 792 1272
rect 808 1208 872 1272
rect 888 1208 952 1272
rect 968 1208 1032 1272
rect 1048 1208 1112 1272
rect 1128 1208 1192 1272
rect 1208 1208 1272 1272
rect 1288 1208 1352 1272
rect 1368 1208 1432 1272
rect 1448 1208 1512 1272
rect 1528 1208 1592 1272
rect 1608 1208 1672 1272
rect 1688 1208 1752 1272
rect 1768 1208 1832 1272
rect 1848 1208 1912 1272
rect 1928 1208 1992 1272
rect 2008 1208 2072 1272
rect 2088 1208 2152 1272
rect 2168 1208 2232 1272
rect 2248 1208 2312 1272
rect 2328 1208 2392 1272
rect 2408 1208 2472 1272
rect 2488 1208 2552 1272
rect 2568 1208 2632 1272
rect 2648 1208 2712 1272
rect 2728 1208 2792 1272
rect 2808 1208 2872 1272
rect 2888 1208 2952 1272
rect 2968 1208 3032 1272
rect 3048 1208 3112 1272
rect 3128 1208 3192 1272
rect 3208 1208 3272 1272
rect 3288 1208 3352 1272
rect 3368 1208 3432 1272
rect 3448 1208 3512 1272
rect 3528 1208 3592 1272
rect 3608 1208 3672 1272
rect 3688 1208 3752 1272
rect 3768 1208 3832 1272
rect 3848 1208 3912 1272
rect 3928 1208 3992 1272
rect 19112 1208 19176 1272
rect 19192 1208 19256 1272
rect 19272 1208 19336 1272
rect 19352 1208 19416 1272
rect 29112 1208 29176 1272
rect 29192 1208 29256 1272
rect 29272 1208 29336 1272
rect 29352 1208 29416 1272
rect 41376 1208 41440 1272
rect 41456 1208 41520 1272
rect 41536 1208 41600 1272
rect 41616 1208 41680 1272
rect 41696 1208 41760 1272
rect 41776 1208 41840 1272
rect 41856 1208 41920 1272
rect 41936 1208 42000 1272
rect 42016 1208 42080 1272
rect 42096 1208 42160 1272
rect 42176 1208 42240 1272
rect 42256 1208 42320 1272
rect 42336 1208 42400 1272
rect 42416 1208 42480 1272
rect 42496 1208 42560 1272
rect 42576 1208 42640 1272
rect 42656 1208 42720 1272
rect 42736 1208 42800 1272
rect 42816 1208 42880 1272
rect 42896 1208 42960 1272
rect 42976 1208 43040 1272
rect 43056 1208 43120 1272
rect 43136 1208 43200 1272
rect 43216 1208 43280 1272
rect 43296 1208 43360 1272
rect 43376 1208 43440 1272
rect 43456 1208 43520 1272
rect 43536 1208 43600 1272
rect 43616 1208 43680 1272
rect 43696 1208 43760 1272
rect 43776 1208 43840 1272
rect 43856 1208 43920 1272
rect 43936 1208 44000 1272
rect 44016 1208 44080 1272
rect 44096 1208 44160 1272
rect 44176 1208 44240 1272
rect 44256 1208 44320 1272
rect 44336 1208 44400 1272
rect 44416 1208 44480 1272
rect 44496 1208 44560 1272
rect 44576 1208 44640 1272
rect 44656 1208 44720 1272
rect 44736 1208 44800 1272
rect 44816 1208 44880 1272
rect 44896 1208 44960 1272
rect 44976 1208 45040 1272
rect 45056 1208 45120 1272
rect 45136 1208 45200 1272
rect 45216 1208 45280 1272
rect 45296 1208 45360 1272
rect 8 1128 72 1192
rect 88 1128 152 1192
rect 168 1128 232 1192
rect 248 1128 312 1192
rect 328 1128 392 1192
rect 408 1128 472 1192
rect 488 1128 552 1192
rect 568 1128 632 1192
rect 648 1128 712 1192
rect 728 1128 792 1192
rect 808 1128 872 1192
rect 888 1128 952 1192
rect 968 1128 1032 1192
rect 1048 1128 1112 1192
rect 1128 1128 1192 1192
rect 1208 1128 1272 1192
rect 1288 1128 1352 1192
rect 1368 1128 1432 1192
rect 1448 1128 1512 1192
rect 1528 1128 1592 1192
rect 1608 1128 1672 1192
rect 1688 1128 1752 1192
rect 1768 1128 1832 1192
rect 1848 1128 1912 1192
rect 1928 1128 1992 1192
rect 2008 1128 2072 1192
rect 2088 1128 2152 1192
rect 2168 1128 2232 1192
rect 2248 1128 2312 1192
rect 2328 1128 2392 1192
rect 2408 1128 2472 1192
rect 2488 1128 2552 1192
rect 2568 1128 2632 1192
rect 2648 1128 2712 1192
rect 2728 1128 2792 1192
rect 2808 1128 2872 1192
rect 2888 1128 2952 1192
rect 2968 1128 3032 1192
rect 3048 1128 3112 1192
rect 3128 1128 3192 1192
rect 3208 1128 3272 1192
rect 3288 1128 3352 1192
rect 3368 1128 3432 1192
rect 3448 1128 3512 1192
rect 3528 1128 3592 1192
rect 3608 1128 3672 1192
rect 3688 1128 3752 1192
rect 3768 1128 3832 1192
rect 3848 1128 3912 1192
rect 3928 1128 3992 1192
rect 19112 1128 19176 1192
rect 19192 1128 19256 1192
rect 19272 1128 19336 1192
rect 19352 1128 19416 1192
rect 29112 1128 29176 1192
rect 29192 1128 29256 1192
rect 29272 1128 29336 1192
rect 29352 1128 29416 1192
rect 41376 1128 41440 1192
rect 41456 1128 41520 1192
rect 41536 1128 41600 1192
rect 41616 1128 41680 1192
rect 41696 1128 41760 1192
rect 41776 1128 41840 1192
rect 41856 1128 41920 1192
rect 41936 1128 42000 1192
rect 42016 1128 42080 1192
rect 42096 1128 42160 1192
rect 42176 1128 42240 1192
rect 42256 1128 42320 1192
rect 42336 1128 42400 1192
rect 42416 1128 42480 1192
rect 42496 1128 42560 1192
rect 42576 1128 42640 1192
rect 42656 1128 42720 1192
rect 42736 1128 42800 1192
rect 42816 1128 42880 1192
rect 42896 1128 42960 1192
rect 42976 1128 43040 1192
rect 43056 1128 43120 1192
rect 43136 1128 43200 1192
rect 43216 1128 43280 1192
rect 43296 1128 43360 1192
rect 43376 1128 43440 1192
rect 43456 1128 43520 1192
rect 43536 1128 43600 1192
rect 43616 1128 43680 1192
rect 43696 1128 43760 1192
rect 43776 1128 43840 1192
rect 43856 1128 43920 1192
rect 43936 1128 44000 1192
rect 44016 1128 44080 1192
rect 44096 1128 44160 1192
rect 44176 1128 44240 1192
rect 44256 1128 44320 1192
rect 44336 1128 44400 1192
rect 44416 1128 44480 1192
rect 44496 1128 44560 1192
rect 44576 1128 44640 1192
rect 44656 1128 44720 1192
rect 44736 1128 44800 1192
rect 44816 1128 44880 1192
rect 44896 1128 44960 1192
rect 44976 1128 45040 1192
rect 45056 1128 45120 1192
rect 45136 1128 45200 1192
rect 45216 1128 45280 1192
rect 45296 1128 45360 1192
rect 8 1048 72 1112
rect 88 1048 152 1112
rect 168 1048 232 1112
rect 248 1048 312 1112
rect 328 1048 392 1112
rect 408 1048 472 1112
rect 488 1048 552 1112
rect 568 1048 632 1112
rect 648 1048 712 1112
rect 728 1048 792 1112
rect 808 1048 872 1112
rect 888 1048 952 1112
rect 968 1048 1032 1112
rect 1048 1048 1112 1112
rect 1128 1048 1192 1112
rect 1208 1048 1272 1112
rect 1288 1048 1352 1112
rect 1368 1048 1432 1112
rect 1448 1048 1512 1112
rect 1528 1048 1592 1112
rect 1608 1048 1672 1112
rect 1688 1048 1752 1112
rect 1768 1048 1832 1112
rect 1848 1048 1912 1112
rect 1928 1048 1992 1112
rect 2008 1048 2072 1112
rect 2088 1048 2152 1112
rect 2168 1048 2232 1112
rect 2248 1048 2312 1112
rect 2328 1048 2392 1112
rect 2408 1048 2472 1112
rect 2488 1048 2552 1112
rect 2568 1048 2632 1112
rect 2648 1048 2712 1112
rect 2728 1048 2792 1112
rect 2808 1048 2872 1112
rect 2888 1048 2952 1112
rect 2968 1048 3032 1112
rect 3048 1048 3112 1112
rect 3128 1048 3192 1112
rect 3208 1048 3272 1112
rect 3288 1048 3352 1112
rect 3368 1048 3432 1112
rect 3448 1048 3512 1112
rect 3528 1048 3592 1112
rect 3608 1048 3672 1112
rect 3688 1048 3752 1112
rect 3768 1048 3832 1112
rect 3848 1048 3912 1112
rect 3928 1048 3992 1112
rect 19112 1048 19176 1112
rect 19192 1048 19256 1112
rect 19272 1048 19336 1112
rect 19352 1048 19416 1112
rect 29112 1048 29176 1112
rect 29192 1048 29256 1112
rect 29272 1048 29336 1112
rect 29352 1048 29416 1112
rect 41376 1048 41440 1112
rect 41456 1048 41520 1112
rect 41536 1048 41600 1112
rect 41616 1048 41680 1112
rect 41696 1048 41760 1112
rect 41776 1048 41840 1112
rect 41856 1048 41920 1112
rect 41936 1048 42000 1112
rect 42016 1048 42080 1112
rect 42096 1048 42160 1112
rect 42176 1048 42240 1112
rect 42256 1048 42320 1112
rect 42336 1048 42400 1112
rect 42416 1048 42480 1112
rect 42496 1048 42560 1112
rect 42576 1048 42640 1112
rect 42656 1048 42720 1112
rect 42736 1048 42800 1112
rect 42816 1048 42880 1112
rect 42896 1048 42960 1112
rect 42976 1048 43040 1112
rect 43056 1048 43120 1112
rect 43136 1048 43200 1112
rect 43216 1048 43280 1112
rect 43296 1048 43360 1112
rect 43376 1048 43440 1112
rect 43456 1048 43520 1112
rect 43536 1048 43600 1112
rect 43616 1048 43680 1112
rect 43696 1048 43760 1112
rect 43776 1048 43840 1112
rect 43856 1048 43920 1112
rect 43936 1048 44000 1112
rect 44016 1048 44080 1112
rect 44096 1048 44160 1112
rect 44176 1048 44240 1112
rect 44256 1048 44320 1112
rect 44336 1048 44400 1112
rect 44416 1048 44480 1112
rect 44496 1048 44560 1112
rect 44576 1048 44640 1112
rect 44656 1048 44720 1112
rect 44736 1048 44800 1112
rect 44816 1048 44880 1112
rect 44896 1048 44960 1112
rect 44976 1048 45040 1112
rect 45056 1048 45120 1112
rect 45136 1048 45200 1112
rect 45216 1048 45280 1112
rect 45296 1048 45360 1112
rect 8 968 72 1032
rect 88 968 152 1032
rect 168 968 232 1032
rect 248 968 312 1032
rect 328 968 392 1032
rect 408 968 472 1032
rect 488 968 552 1032
rect 568 968 632 1032
rect 648 968 712 1032
rect 728 968 792 1032
rect 808 968 872 1032
rect 888 968 952 1032
rect 968 968 1032 1032
rect 1048 968 1112 1032
rect 1128 968 1192 1032
rect 1208 968 1272 1032
rect 1288 968 1352 1032
rect 1368 968 1432 1032
rect 1448 968 1512 1032
rect 1528 968 1592 1032
rect 1608 968 1672 1032
rect 1688 968 1752 1032
rect 1768 968 1832 1032
rect 1848 968 1912 1032
rect 1928 968 1992 1032
rect 2008 968 2072 1032
rect 2088 968 2152 1032
rect 2168 968 2232 1032
rect 2248 968 2312 1032
rect 2328 968 2392 1032
rect 2408 968 2472 1032
rect 2488 968 2552 1032
rect 2568 968 2632 1032
rect 2648 968 2712 1032
rect 2728 968 2792 1032
rect 2808 968 2872 1032
rect 2888 968 2952 1032
rect 2968 968 3032 1032
rect 3048 968 3112 1032
rect 3128 968 3192 1032
rect 3208 968 3272 1032
rect 3288 968 3352 1032
rect 3368 968 3432 1032
rect 3448 968 3512 1032
rect 3528 968 3592 1032
rect 3608 968 3672 1032
rect 3688 968 3752 1032
rect 3768 968 3832 1032
rect 3848 968 3912 1032
rect 3928 968 3992 1032
rect 19112 968 19176 1032
rect 19192 968 19256 1032
rect 19272 968 19336 1032
rect 19352 968 19416 1032
rect 29112 968 29176 1032
rect 29192 968 29256 1032
rect 29272 968 29336 1032
rect 29352 968 29416 1032
rect 41376 968 41440 1032
rect 41456 968 41520 1032
rect 41536 968 41600 1032
rect 41616 968 41680 1032
rect 41696 968 41760 1032
rect 41776 968 41840 1032
rect 41856 968 41920 1032
rect 41936 968 42000 1032
rect 42016 968 42080 1032
rect 42096 968 42160 1032
rect 42176 968 42240 1032
rect 42256 968 42320 1032
rect 42336 968 42400 1032
rect 42416 968 42480 1032
rect 42496 968 42560 1032
rect 42576 968 42640 1032
rect 42656 968 42720 1032
rect 42736 968 42800 1032
rect 42816 968 42880 1032
rect 42896 968 42960 1032
rect 42976 968 43040 1032
rect 43056 968 43120 1032
rect 43136 968 43200 1032
rect 43216 968 43280 1032
rect 43296 968 43360 1032
rect 43376 968 43440 1032
rect 43456 968 43520 1032
rect 43536 968 43600 1032
rect 43616 968 43680 1032
rect 43696 968 43760 1032
rect 43776 968 43840 1032
rect 43856 968 43920 1032
rect 43936 968 44000 1032
rect 44016 968 44080 1032
rect 44096 968 44160 1032
rect 44176 968 44240 1032
rect 44256 968 44320 1032
rect 44336 968 44400 1032
rect 44416 968 44480 1032
rect 44496 968 44560 1032
rect 44576 968 44640 1032
rect 44656 968 44720 1032
rect 44736 968 44800 1032
rect 44816 968 44880 1032
rect 44896 968 44960 1032
rect 44976 968 45040 1032
rect 45056 968 45120 1032
rect 45136 968 45200 1032
rect 45216 968 45280 1032
rect 45296 968 45360 1032
rect 8 888 72 952
rect 88 888 152 952
rect 168 888 232 952
rect 248 888 312 952
rect 328 888 392 952
rect 408 888 472 952
rect 488 888 552 952
rect 568 888 632 952
rect 648 888 712 952
rect 728 888 792 952
rect 808 888 872 952
rect 888 888 952 952
rect 968 888 1032 952
rect 1048 888 1112 952
rect 1128 888 1192 952
rect 1208 888 1272 952
rect 1288 888 1352 952
rect 1368 888 1432 952
rect 1448 888 1512 952
rect 1528 888 1592 952
rect 1608 888 1672 952
rect 1688 888 1752 952
rect 1768 888 1832 952
rect 1848 888 1912 952
rect 1928 888 1992 952
rect 2008 888 2072 952
rect 2088 888 2152 952
rect 2168 888 2232 952
rect 2248 888 2312 952
rect 2328 888 2392 952
rect 2408 888 2472 952
rect 2488 888 2552 952
rect 2568 888 2632 952
rect 2648 888 2712 952
rect 2728 888 2792 952
rect 2808 888 2872 952
rect 2888 888 2952 952
rect 2968 888 3032 952
rect 3048 888 3112 952
rect 3128 888 3192 952
rect 3208 888 3272 952
rect 3288 888 3352 952
rect 3368 888 3432 952
rect 3448 888 3512 952
rect 3528 888 3592 952
rect 3608 888 3672 952
rect 3688 888 3752 952
rect 3768 888 3832 952
rect 3848 888 3912 952
rect 3928 888 3992 952
rect 19112 888 19176 952
rect 19192 888 19256 952
rect 19272 888 19336 952
rect 19352 888 19416 952
rect 29112 888 29176 952
rect 29192 888 29256 952
rect 29272 888 29336 952
rect 29352 888 29416 952
rect 41376 888 41440 952
rect 41456 888 41520 952
rect 41536 888 41600 952
rect 41616 888 41680 952
rect 41696 888 41760 952
rect 41776 888 41840 952
rect 41856 888 41920 952
rect 41936 888 42000 952
rect 42016 888 42080 952
rect 42096 888 42160 952
rect 42176 888 42240 952
rect 42256 888 42320 952
rect 42336 888 42400 952
rect 42416 888 42480 952
rect 42496 888 42560 952
rect 42576 888 42640 952
rect 42656 888 42720 952
rect 42736 888 42800 952
rect 42816 888 42880 952
rect 42896 888 42960 952
rect 42976 888 43040 952
rect 43056 888 43120 952
rect 43136 888 43200 952
rect 43216 888 43280 952
rect 43296 888 43360 952
rect 43376 888 43440 952
rect 43456 888 43520 952
rect 43536 888 43600 952
rect 43616 888 43680 952
rect 43696 888 43760 952
rect 43776 888 43840 952
rect 43856 888 43920 952
rect 43936 888 44000 952
rect 44016 888 44080 952
rect 44096 888 44160 952
rect 44176 888 44240 952
rect 44256 888 44320 952
rect 44336 888 44400 952
rect 44416 888 44480 952
rect 44496 888 44560 952
rect 44576 888 44640 952
rect 44656 888 44720 952
rect 44736 888 44800 952
rect 44816 888 44880 952
rect 44896 888 44960 952
rect 44976 888 45040 952
rect 45056 888 45120 952
rect 45136 888 45200 952
rect 45216 888 45280 952
rect 45296 888 45360 952
rect 8 808 72 872
rect 88 808 152 872
rect 168 808 232 872
rect 248 808 312 872
rect 328 808 392 872
rect 408 808 472 872
rect 488 808 552 872
rect 568 808 632 872
rect 648 808 712 872
rect 728 808 792 872
rect 808 808 872 872
rect 888 808 952 872
rect 968 808 1032 872
rect 1048 808 1112 872
rect 1128 808 1192 872
rect 1208 808 1272 872
rect 1288 808 1352 872
rect 1368 808 1432 872
rect 1448 808 1512 872
rect 1528 808 1592 872
rect 1608 808 1672 872
rect 1688 808 1752 872
rect 1768 808 1832 872
rect 1848 808 1912 872
rect 1928 808 1992 872
rect 2008 808 2072 872
rect 2088 808 2152 872
rect 2168 808 2232 872
rect 2248 808 2312 872
rect 2328 808 2392 872
rect 2408 808 2472 872
rect 2488 808 2552 872
rect 2568 808 2632 872
rect 2648 808 2712 872
rect 2728 808 2792 872
rect 2808 808 2872 872
rect 2888 808 2952 872
rect 2968 808 3032 872
rect 3048 808 3112 872
rect 3128 808 3192 872
rect 3208 808 3272 872
rect 3288 808 3352 872
rect 3368 808 3432 872
rect 3448 808 3512 872
rect 3528 808 3592 872
rect 3608 808 3672 872
rect 3688 808 3752 872
rect 3768 808 3832 872
rect 3848 808 3912 872
rect 3928 808 3992 872
rect 19112 808 19176 872
rect 19192 808 19256 872
rect 19272 808 19336 872
rect 19352 808 19416 872
rect 29112 808 29176 872
rect 29192 808 29256 872
rect 29272 808 29336 872
rect 29352 808 29416 872
rect 41376 808 41440 872
rect 41456 808 41520 872
rect 41536 808 41600 872
rect 41616 808 41680 872
rect 41696 808 41760 872
rect 41776 808 41840 872
rect 41856 808 41920 872
rect 41936 808 42000 872
rect 42016 808 42080 872
rect 42096 808 42160 872
rect 42176 808 42240 872
rect 42256 808 42320 872
rect 42336 808 42400 872
rect 42416 808 42480 872
rect 42496 808 42560 872
rect 42576 808 42640 872
rect 42656 808 42720 872
rect 42736 808 42800 872
rect 42816 808 42880 872
rect 42896 808 42960 872
rect 42976 808 43040 872
rect 43056 808 43120 872
rect 43136 808 43200 872
rect 43216 808 43280 872
rect 43296 808 43360 872
rect 43376 808 43440 872
rect 43456 808 43520 872
rect 43536 808 43600 872
rect 43616 808 43680 872
rect 43696 808 43760 872
rect 43776 808 43840 872
rect 43856 808 43920 872
rect 43936 808 44000 872
rect 44016 808 44080 872
rect 44096 808 44160 872
rect 44176 808 44240 872
rect 44256 808 44320 872
rect 44336 808 44400 872
rect 44416 808 44480 872
rect 44496 808 44560 872
rect 44576 808 44640 872
rect 44656 808 44720 872
rect 44736 808 44800 872
rect 44816 808 44880 872
rect 44896 808 44960 872
rect 44976 808 45040 872
rect 45056 808 45120 872
rect 45136 808 45200 872
rect 45216 808 45280 872
rect 45296 808 45360 872
rect 8 728 72 792
rect 88 728 152 792
rect 168 728 232 792
rect 248 728 312 792
rect 328 728 392 792
rect 408 728 472 792
rect 488 728 552 792
rect 568 728 632 792
rect 648 728 712 792
rect 728 728 792 792
rect 808 728 872 792
rect 888 728 952 792
rect 968 728 1032 792
rect 1048 728 1112 792
rect 1128 728 1192 792
rect 1208 728 1272 792
rect 1288 728 1352 792
rect 1368 728 1432 792
rect 1448 728 1512 792
rect 1528 728 1592 792
rect 1608 728 1672 792
rect 1688 728 1752 792
rect 1768 728 1832 792
rect 1848 728 1912 792
rect 1928 728 1992 792
rect 2008 728 2072 792
rect 2088 728 2152 792
rect 2168 728 2232 792
rect 2248 728 2312 792
rect 2328 728 2392 792
rect 2408 728 2472 792
rect 2488 728 2552 792
rect 2568 728 2632 792
rect 2648 728 2712 792
rect 2728 728 2792 792
rect 2808 728 2872 792
rect 2888 728 2952 792
rect 2968 728 3032 792
rect 3048 728 3112 792
rect 3128 728 3192 792
rect 3208 728 3272 792
rect 3288 728 3352 792
rect 3368 728 3432 792
rect 3448 728 3512 792
rect 3528 728 3592 792
rect 3608 728 3672 792
rect 3688 728 3752 792
rect 3768 728 3832 792
rect 3848 728 3912 792
rect 3928 728 3992 792
rect 19112 728 19176 792
rect 19192 728 19256 792
rect 19272 728 19336 792
rect 19352 728 19416 792
rect 29112 728 29176 792
rect 29192 728 29256 792
rect 29272 728 29336 792
rect 29352 728 29416 792
rect 41376 728 41440 792
rect 41456 728 41520 792
rect 41536 728 41600 792
rect 41616 728 41680 792
rect 41696 728 41760 792
rect 41776 728 41840 792
rect 41856 728 41920 792
rect 41936 728 42000 792
rect 42016 728 42080 792
rect 42096 728 42160 792
rect 42176 728 42240 792
rect 42256 728 42320 792
rect 42336 728 42400 792
rect 42416 728 42480 792
rect 42496 728 42560 792
rect 42576 728 42640 792
rect 42656 728 42720 792
rect 42736 728 42800 792
rect 42816 728 42880 792
rect 42896 728 42960 792
rect 42976 728 43040 792
rect 43056 728 43120 792
rect 43136 728 43200 792
rect 43216 728 43280 792
rect 43296 728 43360 792
rect 43376 728 43440 792
rect 43456 728 43520 792
rect 43536 728 43600 792
rect 43616 728 43680 792
rect 43696 728 43760 792
rect 43776 728 43840 792
rect 43856 728 43920 792
rect 43936 728 44000 792
rect 44016 728 44080 792
rect 44096 728 44160 792
rect 44176 728 44240 792
rect 44256 728 44320 792
rect 44336 728 44400 792
rect 44416 728 44480 792
rect 44496 728 44560 792
rect 44576 728 44640 792
rect 44656 728 44720 792
rect 44736 728 44800 792
rect 44816 728 44880 792
rect 44896 728 44960 792
rect 44976 728 45040 792
rect 45056 728 45120 792
rect 45136 728 45200 792
rect 45216 728 45280 792
rect 45296 728 45360 792
rect 8 648 72 712
rect 88 648 152 712
rect 168 648 232 712
rect 248 648 312 712
rect 328 648 392 712
rect 408 648 472 712
rect 488 648 552 712
rect 568 648 632 712
rect 648 648 712 712
rect 728 648 792 712
rect 808 648 872 712
rect 888 648 952 712
rect 968 648 1032 712
rect 1048 648 1112 712
rect 1128 648 1192 712
rect 1208 648 1272 712
rect 1288 648 1352 712
rect 1368 648 1432 712
rect 1448 648 1512 712
rect 1528 648 1592 712
rect 1608 648 1672 712
rect 1688 648 1752 712
rect 1768 648 1832 712
rect 1848 648 1912 712
rect 1928 648 1992 712
rect 2008 648 2072 712
rect 2088 648 2152 712
rect 2168 648 2232 712
rect 2248 648 2312 712
rect 2328 648 2392 712
rect 2408 648 2472 712
rect 2488 648 2552 712
rect 2568 648 2632 712
rect 2648 648 2712 712
rect 2728 648 2792 712
rect 2808 648 2872 712
rect 2888 648 2952 712
rect 2968 648 3032 712
rect 3048 648 3112 712
rect 3128 648 3192 712
rect 3208 648 3272 712
rect 3288 648 3352 712
rect 3368 648 3432 712
rect 3448 648 3512 712
rect 3528 648 3592 712
rect 3608 648 3672 712
rect 3688 648 3752 712
rect 3768 648 3832 712
rect 3848 648 3912 712
rect 3928 648 3992 712
rect 19112 648 19176 712
rect 19192 648 19256 712
rect 19272 648 19336 712
rect 19352 648 19416 712
rect 29112 648 29176 712
rect 29192 648 29256 712
rect 29272 648 29336 712
rect 29352 648 29416 712
rect 41376 648 41440 712
rect 41456 648 41520 712
rect 41536 648 41600 712
rect 41616 648 41680 712
rect 41696 648 41760 712
rect 41776 648 41840 712
rect 41856 648 41920 712
rect 41936 648 42000 712
rect 42016 648 42080 712
rect 42096 648 42160 712
rect 42176 648 42240 712
rect 42256 648 42320 712
rect 42336 648 42400 712
rect 42416 648 42480 712
rect 42496 648 42560 712
rect 42576 648 42640 712
rect 42656 648 42720 712
rect 42736 648 42800 712
rect 42816 648 42880 712
rect 42896 648 42960 712
rect 42976 648 43040 712
rect 43056 648 43120 712
rect 43136 648 43200 712
rect 43216 648 43280 712
rect 43296 648 43360 712
rect 43376 648 43440 712
rect 43456 648 43520 712
rect 43536 648 43600 712
rect 43616 648 43680 712
rect 43696 648 43760 712
rect 43776 648 43840 712
rect 43856 648 43920 712
rect 43936 648 44000 712
rect 44016 648 44080 712
rect 44096 648 44160 712
rect 44176 648 44240 712
rect 44256 648 44320 712
rect 44336 648 44400 712
rect 44416 648 44480 712
rect 44496 648 44560 712
rect 44576 648 44640 712
rect 44656 648 44720 712
rect 44736 648 44800 712
rect 44816 648 44880 712
rect 44896 648 44960 712
rect 44976 648 45040 712
rect 45056 648 45120 712
rect 45136 648 45200 712
rect 45216 648 45280 712
rect 45296 648 45360 712
rect 8 568 72 632
rect 88 568 152 632
rect 168 568 232 632
rect 248 568 312 632
rect 328 568 392 632
rect 408 568 472 632
rect 488 568 552 632
rect 568 568 632 632
rect 648 568 712 632
rect 728 568 792 632
rect 808 568 872 632
rect 888 568 952 632
rect 968 568 1032 632
rect 1048 568 1112 632
rect 1128 568 1192 632
rect 1208 568 1272 632
rect 1288 568 1352 632
rect 1368 568 1432 632
rect 1448 568 1512 632
rect 1528 568 1592 632
rect 1608 568 1672 632
rect 1688 568 1752 632
rect 1768 568 1832 632
rect 1848 568 1912 632
rect 1928 568 1992 632
rect 2008 568 2072 632
rect 2088 568 2152 632
rect 2168 568 2232 632
rect 2248 568 2312 632
rect 2328 568 2392 632
rect 2408 568 2472 632
rect 2488 568 2552 632
rect 2568 568 2632 632
rect 2648 568 2712 632
rect 2728 568 2792 632
rect 2808 568 2872 632
rect 2888 568 2952 632
rect 2968 568 3032 632
rect 3048 568 3112 632
rect 3128 568 3192 632
rect 3208 568 3272 632
rect 3288 568 3352 632
rect 3368 568 3432 632
rect 3448 568 3512 632
rect 3528 568 3592 632
rect 3608 568 3672 632
rect 3688 568 3752 632
rect 3768 568 3832 632
rect 3848 568 3912 632
rect 3928 568 3992 632
rect 19112 568 19176 632
rect 19192 568 19256 632
rect 19272 568 19336 632
rect 19352 568 19416 632
rect 29112 568 29176 632
rect 29192 568 29256 632
rect 29272 568 29336 632
rect 29352 568 29416 632
rect 41376 568 41440 632
rect 41456 568 41520 632
rect 41536 568 41600 632
rect 41616 568 41680 632
rect 41696 568 41760 632
rect 41776 568 41840 632
rect 41856 568 41920 632
rect 41936 568 42000 632
rect 42016 568 42080 632
rect 42096 568 42160 632
rect 42176 568 42240 632
rect 42256 568 42320 632
rect 42336 568 42400 632
rect 42416 568 42480 632
rect 42496 568 42560 632
rect 42576 568 42640 632
rect 42656 568 42720 632
rect 42736 568 42800 632
rect 42816 568 42880 632
rect 42896 568 42960 632
rect 42976 568 43040 632
rect 43056 568 43120 632
rect 43136 568 43200 632
rect 43216 568 43280 632
rect 43296 568 43360 632
rect 43376 568 43440 632
rect 43456 568 43520 632
rect 43536 568 43600 632
rect 43616 568 43680 632
rect 43696 568 43760 632
rect 43776 568 43840 632
rect 43856 568 43920 632
rect 43936 568 44000 632
rect 44016 568 44080 632
rect 44096 568 44160 632
rect 44176 568 44240 632
rect 44256 568 44320 632
rect 44336 568 44400 632
rect 44416 568 44480 632
rect 44496 568 44560 632
rect 44576 568 44640 632
rect 44656 568 44720 632
rect 44736 568 44800 632
rect 44816 568 44880 632
rect 44896 568 44960 632
rect 44976 568 45040 632
rect 45056 568 45120 632
rect 45136 568 45200 632
rect 45216 568 45280 632
rect 45296 568 45360 632
rect 8 488 72 552
rect 88 488 152 552
rect 168 488 232 552
rect 248 488 312 552
rect 328 488 392 552
rect 408 488 472 552
rect 488 488 552 552
rect 568 488 632 552
rect 648 488 712 552
rect 728 488 792 552
rect 808 488 872 552
rect 888 488 952 552
rect 968 488 1032 552
rect 1048 488 1112 552
rect 1128 488 1192 552
rect 1208 488 1272 552
rect 1288 488 1352 552
rect 1368 488 1432 552
rect 1448 488 1512 552
rect 1528 488 1592 552
rect 1608 488 1672 552
rect 1688 488 1752 552
rect 1768 488 1832 552
rect 1848 488 1912 552
rect 1928 488 1992 552
rect 2008 488 2072 552
rect 2088 488 2152 552
rect 2168 488 2232 552
rect 2248 488 2312 552
rect 2328 488 2392 552
rect 2408 488 2472 552
rect 2488 488 2552 552
rect 2568 488 2632 552
rect 2648 488 2712 552
rect 2728 488 2792 552
rect 2808 488 2872 552
rect 2888 488 2952 552
rect 2968 488 3032 552
rect 3048 488 3112 552
rect 3128 488 3192 552
rect 3208 488 3272 552
rect 3288 488 3352 552
rect 3368 488 3432 552
rect 3448 488 3512 552
rect 3528 488 3592 552
rect 3608 488 3672 552
rect 3688 488 3752 552
rect 3768 488 3832 552
rect 3848 488 3912 552
rect 3928 488 3992 552
rect 19112 488 19176 552
rect 19192 488 19256 552
rect 19272 488 19336 552
rect 19352 488 19416 552
rect 29112 488 29176 552
rect 29192 488 29256 552
rect 29272 488 29336 552
rect 29352 488 29416 552
rect 41376 488 41440 552
rect 41456 488 41520 552
rect 41536 488 41600 552
rect 41616 488 41680 552
rect 41696 488 41760 552
rect 41776 488 41840 552
rect 41856 488 41920 552
rect 41936 488 42000 552
rect 42016 488 42080 552
rect 42096 488 42160 552
rect 42176 488 42240 552
rect 42256 488 42320 552
rect 42336 488 42400 552
rect 42416 488 42480 552
rect 42496 488 42560 552
rect 42576 488 42640 552
rect 42656 488 42720 552
rect 42736 488 42800 552
rect 42816 488 42880 552
rect 42896 488 42960 552
rect 42976 488 43040 552
rect 43056 488 43120 552
rect 43136 488 43200 552
rect 43216 488 43280 552
rect 43296 488 43360 552
rect 43376 488 43440 552
rect 43456 488 43520 552
rect 43536 488 43600 552
rect 43616 488 43680 552
rect 43696 488 43760 552
rect 43776 488 43840 552
rect 43856 488 43920 552
rect 43936 488 44000 552
rect 44016 488 44080 552
rect 44096 488 44160 552
rect 44176 488 44240 552
rect 44256 488 44320 552
rect 44336 488 44400 552
rect 44416 488 44480 552
rect 44496 488 44560 552
rect 44576 488 44640 552
rect 44656 488 44720 552
rect 44736 488 44800 552
rect 44816 488 44880 552
rect 44896 488 44960 552
rect 44976 488 45040 552
rect 45056 488 45120 552
rect 45136 488 45200 552
rect 45216 488 45280 552
rect 45296 488 45360 552
rect 8 408 72 472
rect 88 408 152 472
rect 168 408 232 472
rect 248 408 312 472
rect 328 408 392 472
rect 408 408 472 472
rect 488 408 552 472
rect 568 408 632 472
rect 648 408 712 472
rect 728 408 792 472
rect 808 408 872 472
rect 888 408 952 472
rect 968 408 1032 472
rect 1048 408 1112 472
rect 1128 408 1192 472
rect 1208 408 1272 472
rect 1288 408 1352 472
rect 1368 408 1432 472
rect 1448 408 1512 472
rect 1528 408 1592 472
rect 1608 408 1672 472
rect 1688 408 1752 472
rect 1768 408 1832 472
rect 1848 408 1912 472
rect 1928 408 1992 472
rect 2008 408 2072 472
rect 2088 408 2152 472
rect 2168 408 2232 472
rect 2248 408 2312 472
rect 2328 408 2392 472
rect 2408 408 2472 472
rect 2488 408 2552 472
rect 2568 408 2632 472
rect 2648 408 2712 472
rect 2728 408 2792 472
rect 2808 408 2872 472
rect 2888 408 2952 472
rect 2968 408 3032 472
rect 3048 408 3112 472
rect 3128 408 3192 472
rect 3208 408 3272 472
rect 3288 408 3352 472
rect 3368 408 3432 472
rect 3448 408 3512 472
rect 3528 408 3592 472
rect 3608 408 3672 472
rect 3688 408 3752 472
rect 3768 408 3832 472
rect 3848 408 3912 472
rect 3928 408 3992 472
rect 19112 408 19176 472
rect 19192 408 19256 472
rect 19272 408 19336 472
rect 19352 408 19416 472
rect 29112 408 29176 472
rect 29192 408 29256 472
rect 29272 408 29336 472
rect 29352 408 29416 472
rect 41376 408 41440 472
rect 41456 408 41520 472
rect 41536 408 41600 472
rect 41616 408 41680 472
rect 41696 408 41760 472
rect 41776 408 41840 472
rect 41856 408 41920 472
rect 41936 408 42000 472
rect 42016 408 42080 472
rect 42096 408 42160 472
rect 42176 408 42240 472
rect 42256 408 42320 472
rect 42336 408 42400 472
rect 42416 408 42480 472
rect 42496 408 42560 472
rect 42576 408 42640 472
rect 42656 408 42720 472
rect 42736 408 42800 472
rect 42816 408 42880 472
rect 42896 408 42960 472
rect 42976 408 43040 472
rect 43056 408 43120 472
rect 43136 408 43200 472
rect 43216 408 43280 472
rect 43296 408 43360 472
rect 43376 408 43440 472
rect 43456 408 43520 472
rect 43536 408 43600 472
rect 43616 408 43680 472
rect 43696 408 43760 472
rect 43776 408 43840 472
rect 43856 408 43920 472
rect 43936 408 44000 472
rect 44016 408 44080 472
rect 44096 408 44160 472
rect 44176 408 44240 472
rect 44256 408 44320 472
rect 44336 408 44400 472
rect 44416 408 44480 472
rect 44496 408 44560 472
rect 44576 408 44640 472
rect 44656 408 44720 472
rect 44736 408 44800 472
rect 44816 408 44880 472
rect 44896 408 44960 472
rect 44976 408 45040 472
rect 45056 408 45120 472
rect 45136 408 45200 472
rect 45216 408 45280 472
rect 45296 408 45360 472
rect 8 328 72 392
rect 88 328 152 392
rect 168 328 232 392
rect 248 328 312 392
rect 328 328 392 392
rect 408 328 472 392
rect 488 328 552 392
rect 568 328 632 392
rect 648 328 712 392
rect 728 328 792 392
rect 808 328 872 392
rect 888 328 952 392
rect 968 328 1032 392
rect 1048 328 1112 392
rect 1128 328 1192 392
rect 1208 328 1272 392
rect 1288 328 1352 392
rect 1368 328 1432 392
rect 1448 328 1512 392
rect 1528 328 1592 392
rect 1608 328 1672 392
rect 1688 328 1752 392
rect 1768 328 1832 392
rect 1848 328 1912 392
rect 1928 328 1992 392
rect 2008 328 2072 392
rect 2088 328 2152 392
rect 2168 328 2232 392
rect 2248 328 2312 392
rect 2328 328 2392 392
rect 2408 328 2472 392
rect 2488 328 2552 392
rect 2568 328 2632 392
rect 2648 328 2712 392
rect 2728 328 2792 392
rect 2808 328 2872 392
rect 2888 328 2952 392
rect 2968 328 3032 392
rect 3048 328 3112 392
rect 3128 328 3192 392
rect 3208 328 3272 392
rect 3288 328 3352 392
rect 3368 328 3432 392
rect 3448 328 3512 392
rect 3528 328 3592 392
rect 3608 328 3672 392
rect 3688 328 3752 392
rect 3768 328 3832 392
rect 3848 328 3912 392
rect 3928 328 3992 392
rect 19112 328 19176 392
rect 19192 328 19256 392
rect 19272 328 19336 392
rect 19352 328 19416 392
rect 29112 328 29176 392
rect 29192 328 29256 392
rect 29272 328 29336 392
rect 29352 328 29416 392
rect 41376 328 41440 392
rect 41456 328 41520 392
rect 41536 328 41600 392
rect 41616 328 41680 392
rect 41696 328 41760 392
rect 41776 328 41840 392
rect 41856 328 41920 392
rect 41936 328 42000 392
rect 42016 328 42080 392
rect 42096 328 42160 392
rect 42176 328 42240 392
rect 42256 328 42320 392
rect 42336 328 42400 392
rect 42416 328 42480 392
rect 42496 328 42560 392
rect 42576 328 42640 392
rect 42656 328 42720 392
rect 42736 328 42800 392
rect 42816 328 42880 392
rect 42896 328 42960 392
rect 42976 328 43040 392
rect 43056 328 43120 392
rect 43136 328 43200 392
rect 43216 328 43280 392
rect 43296 328 43360 392
rect 43376 328 43440 392
rect 43456 328 43520 392
rect 43536 328 43600 392
rect 43616 328 43680 392
rect 43696 328 43760 392
rect 43776 328 43840 392
rect 43856 328 43920 392
rect 43936 328 44000 392
rect 44016 328 44080 392
rect 44096 328 44160 392
rect 44176 328 44240 392
rect 44256 328 44320 392
rect 44336 328 44400 392
rect 44416 328 44480 392
rect 44496 328 44560 392
rect 44576 328 44640 392
rect 44656 328 44720 392
rect 44736 328 44800 392
rect 44816 328 44880 392
rect 44896 328 44960 392
rect 44976 328 45040 392
rect 45056 328 45120 392
rect 45136 328 45200 392
rect 45216 328 45280 392
rect 45296 328 45360 392
rect 8 248 72 312
rect 88 248 152 312
rect 168 248 232 312
rect 248 248 312 312
rect 328 248 392 312
rect 408 248 472 312
rect 488 248 552 312
rect 568 248 632 312
rect 648 248 712 312
rect 728 248 792 312
rect 808 248 872 312
rect 888 248 952 312
rect 968 248 1032 312
rect 1048 248 1112 312
rect 1128 248 1192 312
rect 1208 248 1272 312
rect 1288 248 1352 312
rect 1368 248 1432 312
rect 1448 248 1512 312
rect 1528 248 1592 312
rect 1608 248 1672 312
rect 1688 248 1752 312
rect 1768 248 1832 312
rect 1848 248 1912 312
rect 1928 248 1992 312
rect 2008 248 2072 312
rect 2088 248 2152 312
rect 2168 248 2232 312
rect 2248 248 2312 312
rect 2328 248 2392 312
rect 2408 248 2472 312
rect 2488 248 2552 312
rect 2568 248 2632 312
rect 2648 248 2712 312
rect 2728 248 2792 312
rect 2808 248 2872 312
rect 2888 248 2952 312
rect 2968 248 3032 312
rect 3048 248 3112 312
rect 3128 248 3192 312
rect 3208 248 3272 312
rect 3288 248 3352 312
rect 3368 248 3432 312
rect 3448 248 3512 312
rect 3528 248 3592 312
rect 3608 248 3672 312
rect 3688 248 3752 312
rect 3768 248 3832 312
rect 3848 248 3912 312
rect 3928 248 3992 312
rect 19112 248 19176 312
rect 19192 248 19256 312
rect 19272 248 19336 312
rect 19352 248 19416 312
rect 29112 248 29176 312
rect 29192 248 29256 312
rect 29272 248 29336 312
rect 29352 248 29416 312
rect 41376 248 41440 312
rect 41456 248 41520 312
rect 41536 248 41600 312
rect 41616 248 41680 312
rect 41696 248 41760 312
rect 41776 248 41840 312
rect 41856 248 41920 312
rect 41936 248 42000 312
rect 42016 248 42080 312
rect 42096 248 42160 312
rect 42176 248 42240 312
rect 42256 248 42320 312
rect 42336 248 42400 312
rect 42416 248 42480 312
rect 42496 248 42560 312
rect 42576 248 42640 312
rect 42656 248 42720 312
rect 42736 248 42800 312
rect 42816 248 42880 312
rect 42896 248 42960 312
rect 42976 248 43040 312
rect 43056 248 43120 312
rect 43136 248 43200 312
rect 43216 248 43280 312
rect 43296 248 43360 312
rect 43376 248 43440 312
rect 43456 248 43520 312
rect 43536 248 43600 312
rect 43616 248 43680 312
rect 43696 248 43760 312
rect 43776 248 43840 312
rect 43856 248 43920 312
rect 43936 248 44000 312
rect 44016 248 44080 312
rect 44096 248 44160 312
rect 44176 248 44240 312
rect 44256 248 44320 312
rect 44336 248 44400 312
rect 44416 248 44480 312
rect 44496 248 44560 312
rect 44576 248 44640 312
rect 44656 248 44720 312
rect 44736 248 44800 312
rect 44816 248 44880 312
rect 44896 248 44960 312
rect 44976 248 45040 312
rect 45056 248 45120 312
rect 45136 248 45200 312
rect 45216 248 45280 312
rect 45296 248 45360 312
rect 8 168 72 232
rect 88 168 152 232
rect 168 168 232 232
rect 248 168 312 232
rect 328 168 392 232
rect 408 168 472 232
rect 488 168 552 232
rect 568 168 632 232
rect 648 168 712 232
rect 728 168 792 232
rect 808 168 872 232
rect 888 168 952 232
rect 968 168 1032 232
rect 1048 168 1112 232
rect 1128 168 1192 232
rect 1208 168 1272 232
rect 1288 168 1352 232
rect 1368 168 1432 232
rect 1448 168 1512 232
rect 1528 168 1592 232
rect 1608 168 1672 232
rect 1688 168 1752 232
rect 1768 168 1832 232
rect 1848 168 1912 232
rect 1928 168 1992 232
rect 2008 168 2072 232
rect 2088 168 2152 232
rect 2168 168 2232 232
rect 2248 168 2312 232
rect 2328 168 2392 232
rect 2408 168 2472 232
rect 2488 168 2552 232
rect 2568 168 2632 232
rect 2648 168 2712 232
rect 2728 168 2792 232
rect 2808 168 2872 232
rect 2888 168 2952 232
rect 2968 168 3032 232
rect 3048 168 3112 232
rect 3128 168 3192 232
rect 3208 168 3272 232
rect 3288 168 3352 232
rect 3368 168 3432 232
rect 3448 168 3512 232
rect 3528 168 3592 232
rect 3608 168 3672 232
rect 3688 168 3752 232
rect 3768 168 3832 232
rect 3848 168 3912 232
rect 3928 168 3992 232
rect 19112 168 19176 232
rect 19192 168 19256 232
rect 19272 168 19336 232
rect 19352 168 19416 232
rect 29112 168 29176 232
rect 29192 168 29256 232
rect 29272 168 29336 232
rect 29352 168 29416 232
rect 41376 168 41440 232
rect 41456 168 41520 232
rect 41536 168 41600 232
rect 41616 168 41680 232
rect 41696 168 41760 232
rect 41776 168 41840 232
rect 41856 168 41920 232
rect 41936 168 42000 232
rect 42016 168 42080 232
rect 42096 168 42160 232
rect 42176 168 42240 232
rect 42256 168 42320 232
rect 42336 168 42400 232
rect 42416 168 42480 232
rect 42496 168 42560 232
rect 42576 168 42640 232
rect 42656 168 42720 232
rect 42736 168 42800 232
rect 42816 168 42880 232
rect 42896 168 42960 232
rect 42976 168 43040 232
rect 43056 168 43120 232
rect 43136 168 43200 232
rect 43216 168 43280 232
rect 43296 168 43360 232
rect 43376 168 43440 232
rect 43456 168 43520 232
rect 43536 168 43600 232
rect 43616 168 43680 232
rect 43696 168 43760 232
rect 43776 168 43840 232
rect 43856 168 43920 232
rect 43936 168 44000 232
rect 44016 168 44080 232
rect 44096 168 44160 232
rect 44176 168 44240 232
rect 44256 168 44320 232
rect 44336 168 44400 232
rect 44416 168 44480 232
rect 44496 168 44560 232
rect 44576 168 44640 232
rect 44656 168 44720 232
rect 44736 168 44800 232
rect 44816 168 44880 232
rect 44896 168 44960 232
rect 44976 168 45040 232
rect 45056 168 45120 232
rect 45136 168 45200 232
rect 45216 168 45280 232
rect 45296 168 45360 232
rect 8 88 72 152
rect 88 88 152 152
rect 168 88 232 152
rect 248 88 312 152
rect 328 88 392 152
rect 408 88 472 152
rect 488 88 552 152
rect 568 88 632 152
rect 648 88 712 152
rect 728 88 792 152
rect 808 88 872 152
rect 888 88 952 152
rect 968 88 1032 152
rect 1048 88 1112 152
rect 1128 88 1192 152
rect 1208 88 1272 152
rect 1288 88 1352 152
rect 1368 88 1432 152
rect 1448 88 1512 152
rect 1528 88 1592 152
rect 1608 88 1672 152
rect 1688 88 1752 152
rect 1768 88 1832 152
rect 1848 88 1912 152
rect 1928 88 1992 152
rect 2008 88 2072 152
rect 2088 88 2152 152
rect 2168 88 2232 152
rect 2248 88 2312 152
rect 2328 88 2392 152
rect 2408 88 2472 152
rect 2488 88 2552 152
rect 2568 88 2632 152
rect 2648 88 2712 152
rect 2728 88 2792 152
rect 2808 88 2872 152
rect 2888 88 2952 152
rect 2968 88 3032 152
rect 3048 88 3112 152
rect 3128 88 3192 152
rect 3208 88 3272 152
rect 3288 88 3352 152
rect 3368 88 3432 152
rect 3448 88 3512 152
rect 3528 88 3592 152
rect 3608 88 3672 152
rect 3688 88 3752 152
rect 3768 88 3832 152
rect 3848 88 3912 152
rect 3928 88 3992 152
rect 19112 88 19176 152
rect 19192 88 19256 152
rect 19272 88 19336 152
rect 19352 88 19416 152
rect 29112 88 29176 152
rect 29192 88 29256 152
rect 29272 88 29336 152
rect 29352 88 29416 152
rect 41376 88 41440 152
rect 41456 88 41520 152
rect 41536 88 41600 152
rect 41616 88 41680 152
rect 41696 88 41760 152
rect 41776 88 41840 152
rect 41856 88 41920 152
rect 41936 88 42000 152
rect 42016 88 42080 152
rect 42096 88 42160 152
rect 42176 88 42240 152
rect 42256 88 42320 152
rect 42336 88 42400 152
rect 42416 88 42480 152
rect 42496 88 42560 152
rect 42576 88 42640 152
rect 42656 88 42720 152
rect 42736 88 42800 152
rect 42816 88 42880 152
rect 42896 88 42960 152
rect 42976 88 43040 152
rect 43056 88 43120 152
rect 43136 88 43200 152
rect 43216 88 43280 152
rect 43296 88 43360 152
rect 43376 88 43440 152
rect 43456 88 43520 152
rect 43536 88 43600 152
rect 43616 88 43680 152
rect 43696 88 43760 152
rect 43776 88 43840 152
rect 43856 88 43920 152
rect 43936 88 44000 152
rect 44016 88 44080 152
rect 44096 88 44160 152
rect 44176 88 44240 152
rect 44256 88 44320 152
rect 44336 88 44400 152
rect 44416 88 44480 152
rect 44496 88 44560 152
rect 44576 88 44640 152
rect 44656 88 44720 152
rect 44736 88 44800 152
rect 44816 88 44880 152
rect 44896 88 44960 152
rect 44976 88 45040 152
rect 45056 88 45120 152
rect 45136 88 45200 152
rect 45216 88 45280 152
rect 45296 88 45360 152
rect 8 8 72 72
rect 88 8 152 72
rect 168 8 232 72
rect 248 8 312 72
rect 328 8 392 72
rect 408 8 472 72
rect 488 8 552 72
rect 568 8 632 72
rect 648 8 712 72
rect 728 8 792 72
rect 808 8 872 72
rect 888 8 952 72
rect 968 8 1032 72
rect 1048 8 1112 72
rect 1128 8 1192 72
rect 1208 8 1272 72
rect 1288 8 1352 72
rect 1368 8 1432 72
rect 1448 8 1512 72
rect 1528 8 1592 72
rect 1608 8 1672 72
rect 1688 8 1752 72
rect 1768 8 1832 72
rect 1848 8 1912 72
rect 1928 8 1992 72
rect 2008 8 2072 72
rect 2088 8 2152 72
rect 2168 8 2232 72
rect 2248 8 2312 72
rect 2328 8 2392 72
rect 2408 8 2472 72
rect 2488 8 2552 72
rect 2568 8 2632 72
rect 2648 8 2712 72
rect 2728 8 2792 72
rect 2808 8 2872 72
rect 2888 8 2952 72
rect 2968 8 3032 72
rect 3048 8 3112 72
rect 3128 8 3192 72
rect 3208 8 3272 72
rect 3288 8 3352 72
rect 3368 8 3432 72
rect 3448 8 3512 72
rect 3528 8 3592 72
rect 3608 8 3672 72
rect 3688 8 3752 72
rect 3768 8 3832 72
rect 3848 8 3912 72
rect 3928 8 3992 72
rect 19112 8 19176 72
rect 19192 8 19256 72
rect 19272 8 19336 72
rect 19352 8 19416 72
rect 29112 8 29176 72
rect 29192 8 29256 72
rect 29272 8 29336 72
rect 29352 8 29416 72
rect 41376 8 41440 72
rect 41456 8 41520 72
rect 41536 8 41600 72
rect 41616 8 41680 72
rect 41696 8 41760 72
rect 41776 8 41840 72
rect 41856 8 41920 72
rect 41936 8 42000 72
rect 42016 8 42080 72
rect 42096 8 42160 72
rect 42176 8 42240 72
rect 42256 8 42320 72
rect 42336 8 42400 72
rect 42416 8 42480 72
rect 42496 8 42560 72
rect 42576 8 42640 72
rect 42656 8 42720 72
rect 42736 8 42800 72
rect 42816 8 42880 72
rect 42896 8 42960 72
rect 42976 8 43040 72
rect 43056 8 43120 72
rect 43136 8 43200 72
rect 43216 8 43280 72
rect 43296 8 43360 72
rect 43376 8 43440 72
rect 43456 8 43520 72
rect 43536 8 43600 72
rect 43616 8 43680 72
rect 43696 8 43760 72
rect 43776 8 43840 72
rect 43856 8 43920 72
rect 43936 8 44000 72
rect 44016 8 44080 72
rect 44096 8 44160 72
rect 44176 8 44240 72
rect 44256 8 44320 72
rect 44336 8 44400 72
rect 44416 8 44480 72
rect 44496 8 44560 72
rect 44576 8 44640 72
rect 44656 8 44720 72
rect 44736 8 44800 72
rect 44816 8 44880 72
rect 44896 8 44960 72
rect 44976 8 45040 72
rect 45056 8 45120 72
rect 45136 8 45200 72
rect 45216 8 45280 72
rect 45296 8 45360 72
<< metal4 >>
rect 0 45384 4000 45392
rect 0 45320 8 45384
rect 72 45320 88 45384
rect 152 45320 168 45384
rect 232 45320 248 45384
rect 312 45320 328 45384
rect 392 45320 408 45384
rect 472 45320 488 45384
rect 552 45320 568 45384
rect 632 45320 648 45384
rect 712 45320 728 45384
rect 792 45320 808 45384
rect 872 45320 888 45384
rect 952 45320 968 45384
rect 1032 45320 1048 45384
rect 1112 45320 1128 45384
rect 1192 45320 1208 45384
rect 1272 45320 1288 45384
rect 1352 45320 1368 45384
rect 1432 45320 1448 45384
rect 1512 45320 1528 45384
rect 1592 45320 1608 45384
rect 1672 45320 1688 45384
rect 1752 45320 1768 45384
rect 1832 45320 1848 45384
rect 1912 45320 1928 45384
rect 1992 45320 2008 45384
rect 2072 45320 2088 45384
rect 2152 45320 2168 45384
rect 2232 45320 2248 45384
rect 2312 45320 2328 45384
rect 2392 45320 2408 45384
rect 2472 45320 2488 45384
rect 2552 45320 2568 45384
rect 2632 45320 2648 45384
rect 2712 45320 2728 45384
rect 2792 45320 2808 45384
rect 2872 45320 2888 45384
rect 2952 45320 2968 45384
rect 3032 45320 3048 45384
rect 3112 45320 3128 45384
rect 3192 45320 3208 45384
rect 3272 45320 3288 45384
rect 3352 45320 3368 45384
rect 3432 45320 3448 45384
rect 3512 45320 3528 45384
rect 3592 45320 3608 45384
rect 3672 45320 3688 45384
rect 3752 45320 3768 45384
rect 3832 45320 3848 45384
rect 3912 45320 3928 45384
rect 3992 45320 4000 45384
rect 0 45304 4000 45320
rect 0 45240 8 45304
rect 72 45240 88 45304
rect 152 45240 168 45304
rect 232 45240 248 45304
rect 312 45240 328 45304
rect 392 45240 408 45304
rect 472 45240 488 45304
rect 552 45240 568 45304
rect 632 45240 648 45304
rect 712 45240 728 45304
rect 792 45240 808 45304
rect 872 45240 888 45304
rect 952 45240 968 45304
rect 1032 45240 1048 45304
rect 1112 45240 1128 45304
rect 1192 45240 1208 45304
rect 1272 45240 1288 45304
rect 1352 45240 1368 45304
rect 1432 45240 1448 45304
rect 1512 45240 1528 45304
rect 1592 45240 1608 45304
rect 1672 45240 1688 45304
rect 1752 45240 1768 45304
rect 1832 45240 1848 45304
rect 1912 45240 1928 45304
rect 1992 45240 2008 45304
rect 2072 45240 2088 45304
rect 2152 45240 2168 45304
rect 2232 45240 2248 45304
rect 2312 45240 2328 45304
rect 2392 45240 2408 45304
rect 2472 45240 2488 45304
rect 2552 45240 2568 45304
rect 2632 45240 2648 45304
rect 2712 45240 2728 45304
rect 2792 45240 2808 45304
rect 2872 45240 2888 45304
rect 2952 45240 2968 45304
rect 3032 45240 3048 45304
rect 3112 45240 3128 45304
rect 3192 45240 3208 45304
rect 3272 45240 3288 45304
rect 3352 45240 3368 45304
rect 3432 45240 3448 45304
rect 3512 45240 3528 45304
rect 3592 45240 3608 45304
rect 3672 45240 3688 45304
rect 3752 45240 3768 45304
rect 3832 45240 3848 45304
rect 3912 45240 3928 45304
rect 3992 45240 4000 45304
rect 0 45224 4000 45240
rect 0 45160 8 45224
rect 72 45160 88 45224
rect 152 45160 168 45224
rect 232 45160 248 45224
rect 312 45160 328 45224
rect 392 45160 408 45224
rect 472 45160 488 45224
rect 552 45160 568 45224
rect 632 45160 648 45224
rect 712 45160 728 45224
rect 792 45160 808 45224
rect 872 45160 888 45224
rect 952 45160 968 45224
rect 1032 45160 1048 45224
rect 1112 45160 1128 45224
rect 1192 45160 1208 45224
rect 1272 45160 1288 45224
rect 1352 45160 1368 45224
rect 1432 45160 1448 45224
rect 1512 45160 1528 45224
rect 1592 45160 1608 45224
rect 1672 45160 1688 45224
rect 1752 45160 1768 45224
rect 1832 45160 1848 45224
rect 1912 45160 1928 45224
rect 1992 45160 2008 45224
rect 2072 45160 2088 45224
rect 2152 45160 2168 45224
rect 2232 45160 2248 45224
rect 2312 45160 2328 45224
rect 2392 45160 2408 45224
rect 2472 45160 2488 45224
rect 2552 45160 2568 45224
rect 2632 45160 2648 45224
rect 2712 45160 2728 45224
rect 2792 45160 2808 45224
rect 2872 45160 2888 45224
rect 2952 45160 2968 45224
rect 3032 45160 3048 45224
rect 3112 45160 3128 45224
rect 3192 45160 3208 45224
rect 3272 45160 3288 45224
rect 3352 45160 3368 45224
rect 3432 45160 3448 45224
rect 3512 45160 3528 45224
rect 3592 45160 3608 45224
rect 3672 45160 3688 45224
rect 3752 45160 3768 45224
rect 3832 45160 3848 45224
rect 3912 45160 3928 45224
rect 3992 45160 4000 45224
rect 0 45144 4000 45160
rect 0 45080 8 45144
rect 72 45080 88 45144
rect 152 45080 168 45144
rect 232 45080 248 45144
rect 312 45080 328 45144
rect 392 45080 408 45144
rect 472 45080 488 45144
rect 552 45080 568 45144
rect 632 45080 648 45144
rect 712 45080 728 45144
rect 792 45080 808 45144
rect 872 45080 888 45144
rect 952 45080 968 45144
rect 1032 45080 1048 45144
rect 1112 45080 1128 45144
rect 1192 45080 1208 45144
rect 1272 45080 1288 45144
rect 1352 45080 1368 45144
rect 1432 45080 1448 45144
rect 1512 45080 1528 45144
rect 1592 45080 1608 45144
rect 1672 45080 1688 45144
rect 1752 45080 1768 45144
rect 1832 45080 1848 45144
rect 1912 45080 1928 45144
rect 1992 45080 2008 45144
rect 2072 45080 2088 45144
rect 2152 45080 2168 45144
rect 2232 45080 2248 45144
rect 2312 45080 2328 45144
rect 2392 45080 2408 45144
rect 2472 45080 2488 45144
rect 2552 45080 2568 45144
rect 2632 45080 2648 45144
rect 2712 45080 2728 45144
rect 2792 45080 2808 45144
rect 2872 45080 2888 45144
rect 2952 45080 2968 45144
rect 3032 45080 3048 45144
rect 3112 45080 3128 45144
rect 3192 45080 3208 45144
rect 3272 45080 3288 45144
rect 3352 45080 3368 45144
rect 3432 45080 3448 45144
rect 3512 45080 3528 45144
rect 3592 45080 3608 45144
rect 3672 45080 3688 45144
rect 3752 45080 3768 45144
rect 3832 45080 3848 45144
rect 3912 45080 3928 45144
rect 3992 45080 4000 45144
rect 0 45064 4000 45080
rect 0 45000 8 45064
rect 72 45000 88 45064
rect 152 45000 168 45064
rect 232 45000 248 45064
rect 312 45000 328 45064
rect 392 45000 408 45064
rect 472 45000 488 45064
rect 552 45000 568 45064
rect 632 45000 648 45064
rect 712 45000 728 45064
rect 792 45000 808 45064
rect 872 45000 888 45064
rect 952 45000 968 45064
rect 1032 45000 1048 45064
rect 1112 45000 1128 45064
rect 1192 45000 1208 45064
rect 1272 45000 1288 45064
rect 1352 45000 1368 45064
rect 1432 45000 1448 45064
rect 1512 45000 1528 45064
rect 1592 45000 1608 45064
rect 1672 45000 1688 45064
rect 1752 45000 1768 45064
rect 1832 45000 1848 45064
rect 1912 45000 1928 45064
rect 1992 45000 2008 45064
rect 2072 45000 2088 45064
rect 2152 45000 2168 45064
rect 2232 45000 2248 45064
rect 2312 45000 2328 45064
rect 2392 45000 2408 45064
rect 2472 45000 2488 45064
rect 2552 45000 2568 45064
rect 2632 45000 2648 45064
rect 2712 45000 2728 45064
rect 2792 45000 2808 45064
rect 2872 45000 2888 45064
rect 2952 45000 2968 45064
rect 3032 45000 3048 45064
rect 3112 45000 3128 45064
rect 3192 45000 3208 45064
rect 3272 45000 3288 45064
rect 3352 45000 3368 45064
rect 3432 45000 3448 45064
rect 3512 45000 3528 45064
rect 3592 45000 3608 45064
rect 3672 45000 3688 45064
rect 3752 45000 3768 45064
rect 3832 45000 3848 45064
rect 3912 45000 3928 45064
rect 3992 45000 4000 45064
rect 0 44984 4000 45000
rect 0 44920 8 44984
rect 72 44920 88 44984
rect 152 44920 168 44984
rect 232 44920 248 44984
rect 312 44920 328 44984
rect 392 44920 408 44984
rect 472 44920 488 44984
rect 552 44920 568 44984
rect 632 44920 648 44984
rect 712 44920 728 44984
rect 792 44920 808 44984
rect 872 44920 888 44984
rect 952 44920 968 44984
rect 1032 44920 1048 44984
rect 1112 44920 1128 44984
rect 1192 44920 1208 44984
rect 1272 44920 1288 44984
rect 1352 44920 1368 44984
rect 1432 44920 1448 44984
rect 1512 44920 1528 44984
rect 1592 44920 1608 44984
rect 1672 44920 1688 44984
rect 1752 44920 1768 44984
rect 1832 44920 1848 44984
rect 1912 44920 1928 44984
rect 1992 44920 2008 44984
rect 2072 44920 2088 44984
rect 2152 44920 2168 44984
rect 2232 44920 2248 44984
rect 2312 44920 2328 44984
rect 2392 44920 2408 44984
rect 2472 44920 2488 44984
rect 2552 44920 2568 44984
rect 2632 44920 2648 44984
rect 2712 44920 2728 44984
rect 2792 44920 2808 44984
rect 2872 44920 2888 44984
rect 2952 44920 2968 44984
rect 3032 44920 3048 44984
rect 3112 44920 3128 44984
rect 3192 44920 3208 44984
rect 3272 44920 3288 44984
rect 3352 44920 3368 44984
rect 3432 44920 3448 44984
rect 3512 44920 3528 44984
rect 3592 44920 3608 44984
rect 3672 44920 3688 44984
rect 3752 44920 3768 44984
rect 3832 44920 3848 44984
rect 3912 44920 3928 44984
rect 3992 44920 4000 44984
rect 0 44904 4000 44920
rect 0 44840 8 44904
rect 72 44840 88 44904
rect 152 44840 168 44904
rect 232 44840 248 44904
rect 312 44840 328 44904
rect 392 44840 408 44904
rect 472 44840 488 44904
rect 552 44840 568 44904
rect 632 44840 648 44904
rect 712 44840 728 44904
rect 792 44840 808 44904
rect 872 44840 888 44904
rect 952 44840 968 44904
rect 1032 44840 1048 44904
rect 1112 44840 1128 44904
rect 1192 44840 1208 44904
rect 1272 44840 1288 44904
rect 1352 44840 1368 44904
rect 1432 44840 1448 44904
rect 1512 44840 1528 44904
rect 1592 44840 1608 44904
rect 1672 44840 1688 44904
rect 1752 44840 1768 44904
rect 1832 44840 1848 44904
rect 1912 44840 1928 44904
rect 1992 44840 2008 44904
rect 2072 44840 2088 44904
rect 2152 44840 2168 44904
rect 2232 44840 2248 44904
rect 2312 44840 2328 44904
rect 2392 44840 2408 44904
rect 2472 44840 2488 44904
rect 2552 44840 2568 44904
rect 2632 44840 2648 44904
rect 2712 44840 2728 44904
rect 2792 44840 2808 44904
rect 2872 44840 2888 44904
rect 2952 44840 2968 44904
rect 3032 44840 3048 44904
rect 3112 44840 3128 44904
rect 3192 44840 3208 44904
rect 3272 44840 3288 44904
rect 3352 44840 3368 44904
rect 3432 44840 3448 44904
rect 3512 44840 3528 44904
rect 3592 44840 3608 44904
rect 3672 44840 3688 44904
rect 3752 44840 3768 44904
rect 3832 44840 3848 44904
rect 3912 44840 3928 44904
rect 3992 44840 4000 44904
rect 0 44824 4000 44840
rect 0 44760 8 44824
rect 72 44760 88 44824
rect 152 44760 168 44824
rect 232 44760 248 44824
rect 312 44760 328 44824
rect 392 44760 408 44824
rect 472 44760 488 44824
rect 552 44760 568 44824
rect 632 44760 648 44824
rect 712 44760 728 44824
rect 792 44760 808 44824
rect 872 44760 888 44824
rect 952 44760 968 44824
rect 1032 44760 1048 44824
rect 1112 44760 1128 44824
rect 1192 44760 1208 44824
rect 1272 44760 1288 44824
rect 1352 44760 1368 44824
rect 1432 44760 1448 44824
rect 1512 44760 1528 44824
rect 1592 44760 1608 44824
rect 1672 44760 1688 44824
rect 1752 44760 1768 44824
rect 1832 44760 1848 44824
rect 1912 44760 1928 44824
rect 1992 44760 2008 44824
rect 2072 44760 2088 44824
rect 2152 44760 2168 44824
rect 2232 44760 2248 44824
rect 2312 44760 2328 44824
rect 2392 44760 2408 44824
rect 2472 44760 2488 44824
rect 2552 44760 2568 44824
rect 2632 44760 2648 44824
rect 2712 44760 2728 44824
rect 2792 44760 2808 44824
rect 2872 44760 2888 44824
rect 2952 44760 2968 44824
rect 3032 44760 3048 44824
rect 3112 44760 3128 44824
rect 3192 44760 3208 44824
rect 3272 44760 3288 44824
rect 3352 44760 3368 44824
rect 3432 44760 3448 44824
rect 3512 44760 3528 44824
rect 3592 44760 3608 44824
rect 3672 44760 3688 44824
rect 3752 44760 3768 44824
rect 3832 44760 3848 44824
rect 3912 44760 3928 44824
rect 3992 44760 4000 44824
rect 0 44744 4000 44760
rect 0 44680 8 44744
rect 72 44680 88 44744
rect 152 44680 168 44744
rect 232 44680 248 44744
rect 312 44680 328 44744
rect 392 44680 408 44744
rect 472 44680 488 44744
rect 552 44680 568 44744
rect 632 44680 648 44744
rect 712 44680 728 44744
rect 792 44680 808 44744
rect 872 44680 888 44744
rect 952 44680 968 44744
rect 1032 44680 1048 44744
rect 1112 44680 1128 44744
rect 1192 44680 1208 44744
rect 1272 44680 1288 44744
rect 1352 44680 1368 44744
rect 1432 44680 1448 44744
rect 1512 44680 1528 44744
rect 1592 44680 1608 44744
rect 1672 44680 1688 44744
rect 1752 44680 1768 44744
rect 1832 44680 1848 44744
rect 1912 44680 1928 44744
rect 1992 44680 2008 44744
rect 2072 44680 2088 44744
rect 2152 44680 2168 44744
rect 2232 44680 2248 44744
rect 2312 44680 2328 44744
rect 2392 44680 2408 44744
rect 2472 44680 2488 44744
rect 2552 44680 2568 44744
rect 2632 44680 2648 44744
rect 2712 44680 2728 44744
rect 2792 44680 2808 44744
rect 2872 44680 2888 44744
rect 2952 44680 2968 44744
rect 3032 44680 3048 44744
rect 3112 44680 3128 44744
rect 3192 44680 3208 44744
rect 3272 44680 3288 44744
rect 3352 44680 3368 44744
rect 3432 44680 3448 44744
rect 3512 44680 3528 44744
rect 3592 44680 3608 44744
rect 3672 44680 3688 44744
rect 3752 44680 3768 44744
rect 3832 44680 3848 44744
rect 3912 44680 3928 44744
rect 3992 44680 4000 44744
rect 0 44664 4000 44680
rect 0 44600 8 44664
rect 72 44600 88 44664
rect 152 44600 168 44664
rect 232 44600 248 44664
rect 312 44600 328 44664
rect 392 44600 408 44664
rect 472 44600 488 44664
rect 552 44600 568 44664
rect 632 44600 648 44664
rect 712 44600 728 44664
rect 792 44600 808 44664
rect 872 44600 888 44664
rect 952 44600 968 44664
rect 1032 44600 1048 44664
rect 1112 44600 1128 44664
rect 1192 44600 1208 44664
rect 1272 44600 1288 44664
rect 1352 44600 1368 44664
rect 1432 44600 1448 44664
rect 1512 44600 1528 44664
rect 1592 44600 1608 44664
rect 1672 44600 1688 44664
rect 1752 44600 1768 44664
rect 1832 44600 1848 44664
rect 1912 44600 1928 44664
rect 1992 44600 2008 44664
rect 2072 44600 2088 44664
rect 2152 44600 2168 44664
rect 2232 44600 2248 44664
rect 2312 44600 2328 44664
rect 2392 44600 2408 44664
rect 2472 44600 2488 44664
rect 2552 44600 2568 44664
rect 2632 44600 2648 44664
rect 2712 44600 2728 44664
rect 2792 44600 2808 44664
rect 2872 44600 2888 44664
rect 2952 44600 2968 44664
rect 3032 44600 3048 44664
rect 3112 44600 3128 44664
rect 3192 44600 3208 44664
rect 3272 44600 3288 44664
rect 3352 44600 3368 44664
rect 3432 44600 3448 44664
rect 3512 44600 3528 44664
rect 3592 44600 3608 44664
rect 3672 44600 3688 44664
rect 3752 44600 3768 44664
rect 3832 44600 3848 44664
rect 3912 44600 3928 44664
rect 3992 44600 4000 44664
rect 0 44584 4000 44600
rect 0 44520 8 44584
rect 72 44520 88 44584
rect 152 44520 168 44584
rect 232 44520 248 44584
rect 312 44520 328 44584
rect 392 44520 408 44584
rect 472 44520 488 44584
rect 552 44520 568 44584
rect 632 44520 648 44584
rect 712 44520 728 44584
rect 792 44520 808 44584
rect 872 44520 888 44584
rect 952 44520 968 44584
rect 1032 44520 1048 44584
rect 1112 44520 1128 44584
rect 1192 44520 1208 44584
rect 1272 44520 1288 44584
rect 1352 44520 1368 44584
rect 1432 44520 1448 44584
rect 1512 44520 1528 44584
rect 1592 44520 1608 44584
rect 1672 44520 1688 44584
rect 1752 44520 1768 44584
rect 1832 44520 1848 44584
rect 1912 44520 1928 44584
rect 1992 44520 2008 44584
rect 2072 44520 2088 44584
rect 2152 44520 2168 44584
rect 2232 44520 2248 44584
rect 2312 44520 2328 44584
rect 2392 44520 2408 44584
rect 2472 44520 2488 44584
rect 2552 44520 2568 44584
rect 2632 44520 2648 44584
rect 2712 44520 2728 44584
rect 2792 44520 2808 44584
rect 2872 44520 2888 44584
rect 2952 44520 2968 44584
rect 3032 44520 3048 44584
rect 3112 44520 3128 44584
rect 3192 44520 3208 44584
rect 3272 44520 3288 44584
rect 3352 44520 3368 44584
rect 3432 44520 3448 44584
rect 3512 44520 3528 44584
rect 3592 44520 3608 44584
rect 3672 44520 3688 44584
rect 3752 44520 3768 44584
rect 3832 44520 3848 44584
rect 3912 44520 3928 44584
rect 3992 44520 4000 44584
rect 0 44504 4000 44520
rect 0 44440 8 44504
rect 72 44440 88 44504
rect 152 44440 168 44504
rect 232 44440 248 44504
rect 312 44440 328 44504
rect 392 44440 408 44504
rect 472 44440 488 44504
rect 552 44440 568 44504
rect 632 44440 648 44504
rect 712 44440 728 44504
rect 792 44440 808 44504
rect 872 44440 888 44504
rect 952 44440 968 44504
rect 1032 44440 1048 44504
rect 1112 44440 1128 44504
rect 1192 44440 1208 44504
rect 1272 44440 1288 44504
rect 1352 44440 1368 44504
rect 1432 44440 1448 44504
rect 1512 44440 1528 44504
rect 1592 44440 1608 44504
rect 1672 44440 1688 44504
rect 1752 44440 1768 44504
rect 1832 44440 1848 44504
rect 1912 44440 1928 44504
rect 1992 44440 2008 44504
rect 2072 44440 2088 44504
rect 2152 44440 2168 44504
rect 2232 44440 2248 44504
rect 2312 44440 2328 44504
rect 2392 44440 2408 44504
rect 2472 44440 2488 44504
rect 2552 44440 2568 44504
rect 2632 44440 2648 44504
rect 2712 44440 2728 44504
rect 2792 44440 2808 44504
rect 2872 44440 2888 44504
rect 2952 44440 2968 44504
rect 3032 44440 3048 44504
rect 3112 44440 3128 44504
rect 3192 44440 3208 44504
rect 3272 44440 3288 44504
rect 3352 44440 3368 44504
rect 3432 44440 3448 44504
rect 3512 44440 3528 44504
rect 3592 44440 3608 44504
rect 3672 44440 3688 44504
rect 3752 44440 3768 44504
rect 3832 44440 3848 44504
rect 3912 44440 3928 44504
rect 3992 44440 4000 44504
rect 0 44424 4000 44440
rect 0 44360 8 44424
rect 72 44360 88 44424
rect 152 44360 168 44424
rect 232 44360 248 44424
rect 312 44360 328 44424
rect 392 44360 408 44424
rect 472 44360 488 44424
rect 552 44360 568 44424
rect 632 44360 648 44424
rect 712 44360 728 44424
rect 792 44360 808 44424
rect 872 44360 888 44424
rect 952 44360 968 44424
rect 1032 44360 1048 44424
rect 1112 44360 1128 44424
rect 1192 44360 1208 44424
rect 1272 44360 1288 44424
rect 1352 44360 1368 44424
rect 1432 44360 1448 44424
rect 1512 44360 1528 44424
rect 1592 44360 1608 44424
rect 1672 44360 1688 44424
rect 1752 44360 1768 44424
rect 1832 44360 1848 44424
rect 1912 44360 1928 44424
rect 1992 44360 2008 44424
rect 2072 44360 2088 44424
rect 2152 44360 2168 44424
rect 2232 44360 2248 44424
rect 2312 44360 2328 44424
rect 2392 44360 2408 44424
rect 2472 44360 2488 44424
rect 2552 44360 2568 44424
rect 2632 44360 2648 44424
rect 2712 44360 2728 44424
rect 2792 44360 2808 44424
rect 2872 44360 2888 44424
rect 2952 44360 2968 44424
rect 3032 44360 3048 44424
rect 3112 44360 3128 44424
rect 3192 44360 3208 44424
rect 3272 44360 3288 44424
rect 3352 44360 3368 44424
rect 3432 44360 3448 44424
rect 3512 44360 3528 44424
rect 3592 44360 3608 44424
rect 3672 44360 3688 44424
rect 3752 44360 3768 44424
rect 3832 44360 3848 44424
rect 3912 44360 3928 44424
rect 3992 44360 4000 44424
rect 0 44344 4000 44360
rect 0 44280 8 44344
rect 72 44280 88 44344
rect 152 44280 168 44344
rect 232 44280 248 44344
rect 312 44280 328 44344
rect 392 44280 408 44344
rect 472 44280 488 44344
rect 552 44280 568 44344
rect 632 44280 648 44344
rect 712 44280 728 44344
rect 792 44280 808 44344
rect 872 44280 888 44344
rect 952 44280 968 44344
rect 1032 44280 1048 44344
rect 1112 44280 1128 44344
rect 1192 44280 1208 44344
rect 1272 44280 1288 44344
rect 1352 44280 1368 44344
rect 1432 44280 1448 44344
rect 1512 44280 1528 44344
rect 1592 44280 1608 44344
rect 1672 44280 1688 44344
rect 1752 44280 1768 44344
rect 1832 44280 1848 44344
rect 1912 44280 1928 44344
rect 1992 44280 2008 44344
rect 2072 44280 2088 44344
rect 2152 44280 2168 44344
rect 2232 44280 2248 44344
rect 2312 44280 2328 44344
rect 2392 44280 2408 44344
rect 2472 44280 2488 44344
rect 2552 44280 2568 44344
rect 2632 44280 2648 44344
rect 2712 44280 2728 44344
rect 2792 44280 2808 44344
rect 2872 44280 2888 44344
rect 2952 44280 2968 44344
rect 3032 44280 3048 44344
rect 3112 44280 3128 44344
rect 3192 44280 3208 44344
rect 3272 44280 3288 44344
rect 3352 44280 3368 44344
rect 3432 44280 3448 44344
rect 3512 44280 3528 44344
rect 3592 44280 3608 44344
rect 3672 44280 3688 44344
rect 3752 44280 3768 44344
rect 3832 44280 3848 44344
rect 3912 44280 3928 44344
rect 3992 44280 4000 44344
rect 0 44264 4000 44280
rect 0 44200 8 44264
rect 72 44200 88 44264
rect 152 44200 168 44264
rect 232 44200 248 44264
rect 312 44200 328 44264
rect 392 44200 408 44264
rect 472 44200 488 44264
rect 552 44200 568 44264
rect 632 44200 648 44264
rect 712 44200 728 44264
rect 792 44200 808 44264
rect 872 44200 888 44264
rect 952 44200 968 44264
rect 1032 44200 1048 44264
rect 1112 44200 1128 44264
rect 1192 44200 1208 44264
rect 1272 44200 1288 44264
rect 1352 44200 1368 44264
rect 1432 44200 1448 44264
rect 1512 44200 1528 44264
rect 1592 44200 1608 44264
rect 1672 44200 1688 44264
rect 1752 44200 1768 44264
rect 1832 44200 1848 44264
rect 1912 44200 1928 44264
rect 1992 44200 2008 44264
rect 2072 44200 2088 44264
rect 2152 44200 2168 44264
rect 2232 44200 2248 44264
rect 2312 44200 2328 44264
rect 2392 44200 2408 44264
rect 2472 44200 2488 44264
rect 2552 44200 2568 44264
rect 2632 44200 2648 44264
rect 2712 44200 2728 44264
rect 2792 44200 2808 44264
rect 2872 44200 2888 44264
rect 2952 44200 2968 44264
rect 3032 44200 3048 44264
rect 3112 44200 3128 44264
rect 3192 44200 3208 44264
rect 3272 44200 3288 44264
rect 3352 44200 3368 44264
rect 3432 44200 3448 44264
rect 3512 44200 3528 44264
rect 3592 44200 3608 44264
rect 3672 44200 3688 44264
rect 3752 44200 3768 44264
rect 3832 44200 3848 44264
rect 3912 44200 3928 44264
rect 3992 44200 4000 44264
rect 0 44184 4000 44200
rect 0 44120 8 44184
rect 72 44120 88 44184
rect 152 44120 168 44184
rect 232 44120 248 44184
rect 312 44120 328 44184
rect 392 44120 408 44184
rect 472 44120 488 44184
rect 552 44120 568 44184
rect 632 44120 648 44184
rect 712 44120 728 44184
rect 792 44120 808 44184
rect 872 44120 888 44184
rect 952 44120 968 44184
rect 1032 44120 1048 44184
rect 1112 44120 1128 44184
rect 1192 44120 1208 44184
rect 1272 44120 1288 44184
rect 1352 44120 1368 44184
rect 1432 44120 1448 44184
rect 1512 44120 1528 44184
rect 1592 44120 1608 44184
rect 1672 44120 1688 44184
rect 1752 44120 1768 44184
rect 1832 44120 1848 44184
rect 1912 44120 1928 44184
rect 1992 44120 2008 44184
rect 2072 44120 2088 44184
rect 2152 44120 2168 44184
rect 2232 44120 2248 44184
rect 2312 44120 2328 44184
rect 2392 44120 2408 44184
rect 2472 44120 2488 44184
rect 2552 44120 2568 44184
rect 2632 44120 2648 44184
rect 2712 44120 2728 44184
rect 2792 44120 2808 44184
rect 2872 44120 2888 44184
rect 2952 44120 2968 44184
rect 3032 44120 3048 44184
rect 3112 44120 3128 44184
rect 3192 44120 3208 44184
rect 3272 44120 3288 44184
rect 3352 44120 3368 44184
rect 3432 44120 3448 44184
rect 3512 44120 3528 44184
rect 3592 44120 3608 44184
rect 3672 44120 3688 44184
rect 3752 44120 3768 44184
rect 3832 44120 3848 44184
rect 3912 44120 3928 44184
rect 3992 44120 4000 44184
rect 0 44104 4000 44120
rect 0 44040 8 44104
rect 72 44040 88 44104
rect 152 44040 168 44104
rect 232 44040 248 44104
rect 312 44040 328 44104
rect 392 44040 408 44104
rect 472 44040 488 44104
rect 552 44040 568 44104
rect 632 44040 648 44104
rect 712 44040 728 44104
rect 792 44040 808 44104
rect 872 44040 888 44104
rect 952 44040 968 44104
rect 1032 44040 1048 44104
rect 1112 44040 1128 44104
rect 1192 44040 1208 44104
rect 1272 44040 1288 44104
rect 1352 44040 1368 44104
rect 1432 44040 1448 44104
rect 1512 44040 1528 44104
rect 1592 44040 1608 44104
rect 1672 44040 1688 44104
rect 1752 44040 1768 44104
rect 1832 44040 1848 44104
rect 1912 44040 1928 44104
rect 1992 44040 2008 44104
rect 2072 44040 2088 44104
rect 2152 44040 2168 44104
rect 2232 44040 2248 44104
rect 2312 44040 2328 44104
rect 2392 44040 2408 44104
rect 2472 44040 2488 44104
rect 2552 44040 2568 44104
rect 2632 44040 2648 44104
rect 2712 44040 2728 44104
rect 2792 44040 2808 44104
rect 2872 44040 2888 44104
rect 2952 44040 2968 44104
rect 3032 44040 3048 44104
rect 3112 44040 3128 44104
rect 3192 44040 3208 44104
rect 3272 44040 3288 44104
rect 3352 44040 3368 44104
rect 3432 44040 3448 44104
rect 3512 44040 3528 44104
rect 3592 44040 3608 44104
rect 3672 44040 3688 44104
rect 3752 44040 3768 44104
rect 3832 44040 3848 44104
rect 3912 44040 3928 44104
rect 3992 44040 4000 44104
rect 0 44024 4000 44040
rect 0 43960 8 44024
rect 72 43960 88 44024
rect 152 43960 168 44024
rect 232 43960 248 44024
rect 312 43960 328 44024
rect 392 43960 408 44024
rect 472 43960 488 44024
rect 552 43960 568 44024
rect 632 43960 648 44024
rect 712 43960 728 44024
rect 792 43960 808 44024
rect 872 43960 888 44024
rect 952 43960 968 44024
rect 1032 43960 1048 44024
rect 1112 43960 1128 44024
rect 1192 43960 1208 44024
rect 1272 43960 1288 44024
rect 1352 43960 1368 44024
rect 1432 43960 1448 44024
rect 1512 43960 1528 44024
rect 1592 43960 1608 44024
rect 1672 43960 1688 44024
rect 1752 43960 1768 44024
rect 1832 43960 1848 44024
rect 1912 43960 1928 44024
rect 1992 43960 2008 44024
rect 2072 43960 2088 44024
rect 2152 43960 2168 44024
rect 2232 43960 2248 44024
rect 2312 43960 2328 44024
rect 2392 43960 2408 44024
rect 2472 43960 2488 44024
rect 2552 43960 2568 44024
rect 2632 43960 2648 44024
rect 2712 43960 2728 44024
rect 2792 43960 2808 44024
rect 2872 43960 2888 44024
rect 2952 43960 2968 44024
rect 3032 43960 3048 44024
rect 3112 43960 3128 44024
rect 3192 43960 3208 44024
rect 3272 43960 3288 44024
rect 3352 43960 3368 44024
rect 3432 43960 3448 44024
rect 3512 43960 3528 44024
rect 3592 43960 3608 44024
rect 3672 43960 3688 44024
rect 3752 43960 3768 44024
rect 3832 43960 3848 44024
rect 3912 43960 3928 44024
rect 3992 43960 4000 44024
rect 0 43944 4000 43960
rect 0 43880 8 43944
rect 72 43880 88 43944
rect 152 43880 168 43944
rect 232 43880 248 43944
rect 312 43880 328 43944
rect 392 43880 408 43944
rect 472 43880 488 43944
rect 552 43880 568 43944
rect 632 43880 648 43944
rect 712 43880 728 43944
rect 792 43880 808 43944
rect 872 43880 888 43944
rect 952 43880 968 43944
rect 1032 43880 1048 43944
rect 1112 43880 1128 43944
rect 1192 43880 1208 43944
rect 1272 43880 1288 43944
rect 1352 43880 1368 43944
rect 1432 43880 1448 43944
rect 1512 43880 1528 43944
rect 1592 43880 1608 43944
rect 1672 43880 1688 43944
rect 1752 43880 1768 43944
rect 1832 43880 1848 43944
rect 1912 43880 1928 43944
rect 1992 43880 2008 43944
rect 2072 43880 2088 43944
rect 2152 43880 2168 43944
rect 2232 43880 2248 43944
rect 2312 43880 2328 43944
rect 2392 43880 2408 43944
rect 2472 43880 2488 43944
rect 2552 43880 2568 43944
rect 2632 43880 2648 43944
rect 2712 43880 2728 43944
rect 2792 43880 2808 43944
rect 2872 43880 2888 43944
rect 2952 43880 2968 43944
rect 3032 43880 3048 43944
rect 3112 43880 3128 43944
rect 3192 43880 3208 43944
rect 3272 43880 3288 43944
rect 3352 43880 3368 43944
rect 3432 43880 3448 43944
rect 3512 43880 3528 43944
rect 3592 43880 3608 43944
rect 3672 43880 3688 43944
rect 3752 43880 3768 43944
rect 3832 43880 3848 43944
rect 3912 43880 3928 43944
rect 3992 43880 4000 43944
rect 0 43864 4000 43880
rect 0 43800 8 43864
rect 72 43800 88 43864
rect 152 43800 168 43864
rect 232 43800 248 43864
rect 312 43800 328 43864
rect 392 43800 408 43864
rect 472 43800 488 43864
rect 552 43800 568 43864
rect 632 43800 648 43864
rect 712 43800 728 43864
rect 792 43800 808 43864
rect 872 43800 888 43864
rect 952 43800 968 43864
rect 1032 43800 1048 43864
rect 1112 43800 1128 43864
rect 1192 43800 1208 43864
rect 1272 43800 1288 43864
rect 1352 43800 1368 43864
rect 1432 43800 1448 43864
rect 1512 43800 1528 43864
rect 1592 43800 1608 43864
rect 1672 43800 1688 43864
rect 1752 43800 1768 43864
rect 1832 43800 1848 43864
rect 1912 43800 1928 43864
rect 1992 43800 2008 43864
rect 2072 43800 2088 43864
rect 2152 43800 2168 43864
rect 2232 43800 2248 43864
rect 2312 43800 2328 43864
rect 2392 43800 2408 43864
rect 2472 43800 2488 43864
rect 2552 43800 2568 43864
rect 2632 43800 2648 43864
rect 2712 43800 2728 43864
rect 2792 43800 2808 43864
rect 2872 43800 2888 43864
rect 2952 43800 2968 43864
rect 3032 43800 3048 43864
rect 3112 43800 3128 43864
rect 3192 43800 3208 43864
rect 3272 43800 3288 43864
rect 3352 43800 3368 43864
rect 3432 43800 3448 43864
rect 3512 43800 3528 43864
rect 3592 43800 3608 43864
rect 3672 43800 3688 43864
rect 3752 43800 3768 43864
rect 3832 43800 3848 43864
rect 3912 43800 3928 43864
rect 3992 43800 4000 43864
rect 0 43784 4000 43800
rect 0 43720 8 43784
rect 72 43720 88 43784
rect 152 43720 168 43784
rect 232 43720 248 43784
rect 312 43720 328 43784
rect 392 43720 408 43784
rect 472 43720 488 43784
rect 552 43720 568 43784
rect 632 43720 648 43784
rect 712 43720 728 43784
rect 792 43720 808 43784
rect 872 43720 888 43784
rect 952 43720 968 43784
rect 1032 43720 1048 43784
rect 1112 43720 1128 43784
rect 1192 43720 1208 43784
rect 1272 43720 1288 43784
rect 1352 43720 1368 43784
rect 1432 43720 1448 43784
rect 1512 43720 1528 43784
rect 1592 43720 1608 43784
rect 1672 43720 1688 43784
rect 1752 43720 1768 43784
rect 1832 43720 1848 43784
rect 1912 43720 1928 43784
rect 1992 43720 2008 43784
rect 2072 43720 2088 43784
rect 2152 43720 2168 43784
rect 2232 43720 2248 43784
rect 2312 43720 2328 43784
rect 2392 43720 2408 43784
rect 2472 43720 2488 43784
rect 2552 43720 2568 43784
rect 2632 43720 2648 43784
rect 2712 43720 2728 43784
rect 2792 43720 2808 43784
rect 2872 43720 2888 43784
rect 2952 43720 2968 43784
rect 3032 43720 3048 43784
rect 3112 43720 3128 43784
rect 3192 43720 3208 43784
rect 3272 43720 3288 43784
rect 3352 43720 3368 43784
rect 3432 43720 3448 43784
rect 3512 43720 3528 43784
rect 3592 43720 3608 43784
rect 3672 43720 3688 43784
rect 3752 43720 3768 43784
rect 3832 43720 3848 43784
rect 3912 43720 3928 43784
rect 3992 43720 4000 43784
rect 0 43704 4000 43720
rect 0 43640 8 43704
rect 72 43640 88 43704
rect 152 43640 168 43704
rect 232 43640 248 43704
rect 312 43640 328 43704
rect 392 43640 408 43704
rect 472 43640 488 43704
rect 552 43640 568 43704
rect 632 43640 648 43704
rect 712 43640 728 43704
rect 792 43640 808 43704
rect 872 43640 888 43704
rect 952 43640 968 43704
rect 1032 43640 1048 43704
rect 1112 43640 1128 43704
rect 1192 43640 1208 43704
rect 1272 43640 1288 43704
rect 1352 43640 1368 43704
rect 1432 43640 1448 43704
rect 1512 43640 1528 43704
rect 1592 43640 1608 43704
rect 1672 43640 1688 43704
rect 1752 43640 1768 43704
rect 1832 43640 1848 43704
rect 1912 43640 1928 43704
rect 1992 43640 2008 43704
rect 2072 43640 2088 43704
rect 2152 43640 2168 43704
rect 2232 43640 2248 43704
rect 2312 43640 2328 43704
rect 2392 43640 2408 43704
rect 2472 43640 2488 43704
rect 2552 43640 2568 43704
rect 2632 43640 2648 43704
rect 2712 43640 2728 43704
rect 2792 43640 2808 43704
rect 2872 43640 2888 43704
rect 2952 43640 2968 43704
rect 3032 43640 3048 43704
rect 3112 43640 3128 43704
rect 3192 43640 3208 43704
rect 3272 43640 3288 43704
rect 3352 43640 3368 43704
rect 3432 43640 3448 43704
rect 3512 43640 3528 43704
rect 3592 43640 3608 43704
rect 3672 43640 3688 43704
rect 3752 43640 3768 43704
rect 3832 43640 3848 43704
rect 3912 43640 3928 43704
rect 3992 43640 4000 43704
rect 0 43624 4000 43640
rect 0 43560 8 43624
rect 72 43560 88 43624
rect 152 43560 168 43624
rect 232 43560 248 43624
rect 312 43560 328 43624
rect 392 43560 408 43624
rect 472 43560 488 43624
rect 552 43560 568 43624
rect 632 43560 648 43624
rect 712 43560 728 43624
rect 792 43560 808 43624
rect 872 43560 888 43624
rect 952 43560 968 43624
rect 1032 43560 1048 43624
rect 1112 43560 1128 43624
rect 1192 43560 1208 43624
rect 1272 43560 1288 43624
rect 1352 43560 1368 43624
rect 1432 43560 1448 43624
rect 1512 43560 1528 43624
rect 1592 43560 1608 43624
rect 1672 43560 1688 43624
rect 1752 43560 1768 43624
rect 1832 43560 1848 43624
rect 1912 43560 1928 43624
rect 1992 43560 2008 43624
rect 2072 43560 2088 43624
rect 2152 43560 2168 43624
rect 2232 43560 2248 43624
rect 2312 43560 2328 43624
rect 2392 43560 2408 43624
rect 2472 43560 2488 43624
rect 2552 43560 2568 43624
rect 2632 43560 2648 43624
rect 2712 43560 2728 43624
rect 2792 43560 2808 43624
rect 2872 43560 2888 43624
rect 2952 43560 2968 43624
rect 3032 43560 3048 43624
rect 3112 43560 3128 43624
rect 3192 43560 3208 43624
rect 3272 43560 3288 43624
rect 3352 43560 3368 43624
rect 3432 43560 3448 43624
rect 3512 43560 3528 43624
rect 3592 43560 3608 43624
rect 3672 43560 3688 43624
rect 3752 43560 3768 43624
rect 3832 43560 3848 43624
rect 3912 43560 3928 43624
rect 3992 43560 4000 43624
rect 0 43544 4000 43560
rect 0 43480 8 43544
rect 72 43480 88 43544
rect 152 43480 168 43544
rect 232 43480 248 43544
rect 312 43480 328 43544
rect 392 43480 408 43544
rect 472 43480 488 43544
rect 552 43480 568 43544
rect 632 43480 648 43544
rect 712 43480 728 43544
rect 792 43480 808 43544
rect 872 43480 888 43544
rect 952 43480 968 43544
rect 1032 43480 1048 43544
rect 1112 43480 1128 43544
rect 1192 43480 1208 43544
rect 1272 43480 1288 43544
rect 1352 43480 1368 43544
rect 1432 43480 1448 43544
rect 1512 43480 1528 43544
rect 1592 43480 1608 43544
rect 1672 43480 1688 43544
rect 1752 43480 1768 43544
rect 1832 43480 1848 43544
rect 1912 43480 1928 43544
rect 1992 43480 2008 43544
rect 2072 43480 2088 43544
rect 2152 43480 2168 43544
rect 2232 43480 2248 43544
rect 2312 43480 2328 43544
rect 2392 43480 2408 43544
rect 2472 43480 2488 43544
rect 2552 43480 2568 43544
rect 2632 43480 2648 43544
rect 2712 43480 2728 43544
rect 2792 43480 2808 43544
rect 2872 43480 2888 43544
rect 2952 43480 2968 43544
rect 3032 43480 3048 43544
rect 3112 43480 3128 43544
rect 3192 43480 3208 43544
rect 3272 43480 3288 43544
rect 3352 43480 3368 43544
rect 3432 43480 3448 43544
rect 3512 43480 3528 43544
rect 3592 43480 3608 43544
rect 3672 43480 3688 43544
rect 3752 43480 3768 43544
rect 3832 43480 3848 43544
rect 3912 43480 3928 43544
rect 3992 43480 4000 43544
rect 0 43464 4000 43480
rect 0 43400 8 43464
rect 72 43400 88 43464
rect 152 43400 168 43464
rect 232 43400 248 43464
rect 312 43400 328 43464
rect 392 43400 408 43464
rect 472 43400 488 43464
rect 552 43400 568 43464
rect 632 43400 648 43464
rect 712 43400 728 43464
rect 792 43400 808 43464
rect 872 43400 888 43464
rect 952 43400 968 43464
rect 1032 43400 1048 43464
rect 1112 43400 1128 43464
rect 1192 43400 1208 43464
rect 1272 43400 1288 43464
rect 1352 43400 1368 43464
rect 1432 43400 1448 43464
rect 1512 43400 1528 43464
rect 1592 43400 1608 43464
rect 1672 43400 1688 43464
rect 1752 43400 1768 43464
rect 1832 43400 1848 43464
rect 1912 43400 1928 43464
rect 1992 43400 2008 43464
rect 2072 43400 2088 43464
rect 2152 43400 2168 43464
rect 2232 43400 2248 43464
rect 2312 43400 2328 43464
rect 2392 43400 2408 43464
rect 2472 43400 2488 43464
rect 2552 43400 2568 43464
rect 2632 43400 2648 43464
rect 2712 43400 2728 43464
rect 2792 43400 2808 43464
rect 2872 43400 2888 43464
rect 2952 43400 2968 43464
rect 3032 43400 3048 43464
rect 3112 43400 3128 43464
rect 3192 43400 3208 43464
rect 3272 43400 3288 43464
rect 3352 43400 3368 43464
rect 3432 43400 3448 43464
rect 3512 43400 3528 43464
rect 3592 43400 3608 43464
rect 3672 43400 3688 43464
rect 3752 43400 3768 43464
rect 3832 43400 3848 43464
rect 3912 43400 3928 43464
rect 3992 43400 4000 43464
rect 0 43384 4000 43400
rect 0 43320 8 43384
rect 72 43320 88 43384
rect 152 43320 168 43384
rect 232 43320 248 43384
rect 312 43320 328 43384
rect 392 43320 408 43384
rect 472 43320 488 43384
rect 552 43320 568 43384
rect 632 43320 648 43384
rect 712 43320 728 43384
rect 792 43320 808 43384
rect 872 43320 888 43384
rect 952 43320 968 43384
rect 1032 43320 1048 43384
rect 1112 43320 1128 43384
rect 1192 43320 1208 43384
rect 1272 43320 1288 43384
rect 1352 43320 1368 43384
rect 1432 43320 1448 43384
rect 1512 43320 1528 43384
rect 1592 43320 1608 43384
rect 1672 43320 1688 43384
rect 1752 43320 1768 43384
rect 1832 43320 1848 43384
rect 1912 43320 1928 43384
rect 1992 43320 2008 43384
rect 2072 43320 2088 43384
rect 2152 43320 2168 43384
rect 2232 43320 2248 43384
rect 2312 43320 2328 43384
rect 2392 43320 2408 43384
rect 2472 43320 2488 43384
rect 2552 43320 2568 43384
rect 2632 43320 2648 43384
rect 2712 43320 2728 43384
rect 2792 43320 2808 43384
rect 2872 43320 2888 43384
rect 2952 43320 2968 43384
rect 3032 43320 3048 43384
rect 3112 43320 3128 43384
rect 3192 43320 3208 43384
rect 3272 43320 3288 43384
rect 3352 43320 3368 43384
rect 3432 43320 3448 43384
rect 3512 43320 3528 43384
rect 3592 43320 3608 43384
rect 3672 43320 3688 43384
rect 3752 43320 3768 43384
rect 3832 43320 3848 43384
rect 3912 43320 3928 43384
rect 3992 43320 4000 43384
rect 0 43304 4000 43320
rect 0 43240 8 43304
rect 72 43240 88 43304
rect 152 43240 168 43304
rect 232 43240 248 43304
rect 312 43240 328 43304
rect 392 43240 408 43304
rect 472 43240 488 43304
rect 552 43240 568 43304
rect 632 43240 648 43304
rect 712 43240 728 43304
rect 792 43240 808 43304
rect 872 43240 888 43304
rect 952 43240 968 43304
rect 1032 43240 1048 43304
rect 1112 43240 1128 43304
rect 1192 43240 1208 43304
rect 1272 43240 1288 43304
rect 1352 43240 1368 43304
rect 1432 43240 1448 43304
rect 1512 43240 1528 43304
rect 1592 43240 1608 43304
rect 1672 43240 1688 43304
rect 1752 43240 1768 43304
rect 1832 43240 1848 43304
rect 1912 43240 1928 43304
rect 1992 43240 2008 43304
rect 2072 43240 2088 43304
rect 2152 43240 2168 43304
rect 2232 43240 2248 43304
rect 2312 43240 2328 43304
rect 2392 43240 2408 43304
rect 2472 43240 2488 43304
rect 2552 43240 2568 43304
rect 2632 43240 2648 43304
rect 2712 43240 2728 43304
rect 2792 43240 2808 43304
rect 2872 43240 2888 43304
rect 2952 43240 2968 43304
rect 3032 43240 3048 43304
rect 3112 43240 3128 43304
rect 3192 43240 3208 43304
rect 3272 43240 3288 43304
rect 3352 43240 3368 43304
rect 3432 43240 3448 43304
rect 3512 43240 3528 43304
rect 3592 43240 3608 43304
rect 3672 43240 3688 43304
rect 3752 43240 3768 43304
rect 3832 43240 3848 43304
rect 3912 43240 3928 43304
rect 3992 43240 4000 43304
rect 0 43224 4000 43240
rect 0 43160 8 43224
rect 72 43160 88 43224
rect 152 43160 168 43224
rect 232 43160 248 43224
rect 312 43160 328 43224
rect 392 43160 408 43224
rect 472 43160 488 43224
rect 552 43160 568 43224
rect 632 43160 648 43224
rect 712 43160 728 43224
rect 792 43160 808 43224
rect 872 43160 888 43224
rect 952 43160 968 43224
rect 1032 43160 1048 43224
rect 1112 43160 1128 43224
rect 1192 43160 1208 43224
rect 1272 43160 1288 43224
rect 1352 43160 1368 43224
rect 1432 43160 1448 43224
rect 1512 43160 1528 43224
rect 1592 43160 1608 43224
rect 1672 43160 1688 43224
rect 1752 43160 1768 43224
rect 1832 43160 1848 43224
rect 1912 43160 1928 43224
rect 1992 43160 2008 43224
rect 2072 43160 2088 43224
rect 2152 43160 2168 43224
rect 2232 43160 2248 43224
rect 2312 43160 2328 43224
rect 2392 43160 2408 43224
rect 2472 43160 2488 43224
rect 2552 43160 2568 43224
rect 2632 43160 2648 43224
rect 2712 43160 2728 43224
rect 2792 43160 2808 43224
rect 2872 43160 2888 43224
rect 2952 43160 2968 43224
rect 3032 43160 3048 43224
rect 3112 43160 3128 43224
rect 3192 43160 3208 43224
rect 3272 43160 3288 43224
rect 3352 43160 3368 43224
rect 3432 43160 3448 43224
rect 3512 43160 3528 43224
rect 3592 43160 3608 43224
rect 3672 43160 3688 43224
rect 3752 43160 3768 43224
rect 3832 43160 3848 43224
rect 3912 43160 3928 43224
rect 3992 43160 4000 43224
rect 0 43144 4000 43160
rect 0 43080 8 43144
rect 72 43080 88 43144
rect 152 43080 168 43144
rect 232 43080 248 43144
rect 312 43080 328 43144
rect 392 43080 408 43144
rect 472 43080 488 43144
rect 552 43080 568 43144
rect 632 43080 648 43144
rect 712 43080 728 43144
rect 792 43080 808 43144
rect 872 43080 888 43144
rect 952 43080 968 43144
rect 1032 43080 1048 43144
rect 1112 43080 1128 43144
rect 1192 43080 1208 43144
rect 1272 43080 1288 43144
rect 1352 43080 1368 43144
rect 1432 43080 1448 43144
rect 1512 43080 1528 43144
rect 1592 43080 1608 43144
rect 1672 43080 1688 43144
rect 1752 43080 1768 43144
rect 1832 43080 1848 43144
rect 1912 43080 1928 43144
rect 1992 43080 2008 43144
rect 2072 43080 2088 43144
rect 2152 43080 2168 43144
rect 2232 43080 2248 43144
rect 2312 43080 2328 43144
rect 2392 43080 2408 43144
rect 2472 43080 2488 43144
rect 2552 43080 2568 43144
rect 2632 43080 2648 43144
rect 2712 43080 2728 43144
rect 2792 43080 2808 43144
rect 2872 43080 2888 43144
rect 2952 43080 2968 43144
rect 3032 43080 3048 43144
rect 3112 43080 3128 43144
rect 3192 43080 3208 43144
rect 3272 43080 3288 43144
rect 3352 43080 3368 43144
rect 3432 43080 3448 43144
rect 3512 43080 3528 43144
rect 3592 43080 3608 43144
rect 3672 43080 3688 43144
rect 3752 43080 3768 43144
rect 3832 43080 3848 43144
rect 3912 43080 3928 43144
rect 3992 43080 4000 43144
rect 0 43064 4000 43080
rect 0 43000 8 43064
rect 72 43000 88 43064
rect 152 43000 168 43064
rect 232 43000 248 43064
rect 312 43000 328 43064
rect 392 43000 408 43064
rect 472 43000 488 43064
rect 552 43000 568 43064
rect 632 43000 648 43064
rect 712 43000 728 43064
rect 792 43000 808 43064
rect 872 43000 888 43064
rect 952 43000 968 43064
rect 1032 43000 1048 43064
rect 1112 43000 1128 43064
rect 1192 43000 1208 43064
rect 1272 43000 1288 43064
rect 1352 43000 1368 43064
rect 1432 43000 1448 43064
rect 1512 43000 1528 43064
rect 1592 43000 1608 43064
rect 1672 43000 1688 43064
rect 1752 43000 1768 43064
rect 1832 43000 1848 43064
rect 1912 43000 1928 43064
rect 1992 43000 2008 43064
rect 2072 43000 2088 43064
rect 2152 43000 2168 43064
rect 2232 43000 2248 43064
rect 2312 43000 2328 43064
rect 2392 43000 2408 43064
rect 2472 43000 2488 43064
rect 2552 43000 2568 43064
rect 2632 43000 2648 43064
rect 2712 43000 2728 43064
rect 2792 43000 2808 43064
rect 2872 43000 2888 43064
rect 2952 43000 2968 43064
rect 3032 43000 3048 43064
rect 3112 43000 3128 43064
rect 3192 43000 3208 43064
rect 3272 43000 3288 43064
rect 3352 43000 3368 43064
rect 3432 43000 3448 43064
rect 3512 43000 3528 43064
rect 3592 43000 3608 43064
rect 3672 43000 3688 43064
rect 3752 43000 3768 43064
rect 3832 43000 3848 43064
rect 3912 43000 3928 43064
rect 3992 43000 4000 43064
rect 0 42984 4000 43000
rect 0 42920 8 42984
rect 72 42920 88 42984
rect 152 42920 168 42984
rect 232 42920 248 42984
rect 312 42920 328 42984
rect 392 42920 408 42984
rect 472 42920 488 42984
rect 552 42920 568 42984
rect 632 42920 648 42984
rect 712 42920 728 42984
rect 792 42920 808 42984
rect 872 42920 888 42984
rect 952 42920 968 42984
rect 1032 42920 1048 42984
rect 1112 42920 1128 42984
rect 1192 42920 1208 42984
rect 1272 42920 1288 42984
rect 1352 42920 1368 42984
rect 1432 42920 1448 42984
rect 1512 42920 1528 42984
rect 1592 42920 1608 42984
rect 1672 42920 1688 42984
rect 1752 42920 1768 42984
rect 1832 42920 1848 42984
rect 1912 42920 1928 42984
rect 1992 42920 2008 42984
rect 2072 42920 2088 42984
rect 2152 42920 2168 42984
rect 2232 42920 2248 42984
rect 2312 42920 2328 42984
rect 2392 42920 2408 42984
rect 2472 42920 2488 42984
rect 2552 42920 2568 42984
rect 2632 42920 2648 42984
rect 2712 42920 2728 42984
rect 2792 42920 2808 42984
rect 2872 42920 2888 42984
rect 2952 42920 2968 42984
rect 3032 42920 3048 42984
rect 3112 42920 3128 42984
rect 3192 42920 3208 42984
rect 3272 42920 3288 42984
rect 3352 42920 3368 42984
rect 3432 42920 3448 42984
rect 3512 42920 3528 42984
rect 3592 42920 3608 42984
rect 3672 42920 3688 42984
rect 3752 42920 3768 42984
rect 3832 42920 3848 42984
rect 3912 42920 3928 42984
rect 3992 42920 4000 42984
rect 0 42904 4000 42920
rect 0 42840 8 42904
rect 72 42840 88 42904
rect 152 42840 168 42904
rect 232 42840 248 42904
rect 312 42840 328 42904
rect 392 42840 408 42904
rect 472 42840 488 42904
rect 552 42840 568 42904
rect 632 42840 648 42904
rect 712 42840 728 42904
rect 792 42840 808 42904
rect 872 42840 888 42904
rect 952 42840 968 42904
rect 1032 42840 1048 42904
rect 1112 42840 1128 42904
rect 1192 42840 1208 42904
rect 1272 42840 1288 42904
rect 1352 42840 1368 42904
rect 1432 42840 1448 42904
rect 1512 42840 1528 42904
rect 1592 42840 1608 42904
rect 1672 42840 1688 42904
rect 1752 42840 1768 42904
rect 1832 42840 1848 42904
rect 1912 42840 1928 42904
rect 1992 42840 2008 42904
rect 2072 42840 2088 42904
rect 2152 42840 2168 42904
rect 2232 42840 2248 42904
rect 2312 42840 2328 42904
rect 2392 42840 2408 42904
rect 2472 42840 2488 42904
rect 2552 42840 2568 42904
rect 2632 42840 2648 42904
rect 2712 42840 2728 42904
rect 2792 42840 2808 42904
rect 2872 42840 2888 42904
rect 2952 42840 2968 42904
rect 3032 42840 3048 42904
rect 3112 42840 3128 42904
rect 3192 42840 3208 42904
rect 3272 42840 3288 42904
rect 3352 42840 3368 42904
rect 3432 42840 3448 42904
rect 3512 42840 3528 42904
rect 3592 42840 3608 42904
rect 3672 42840 3688 42904
rect 3752 42840 3768 42904
rect 3832 42840 3848 42904
rect 3912 42840 3928 42904
rect 3992 42840 4000 42904
rect 0 42824 4000 42840
rect 0 42760 8 42824
rect 72 42760 88 42824
rect 152 42760 168 42824
rect 232 42760 248 42824
rect 312 42760 328 42824
rect 392 42760 408 42824
rect 472 42760 488 42824
rect 552 42760 568 42824
rect 632 42760 648 42824
rect 712 42760 728 42824
rect 792 42760 808 42824
rect 872 42760 888 42824
rect 952 42760 968 42824
rect 1032 42760 1048 42824
rect 1112 42760 1128 42824
rect 1192 42760 1208 42824
rect 1272 42760 1288 42824
rect 1352 42760 1368 42824
rect 1432 42760 1448 42824
rect 1512 42760 1528 42824
rect 1592 42760 1608 42824
rect 1672 42760 1688 42824
rect 1752 42760 1768 42824
rect 1832 42760 1848 42824
rect 1912 42760 1928 42824
rect 1992 42760 2008 42824
rect 2072 42760 2088 42824
rect 2152 42760 2168 42824
rect 2232 42760 2248 42824
rect 2312 42760 2328 42824
rect 2392 42760 2408 42824
rect 2472 42760 2488 42824
rect 2552 42760 2568 42824
rect 2632 42760 2648 42824
rect 2712 42760 2728 42824
rect 2792 42760 2808 42824
rect 2872 42760 2888 42824
rect 2952 42760 2968 42824
rect 3032 42760 3048 42824
rect 3112 42760 3128 42824
rect 3192 42760 3208 42824
rect 3272 42760 3288 42824
rect 3352 42760 3368 42824
rect 3432 42760 3448 42824
rect 3512 42760 3528 42824
rect 3592 42760 3608 42824
rect 3672 42760 3688 42824
rect 3752 42760 3768 42824
rect 3832 42760 3848 42824
rect 3912 42760 3928 42824
rect 3992 42760 4000 42824
rect 0 42744 4000 42760
rect 0 42680 8 42744
rect 72 42680 88 42744
rect 152 42680 168 42744
rect 232 42680 248 42744
rect 312 42680 328 42744
rect 392 42680 408 42744
rect 472 42680 488 42744
rect 552 42680 568 42744
rect 632 42680 648 42744
rect 712 42680 728 42744
rect 792 42680 808 42744
rect 872 42680 888 42744
rect 952 42680 968 42744
rect 1032 42680 1048 42744
rect 1112 42680 1128 42744
rect 1192 42680 1208 42744
rect 1272 42680 1288 42744
rect 1352 42680 1368 42744
rect 1432 42680 1448 42744
rect 1512 42680 1528 42744
rect 1592 42680 1608 42744
rect 1672 42680 1688 42744
rect 1752 42680 1768 42744
rect 1832 42680 1848 42744
rect 1912 42680 1928 42744
rect 1992 42680 2008 42744
rect 2072 42680 2088 42744
rect 2152 42680 2168 42744
rect 2232 42680 2248 42744
rect 2312 42680 2328 42744
rect 2392 42680 2408 42744
rect 2472 42680 2488 42744
rect 2552 42680 2568 42744
rect 2632 42680 2648 42744
rect 2712 42680 2728 42744
rect 2792 42680 2808 42744
rect 2872 42680 2888 42744
rect 2952 42680 2968 42744
rect 3032 42680 3048 42744
rect 3112 42680 3128 42744
rect 3192 42680 3208 42744
rect 3272 42680 3288 42744
rect 3352 42680 3368 42744
rect 3432 42680 3448 42744
rect 3512 42680 3528 42744
rect 3592 42680 3608 42744
rect 3672 42680 3688 42744
rect 3752 42680 3768 42744
rect 3832 42680 3848 42744
rect 3912 42680 3928 42744
rect 3992 42680 4000 42744
rect 0 42664 4000 42680
rect 0 42600 8 42664
rect 72 42600 88 42664
rect 152 42600 168 42664
rect 232 42600 248 42664
rect 312 42600 328 42664
rect 392 42600 408 42664
rect 472 42600 488 42664
rect 552 42600 568 42664
rect 632 42600 648 42664
rect 712 42600 728 42664
rect 792 42600 808 42664
rect 872 42600 888 42664
rect 952 42600 968 42664
rect 1032 42600 1048 42664
rect 1112 42600 1128 42664
rect 1192 42600 1208 42664
rect 1272 42600 1288 42664
rect 1352 42600 1368 42664
rect 1432 42600 1448 42664
rect 1512 42600 1528 42664
rect 1592 42600 1608 42664
rect 1672 42600 1688 42664
rect 1752 42600 1768 42664
rect 1832 42600 1848 42664
rect 1912 42600 1928 42664
rect 1992 42600 2008 42664
rect 2072 42600 2088 42664
rect 2152 42600 2168 42664
rect 2232 42600 2248 42664
rect 2312 42600 2328 42664
rect 2392 42600 2408 42664
rect 2472 42600 2488 42664
rect 2552 42600 2568 42664
rect 2632 42600 2648 42664
rect 2712 42600 2728 42664
rect 2792 42600 2808 42664
rect 2872 42600 2888 42664
rect 2952 42600 2968 42664
rect 3032 42600 3048 42664
rect 3112 42600 3128 42664
rect 3192 42600 3208 42664
rect 3272 42600 3288 42664
rect 3352 42600 3368 42664
rect 3432 42600 3448 42664
rect 3512 42600 3528 42664
rect 3592 42600 3608 42664
rect 3672 42600 3688 42664
rect 3752 42600 3768 42664
rect 3832 42600 3848 42664
rect 3912 42600 3928 42664
rect 3992 42600 4000 42664
rect 0 42584 4000 42600
rect 0 42520 8 42584
rect 72 42520 88 42584
rect 152 42520 168 42584
rect 232 42520 248 42584
rect 312 42520 328 42584
rect 392 42520 408 42584
rect 472 42520 488 42584
rect 552 42520 568 42584
rect 632 42520 648 42584
rect 712 42520 728 42584
rect 792 42520 808 42584
rect 872 42520 888 42584
rect 952 42520 968 42584
rect 1032 42520 1048 42584
rect 1112 42520 1128 42584
rect 1192 42520 1208 42584
rect 1272 42520 1288 42584
rect 1352 42520 1368 42584
rect 1432 42520 1448 42584
rect 1512 42520 1528 42584
rect 1592 42520 1608 42584
rect 1672 42520 1688 42584
rect 1752 42520 1768 42584
rect 1832 42520 1848 42584
rect 1912 42520 1928 42584
rect 1992 42520 2008 42584
rect 2072 42520 2088 42584
rect 2152 42520 2168 42584
rect 2232 42520 2248 42584
rect 2312 42520 2328 42584
rect 2392 42520 2408 42584
rect 2472 42520 2488 42584
rect 2552 42520 2568 42584
rect 2632 42520 2648 42584
rect 2712 42520 2728 42584
rect 2792 42520 2808 42584
rect 2872 42520 2888 42584
rect 2952 42520 2968 42584
rect 3032 42520 3048 42584
rect 3112 42520 3128 42584
rect 3192 42520 3208 42584
rect 3272 42520 3288 42584
rect 3352 42520 3368 42584
rect 3432 42520 3448 42584
rect 3512 42520 3528 42584
rect 3592 42520 3608 42584
rect 3672 42520 3688 42584
rect 3752 42520 3768 42584
rect 3832 42520 3848 42584
rect 3912 42520 3928 42584
rect 3992 42520 4000 42584
rect 0 42504 4000 42520
rect 0 42440 8 42504
rect 72 42440 88 42504
rect 152 42440 168 42504
rect 232 42440 248 42504
rect 312 42440 328 42504
rect 392 42440 408 42504
rect 472 42440 488 42504
rect 552 42440 568 42504
rect 632 42440 648 42504
rect 712 42440 728 42504
rect 792 42440 808 42504
rect 872 42440 888 42504
rect 952 42440 968 42504
rect 1032 42440 1048 42504
rect 1112 42440 1128 42504
rect 1192 42440 1208 42504
rect 1272 42440 1288 42504
rect 1352 42440 1368 42504
rect 1432 42440 1448 42504
rect 1512 42440 1528 42504
rect 1592 42440 1608 42504
rect 1672 42440 1688 42504
rect 1752 42440 1768 42504
rect 1832 42440 1848 42504
rect 1912 42440 1928 42504
rect 1992 42440 2008 42504
rect 2072 42440 2088 42504
rect 2152 42440 2168 42504
rect 2232 42440 2248 42504
rect 2312 42440 2328 42504
rect 2392 42440 2408 42504
rect 2472 42440 2488 42504
rect 2552 42440 2568 42504
rect 2632 42440 2648 42504
rect 2712 42440 2728 42504
rect 2792 42440 2808 42504
rect 2872 42440 2888 42504
rect 2952 42440 2968 42504
rect 3032 42440 3048 42504
rect 3112 42440 3128 42504
rect 3192 42440 3208 42504
rect 3272 42440 3288 42504
rect 3352 42440 3368 42504
rect 3432 42440 3448 42504
rect 3512 42440 3528 42504
rect 3592 42440 3608 42504
rect 3672 42440 3688 42504
rect 3752 42440 3768 42504
rect 3832 42440 3848 42504
rect 3912 42440 3928 42504
rect 3992 42440 4000 42504
rect 0 42424 4000 42440
rect 0 42360 8 42424
rect 72 42360 88 42424
rect 152 42360 168 42424
rect 232 42360 248 42424
rect 312 42360 328 42424
rect 392 42360 408 42424
rect 472 42360 488 42424
rect 552 42360 568 42424
rect 632 42360 648 42424
rect 712 42360 728 42424
rect 792 42360 808 42424
rect 872 42360 888 42424
rect 952 42360 968 42424
rect 1032 42360 1048 42424
rect 1112 42360 1128 42424
rect 1192 42360 1208 42424
rect 1272 42360 1288 42424
rect 1352 42360 1368 42424
rect 1432 42360 1448 42424
rect 1512 42360 1528 42424
rect 1592 42360 1608 42424
rect 1672 42360 1688 42424
rect 1752 42360 1768 42424
rect 1832 42360 1848 42424
rect 1912 42360 1928 42424
rect 1992 42360 2008 42424
rect 2072 42360 2088 42424
rect 2152 42360 2168 42424
rect 2232 42360 2248 42424
rect 2312 42360 2328 42424
rect 2392 42360 2408 42424
rect 2472 42360 2488 42424
rect 2552 42360 2568 42424
rect 2632 42360 2648 42424
rect 2712 42360 2728 42424
rect 2792 42360 2808 42424
rect 2872 42360 2888 42424
rect 2952 42360 2968 42424
rect 3032 42360 3048 42424
rect 3112 42360 3128 42424
rect 3192 42360 3208 42424
rect 3272 42360 3288 42424
rect 3352 42360 3368 42424
rect 3432 42360 3448 42424
rect 3512 42360 3528 42424
rect 3592 42360 3608 42424
rect 3672 42360 3688 42424
rect 3752 42360 3768 42424
rect 3832 42360 3848 42424
rect 3912 42360 3928 42424
rect 3992 42360 4000 42424
rect 0 42344 4000 42360
rect 0 42280 8 42344
rect 72 42280 88 42344
rect 152 42280 168 42344
rect 232 42280 248 42344
rect 312 42280 328 42344
rect 392 42280 408 42344
rect 472 42280 488 42344
rect 552 42280 568 42344
rect 632 42280 648 42344
rect 712 42280 728 42344
rect 792 42280 808 42344
rect 872 42280 888 42344
rect 952 42280 968 42344
rect 1032 42280 1048 42344
rect 1112 42280 1128 42344
rect 1192 42280 1208 42344
rect 1272 42280 1288 42344
rect 1352 42280 1368 42344
rect 1432 42280 1448 42344
rect 1512 42280 1528 42344
rect 1592 42280 1608 42344
rect 1672 42280 1688 42344
rect 1752 42280 1768 42344
rect 1832 42280 1848 42344
rect 1912 42280 1928 42344
rect 1992 42280 2008 42344
rect 2072 42280 2088 42344
rect 2152 42280 2168 42344
rect 2232 42280 2248 42344
rect 2312 42280 2328 42344
rect 2392 42280 2408 42344
rect 2472 42280 2488 42344
rect 2552 42280 2568 42344
rect 2632 42280 2648 42344
rect 2712 42280 2728 42344
rect 2792 42280 2808 42344
rect 2872 42280 2888 42344
rect 2952 42280 2968 42344
rect 3032 42280 3048 42344
rect 3112 42280 3128 42344
rect 3192 42280 3208 42344
rect 3272 42280 3288 42344
rect 3352 42280 3368 42344
rect 3432 42280 3448 42344
rect 3512 42280 3528 42344
rect 3592 42280 3608 42344
rect 3672 42280 3688 42344
rect 3752 42280 3768 42344
rect 3832 42280 3848 42344
rect 3912 42280 3928 42344
rect 3992 42280 4000 42344
rect 0 42264 4000 42280
rect 0 42200 8 42264
rect 72 42200 88 42264
rect 152 42200 168 42264
rect 232 42200 248 42264
rect 312 42200 328 42264
rect 392 42200 408 42264
rect 472 42200 488 42264
rect 552 42200 568 42264
rect 632 42200 648 42264
rect 712 42200 728 42264
rect 792 42200 808 42264
rect 872 42200 888 42264
rect 952 42200 968 42264
rect 1032 42200 1048 42264
rect 1112 42200 1128 42264
rect 1192 42200 1208 42264
rect 1272 42200 1288 42264
rect 1352 42200 1368 42264
rect 1432 42200 1448 42264
rect 1512 42200 1528 42264
rect 1592 42200 1608 42264
rect 1672 42200 1688 42264
rect 1752 42200 1768 42264
rect 1832 42200 1848 42264
rect 1912 42200 1928 42264
rect 1992 42200 2008 42264
rect 2072 42200 2088 42264
rect 2152 42200 2168 42264
rect 2232 42200 2248 42264
rect 2312 42200 2328 42264
rect 2392 42200 2408 42264
rect 2472 42200 2488 42264
rect 2552 42200 2568 42264
rect 2632 42200 2648 42264
rect 2712 42200 2728 42264
rect 2792 42200 2808 42264
rect 2872 42200 2888 42264
rect 2952 42200 2968 42264
rect 3032 42200 3048 42264
rect 3112 42200 3128 42264
rect 3192 42200 3208 42264
rect 3272 42200 3288 42264
rect 3352 42200 3368 42264
rect 3432 42200 3448 42264
rect 3512 42200 3528 42264
rect 3592 42200 3608 42264
rect 3672 42200 3688 42264
rect 3752 42200 3768 42264
rect 3832 42200 3848 42264
rect 3912 42200 3928 42264
rect 3992 42200 4000 42264
rect 0 42184 4000 42200
rect 0 42120 8 42184
rect 72 42120 88 42184
rect 152 42120 168 42184
rect 232 42120 248 42184
rect 312 42120 328 42184
rect 392 42120 408 42184
rect 472 42120 488 42184
rect 552 42120 568 42184
rect 632 42120 648 42184
rect 712 42120 728 42184
rect 792 42120 808 42184
rect 872 42120 888 42184
rect 952 42120 968 42184
rect 1032 42120 1048 42184
rect 1112 42120 1128 42184
rect 1192 42120 1208 42184
rect 1272 42120 1288 42184
rect 1352 42120 1368 42184
rect 1432 42120 1448 42184
rect 1512 42120 1528 42184
rect 1592 42120 1608 42184
rect 1672 42120 1688 42184
rect 1752 42120 1768 42184
rect 1832 42120 1848 42184
rect 1912 42120 1928 42184
rect 1992 42120 2008 42184
rect 2072 42120 2088 42184
rect 2152 42120 2168 42184
rect 2232 42120 2248 42184
rect 2312 42120 2328 42184
rect 2392 42120 2408 42184
rect 2472 42120 2488 42184
rect 2552 42120 2568 42184
rect 2632 42120 2648 42184
rect 2712 42120 2728 42184
rect 2792 42120 2808 42184
rect 2872 42120 2888 42184
rect 2952 42120 2968 42184
rect 3032 42120 3048 42184
rect 3112 42120 3128 42184
rect 3192 42120 3208 42184
rect 3272 42120 3288 42184
rect 3352 42120 3368 42184
rect 3432 42120 3448 42184
rect 3512 42120 3528 42184
rect 3592 42120 3608 42184
rect 3672 42120 3688 42184
rect 3752 42120 3768 42184
rect 3832 42120 3848 42184
rect 3912 42120 3928 42184
rect 3992 42120 4000 42184
rect 0 42104 4000 42120
rect 0 42040 8 42104
rect 72 42040 88 42104
rect 152 42040 168 42104
rect 232 42040 248 42104
rect 312 42040 328 42104
rect 392 42040 408 42104
rect 472 42040 488 42104
rect 552 42040 568 42104
rect 632 42040 648 42104
rect 712 42040 728 42104
rect 792 42040 808 42104
rect 872 42040 888 42104
rect 952 42040 968 42104
rect 1032 42040 1048 42104
rect 1112 42040 1128 42104
rect 1192 42040 1208 42104
rect 1272 42040 1288 42104
rect 1352 42040 1368 42104
rect 1432 42040 1448 42104
rect 1512 42040 1528 42104
rect 1592 42040 1608 42104
rect 1672 42040 1688 42104
rect 1752 42040 1768 42104
rect 1832 42040 1848 42104
rect 1912 42040 1928 42104
rect 1992 42040 2008 42104
rect 2072 42040 2088 42104
rect 2152 42040 2168 42104
rect 2232 42040 2248 42104
rect 2312 42040 2328 42104
rect 2392 42040 2408 42104
rect 2472 42040 2488 42104
rect 2552 42040 2568 42104
rect 2632 42040 2648 42104
rect 2712 42040 2728 42104
rect 2792 42040 2808 42104
rect 2872 42040 2888 42104
rect 2952 42040 2968 42104
rect 3032 42040 3048 42104
rect 3112 42040 3128 42104
rect 3192 42040 3208 42104
rect 3272 42040 3288 42104
rect 3352 42040 3368 42104
rect 3432 42040 3448 42104
rect 3512 42040 3528 42104
rect 3592 42040 3608 42104
rect 3672 42040 3688 42104
rect 3752 42040 3768 42104
rect 3832 42040 3848 42104
rect 3912 42040 3928 42104
rect 3992 42040 4000 42104
rect 0 42024 4000 42040
rect 0 41960 8 42024
rect 72 41960 88 42024
rect 152 41960 168 42024
rect 232 41960 248 42024
rect 312 41960 328 42024
rect 392 41960 408 42024
rect 472 41960 488 42024
rect 552 41960 568 42024
rect 632 41960 648 42024
rect 712 41960 728 42024
rect 792 41960 808 42024
rect 872 41960 888 42024
rect 952 41960 968 42024
rect 1032 41960 1048 42024
rect 1112 41960 1128 42024
rect 1192 41960 1208 42024
rect 1272 41960 1288 42024
rect 1352 41960 1368 42024
rect 1432 41960 1448 42024
rect 1512 41960 1528 42024
rect 1592 41960 1608 42024
rect 1672 41960 1688 42024
rect 1752 41960 1768 42024
rect 1832 41960 1848 42024
rect 1912 41960 1928 42024
rect 1992 41960 2008 42024
rect 2072 41960 2088 42024
rect 2152 41960 2168 42024
rect 2232 41960 2248 42024
rect 2312 41960 2328 42024
rect 2392 41960 2408 42024
rect 2472 41960 2488 42024
rect 2552 41960 2568 42024
rect 2632 41960 2648 42024
rect 2712 41960 2728 42024
rect 2792 41960 2808 42024
rect 2872 41960 2888 42024
rect 2952 41960 2968 42024
rect 3032 41960 3048 42024
rect 3112 41960 3128 42024
rect 3192 41960 3208 42024
rect 3272 41960 3288 42024
rect 3352 41960 3368 42024
rect 3432 41960 3448 42024
rect 3512 41960 3528 42024
rect 3592 41960 3608 42024
rect 3672 41960 3688 42024
rect 3752 41960 3768 42024
rect 3832 41960 3848 42024
rect 3912 41960 3928 42024
rect 3992 41960 4000 42024
rect 0 41944 4000 41960
rect 0 41880 8 41944
rect 72 41880 88 41944
rect 152 41880 168 41944
rect 232 41880 248 41944
rect 312 41880 328 41944
rect 392 41880 408 41944
rect 472 41880 488 41944
rect 552 41880 568 41944
rect 632 41880 648 41944
rect 712 41880 728 41944
rect 792 41880 808 41944
rect 872 41880 888 41944
rect 952 41880 968 41944
rect 1032 41880 1048 41944
rect 1112 41880 1128 41944
rect 1192 41880 1208 41944
rect 1272 41880 1288 41944
rect 1352 41880 1368 41944
rect 1432 41880 1448 41944
rect 1512 41880 1528 41944
rect 1592 41880 1608 41944
rect 1672 41880 1688 41944
rect 1752 41880 1768 41944
rect 1832 41880 1848 41944
rect 1912 41880 1928 41944
rect 1992 41880 2008 41944
rect 2072 41880 2088 41944
rect 2152 41880 2168 41944
rect 2232 41880 2248 41944
rect 2312 41880 2328 41944
rect 2392 41880 2408 41944
rect 2472 41880 2488 41944
rect 2552 41880 2568 41944
rect 2632 41880 2648 41944
rect 2712 41880 2728 41944
rect 2792 41880 2808 41944
rect 2872 41880 2888 41944
rect 2952 41880 2968 41944
rect 3032 41880 3048 41944
rect 3112 41880 3128 41944
rect 3192 41880 3208 41944
rect 3272 41880 3288 41944
rect 3352 41880 3368 41944
rect 3432 41880 3448 41944
rect 3512 41880 3528 41944
rect 3592 41880 3608 41944
rect 3672 41880 3688 41944
rect 3752 41880 3768 41944
rect 3832 41880 3848 41944
rect 3912 41880 3928 41944
rect 3992 41880 4000 41944
rect 0 41864 4000 41880
rect 0 41800 8 41864
rect 72 41800 88 41864
rect 152 41800 168 41864
rect 232 41800 248 41864
rect 312 41800 328 41864
rect 392 41800 408 41864
rect 472 41800 488 41864
rect 552 41800 568 41864
rect 632 41800 648 41864
rect 712 41800 728 41864
rect 792 41800 808 41864
rect 872 41800 888 41864
rect 952 41800 968 41864
rect 1032 41800 1048 41864
rect 1112 41800 1128 41864
rect 1192 41800 1208 41864
rect 1272 41800 1288 41864
rect 1352 41800 1368 41864
rect 1432 41800 1448 41864
rect 1512 41800 1528 41864
rect 1592 41800 1608 41864
rect 1672 41800 1688 41864
rect 1752 41800 1768 41864
rect 1832 41800 1848 41864
rect 1912 41800 1928 41864
rect 1992 41800 2008 41864
rect 2072 41800 2088 41864
rect 2152 41800 2168 41864
rect 2232 41800 2248 41864
rect 2312 41800 2328 41864
rect 2392 41800 2408 41864
rect 2472 41800 2488 41864
rect 2552 41800 2568 41864
rect 2632 41800 2648 41864
rect 2712 41800 2728 41864
rect 2792 41800 2808 41864
rect 2872 41800 2888 41864
rect 2952 41800 2968 41864
rect 3032 41800 3048 41864
rect 3112 41800 3128 41864
rect 3192 41800 3208 41864
rect 3272 41800 3288 41864
rect 3352 41800 3368 41864
rect 3432 41800 3448 41864
rect 3512 41800 3528 41864
rect 3592 41800 3608 41864
rect 3672 41800 3688 41864
rect 3752 41800 3768 41864
rect 3832 41800 3848 41864
rect 3912 41800 3928 41864
rect 3992 41800 4000 41864
rect 0 41784 4000 41800
rect 0 41720 8 41784
rect 72 41720 88 41784
rect 152 41720 168 41784
rect 232 41720 248 41784
rect 312 41720 328 41784
rect 392 41720 408 41784
rect 472 41720 488 41784
rect 552 41720 568 41784
rect 632 41720 648 41784
rect 712 41720 728 41784
rect 792 41720 808 41784
rect 872 41720 888 41784
rect 952 41720 968 41784
rect 1032 41720 1048 41784
rect 1112 41720 1128 41784
rect 1192 41720 1208 41784
rect 1272 41720 1288 41784
rect 1352 41720 1368 41784
rect 1432 41720 1448 41784
rect 1512 41720 1528 41784
rect 1592 41720 1608 41784
rect 1672 41720 1688 41784
rect 1752 41720 1768 41784
rect 1832 41720 1848 41784
rect 1912 41720 1928 41784
rect 1992 41720 2008 41784
rect 2072 41720 2088 41784
rect 2152 41720 2168 41784
rect 2232 41720 2248 41784
rect 2312 41720 2328 41784
rect 2392 41720 2408 41784
rect 2472 41720 2488 41784
rect 2552 41720 2568 41784
rect 2632 41720 2648 41784
rect 2712 41720 2728 41784
rect 2792 41720 2808 41784
rect 2872 41720 2888 41784
rect 2952 41720 2968 41784
rect 3032 41720 3048 41784
rect 3112 41720 3128 41784
rect 3192 41720 3208 41784
rect 3272 41720 3288 41784
rect 3352 41720 3368 41784
rect 3432 41720 3448 41784
rect 3512 41720 3528 41784
rect 3592 41720 3608 41784
rect 3672 41720 3688 41784
rect 3752 41720 3768 41784
rect 3832 41720 3848 41784
rect 3912 41720 3928 41784
rect 3992 41720 4000 41784
rect 0 41704 4000 41720
rect 0 41640 8 41704
rect 72 41640 88 41704
rect 152 41640 168 41704
rect 232 41640 248 41704
rect 312 41640 328 41704
rect 392 41640 408 41704
rect 472 41640 488 41704
rect 552 41640 568 41704
rect 632 41640 648 41704
rect 712 41640 728 41704
rect 792 41640 808 41704
rect 872 41640 888 41704
rect 952 41640 968 41704
rect 1032 41640 1048 41704
rect 1112 41640 1128 41704
rect 1192 41640 1208 41704
rect 1272 41640 1288 41704
rect 1352 41640 1368 41704
rect 1432 41640 1448 41704
rect 1512 41640 1528 41704
rect 1592 41640 1608 41704
rect 1672 41640 1688 41704
rect 1752 41640 1768 41704
rect 1832 41640 1848 41704
rect 1912 41640 1928 41704
rect 1992 41640 2008 41704
rect 2072 41640 2088 41704
rect 2152 41640 2168 41704
rect 2232 41640 2248 41704
rect 2312 41640 2328 41704
rect 2392 41640 2408 41704
rect 2472 41640 2488 41704
rect 2552 41640 2568 41704
rect 2632 41640 2648 41704
rect 2712 41640 2728 41704
rect 2792 41640 2808 41704
rect 2872 41640 2888 41704
rect 2952 41640 2968 41704
rect 3032 41640 3048 41704
rect 3112 41640 3128 41704
rect 3192 41640 3208 41704
rect 3272 41640 3288 41704
rect 3352 41640 3368 41704
rect 3432 41640 3448 41704
rect 3512 41640 3528 41704
rect 3592 41640 3608 41704
rect 3672 41640 3688 41704
rect 3752 41640 3768 41704
rect 3832 41640 3848 41704
rect 3912 41640 3928 41704
rect 3992 41640 4000 41704
rect 0 41624 4000 41640
rect 0 41560 8 41624
rect 72 41560 88 41624
rect 152 41560 168 41624
rect 232 41560 248 41624
rect 312 41560 328 41624
rect 392 41560 408 41624
rect 472 41560 488 41624
rect 552 41560 568 41624
rect 632 41560 648 41624
rect 712 41560 728 41624
rect 792 41560 808 41624
rect 872 41560 888 41624
rect 952 41560 968 41624
rect 1032 41560 1048 41624
rect 1112 41560 1128 41624
rect 1192 41560 1208 41624
rect 1272 41560 1288 41624
rect 1352 41560 1368 41624
rect 1432 41560 1448 41624
rect 1512 41560 1528 41624
rect 1592 41560 1608 41624
rect 1672 41560 1688 41624
rect 1752 41560 1768 41624
rect 1832 41560 1848 41624
rect 1912 41560 1928 41624
rect 1992 41560 2008 41624
rect 2072 41560 2088 41624
rect 2152 41560 2168 41624
rect 2232 41560 2248 41624
rect 2312 41560 2328 41624
rect 2392 41560 2408 41624
rect 2472 41560 2488 41624
rect 2552 41560 2568 41624
rect 2632 41560 2648 41624
rect 2712 41560 2728 41624
rect 2792 41560 2808 41624
rect 2872 41560 2888 41624
rect 2952 41560 2968 41624
rect 3032 41560 3048 41624
rect 3112 41560 3128 41624
rect 3192 41560 3208 41624
rect 3272 41560 3288 41624
rect 3352 41560 3368 41624
rect 3432 41560 3448 41624
rect 3512 41560 3528 41624
rect 3592 41560 3608 41624
rect 3672 41560 3688 41624
rect 3752 41560 3768 41624
rect 3832 41560 3848 41624
rect 3912 41560 3928 41624
rect 3992 41560 4000 41624
rect 0 41544 4000 41560
rect 0 41480 8 41544
rect 72 41480 88 41544
rect 152 41480 168 41544
rect 232 41480 248 41544
rect 312 41480 328 41544
rect 392 41480 408 41544
rect 472 41480 488 41544
rect 552 41480 568 41544
rect 632 41480 648 41544
rect 712 41480 728 41544
rect 792 41480 808 41544
rect 872 41480 888 41544
rect 952 41480 968 41544
rect 1032 41480 1048 41544
rect 1112 41480 1128 41544
rect 1192 41480 1208 41544
rect 1272 41480 1288 41544
rect 1352 41480 1368 41544
rect 1432 41480 1448 41544
rect 1512 41480 1528 41544
rect 1592 41480 1608 41544
rect 1672 41480 1688 41544
rect 1752 41480 1768 41544
rect 1832 41480 1848 41544
rect 1912 41480 1928 41544
rect 1992 41480 2008 41544
rect 2072 41480 2088 41544
rect 2152 41480 2168 41544
rect 2232 41480 2248 41544
rect 2312 41480 2328 41544
rect 2392 41480 2408 41544
rect 2472 41480 2488 41544
rect 2552 41480 2568 41544
rect 2632 41480 2648 41544
rect 2712 41480 2728 41544
rect 2792 41480 2808 41544
rect 2872 41480 2888 41544
rect 2952 41480 2968 41544
rect 3032 41480 3048 41544
rect 3112 41480 3128 41544
rect 3192 41480 3208 41544
rect 3272 41480 3288 41544
rect 3352 41480 3368 41544
rect 3432 41480 3448 41544
rect 3512 41480 3528 41544
rect 3592 41480 3608 41544
rect 3672 41480 3688 41544
rect 3752 41480 3768 41544
rect 3832 41480 3848 41544
rect 3912 41480 3928 41544
rect 3992 41480 4000 41544
rect 0 41464 4000 41480
rect 0 41400 8 41464
rect 72 41400 88 41464
rect 152 41400 168 41464
rect 232 41400 248 41464
rect 312 41400 328 41464
rect 392 41400 408 41464
rect 472 41400 488 41464
rect 552 41400 568 41464
rect 632 41400 648 41464
rect 712 41400 728 41464
rect 792 41400 808 41464
rect 872 41400 888 41464
rect 952 41400 968 41464
rect 1032 41400 1048 41464
rect 1112 41400 1128 41464
rect 1192 41400 1208 41464
rect 1272 41400 1288 41464
rect 1352 41400 1368 41464
rect 1432 41400 1448 41464
rect 1512 41400 1528 41464
rect 1592 41400 1608 41464
rect 1672 41400 1688 41464
rect 1752 41400 1768 41464
rect 1832 41400 1848 41464
rect 1912 41400 1928 41464
rect 1992 41400 2008 41464
rect 2072 41400 2088 41464
rect 2152 41400 2168 41464
rect 2232 41400 2248 41464
rect 2312 41400 2328 41464
rect 2392 41400 2408 41464
rect 2472 41400 2488 41464
rect 2552 41400 2568 41464
rect 2632 41400 2648 41464
rect 2712 41400 2728 41464
rect 2792 41400 2808 41464
rect 2872 41400 2888 41464
rect 2952 41400 2968 41464
rect 3032 41400 3048 41464
rect 3112 41400 3128 41464
rect 3192 41400 3208 41464
rect 3272 41400 3288 41464
rect 3352 41400 3368 41464
rect 3432 41400 3448 41464
rect 3512 41400 3528 41464
rect 3592 41400 3608 41464
rect 3672 41400 3688 41464
rect 3752 41400 3768 41464
rect 3832 41400 3848 41464
rect 3912 41400 3928 41464
rect 3992 41400 4000 41464
rect 0 3992 4000 41400
rect 5000 40384 9000 40392
rect 5000 40320 5008 40384
rect 5072 40320 5088 40384
rect 5152 40320 5168 40384
rect 5232 40320 5248 40384
rect 5312 40320 5328 40384
rect 5392 40320 5408 40384
rect 5472 40320 5488 40384
rect 5552 40320 5568 40384
rect 5632 40320 5648 40384
rect 5712 40320 5728 40384
rect 5792 40320 5808 40384
rect 5872 40320 5888 40384
rect 5952 40320 5968 40384
rect 6032 40320 6048 40384
rect 6112 40320 6128 40384
rect 6192 40320 6208 40384
rect 6272 40320 6288 40384
rect 6352 40320 6368 40384
rect 6432 40320 6448 40384
rect 6512 40320 6528 40384
rect 6592 40320 6608 40384
rect 6672 40320 6688 40384
rect 6752 40320 6768 40384
rect 6832 40320 6848 40384
rect 6912 40320 6928 40384
rect 6992 40320 7008 40384
rect 7072 40320 7088 40384
rect 7152 40320 7168 40384
rect 7232 40320 7248 40384
rect 7312 40320 7328 40384
rect 7392 40320 7408 40384
rect 7472 40320 7488 40384
rect 7552 40320 7568 40384
rect 7632 40320 7648 40384
rect 7712 40320 7728 40384
rect 7792 40320 7808 40384
rect 7872 40320 7888 40384
rect 7952 40320 7968 40384
rect 8032 40320 8048 40384
rect 8112 40320 8128 40384
rect 8192 40320 8208 40384
rect 8272 40320 8288 40384
rect 8352 40320 8368 40384
rect 8432 40320 8448 40384
rect 8512 40320 8528 40384
rect 8592 40320 8608 40384
rect 8672 40320 8688 40384
rect 8752 40320 8768 40384
rect 8832 40320 8848 40384
rect 8912 40320 8928 40384
rect 8992 40320 9000 40384
rect 5000 40304 9000 40320
rect 5000 40240 5008 40304
rect 5072 40240 5088 40304
rect 5152 40240 5168 40304
rect 5232 40240 5248 40304
rect 5312 40240 5328 40304
rect 5392 40240 5408 40304
rect 5472 40240 5488 40304
rect 5552 40240 5568 40304
rect 5632 40240 5648 40304
rect 5712 40240 5728 40304
rect 5792 40240 5808 40304
rect 5872 40240 5888 40304
rect 5952 40240 5968 40304
rect 6032 40240 6048 40304
rect 6112 40240 6128 40304
rect 6192 40240 6208 40304
rect 6272 40240 6288 40304
rect 6352 40240 6368 40304
rect 6432 40240 6448 40304
rect 6512 40240 6528 40304
rect 6592 40240 6608 40304
rect 6672 40240 6688 40304
rect 6752 40240 6768 40304
rect 6832 40240 6848 40304
rect 6912 40240 6928 40304
rect 6992 40240 7008 40304
rect 7072 40240 7088 40304
rect 7152 40240 7168 40304
rect 7232 40240 7248 40304
rect 7312 40240 7328 40304
rect 7392 40240 7408 40304
rect 7472 40240 7488 40304
rect 7552 40240 7568 40304
rect 7632 40240 7648 40304
rect 7712 40240 7728 40304
rect 7792 40240 7808 40304
rect 7872 40240 7888 40304
rect 7952 40240 7968 40304
rect 8032 40240 8048 40304
rect 8112 40240 8128 40304
rect 8192 40240 8208 40304
rect 8272 40240 8288 40304
rect 8352 40240 8368 40304
rect 8432 40240 8448 40304
rect 8512 40240 8528 40304
rect 8592 40240 8608 40304
rect 8672 40240 8688 40304
rect 8752 40240 8768 40304
rect 8832 40240 8848 40304
rect 8912 40240 8928 40304
rect 8992 40240 9000 40304
rect 5000 40224 9000 40240
rect 5000 40160 5008 40224
rect 5072 40160 5088 40224
rect 5152 40160 5168 40224
rect 5232 40160 5248 40224
rect 5312 40160 5328 40224
rect 5392 40160 5408 40224
rect 5472 40160 5488 40224
rect 5552 40160 5568 40224
rect 5632 40160 5648 40224
rect 5712 40160 5728 40224
rect 5792 40160 5808 40224
rect 5872 40160 5888 40224
rect 5952 40160 5968 40224
rect 6032 40160 6048 40224
rect 6112 40160 6128 40224
rect 6192 40160 6208 40224
rect 6272 40160 6288 40224
rect 6352 40160 6368 40224
rect 6432 40160 6448 40224
rect 6512 40160 6528 40224
rect 6592 40160 6608 40224
rect 6672 40160 6688 40224
rect 6752 40160 6768 40224
rect 6832 40160 6848 40224
rect 6912 40160 6928 40224
rect 6992 40160 7008 40224
rect 7072 40160 7088 40224
rect 7152 40160 7168 40224
rect 7232 40160 7248 40224
rect 7312 40160 7328 40224
rect 7392 40160 7408 40224
rect 7472 40160 7488 40224
rect 7552 40160 7568 40224
rect 7632 40160 7648 40224
rect 7712 40160 7728 40224
rect 7792 40160 7808 40224
rect 7872 40160 7888 40224
rect 7952 40160 7968 40224
rect 8032 40160 8048 40224
rect 8112 40160 8128 40224
rect 8192 40160 8208 40224
rect 8272 40160 8288 40224
rect 8352 40160 8368 40224
rect 8432 40160 8448 40224
rect 8512 40160 8528 40224
rect 8592 40160 8608 40224
rect 8672 40160 8688 40224
rect 8752 40160 8768 40224
rect 8832 40160 8848 40224
rect 8912 40160 8928 40224
rect 8992 40160 9000 40224
rect 5000 40144 9000 40160
rect 5000 40080 5008 40144
rect 5072 40080 5088 40144
rect 5152 40080 5168 40144
rect 5232 40080 5248 40144
rect 5312 40080 5328 40144
rect 5392 40080 5408 40144
rect 5472 40080 5488 40144
rect 5552 40080 5568 40144
rect 5632 40080 5648 40144
rect 5712 40080 5728 40144
rect 5792 40080 5808 40144
rect 5872 40080 5888 40144
rect 5952 40080 5968 40144
rect 6032 40080 6048 40144
rect 6112 40080 6128 40144
rect 6192 40080 6208 40144
rect 6272 40080 6288 40144
rect 6352 40080 6368 40144
rect 6432 40080 6448 40144
rect 6512 40080 6528 40144
rect 6592 40080 6608 40144
rect 6672 40080 6688 40144
rect 6752 40080 6768 40144
rect 6832 40080 6848 40144
rect 6912 40080 6928 40144
rect 6992 40080 7008 40144
rect 7072 40080 7088 40144
rect 7152 40080 7168 40144
rect 7232 40080 7248 40144
rect 7312 40080 7328 40144
rect 7392 40080 7408 40144
rect 7472 40080 7488 40144
rect 7552 40080 7568 40144
rect 7632 40080 7648 40144
rect 7712 40080 7728 40144
rect 7792 40080 7808 40144
rect 7872 40080 7888 40144
rect 7952 40080 7968 40144
rect 8032 40080 8048 40144
rect 8112 40080 8128 40144
rect 8192 40080 8208 40144
rect 8272 40080 8288 40144
rect 8352 40080 8368 40144
rect 8432 40080 8448 40144
rect 8512 40080 8528 40144
rect 8592 40080 8608 40144
rect 8672 40080 8688 40144
rect 8752 40080 8768 40144
rect 8832 40080 8848 40144
rect 8912 40080 8928 40144
rect 8992 40080 9000 40144
rect 5000 40064 9000 40080
rect 5000 40000 5008 40064
rect 5072 40000 5088 40064
rect 5152 40000 5168 40064
rect 5232 40000 5248 40064
rect 5312 40000 5328 40064
rect 5392 40000 5408 40064
rect 5472 40000 5488 40064
rect 5552 40000 5568 40064
rect 5632 40000 5648 40064
rect 5712 40000 5728 40064
rect 5792 40000 5808 40064
rect 5872 40000 5888 40064
rect 5952 40000 5968 40064
rect 6032 40000 6048 40064
rect 6112 40000 6128 40064
rect 6192 40000 6208 40064
rect 6272 40000 6288 40064
rect 6352 40000 6368 40064
rect 6432 40000 6448 40064
rect 6512 40000 6528 40064
rect 6592 40000 6608 40064
rect 6672 40000 6688 40064
rect 6752 40000 6768 40064
rect 6832 40000 6848 40064
rect 6912 40000 6928 40064
rect 6992 40000 7008 40064
rect 7072 40000 7088 40064
rect 7152 40000 7168 40064
rect 7232 40000 7248 40064
rect 7312 40000 7328 40064
rect 7392 40000 7408 40064
rect 7472 40000 7488 40064
rect 7552 40000 7568 40064
rect 7632 40000 7648 40064
rect 7712 40000 7728 40064
rect 7792 40000 7808 40064
rect 7872 40000 7888 40064
rect 7952 40000 7968 40064
rect 8032 40000 8048 40064
rect 8112 40000 8128 40064
rect 8192 40000 8208 40064
rect 8272 40000 8288 40064
rect 8352 40000 8368 40064
rect 8432 40000 8448 40064
rect 8512 40000 8528 40064
rect 8592 40000 8608 40064
rect 8672 40000 8688 40064
rect 8752 40000 8768 40064
rect 8832 40000 8848 40064
rect 8912 40000 8928 40064
rect 8992 40000 9000 40064
rect 5000 39984 9000 40000
rect 5000 39920 5008 39984
rect 5072 39920 5088 39984
rect 5152 39920 5168 39984
rect 5232 39920 5248 39984
rect 5312 39920 5328 39984
rect 5392 39920 5408 39984
rect 5472 39920 5488 39984
rect 5552 39920 5568 39984
rect 5632 39920 5648 39984
rect 5712 39920 5728 39984
rect 5792 39920 5808 39984
rect 5872 39920 5888 39984
rect 5952 39920 5968 39984
rect 6032 39920 6048 39984
rect 6112 39920 6128 39984
rect 6192 39920 6208 39984
rect 6272 39920 6288 39984
rect 6352 39920 6368 39984
rect 6432 39920 6448 39984
rect 6512 39920 6528 39984
rect 6592 39920 6608 39984
rect 6672 39920 6688 39984
rect 6752 39920 6768 39984
rect 6832 39920 6848 39984
rect 6912 39920 6928 39984
rect 6992 39920 7008 39984
rect 7072 39920 7088 39984
rect 7152 39920 7168 39984
rect 7232 39920 7248 39984
rect 7312 39920 7328 39984
rect 7392 39920 7408 39984
rect 7472 39920 7488 39984
rect 7552 39920 7568 39984
rect 7632 39920 7648 39984
rect 7712 39920 7728 39984
rect 7792 39920 7808 39984
rect 7872 39920 7888 39984
rect 7952 39920 7968 39984
rect 8032 39920 8048 39984
rect 8112 39920 8128 39984
rect 8192 39920 8208 39984
rect 8272 39920 8288 39984
rect 8352 39920 8368 39984
rect 8432 39920 8448 39984
rect 8512 39920 8528 39984
rect 8592 39920 8608 39984
rect 8672 39920 8688 39984
rect 8752 39920 8768 39984
rect 8832 39920 8848 39984
rect 8912 39920 8928 39984
rect 8992 39920 9000 39984
rect 5000 39904 9000 39920
rect 5000 39840 5008 39904
rect 5072 39840 5088 39904
rect 5152 39840 5168 39904
rect 5232 39840 5248 39904
rect 5312 39840 5328 39904
rect 5392 39840 5408 39904
rect 5472 39840 5488 39904
rect 5552 39840 5568 39904
rect 5632 39840 5648 39904
rect 5712 39840 5728 39904
rect 5792 39840 5808 39904
rect 5872 39840 5888 39904
rect 5952 39840 5968 39904
rect 6032 39840 6048 39904
rect 6112 39840 6128 39904
rect 6192 39840 6208 39904
rect 6272 39840 6288 39904
rect 6352 39840 6368 39904
rect 6432 39840 6448 39904
rect 6512 39840 6528 39904
rect 6592 39840 6608 39904
rect 6672 39840 6688 39904
rect 6752 39840 6768 39904
rect 6832 39840 6848 39904
rect 6912 39840 6928 39904
rect 6992 39840 7008 39904
rect 7072 39840 7088 39904
rect 7152 39840 7168 39904
rect 7232 39840 7248 39904
rect 7312 39840 7328 39904
rect 7392 39840 7408 39904
rect 7472 39840 7488 39904
rect 7552 39840 7568 39904
rect 7632 39840 7648 39904
rect 7712 39840 7728 39904
rect 7792 39840 7808 39904
rect 7872 39840 7888 39904
rect 7952 39840 7968 39904
rect 8032 39840 8048 39904
rect 8112 39840 8128 39904
rect 8192 39840 8208 39904
rect 8272 39840 8288 39904
rect 8352 39840 8368 39904
rect 8432 39840 8448 39904
rect 8512 39840 8528 39904
rect 8592 39840 8608 39904
rect 8672 39840 8688 39904
rect 8752 39840 8768 39904
rect 8832 39840 8848 39904
rect 8912 39840 8928 39904
rect 8992 39840 9000 39904
rect 5000 39824 9000 39840
rect 5000 39760 5008 39824
rect 5072 39760 5088 39824
rect 5152 39760 5168 39824
rect 5232 39760 5248 39824
rect 5312 39760 5328 39824
rect 5392 39760 5408 39824
rect 5472 39760 5488 39824
rect 5552 39760 5568 39824
rect 5632 39760 5648 39824
rect 5712 39760 5728 39824
rect 5792 39760 5808 39824
rect 5872 39760 5888 39824
rect 5952 39760 5968 39824
rect 6032 39760 6048 39824
rect 6112 39760 6128 39824
rect 6192 39760 6208 39824
rect 6272 39760 6288 39824
rect 6352 39760 6368 39824
rect 6432 39760 6448 39824
rect 6512 39760 6528 39824
rect 6592 39760 6608 39824
rect 6672 39760 6688 39824
rect 6752 39760 6768 39824
rect 6832 39760 6848 39824
rect 6912 39760 6928 39824
rect 6992 39760 7008 39824
rect 7072 39760 7088 39824
rect 7152 39760 7168 39824
rect 7232 39760 7248 39824
rect 7312 39760 7328 39824
rect 7392 39760 7408 39824
rect 7472 39760 7488 39824
rect 7552 39760 7568 39824
rect 7632 39760 7648 39824
rect 7712 39760 7728 39824
rect 7792 39760 7808 39824
rect 7872 39760 7888 39824
rect 7952 39760 7968 39824
rect 8032 39760 8048 39824
rect 8112 39760 8128 39824
rect 8192 39760 8208 39824
rect 8272 39760 8288 39824
rect 8352 39760 8368 39824
rect 8432 39760 8448 39824
rect 8512 39760 8528 39824
rect 8592 39760 8608 39824
rect 8672 39760 8688 39824
rect 8752 39760 8768 39824
rect 8832 39760 8848 39824
rect 8912 39760 8928 39824
rect 8992 39760 9000 39824
rect 5000 39744 9000 39760
rect 5000 39680 5008 39744
rect 5072 39680 5088 39744
rect 5152 39680 5168 39744
rect 5232 39680 5248 39744
rect 5312 39680 5328 39744
rect 5392 39680 5408 39744
rect 5472 39680 5488 39744
rect 5552 39680 5568 39744
rect 5632 39680 5648 39744
rect 5712 39680 5728 39744
rect 5792 39680 5808 39744
rect 5872 39680 5888 39744
rect 5952 39680 5968 39744
rect 6032 39680 6048 39744
rect 6112 39680 6128 39744
rect 6192 39680 6208 39744
rect 6272 39680 6288 39744
rect 6352 39680 6368 39744
rect 6432 39680 6448 39744
rect 6512 39680 6528 39744
rect 6592 39680 6608 39744
rect 6672 39680 6688 39744
rect 6752 39680 6768 39744
rect 6832 39680 6848 39744
rect 6912 39680 6928 39744
rect 6992 39680 7008 39744
rect 7072 39680 7088 39744
rect 7152 39680 7168 39744
rect 7232 39680 7248 39744
rect 7312 39680 7328 39744
rect 7392 39680 7408 39744
rect 7472 39680 7488 39744
rect 7552 39680 7568 39744
rect 7632 39680 7648 39744
rect 7712 39680 7728 39744
rect 7792 39680 7808 39744
rect 7872 39680 7888 39744
rect 7952 39680 7968 39744
rect 8032 39680 8048 39744
rect 8112 39680 8128 39744
rect 8192 39680 8208 39744
rect 8272 39680 8288 39744
rect 8352 39680 8368 39744
rect 8432 39680 8448 39744
rect 8512 39680 8528 39744
rect 8592 39680 8608 39744
rect 8672 39680 8688 39744
rect 8752 39680 8768 39744
rect 8832 39680 8848 39744
rect 8912 39680 8928 39744
rect 8992 39680 9000 39744
rect 5000 39664 9000 39680
rect 5000 39600 5008 39664
rect 5072 39600 5088 39664
rect 5152 39600 5168 39664
rect 5232 39600 5248 39664
rect 5312 39600 5328 39664
rect 5392 39600 5408 39664
rect 5472 39600 5488 39664
rect 5552 39600 5568 39664
rect 5632 39600 5648 39664
rect 5712 39600 5728 39664
rect 5792 39600 5808 39664
rect 5872 39600 5888 39664
rect 5952 39600 5968 39664
rect 6032 39600 6048 39664
rect 6112 39600 6128 39664
rect 6192 39600 6208 39664
rect 6272 39600 6288 39664
rect 6352 39600 6368 39664
rect 6432 39600 6448 39664
rect 6512 39600 6528 39664
rect 6592 39600 6608 39664
rect 6672 39600 6688 39664
rect 6752 39600 6768 39664
rect 6832 39600 6848 39664
rect 6912 39600 6928 39664
rect 6992 39600 7008 39664
rect 7072 39600 7088 39664
rect 7152 39600 7168 39664
rect 7232 39600 7248 39664
rect 7312 39600 7328 39664
rect 7392 39600 7408 39664
rect 7472 39600 7488 39664
rect 7552 39600 7568 39664
rect 7632 39600 7648 39664
rect 7712 39600 7728 39664
rect 7792 39600 7808 39664
rect 7872 39600 7888 39664
rect 7952 39600 7968 39664
rect 8032 39600 8048 39664
rect 8112 39600 8128 39664
rect 8192 39600 8208 39664
rect 8272 39600 8288 39664
rect 8352 39600 8368 39664
rect 8432 39600 8448 39664
rect 8512 39600 8528 39664
rect 8592 39600 8608 39664
rect 8672 39600 8688 39664
rect 8752 39600 8768 39664
rect 8832 39600 8848 39664
rect 8912 39600 8928 39664
rect 8992 39600 9000 39664
rect 5000 39584 9000 39600
rect 5000 39520 5008 39584
rect 5072 39520 5088 39584
rect 5152 39520 5168 39584
rect 5232 39520 5248 39584
rect 5312 39520 5328 39584
rect 5392 39520 5408 39584
rect 5472 39520 5488 39584
rect 5552 39520 5568 39584
rect 5632 39520 5648 39584
rect 5712 39520 5728 39584
rect 5792 39520 5808 39584
rect 5872 39520 5888 39584
rect 5952 39520 5968 39584
rect 6032 39520 6048 39584
rect 6112 39520 6128 39584
rect 6192 39520 6208 39584
rect 6272 39520 6288 39584
rect 6352 39520 6368 39584
rect 6432 39520 6448 39584
rect 6512 39520 6528 39584
rect 6592 39520 6608 39584
rect 6672 39520 6688 39584
rect 6752 39520 6768 39584
rect 6832 39520 6848 39584
rect 6912 39520 6928 39584
rect 6992 39520 7008 39584
rect 7072 39520 7088 39584
rect 7152 39520 7168 39584
rect 7232 39520 7248 39584
rect 7312 39520 7328 39584
rect 7392 39520 7408 39584
rect 7472 39520 7488 39584
rect 7552 39520 7568 39584
rect 7632 39520 7648 39584
rect 7712 39520 7728 39584
rect 7792 39520 7808 39584
rect 7872 39520 7888 39584
rect 7952 39520 7968 39584
rect 8032 39520 8048 39584
rect 8112 39520 8128 39584
rect 8192 39520 8208 39584
rect 8272 39520 8288 39584
rect 8352 39520 8368 39584
rect 8432 39520 8448 39584
rect 8512 39520 8528 39584
rect 8592 39520 8608 39584
rect 8672 39520 8688 39584
rect 8752 39520 8768 39584
rect 8832 39520 8848 39584
rect 8912 39520 8928 39584
rect 8992 39520 9000 39584
rect 5000 39504 9000 39520
rect 5000 39440 5008 39504
rect 5072 39440 5088 39504
rect 5152 39440 5168 39504
rect 5232 39440 5248 39504
rect 5312 39440 5328 39504
rect 5392 39440 5408 39504
rect 5472 39440 5488 39504
rect 5552 39440 5568 39504
rect 5632 39440 5648 39504
rect 5712 39440 5728 39504
rect 5792 39440 5808 39504
rect 5872 39440 5888 39504
rect 5952 39440 5968 39504
rect 6032 39440 6048 39504
rect 6112 39440 6128 39504
rect 6192 39440 6208 39504
rect 6272 39440 6288 39504
rect 6352 39440 6368 39504
rect 6432 39440 6448 39504
rect 6512 39440 6528 39504
rect 6592 39440 6608 39504
rect 6672 39440 6688 39504
rect 6752 39440 6768 39504
rect 6832 39440 6848 39504
rect 6912 39440 6928 39504
rect 6992 39440 7008 39504
rect 7072 39440 7088 39504
rect 7152 39440 7168 39504
rect 7232 39440 7248 39504
rect 7312 39440 7328 39504
rect 7392 39440 7408 39504
rect 7472 39440 7488 39504
rect 7552 39440 7568 39504
rect 7632 39440 7648 39504
rect 7712 39440 7728 39504
rect 7792 39440 7808 39504
rect 7872 39440 7888 39504
rect 7952 39440 7968 39504
rect 8032 39440 8048 39504
rect 8112 39440 8128 39504
rect 8192 39440 8208 39504
rect 8272 39440 8288 39504
rect 8352 39440 8368 39504
rect 8432 39440 8448 39504
rect 8512 39440 8528 39504
rect 8592 39440 8608 39504
rect 8672 39440 8688 39504
rect 8752 39440 8768 39504
rect 8832 39440 8848 39504
rect 8912 39440 8928 39504
rect 8992 39440 9000 39504
rect 5000 39424 9000 39440
rect 5000 39360 5008 39424
rect 5072 39360 5088 39424
rect 5152 39360 5168 39424
rect 5232 39360 5248 39424
rect 5312 39360 5328 39424
rect 5392 39360 5408 39424
rect 5472 39360 5488 39424
rect 5552 39360 5568 39424
rect 5632 39360 5648 39424
rect 5712 39360 5728 39424
rect 5792 39360 5808 39424
rect 5872 39360 5888 39424
rect 5952 39360 5968 39424
rect 6032 39360 6048 39424
rect 6112 39360 6128 39424
rect 6192 39360 6208 39424
rect 6272 39360 6288 39424
rect 6352 39360 6368 39424
rect 6432 39360 6448 39424
rect 6512 39360 6528 39424
rect 6592 39360 6608 39424
rect 6672 39360 6688 39424
rect 6752 39360 6768 39424
rect 6832 39360 6848 39424
rect 6912 39360 6928 39424
rect 6992 39360 7008 39424
rect 7072 39360 7088 39424
rect 7152 39360 7168 39424
rect 7232 39360 7248 39424
rect 7312 39360 7328 39424
rect 7392 39360 7408 39424
rect 7472 39360 7488 39424
rect 7552 39360 7568 39424
rect 7632 39360 7648 39424
rect 7712 39360 7728 39424
rect 7792 39360 7808 39424
rect 7872 39360 7888 39424
rect 7952 39360 7968 39424
rect 8032 39360 8048 39424
rect 8112 39360 8128 39424
rect 8192 39360 8208 39424
rect 8272 39360 8288 39424
rect 8352 39360 8368 39424
rect 8432 39360 8448 39424
rect 8512 39360 8528 39424
rect 8592 39360 8608 39424
rect 8672 39360 8688 39424
rect 8752 39360 8768 39424
rect 8832 39360 8848 39424
rect 8912 39360 8928 39424
rect 8992 39360 9000 39424
rect 5000 39344 9000 39360
rect 5000 39280 5008 39344
rect 5072 39280 5088 39344
rect 5152 39280 5168 39344
rect 5232 39280 5248 39344
rect 5312 39280 5328 39344
rect 5392 39280 5408 39344
rect 5472 39280 5488 39344
rect 5552 39280 5568 39344
rect 5632 39280 5648 39344
rect 5712 39280 5728 39344
rect 5792 39280 5808 39344
rect 5872 39280 5888 39344
rect 5952 39280 5968 39344
rect 6032 39280 6048 39344
rect 6112 39280 6128 39344
rect 6192 39280 6208 39344
rect 6272 39280 6288 39344
rect 6352 39280 6368 39344
rect 6432 39280 6448 39344
rect 6512 39280 6528 39344
rect 6592 39280 6608 39344
rect 6672 39280 6688 39344
rect 6752 39280 6768 39344
rect 6832 39280 6848 39344
rect 6912 39280 6928 39344
rect 6992 39280 7008 39344
rect 7072 39280 7088 39344
rect 7152 39280 7168 39344
rect 7232 39280 7248 39344
rect 7312 39280 7328 39344
rect 7392 39280 7408 39344
rect 7472 39280 7488 39344
rect 7552 39280 7568 39344
rect 7632 39280 7648 39344
rect 7712 39280 7728 39344
rect 7792 39280 7808 39344
rect 7872 39280 7888 39344
rect 7952 39280 7968 39344
rect 8032 39280 8048 39344
rect 8112 39280 8128 39344
rect 8192 39280 8208 39344
rect 8272 39280 8288 39344
rect 8352 39280 8368 39344
rect 8432 39280 8448 39344
rect 8512 39280 8528 39344
rect 8592 39280 8608 39344
rect 8672 39280 8688 39344
rect 8752 39280 8768 39344
rect 8832 39280 8848 39344
rect 8912 39280 8928 39344
rect 8992 39280 9000 39344
rect 5000 39264 9000 39280
rect 5000 39200 5008 39264
rect 5072 39200 5088 39264
rect 5152 39200 5168 39264
rect 5232 39200 5248 39264
rect 5312 39200 5328 39264
rect 5392 39200 5408 39264
rect 5472 39200 5488 39264
rect 5552 39200 5568 39264
rect 5632 39200 5648 39264
rect 5712 39200 5728 39264
rect 5792 39200 5808 39264
rect 5872 39200 5888 39264
rect 5952 39200 5968 39264
rect 6032 39200 6048 39264
rect 6112 39200 6128 39264
rect 6192 39200 6208 39264
rect 6272 39200 6288 39264
rect 6352 39200 6368 39264
rect 6432 39200 6448 39264
rect 6512 39200 6528 39264
rect 6592 39200 6608 39264
rect 6672 39200 6688 39264
rect 6752 39200 6768 39264
rect 6832 39200 6848 39264
rect 6912 39200 6928 39264
rect 6992 39200 7008 39264
rect 7072 39200 7088 39264
rect 7152 39200 7168 39264
rect 7232 39200 7248 39264
rect 7312 39200 7328 39264
rect 7392 39200 7408 39264
rect 7472 39200 7488 39264
rect 7552 39200 7568 39264
rect 7632 39200 7648 39264
rect 7712 39200 7728 39264
rect 7792 39200 7808 39264
rect 7872 39200 7888 39264
rect 7952 39200 7968 39264
rect 8032 39200 8048 39264
rect 8112 39200 8128 39264
rect 8192 39200 8208 39264
rect 8272 39200 8288 39264
rect 8352 39200 8368 39264
rect 8432 39200 8448 39264
rect 8512 39200 8528 39264
rect 8592 39200 8608 39264
rect 8672 39200 8688 39264
rect 8752 39200 8768 39264
rect 8832 39200 8848 39264
rect 8912 39200 8928 39264
rect 8992 39200 9000 39264
rect 5000 39184 9000 39200
rect 5000 39120 5008 39184
rect 5072 39120 5088 39184
rect 5152 39120 5168 39184
rect 5232 39120 5248 39184
rect 5312 39120 5328 39184
rect 5392 39120 5408 39184
rect 5472 39120 5488 39184
rect 5552 39120 5568 39184
rect 5632 39120 5648 39184
rect 5712 39120 5728 39184
rect 5792 39120 5808 39184
rect 5872 39120 5888 39184
rect 5952 39120 5968 39184
rect 6032 39120 6048 39184
rect 6112 39120 6128 39184
rect 6192 39120 6208 39184
rect 6272 39120 6288 39184
rect 6352 39120 6368 39184
rect 6432 39120 6448 39184
rect 6512 39120 6528 39184
rect 6592 39120 6608 39184
rect 6672 39120 6688 39184
rect 6752 39120 6768 39184
rect 6832 39120 6848 39184
rect 6912 39120 6928 39184
rect 6992 39120 7008 39184
rect 7072 39120 7088 39184
rect 7152 39120 7168 39184
rect 7232 39120 7248 39184
rect 7312 39120 7328 39184
rect 7392 39120 7408 39184
rect 7472 39120 7488 39184
rect 7552 39120 7568 39184
rect 7632 39120 7648 39184
rect 7712 39120 7728 39184
rect 7792 39120 7808 39184
rect 7872 39120 7888 39184
rect 7952 39120 7968 39184
rect 8032 39120 8048 39184
rect 8112 39120 8128 39184
rect 8192 39120 8208 39184
rect 8272 39120 8288 39184
rect 8352 39120 8368 39184
rect 8432 39120 8448 39184
rect 8512 39120 8528 39184
rect 8592 39120 8608 39184
rect 8672 39120 8688 39184
rect 8752 39120 8768 39184
rect 8832 39120 8848 39184
rect 8912 39120 8928 39184
rect 8992 39120 9000 39184
rect 5000 39104 9000 39120
rect 5000 39040 5008 39104
rect 5072 39040 5088 39104
rect 5152 39040 5168 39104
rect 5232 39040 5248 39104
rect 5312 39040 5328 39104
rect 5392 39040 5408 39104
rect 5472 39040 5488 39104
rect 5552 39040 5568 39104
rect 5632 39040 5648 39104
rect 5712 39040 5728 39104
rect 5792 39040 5808 39104
rect 5872 39040 5888 39104
rect 5952 39040 5968 39104
rect 6032 39040 6048 39104
rect 6112 39040 6128 39104
rect 6192 39040 6208 39104
rect 6272 39040 6288 39104
rect 6352 39040 6368 39104
rect 6432 39040 6448 39104
rect 6512 39040 6528 39104
rect 6592 39040 6608 39104
rect 6672 39040 6688 39104
rect 6752 39040 6768 39104
rect 6832 39040 6848 39104
rect 6912 39040 6928 39104
rect 6992 39040 7008 39104
rect 7072 39040 7088 39104
rect 7152 39040 7168 39104
rect 7232 39040 7248 39104
rect 7312 39040 7328 39104
rect 7392 39040 7408 39104
rect 7472 39040 7488 39104
rect 7552 39040 7568 39104
rect 7632 39040 7648 39104
rect 7712 39040 7728 39104
rect 7792 39040 7808 39104
rect 7872 39040 7888 39104
rect 7952 39040 7968 39104
rect 8032 39040 8048 39104
rect 8112 39040 8128 39104
rect 8192 39040 8208 39104
rect 8272 39040 8288 39104
rect 8352 39040 8368 39104
rect 8432 39040 8448 39104
rect 8512 39040 8528 39104
rect 8592 39040 8608 39104
rect 8672 39040 8688 39104
rect 8752 39040 8768 39104
rect 8832 39040 8848 39104
rect 8912 39040 8928 39104
rect 8992 39040 9000 39104
rect 5000 39024 9000 39040
rect 5000 38960 5008 39024
rect 5072 38960 5088 39024
rect 5152 38960 5168 39024
rect 5232 38960 5248 39024
rect 5312 38960 5328 39024
rect 5392 38960 5408 39024
rect 5472 38960 5488 39024
rect 5552 38960 5568 39024
rect 5632 38960 5648 39024
rect 5712 38960 5728 39024
rect 5792 38960 5808 39024
rect 5872 38960 5888 39024
rect 5952 38960 5968 39024
rect 6032 38960 6048 39024
rect 6112 38960 6128 39024
rect 6192 38960 6208 39024
rect 6272 38960 6288 39024
rect 6352 38960 6368 39024
rect 6432 38960 6448 39024
rect 6512 38960 6528 39024
rect 6592 38960 6608 39024
rect 6672 38960 6688 39024
rect 6752 38960 6768 39024
rect 6832 38960 6848 39024
rect 6912 38960 6928 39024
rect 6992 38960 7008 39024
rect 7072 38960 7088 39024
rect 7152 38960 7168 39024
rect 7232 38960 7248 39024
rect 7312 38960 7328 39024
rect 7392 38960 7408 39024
rect 7472 38960 7488 39024
rect 7552 38960 7568 39024
rect 7632 38960 7648 39024
rect 7712 38960 7728 39024
rect 7792 38960 7808 39024
rect 7872 38960 7888 39024
rect 7952 38960 7968 39024
rect 8032 38960 8048 39024
rect 8112 38960 8128 39024
rect 8192 38960 8208 39024
rect 8272 38960 8288 39024
rect 8352 38960 8368 39024
rect 8432 38960 8448 39024
rect 8512 38960 8528 39024
rect 8592 38960 8608 39024
rect 8672 38960 8688 39024
rect 8752 38960 8768 39024
rect 8832 38960 8848 39024
rect 8912 38960 8928 39024
rect 8992 38960 9000 39024
rect 5000 38944 9000 38960
rect 5000 38880 5008 38944
rect 5072 38880 5088 38944
rect 5152 38880 5168 38944
rect 5232 38880 5248 38944
rect 5312 38880 5328 38944
rect 5392 38880 5408 38944
rect 5472 38880 5488 38944
rect 5552 38880 5568 38944
rect 5632 38880 5648 38944
rect 5712 38880 5728 38944
rect 5792 38880 5808 38944
rect 5872 38880 5888 38944
rect 5952 38880 5968 38944
rect 6032 38880 6048 38944
rect 6112 38880 6128 38944
rect 6192 38880 6208 38944
rect 6272 38880 6288 38944
rect 6352 38880 6368 38944
rect 6432 38880 6448 38944
rect 6512 38880 6528 38944
rect 6592 38880 6608 38944
rect 6672 38880 6688 38944
rect 6752 38880 6768 38944
rect 6832 38880 6848 38944
rect 6912 38880 6928 38944
rect 6992 38880 7008 38944
rect 7072 38880 7088 38944
rect 7152 38880 7168 38944
rect 7232 38880 7248 38944
rect 7312 38880 7328 38944
rect 7392 38880 7408 38944
rect 7472 38880 7488 38944
rect 7552 38880 7568 38944
rect 7632 38880 7648 38944
rect 7712 38880 7728 38944
rect 7792 38880 7808 38944
rect 7872 38880 7888 38944
rect 7952 38880 7968 38944
rect 8032 38880 8048 38944
rect 8112 38880 8128 38944
rect 8192 38880 8208 38944
rect 8272 38880 8288 38944
rect 8352 38880 8368 38944
rect 8432 38880 8448 38944
rect 8512 38880 8528 38944
rect 8592 38880 8608 38944
rect 8672 38880 8688 38944
rect 8752 38880 8768 38944
rect 8832 38880 8848 38944
rect 8912 38880 8928 38944
rect 8992 38880 9000 38944
rect 5000 38864 9000 38880
rect 5000 38800 5008 38864
rect 5072 38800 5088 38864
rect 5152 38800 5168 38864
rect 5232 38800 5248 38864
rect 5312 38800 5328 38864
rect 5392 38800 5408 38864
rect 5472 38800 5488 38864
rect 5552 38800 5568 38864
rect 5632 38800 5648 38864
rect 5712 38800 5728 38864
rect 5792 38800 5808 38864
rect 5872 38800 5888 38864
rect 5952 38800 5968 38864
rect 6032 38800 6048 38864
rect 6112 38800 6128 38864
rect 6192 38800 6208 38864
rect 6272 38800 6288 38864
rect 6352 38800 6368 38864
rect 6432 38800 6448 38864
rect 6512 38800 6528 38864
rect 6592 38800 6608 38864
rect 6672 38800 6688 38864
rect 6752 38800 6768 38864
rect 6832 38800 6848 38864
rect 6912 38800 6928 38864
rect 6992 38800 7008 38864
rect 7072 38800 7088 38864
rect 7152 38800 7168 38864
rect 7232 38800 7248 38864
rect 7312 38800 7328 38864
rect 7392 38800 7408 38864
rect 7472 38800 7488 38864
rect 7552 38800 7568 38864
rect 7632 38800 7648 38864
rect 7712 38800 7728 38864
rect 7792 38800 7808 38864
rect 7872 38800 7888 38864
rect 7952 38800 7968 38864
rect 8032 38800 8048 38864
rect 8112 38800 8128 38864
rect 8192 38800 8208 38864
rect 8272 38800 8288 38864
rect 8352 38800 8368 38864
rect 8432 38800 8448 38864
rect 8512 38800 8528 38864
rect 8592 38800 8608 38864
rect 8672 38800 8688 38864
rect 8752 38800 8768 38864
rect 8832 38800 8848 38864
rect 8912 38800 8928 38864
rect 8992 38800 9000 38864
rect 5000 38784 9000 38800
rect 5000 38720 5008 38784
rect 5072 38720 5088 38784
rect 5152 38720 5168 38784
rect 5232 38720 5248 38784
rect 5312 38720 5328 38784
rect 5392 38720 5408 38784
rect 5472 38720 5488 38784
rect 5552 38720 5568 38784
rect 5632 38720 5648 38784
rect 5712 38720 5728 38784
rect 5792 38720 5808 38784
rect 5872 38720 5888 38784
rect 5952 38720 5968 38784
rect 6032 38720 6048 38784
rect 6112 38720 6128 38784
rect 6192 38720 6208 38784
rect 6272 38720 6288 38784
rect 6352 38720 6368 38784
rect 6432 38720 6448 38784
rect 6512 38720 6528 38784
rect 6592 38720 6608 38784
rect 6672 38720 6688 38784
rect 6752 38720 6768 38784
rect 6832 38720 6848 38784
rect 6912 38720 6928 38784
rect 6992 38720 7008 38784
rect 7072 38720 7088 38784
rect 7152 38720 7168 38784
rect 7232 38720 7248 38784
rect 7312 38720 7328 38784
rect 7392 38720 7408 38784
rect 7472 38720 7488 38784
rect 7552 38720 7568 38784
rect 7632 38720 7648 38784
rect 7712 38720 7728 38784
rect 7792 38720 7808 38784
rect 7872 38720 7888 38784
rect 7952 38720 7968 38784
rect 8032 38720 8048 38784
rect 8112 38720 8128 38784
rect 8192 38720 8208 38784
rect 8272 38720 8288 38784
rect 8352 38720 8368 38784
rect 8432 38720 8448 38784
rect 8512 38720 8528 38784
rect 8592 38720 8608 38784
rect 8672 38720 8688 38784
rect 8752 38720 8768 38784
rect 8832 38720 8848 38784
rect 8912 38720 8928 38784
rect 8992 38720 9000 38784
rect 5000 38704 9000 38720
rect 5000 38640 5008 38704
rect 5072 38640 5088 38704
rect 5152 38640 5168 38704
rect 5232 38640 5248 38704
rect 5312 38640 5328 38704
rect 5392 38640 5408 38704
rect 5472 38640 5488 38704
rect 5552 38640 5568 38704
rect 5632 38640 5648 38704
rect 5712 38640 5728 38704
rect 5792 38640 5808 38704
rect 5872 38640 5888 38704
rect 5952 38640 5968 38704
rect 6032 38640 6048 38704
rect 6112 38640 6128 38704
rect 6192 38640 6208 38704
rect 6272 38640 6288 38704
rect 6352 38640 6368 38704
rect 6432 38640 6448 38704
rect 6512 38640 6528 38704
rect 6592 38640 6608 38704
rect 6672 38640 6688 38704
rect 6752 38640 6768 38704
rect 6832 38640 6848 38704
rect 6912 38640 6928 38704
rect 6992 38640 7008 38704
rect 7072 38640 7088 38704
rect 7152 38640 7168 38704
rect 7232 38640 7248 38704
rect 7312 38640 7328 38704
rect 7392 38640 7408 38704
rect 7472 38640 7488 38704
rect 7552 38640 7568 38704
rect 7632 38640 7648 38704
rect 7712 38640 7728 38704
rect 7792 38640 7808 38704
rect 7872 38640 7888 38704
rect 7952 38640 7968 38704
rect 8032 38640 8048 38704
rect 8112 38640 8128 38704
rect 8192 38640 8208 38704
rect 8272 38640 8288 38704
rect 8352 38640 8368 38704
rect 8432 38640 8448 38704
rect 8512 38640 8528 38704
rect 8592 38640 8608 38704
rect 8672 38640 8688 38704
rect 8752 38640 8768 38704
rect 8832 38640 8848 38704
rect 8912 38640 8928 38704
rect 8992 38640 9000 38704
rect 5000 38624 9000 38640
rect 5000 38560 5008 38624
rect 5072 38560 5088 38624
rect 5152 38560 5168 38624
rect 5232 38560 5248 38624
rect 5312 38560 5328 38624
rect 5392 38560 5408 38624
rect 5472 38560 5488 38624
rect 5552 38560 5568 38624
rect 5632 38560 5648 38624
rect 5712 38560 5728 38624
rect 5792 38560 5808 38624
rect 5872 38560 5888 38624
rect 5952 38560 5968 38624
rect 6032 38560 6048 38624
rect 6112 38560 6128 38624
rect 6192 38560 6208 38624
rect 6272 38560 6288 38624
rect 6352 38560 6368 38624
rect 6432 38560 6448 38624
rect 6512 38560 6528 38624
rect 6592 38560 6608 38624
rect 6672 38560 6688 38624
rect 6752 38560 6768 38624
rect 6832 38560 6848 38624
rect 6912 38560 6928 38624
rect 6992 38560 7008 38624
rect 7072 38560 7088 38624
rect 7152 38560 7168 38624
rect 7232 38560 7248 38624
rect 7312 38560 7328 38624
rect 7392 38560 7408 38624
rect 7472 38560 7488 38624
rect 7552 38560 7568 38624
rect 7632 38560 7648 38624
rect 7712 38560 7728 38624
rect 7792 38560 7808 38624
rect 7872 38560 7888 38624
rect 7952 38560 7968 38624
rect 8032 38560 8048 38624
rect 8112 38560 8128 38624
rect 8192 38560 8208 38624
rect 8272 38560 8288 38624
rect 8352 38560 8368 38624
rect 8432 38560 8448 38624
rect 8512 38560 8528 38624
rect 8592 38560 8608 38624
rect 8672 38560 8688 38624
rect 8752 38560 8768 38624
rect 8832 38560 8848 38624
rect 8912 38560 8928 38624
rect 8992 38560 9000 38624
rect 5000 38544 9000 38560
rect 5000 38480 5008 38544
rect 5072 38480 5088 38544
rect 5152 38480 5168 38544
rect 5232 38480 5248 38544
rect 5312 38480 5328 38544
rect 5392 38480 5408 38544
rect 5472 38480 5488 38544
rect 5552 38480 5568 38544
rect 5632 38480 5648 38544
rect 5712 38480 5728 38544
rect 5792 38480 5808 38544
rect 5872 38480 5888 38544
rect 5952 38480 5968 38544
rect 6032 38480 6048 38544
rect 6112 38480 6128 38544
rect 6192 38480 6208 38544
rect 6272 38480 6288 38544
rect 6352 38480 6368 38544
rect 6432 38480 6448 38544
rect 6512 38480 6528 38544
rect 6592 38480 6608 38544
rect 6672 38480 6688 38544
rect 6752 38480 6768 38544
rect 6832 38480 6848 38544
rect 6912 38480 6928 38544
rect 6992 38480 7008 38544
rect 7072 38480 7088 38544
rect 7152 38480 7168 38544
rect 7232 38480 7248 38544
rect 7312 38480 7328 38544
rect 7392 38480 7408 38544
rect 7472 38480 7488 38544
rect 7552 38480 7568 38544
rect 7632 38480 7648 38544
rect 7712 38480 7728 38544
rect 7792 38480 7808 38544
rect 7872 38480 7888 38544
rect 7952 38480 7968 38544
rect 8032 38480 8048 38544
rect 8112 38480 8128 38544
rect 8192 38480 8208 38544
rect 8272 38480 8288 38544
rect 8352 38480 8368 38544
rect 8432 38480 8448 38544
rect 8512 38480 8528 38544
rect 8592 38480 8608 38544
rect 8672 38480 8688 38544
rect 8752 38480 8768 38544
rect 8832 38480 8848 38544
rect 8912 38480 8928 38544
rect 8992 38480 9000 38544
rect 5000 38464 9000 38480
rect 5000 38400 5008 38464
rect 5072 38400 5088 38464
rect 5152 38400 5168 38464
rect 5232 38400 5248 38464
rect 5312 38400 5328 38464
rect 5392 38400 5408 38464
rect 5472 38400 5488 38464
rect 5552 38400 5568 38464
rect 5632 38400 5648 38464
rect 5712 38400 5728 38464
rect 5792 38400 5808 38464
rect 5872 38400 5888 38464
rect 5952 38400 5968 38464
rect 6032 38400 6048 38464
rect 6112 38400 6128 38464
rect 6192 38400 6208 38464
rect 6272 38400 6288 38464
rect 6352 38400 6368 38464
rect 6432 38400 6448 38464
rect 6512 38400 6528 38464
rect 6592 38400 6608 38464
rect 6672 38400 6688 38464
rect 6752 38400 6768 38464
rect 6832 38400 6848 38464
rect 6912 38400 6928 38464
rect 6992 38400 7008 38464
rect 7072 38400 7088 38464
rect 7152 38400 7168 38464
rect 7232 38400 7248 38464
rect 7312 38400 7328 38464
rect 7392 38400 7408 38464
rect 7472 38400 7488 38464
rect 7552 38400 7568 38464
rect 7632 38400 7648 38464
rect 7712 38400 7728 38464
rect 7792 38400 7808 38464
rect 7872 38400 7888 38464
rect 7952 38400 7968 38464
rect 8032 38400 8048 38464
rect 8112 38400 8128 38464
rect 8192 38400 8208 38464
rect 8272 38400 8288 38464
rect 8352 38400 8368 38464
rect 8432 38400 8448 38464
rect 8512 38400 8528 38464
rect 8592 38400 8608 38464
rect 8672 38400 8688 38464
rect 8752 38400 8768 38464
rect 8832 38400 8848 38464
rect 8912 38400 8928 38464
rect 8992 38400 9000 38464
rect 5000 38384 9000 38400
rect 5000 38320 5008 38384
rect 5072 38320 5088 38384
rect 5152 38320 5168 38384
rect 5232 38320 5248 38384
rect 5312 38320 5328 38384
rect 5392 38320 5408 38384
rect 5472 38320 5488 38384
rect 5552 38320 5568 38384
rect 5632 38320 5648 38384
rect 5712 38320 5728 38384
rect 5792 38320 5808 38384
rect 5872 38320 5888 38384
rect 5952 38320 5968 38384
rect 6032 38320 6048 38384
rect 6112 38320 6128 38384
rect 6192 38320 6208 38384
rect 6272 38320 6288 38384
rect 6352 38320 6368 38384
rect 6432 38320 6448 38384
rect 6512 38320 6528 38384
rect 6592 38320 6608 38384
rect 6672 38320 6688 38384
rect 6752 38320 6768 38384
rect 6832 38320 6848 38384
rect 6912 38320 6928 38384
rect 6992 38320 7008 38384
rect 7072 38320 7088 38384
rect 7152 38320 7168 38384
rect 7232 38320 7248 38384
rect 7312 38320 7328 38384
rect 7392 38320 7408 38384
rect 7472 38320 7488 38384
rect 7552 38320 7568 38384
rect 7632 38320 7648 38384
rect 7712 38320 7728 38384
rect 7792 38320 7808 38384
rect 7872 38320 7888 38384
rect 7952 38320 7968 38384
rect 8032 38320 8048 38384
rect 8112 38320 8128 38384
rect 8192 38320 8208 38384
rect 8272 38320 8288 38384
rect 8352 38320 8368 38384
rect 8432 38320 8448 38384
rect 8512 38320 8528 38384
rect 8592 38320 8608 38384
rect 8672 38320 8688 38384
rect 8752 38320 8768 38384
rect 8832 38320 8848 38384
rect 8912 38320 8928 38384
rect 8992 38320 9000 38384
rect 5000 38304 9000 38320
rect 5000 38240 5008 38304
rect 5072 38240 5088 38304
rect 5152 38240 5168 38304
rect 5232 38240 5248 38304
rect 5312 38240 5328 38304
rect 5392 38240 5408 38304
rect 5472 38240 5488 38304
rect 5552 38240 5568 38304
rect 5632 38240 5648 38304
rect 5712 38240 5728 38304
rect 5792 38240 5808 38304
rect 5872 38240 5888 38304
rect 5952 38240 5968 38304
rect 6032 38240 6048 38304
rect 6112 38240 6128 38304
rect 6192 38240 6208 38304
rect 6272 38240 6288 38304
rect 6352 38240 6368 38304
rect 6432 38240 6448 38304
rect 6512 38240 6528 38304
rect 6592 38240 6608 38304
rect 6672 38240 6688 38304
rect 6752 38240 6768 38304
rect 6832 38240 6848 38304
rect 6912 38240 6928 38304
rect 6992 38240 7008 38304
rect 7072 38240 7088 38304
rect 7152 38240 7168 38304
rect 7232 38240 7248 38304
rect 7312 38240 7328 38304
rect 7392 38240 7408 38304
rect 7472 38240 7488 38304
rect 7552 38240 7568 38304
rect 7632 38240 7648 38304
rect 7712 38240 7728 38304
rect 7792 38240 7808 38304
rect 7872 38240 7888 38304
rect 7952 38240 7968 38304
rect 8032 38240 8048 38304
rect 8112 38240 8128 38304
rect 8192 38240 8208 38304
rect 8272 38240 8288 38304
rect 8352 38240 8368 38304
rect 8432 38240 8448 38304
rect 8512 38240 8528 38304
rect 8592 38240 8608 38304
rect 8672 38240 8688 38304
rect 8752 38240 8768 38304
rect 8832 38240 8848 38304
rect 8912 38240 8928 38304
rect 8992 38240 9000 38304
rect 5000 38224 9000 38240
rect 5000 38160 5008 38224
rect 5072 38160 5088 38224
rect 5152 38160 5168 38224
rect 5232 38160 5248 38224
rect 5312 38160 5328 38224
rect 5392 38160 5408 38224
rect 5472 38160 5488 38224
rect 5552 38160 5568 38224
rect 5632 38160 5648 38224
rect 5712 38160 5728 38224
rect 5792 38160 5808 38224
rect 5872 38160 5888 38224
rect 5952 38160 5968 38224
rect 6032 38160 6048 38224
rect 6112 38160 6128 38224
rect 6192 38160 6208 38224
rect 6272 38160 6288 38224
rect 6352 38160 6368 38224
rect 6432 38160 6448 38224
rect 6512 38160 6528 38224
rect 6592 38160 6608 38224
rect 6672 38160 6688 38224
rect 6752 38160 6768 38224
rect 6832 38160 6848 38224
rect 6912 38160 6928 38224
rect 6992 38160 7008 38224
rect 7072 38160 7088 38224
rect 7152 38160 7168 38224
rect 7232 38160 7248 38224
rect 7312 38160 7328 38224
rect 7392 38160 7408 38224
rect 7472 38160 7488 38224
rect 7552 38160 7568 38224
rect 7632 38160 7648 38224
rect 7712 38160 7728 38224
rect 7792 38160 7808 38224
rect 7872 38160 7888 38224
rect 7952 38160 7968 38224
rect 8032 38160 8048 38224
rect 8112 38160 8128 38224
rect 8192 38160 8208 38224
rect 8272 38160 8288 38224
rect 8352 38160 8368 38224
rect 8432 38160 8448 38224
rect 8512 38160 8528 38224
rect 8592 38160 8608 38224
rect 8672 38160 8688 38224
rect 8752 38160 8768 38224
rect 8832 38160 8848 38224
rect 8912 38160 8928 38224
rect 8992 38160 9000 38224
rect 5000 38144 9000 38160
rect 5000 38080 5008 38144
rect 5072 38080 5088 38144
rect 5152 38080 5168 38144
rect 5232 38080 5248 38144
rect 5312 38080 5328 38144
rect 5392 38080 5408 38144
rect 5472 38080 5488 38144
rect 5552 38080 5568 38144
rect 5632 38080 5648 38144
rect 5712 38080 5728 38144
rect 5792 38080 5808 38144
rect 5872 38080 5888 38144
rect 5952 38080 5968 38144
rect 6032 38080 6048 38144
rect 6112 38080 6128 38144
rect 6192 38080 6208 38144
rect 6272 38080 6288 38144
rect 6352 38080 6368 38144
rect 6432 38080 6448 38144
rect 6512 38080 6528 38144
rect 6592 38080 6608 38144
rect 6672 38080 6688 38144
rect 6752 38080 6768 38144
rect 6832 38080 6848 38144
rect 6912 38080 6928 38144
rect 6992 38080 7008 38144
rect 7072 38080 7088 38144
rect 7152 38080 7168 38144
rect 7232 38080 7248 38144
rect 7312 38080 7328 38144
rect 7392 38080 7408 38144
rect 7472 38080 7488 38144
rect 7552 38080 7568 38144
rect 7632 38080 7648 38144
rect 7712 38080 7728 38144
rect 7792 38080 7808 38144
rect 7872 38080 7888 38144
rect 7952 38080 7968 38144
rect 8032 38080 8048 38144
rect 8112 38080 8128 38144
rect 8192 38080 8208 38144
rect 8272 38080 8288 38144
rect 8352 38080 8368 38144
rect 8432 38080 8448 38144
rect 8512 38080 8528 38144
rect 8592 38080 8608 38144
rect 8672 38080 8688 38144
rect 8752 38080 8768 38144
rect 8832 38080 8848 38144
rect 8912 38080 8928 38144
rect 8992 38080 9000 38144
rect 5000 38064 9000 38080
rect 5000 38000 5008 38064
rect 5072 38000 5088 38064
rect 5152 38000 5168 38064
rect 5232 38000 5248 38064
rect 5312 38000 5328 38064
rect 5392 38000 5408 38064
rect 5472 38000 5488 38064
rect 5552 38000 5568 38064
rect 5632 38000 5648 38064
rect 5712 38000 5728 38064
rect 5792 38000 5808 38064
rect 5872 38000 5888 38064
rect 5952 38000 5968 38064
rect 6032 38000 6048 38064
rect 6112 38000 6128 38064
rect 6192 38000 6208 38064
rect 6272 38000 6288 38064
rect 6352 38000 6368 38064
rect 6432 38000 6448 38064
rect 6512 38000 6528 38064
rect 6592 38000 6608 38064
rect 6672 38000 6688 38064
rect 6752 38000 6768 38064
rect 6832 38000 6848 38064
rect 6912 38000 6928 38064
rect 6992 38000 7008 38064
rect 7072 38000 7088 38064
rect 7152 38000 7168 38064
rect 7232 38000 7248 38064
rect 7312 38000 7328 38064
rect 7392 38000 7408 38064
rect 7472 38000 7488 38064
rect 7552 38000 7568 38064
rect 7632 38000 7648 38064
rect 7712 38000 7728 38064
rect 7792 38000 7808 38064
rect 7872 38000 7888 38064
rect 7952 38000 7968 38064
rect 8032 38000 8048 38064
rect 8112 38000 8128 38064
rect 8192 38000 8208 38064
rect 8272 38000 8288 38064
rect 8352 38000 8368 38064
rect 8432 38000 8448 38064
rect 8512 38000 8528 38064
rect 8592 38000 8608 38064
rect 8672 38000 8688 38064
rect 8752 38000 8768 38064
rect 8832 38000 8848 38064
rect 8912 38000 8928 38064
rect 8992 38000 9000 38064
rect 5000 37984 9000 38000
rect 5000 37920 5008 37984
rect 5072 37920 5088 37984
rect 5152 37920 5168 37984
rect 5232 37920 5248 37984
rect 5312 37920 5328 37984
rect 5392 37920 5408 37984
rect 5472 37920 5488 37984
rect 5552 37920 5568 37984
rect 5632 37920 5648 37984
rect 5712 37920 5728 37984
rect 5792 37920 5808 37984
rect 5872 37920 5888 37984
rect 5952 37920 5968 37984
rect 6032 37920 6048 37984
rect 6112 37920 6128 37984
rect 6192 37920 6208 37984
rect 6272 37920 6288 37984
rect 6352 37920 6368 37984
rect 6432 37920 6448 37984
rect 6512 37920 6528 37984
rect 6592 37920 6608 37984
rect 6672 37920 6688 37984
rect 6752 37920 6768 37984
rect 6832 37920 6848 37984
rect 6912 37920 6928 37984
rect 6992 37920 7008 37984
rect 7072 37920 7088 37984
rect 7152 37920 7168 37984
rect 7232 37920 7248 37984
rect 7312 37920 7328 37984
rect 7392 37920 7408 37984
rect 7472 37920 7488 37984
rect 7552 37920 7568 37984
rect 7632 37920 7648 37984
rect 7712 37920 7728 37984
rect 7792 37920 7808 37984
rect 7872 37920 7888 37984
rect 7952 37920 7968 37984
rect 8032 37920 8048 37984
rect 8112 37920 8128 37984
rect 8192 37920 8208 37984
rect 8272 37920 8288 37984
rect 8352 37920 8368 37984
rect 8432 37920 8448 37984
rect 8512 37920 8528 37984
rect 8592 37920 8608 37984
rect 8672 37920 8688 37984
rect 8752 37920 8768 37984
rect 8832 37920 8848 37984
rect 8912 37920 8928 37984
rect 8992 37920 9000 37984
rect 5000 37904 9000 37920
rect 5000 37840 5008 37904
rect 5072 37840 5088 37904
rect 5152 37840 5168 37904
rect 5232 37840 5248 37904
rect 5312 37840 5328 37904
rect 5392 37840 5408 37904
rect 5472 37840 5488 37904
rect 5552 37840 5568 37904
rect 5632 37840 5648 37904
rect 5712 37840 5728 37904
rect 5792 37840 5808 37904
rect 5872 37840 5888 37904
rect 5952 37840 5968 37904
rect 6032 37840 6048 37904
rect 6112 37840 6128 37904
rect 6192 37840 6208 37904
rect 6272 37840 6288 37904
rect 6352 37840 6368 37904
rect 6432 37840 6448 37904
rect 6512 37840 6528 37904
rect 6592 37840 6608 37904
rect 6672 37840 6688 37904
rect 6752 37840 6768 37904
rect 6832 37840 6848 37904
rect 6912 37840 6928 37904
rect 6992 37840 7008 37904
rect 7072 37840 7088 37904
rect 7152 37840 7168 37904
rect 7232 37840 7248 37904
rect 7312 37840 7328 37904
rect 7392 37840 7408 37904
rect 7472 37840 7488 37904
rect 7552 37840 7568 37904
rect 7632 37840 7648 37904
rect 7712 37840 7728 37904
rect 7792 37840 7808 37904
rect 7872 37840 7888 37904
rect 7952 37840 7968 37904
rect 8032 37840 8048 37904
rect 8112 37840 8128 37904
rect 8192 37840 8208 37904
rect 8272 37840 8288 37904
rect 8352 37840 8368 37904
rect 8432 37840 8448 37904
rect 8512 37840 8528 37904
rect 8592 37840 8608 37904
rect 8672 37840 8688 37904
rect 8752 37840 8768 37904
rect 8832 37840 8848 37904
rect 8912 37840 8928 37904
rect 8992 37840 9000 37904
rect 5000 37824 9000 37840
rect 5000 37760 5008 37824
rect 5072 37760 5088 37824
rect 5152 37760 5168 37824
rect 5232 37760 5248 37824
rect 5312 37760 5328 37824
rect 5392 37760 5408 37824
rect 5472 37760 5488 37824
rect 5552 37760 5568 37824
rect 5632 37760 5648 37824
rect 5712 37760 5728 37824
rect 5792 37760 5808 37824
rect 5872 37760 5888 37824
rect 5952 37760 5968 37824
rect 6032 37760 6048 37824
rect 6112 37760 6128 37824
rect 6192 37760 6208 37824
rect 6272 37760 6288 37824
rect 6352 37760 6368 37824
rect 6432 37760 6448 37824
rect 6512 37760 6528 37824
rect 6592 37760 6608 37824
rect 6672 37760 6688 37824
rect 6752 37760 6768 37824
rect 6832 37760 6848 37824
rect 6912 37760 6928 37824
rect 6992 37760 7008 37824
rect 7072 37760 7088 37824
rect 7152 37760 7168 37824
rect 7232 37760 7248 37824
rect 7312 37760 7328 37824
rect 7392 37760 7408 37824
rect 7472 37760 7488 37824
rect 7552 37760 7568 37824
rect 7632 37760 7648 37824
rect 7712 37760 7728 37824
rect 7792 37760 7808 37824
rect 7872 37760 7888 37824
rect 7952 37760 7968 37824
rect 8032 37760 8048 37824
rect 8112 37760 8128 37824
rect 8192 37760 8208 37824
rect 8272 37760 8288 37824
rect 8352 37760 8368 37824
rect 8432 37760 8448 37824
rect 8512 37760 8528 37824
rect 8592 37760 8608 37824
rect 8672 37760 8688 37824
rect 8752 37760 8768 37824
rect 8832 37760 8848 37824
rect 8912 37760 8928 37824
rect 8992 37760 9000 37824
rect 5000 37744 9000 37760
rect 5000 37680 5008 37744
rect 5072 37680 5088 37744
rect 5152 37680 5168 37744
rect 5232 37680 5248 37744
rect 5312 37680 5328 37744
rect 5392 37680 5408 37744
rect 5472 37680 5488 37744
rect 5552 37680 5568 37744
rect 5632 37680 5648 37744
rect 5712 37680 5728 37744
rect 5792 37680 5808 37744
rect 5872 37680 5888 37744
rect 5952 37680 5968 37744
rect 6032 37680 6048 37744
rect 6112 37680 6128 37744
rect 6192 37680 6208 37744
rect 6272 37680 6288 37744
rect 6352 37680 6368 37744
rect 6432 37680 6448 37744
rect 6512 37680 6528 37744
rect 6592 37680 6608 37744
rect 6672 37680 6688 37744
rect 6752 37680 6768 37744
rect 6832 37680 6848 37744
rect 6912 37680 6928 37744
rect 6992 37680 7008 37744
rect 7072 37680 7088 37744
rect 7152 37680 7168 37744
rect 7232 37680 7248 37744
rect 7312 37680 7328 37744
rect 7392 37680 7408 37744
rect 7472 37680 7488 37744
rect 7552 37680 7568 37744
rect 7632 37680 7648 37744
rect 7712 37680 7728 37744
rect 7792 37680 7808 37744
rect 7872 37680 7888 37744
rect 7952 37680 7968 37744
rect 8032 37680 8048 37744
rect 8112 37680 8128 37744
rect 8192 37680 8208 37744
rect 8272 37680 8288 37744
rect 8352 37680 8368 37744
rect 8432 37680 8448 37744
rect 8512 37680 8528 37744
rect 8592 37680 8608 37744
rect 8672 37680 8688 37744
rect 8752 37680 8768 37744
rect 8832 37680 8848 37744
rect 8912 37680 8928 37744
rect 8992 37680 9000 37744
rect 5000 37664 9000 37680
rect 5000 37600 5008 37664
rect 5072 37600 5088 37664
rect 5152 37600 5168 37664
rect 5232 37600 5248 37664
rect 5312 37600 5328 37664
rect 5392 37600 5408 37664
rect 5472 37600 5488 37664
rect 5552 37600 5568 37664
rect 5632 37600 5648 37664
rect 5712 37600 5728 37664
rect 5792 37600 5808 37664
rect 5872 37600 5888 37664
rect 5952 37600 5968 37664
rect 6032 37600 6048 37664
rect 6112 37600 6128 37664
rect 6192 37600 6208 37664
rect 6272 37600 6288 37664
rect 6352 37600 6368 37664
rect 6432 37600 6448 37664
rect 6512 37600 6528 37664
rect 6592 37600 6608 37664
rect 6672 37600 6688 37664
rect 6752 37600 6768 37664
rect 6832 37600 6848 37664
rect 6912 37600 6928 37664
rect 6992 37600 7008 37664
rect 7072 37600 7088 37664
rect 7152 37600 7168 37664
rect 7232 37600 7248 37664
rect 7312 37600 7328 37664
rect 7392 37600 7408 37664
rect 7472 37600 7488 37664
rect 7552 37600 7568 37664
rect 7632 37600 7648 37664
rect 7712 37600 7728 37664
rect 7792 37600 7808 37664
rect 7872 37600 7888 37664
rect 7952 37600 7968 37664
rect 8032 37600 8048 37664
rect 8112 37600 8128 37664
rect 8192 37600 8208 37664
rect 8272 37600 8288 37664
rect 8352 37600 8368 37664
rect 8432 37600 8448 37664
rect 8512 37600 8528 37664
rect 8592 37600 8608 37664
rect 8672 37600 8688 37664
rect 8752 37600 8768 37664
rect 8832 37600 8848 37664
rect 8912 37600 8928 37664
rect 8992 37600 9000 37664
rect 5000 37584 9000 37600
rect 5000 37520 5008 37584
rect 5072 37520 5088 37584
rect 5152 37520 5168 37584
rect 5232 37520 5248 37584
rect 5312 37520 5328 37584
rect 5392 37520 5408 37584
rect 5472 37520 5488 37584
rect 5552 37520 5568 37584
rect 5632 37520 5648 37584
rect 5712 37520 5728 37584
rect 5792 37520 5808 37584
rect 5872 37520 5888 37584
rect 5952 37520 5968 37584
rect 6032 37520 6048 37584
rect 6112 37520 6128 37584
rect 6192 37520 6208 37584
rect 6272 37520 6288 37584
rect 6352 37520 6368 37584
rect 6432 37520 6448 37584
rect 6512 37520 6528 37584
rect 6592 37520 6608 37584
rect 6672 37520 6688 37584
rect 6752 37520 6768 37584
rect 6832 37520 6848 37584
rect 6912 37520 6928 37584
rect 6992 37520 7008 37584
rect 7072 37520 7088 37584
rect 7152 37520 7168 37584
rect 7232 37520 7248 37584
rect 7312 37520 7328 37584
rect 7392 37520 7408 37584
rect 7472 37520 7488 37584
rect 7552 37520 7568 37584
rect 7632 37520 7648 37584
rect 7712 37520 7728 37584
rect 7792 37520 7808 37584
rect 7872 37520 7888 37584
rect 7952 37520 7968 37584
rect 8032 37520 8048 37584
rect 8112 37520 8128 37584
rect 8192 37520 8208 37584
rect 8272 37520 8288 37584
rect 8352 37520 8368 37584
rect 8432 37520 8448 37584
rect 8512 37520 8528 37584
rect 8592 37520 8608 37584
rect 8672 37520 8688 37584
rect 8752 37520 8768 37584
rect 8832 37520 8848 37584
rect 8912 37520 8928 37584
rect 8992 37520 9000 37584
rect 5000 37504 9000 37520
rect 5000 37440 5008 37504
rect 5072 37440 5088 37504
rect 5152 37440 5168 37504
rect 5232 37440 5248 37504
rect 5312 37440 5328 37504
rect 5392 37440 5408 37504
rect 5472 37440 5488 37504
rect 5552 37440 5568 37504
rect 5632 37440 5648 37504
rect 5712 37440 5728 37504
rect 5792 37440 5808 37504
rect 5872 37440 5888 37504
rect 5952 37440 5968 37504
rect 6032 37440 6048 37504
rect 6112 37440 6128 37504
rect 6192 37440 6208 37504
rect 6272 37440 6288 37504
rect 6352 37440 6368 37504
rect 6432 37440 6448 37504
rect 6512 37440 6528 37504
rect 6592 37440 6608 37504
rect 6672 37440 6688 37504
rect 6752 37440 6768 37504
rect 6832 37440 6848 37504
rect 6912 37440 6928 37504
rect 6992 37440 7008 37504
rect 7072 37440 7088 37504
rect 7152 37440 7168 37504
rect 7232 37440 7248 37504
rect 7312 37440 7328 37504
rect 7392 37440 7408 37504
rect 7472 37440 7488 37504
rect 7552 37440 7568 37504
rect 7632 37440 7648 37504
rect 7712 37440 7728 37504
rect 7792 37440 7808 37504
rect 7872 37440 7888 37504
rect 7952 37440 7968 37504
rect 8032 37440 8048 37504
rect 8112 37440 8128 37504
rect 8192 37440 8208 37504
rect 8272 37440 8288 37504
rect 8352 37440 8368 37504
rect 8432 37440 8448 37504
rect 8512 37440 8528 37504
rect 8592 37440 8608 37504
rect 8672 37440 8688 37504
rect 8752 37440 8768 37504
rect 8832 37440 8848 37504
rect 8912 37440 8928 37504
rect 8992 37440 9000 37504
rect 5000 37424 9000 37440
rect 5000 37360 5008 37424
rect 5072 37360 5088 37424
rect 5152 37360 5168 37424
rect 5232 37360 5248 37424
rect 5312 37360 5328 37424
rect 5392 37360 5408 37424
rect 5472 37360 5488 37424
rect 5552 37360 5568 37424
rect 5632 37360 5648 37424
rect 5712 37360 5728 37424
rect 5792 37360 5808 37424
rect 5872 37360 5888 37424
rect 5952 37360 5968 37424
rect 6032 37360 6048 37424
rect 6112 37360 6128 37424
rect 6192 37360 6208 37424
rect 6272 37360 6288 37424
rect 6352 37360 6368 37424
rect 6432 37360 6448 37424
rect 6512 37360 6528 37424
rect 6592 37360 6608 37424
rect 6672 37360 6688 37424
rect 6752 37360 6768 37424
rect 6832 37360 6848 37424
rect 6912 37360 6928 37424
rect 6992 37360 7008 37424
rect 7072 37360 7088 37424
rect 7152 37360 7168 37424
rect 7232 37360 7248 37424
rect 7312 37360 7328 37424
rect 7392 37360 7408 37424
rect 7472 37360 7488 37424
rect 7552 37360 7568 37424
rect 7632 37360 7648 37424
rect 7712 37360 7728 37424
rect 7792 37360 7808 37424
rect 7872 37360 7888 37424
rect 7952 37360 7968 37424
rect 8032 37360 8048 37424
rect 8112 37360 8128 37424
rect 8192 37360 8208 37424
rect 8272 37360 8288 37424
rect 8352 37360 8368 37424
rect 8432 37360 8448 37424
rect 8512 37360 8528 37424
rect 8592 37360 8608 37424
rect 8672 37360 8688 37424
rect 8752 37360 8768 37424
rect 8832 37360 8848 37424
rect 8912 37360 8928 37424
rect 8992 37360 9000 37424
rect 5000 37344 9000 37360
rect 5000 37280 5008 37344
rect 5072 37280 5088 37344
rect 5152 37280 5168 37344
rect 5232 37280 5248 37344
rect 5312 37280 5328 37344
rect 5392 37280 5408 37344
rect 5472 37280 5488 37344
rect 5552 37280 5568 37344
rect 5632 37280 5648 37344
rect 5712 37280 5728 37344
rect 5792 37280 5808 37344
rect 5872 37280 5888 37344
rect 5952 37280 5968 37344
rect 6032 37280 6048 37344
rect 6112 37280 6128 37344
rect 6192 37280 6208 37344
rect 6272 37280 6288 37344
rect 6352 37280 6368 37344
rect 6432 37280 6448 37344
rect 6512 37280 6528 37344
rect 6592 37280 6608 37344
rect 6672 37280 6688 37344
rect 6752 37280 6768 37344
rect 6832 37280 6848 37344
rect 6912 37280 6928 37344
rect 6992 37280 7008 37344
rect 7072 37280 7088 37344
rect 7152 37280 7168 37344
rect 7232 37280 7248 37344
rect 7312 37280 7328 37344
rect 7392 37280 7408 37344
rect 7472 37280 7488 37344
rect 7552 37280 7568 37344
rect 7632 37280 7648 37344
rect 7712 37280 7728 37344
rect 7792 37280 7808 37344
rect 7872 37280 7888 37344
rect 7952 37280 7968 37344
rect 8032 37280 8048 37344
rect 8112 37280 8128 37344
rect 8192 37280 8208 37344
rect 8272 37280 8288 37344
rect 8352 37280 8368 37344
rect 8432 37280 8448 37344
rect 8512 37280 8528 37344
rect 8592 37280 8608 37344
rect 8672 37280 8688 37344
rect 8752 37280 8768 37344
rect 8832 37280 8848 37344
rect 8912 37280 8928 37344
rect 8992 37280 9000 37344
rect 5000 37264 9000 37280
rect 5000 37200 5008 37264
rect 5072 37200 5088 37264
rect 5152 37200 5168 37264
rect 5232 37200 5248 37264
rect 5312 37200 5328 37264
rect 5392 37200 5408 37264
rect 5472 37200 5488 37264
rect 5552 37200 5568 37264
rect 5632 37200 5648 37264
rect 5712 37200 5728 37264
rect 5792 37200 5808 37264
rect 5872 37200 5888 37264
rect 5952 37200 5968 37264
rect 6032 37200 6048 37264
rect 6112 37200 6128 37264
rect 6192 37200 6208 37264
rect 6272 37200 6288 37264
rect 6352 37200 6368 37264
rect 6432 37200 6448 37264
rect 6512 37200 6528 37264
rect 6592 37200 6608 37264
rect 6672 37200 6688 37264
rect 6752 37200 6768 37264
rect 6832 37200 6848 37264
rect 6912 37200 6928 37264
rect 6992 37200 7008 37264
rect 7072 37200 7088 37264
rect 7152 37200 7168 37264
rect 7232 37200 7248 37264
rect 7312 37200 7328 37264
rect 7392 37200 7408 37264
rect 7472 37200 7488 37264
rect 7552 37200 7568 37264
rect 7632 37200 7648 37264
rect 7712 37200 7728 37264
rect 7792 37200 7808 37264
rect 7872 37200 7888 37264
rect 7952 37200 7968 37264
rect 8032 37200 8048 37264
rect 8112 37200 8128 37264
rect 8192 37200 8208 37264
rect 8272 37200 8288 37264
rect 8352 37200 8368 37264
rect 8432 37200 8448 37264
rect 8512 37200 8528 37264
rect 8592 37200 8608 37264
rect 8672 37200 8688 37264
rect 8752 37200 8768 37264
rect 8832 37200 8848 37264
rect 8912 37200 8928 37264
rect 8992 37200 9000 37264
rect 5000 37184 9000 37200
rect 5000 37120 5008 37184
rect 5072 37120 5088 37184
rect 5152 37120 5168 37184
rect 5232 37120 5248 37184
rect 5312 37120 5328 37184
rect 5392 37120 5408 37184
rect 5472 37120 5488 37184
rect 5552 37120 5568 37184
rect 5632 37120 5648 37184
rect 5712 37120 5728 37184
rect 5792 37120 5808 37184
rect 5872 37120 5888 37184
rect 5952 37120 5968 37184
rect 6032 37120 6048 37184
rect 6112 37120 6128 37184
rect 6192 37120 6208 37184
rect 6272 37120 6288 37184
rect 6352 37120 6368 37184
rect 6432 37120 6448 37184
rect 6512 37120 6528 37184
rect 6592 37120 6608 37184
rect 6672 37120 6688 37184
rect 6752 37120 6768 37184
rect 6832 37120 6848 37184
rect 6912 37120 6928 37184
rect 6992 37120 7008 37184
rect 7072 37120 7088 37184
rect 7152 37120 7168 37184
rect 7232 37120 7248 37184
rect 7312 37120 7328 37184
rect 7392 37120 7408 37184
rect 7472 37120 7488 37184
rect 7552 37120 7568 37184
rect 7632 37120 7648 37184
rect 7712 37120 7728 37184
rect 7792 37120 7808 37184
rect 7872 37120 7888 37184
rect 7952 37120 7968 37184
rect 8032 37120 8048 37184
rect 8112 37120 8128 37184
rect 8192 37120 8208 37184
rect 8272 37120 8288 37184
rect 8352 37120 8368 37184
rect 8432 37120 8448 37184
rect 8512 37120 8528 37184
rect 8592 37120 8608 37184
rect 8672 37120 8688 37184
rect 8752 37120 8768 37184
rect 8832 37120 8848 37184
rect 8912 37120 8928 37184
rect 8992 37120 9000 37184
rect 5000 37104 9000 37120
rect 5000 37040 5008 37104
rect 5072 37040 5088 37104
rect 5152 37040 5168 37104
rect 5232 37040 5248 37104
rect 5312 37040 5328 37104
rect 5392 37040 5408 37104
rect 5472 37040 5488 37104
rect 5552 37040 5568 37104
rect 5632 37040 5648 37104
rect 5712 37040 5728 37104
rect 5792 37040 5808 37104
rect 5872 37040 5888 37104
rect 5952 37040 5968 37104
rect 6032 37040 6048 37104
rect 6112 37040 6128 37104
rect 6192 37040 6208 37104
rect 6272 37040 6288 37104
rect 6352 37040 6368 37104
rect 6432 37040 6448 37104
rect 6512 37040 6528 37104
rect 6592 37040 6608 37104
rect 6672 37040 6688 37104
rect 6752 37040 6768 37104
rect 6832 37040 6848 37104
rect 6912 37040 6928 37104
rect 6992 37040 7008 37104
rect 7072 37040 7088 37104
rect 7152 37040 7168 37104
rect 7232 37040 7248 37104
rect 7312 37040 7328 37104
rect 7392 37040 7408 37104
rect 7472 37040 7488 37104
rect 7552 37040 7568 37104
rect 7632 37040 7648 37104
rect 7712 37040 7728 37104
rect 7792 37040 7808 37104
rect 7872 37040 7888 37104
rect 7952 37040 7968 37104
rect 8032 37040 8048 37104
rect 8112 37040 8128 37104
rect 8192 37040 8208 37104
rect 8272 37040 8288 37104
rect 8352 37040 8368 37104
rect 8432 37040 8448 37104
rect 8512 37040 8528 37104
rect 8592 37040 8608 37104
rect 8672 37040 8688 37104
rect 8752 37040 8768 37104
rect 8832 37040 8848 37104
rect 8912 37040 8928 37104
rect 8992 37040 9000 37104
rect 5000 37024 9000 37040
rect 5000 36960 5008 37024
rect 5072 36960 5088 37024
rect 5152 36960 5168 37024
rect 5232 36960 5248 37024
rect 5312 36960 5328 37024
rect 5392 36960 5408 37024
rect 5472 36960 5488 37024
rect 5552 36960 5568 37024
rect 5632 36960 5648 37024
rect 5712 36960 5728 37024
rect 5792 36960 5808 37024
rect 5872 36960 5888 37024
rect 5952 36960 5968 37024
rect 6032 36960 6048 37024
rect 6112 36960 6128 37024
rect 6192 36960 6208 37024
rect 6272 36960 6288 37024
rect 6352 36960 6368 37024
rect 6432 36960 6448 37024
rect 6512 36960 6528 37024
rect 6592 36960 6608 37024
rect 6672 36960 6688 37024
rect 6752 36960 6768 37024
rect 6832 36960 6848 37024
rect 6912 36960 6928 37024
rect 6992 36960 7008 37024
rect 7072 36960 7088 37024
rect 7152 36960 7168 37024
rect 7232 36960 7248 37024
rect 7312 36960 7328 37024
rect 7392 36960 7408 37024
rect 7472 36960 7488 37024
rect 7552 36960 7568 37024
rect 7632 36960 7648 37024
rect 7712 36960 7728 37024
rect 7792 36960 7808 37024
rect 7872 36960 7888 37024
rect 7952 36960 7968 37024
rect 8032 36960 8048 37024
rect 8112 36960 8128 37024
rect 8192 36960 8208 37024
rect 8272 36960 8288 37024
rect 8352 36960 8368 37024
rect 8432 36960 8448 37024
rect 8512 36960 8528 37024
rect 8592 36960 8608 37024
rect 8672 36960 8688 37024
rect 8752 36960 8768 37024
rect 8832 36960 8848 37024
rect 8912 36960 8928 37024
rect 8992 36960 9000 37024
rect 5000 36944 9000 36960
rect 5000 36880 5008 36944
rect 5072 36880 5088 36944
rect 5152 36880 5168 36944
rect 5232 36880 5248 36944
rect 5312 36880 5328 36944
rect 5392 36880 5408 36944
rect 5472 36880 5488 36944
rect 5552 36880 5568 36944
rect 5632 36880 5648 36944
rect 5712 36880 5728 36944
rect 5792 36880 5808 36944
rect 5872 36880 5888 36944
rect 5952 36880 5968 36944
rect 6032 36880 6048 36944
rect 6112 36880 6128 36944
rect 6192 36880 6208 36944
rect 6272 36880 6288 36944
rect 6352 36880 6368 36944
rect 6432 36880 6448 36944
rect 6512 36880 6528 36944
rect 6592 36880 6608 36944
rect 6672 36880 6688 36944
rect 6752 36880 6768 36944
rect 6832 36880 6848 36944
rect 6912 36880 6928 36944
rect 6992 36880 7008 36944
rect 7072 36880 7088 36944
rect 7152 36880 7168 36944
rect 7232 36880 7248 36944
rect 7312 36880 7328 36944
rect 7392 36880 7408 36944
rect 7472 36880 7488 36944
rect 7552 36880 7568 36944
rect 7632 36880 7648 36944
rect 7712 36880 7728 36944
rect 7792 36880 7808 36944
rect 7872 36880 7888 36944
rect 7952 36880 7968 36944
rect 8032 36880 8048 36944
rect 8112 36880 8128 36944
rect 8192 36880 8208 36944
rect 8272 36880 8288 36944
rect 8352 36880 8368 36944
rect 8432 36880 8448 36944
rect 8512 36880 8528 36944
rect 8592 36880 8608 36944
rect 8672 36880 8688 36944
rect 8752 36880 8768 36944
rect 8832 36880 8848 36944
rect 8912 36880 8928 36944
rect 8992 36880 9000 36944
rect 5000 36864 9000 36880
rect 5000 36800 5008 36864
rect 5072 36800 5088 36864
rect 5152 36800 5168 36864
rect 5232 36800 5248 36864
rect 5312 36800 5328 36864
rect 5392 36800 5408 36864
rect 5472 36800 5488 36864
rect 5552 36800 5568 36864
rect 5632 36800 5648 36864
rect 5712 36800 5728 36864
rect 5792 36800 5808 36864
rect 5872 36800 5888 36864
rect 5952 36800 5968 36864
rect 6032 36800 6048 36864
rect 6112 36800 6128 36864
rect 6192 36800 6208 36864
rect 6272 36800 6288 36864
rect 6352 36800 6368 36864
rect 6432 36800 6448 36864
rect 6512 36800 6528 36864
rect 6592 36800 6608 36864
rect 6672 36800 6688 36864
rect 6752 36800 6768 36864
rect 6832 36800 6848 36864
rect 6912 36800 6928 36864
rect 6992 36800 7008 36864
rect 7072 36800 7088 36864
rect 7152 36800 7168 36864
rect 7232 36800 7248 36864
rect 7312 36800 7328 36864
rect 7392 36800 7408 36864
rect 7472 36800 7488 36864
rect 7552 36800 7568 36864
rect 7632 36800 7648 36864
rect 7712 36800 7728 36864
rect 7792 36800 7808 36864
rect 7872 36800 7888 36864
rect 7952 36800 7968 36864
rect 8032 36800 8048 36864
rect 8112 36800 8128 36864
rect 8192 36800 8208 36864
rect 8272 36800 8288 36864
rect 8352 36800 8368 36864
rect 8432 36800 8448 36864
rect 8512 36800 8528 36864
rect 8592 36800 8608 36864
rect 8672 36800 8688 36864
rect 8752 36800 8768 36864
rect 8832 36800 8848 36864
rect 8912 36800 8928 36864
rect 8992 36800 9000 36864
rect 5000 36784 9000 36800
rect 5000 36720 5008 36784
rect 5072 36720 5088 36784
rect 5152 36720 5168 36784
rect 5232 36720 5248 36784
rect 5312 36720 5328 36784
rect 5392 36720 5408 36784
rect 5472 36720 5488 36784
rect 5552 36720 5568 36784
rect 5632 36720 5648 36784
rect 5712 36720 5728 36784
rect 5792 36720 5808 36784
rect 5872 36720 5888 36784
rect 5952 36720 5968 36784
rect 6032 36720 6048 36784
rect 6112 36720 6128 36784
rect 6192 36720 6208 36784
rect 6272 36720 6288 36784
rect 6352 36720 6368 36784
rect 6432 36720 6448 36784
rect 6512 36720 6528 36784
rect 6592 36720 6608 36784
rect 6672 36720 6688 36784
rect 6752 36720 6768 36784
rect 6832 36720 6848 36784
rect 6912 36720 6928 36784
rect 6992 36720 7008 36784
rect 7072 36720 7088 36784
rect 7152 36720 7168 36784
rect 7232 36720 7248 36784
rect 7312 36720 7328 36784
rect 7392 36720 7408 36784
rect 7472 36720 7488 36784
rect 7552 36720 7568 36784
rect 7632 36720 7648 36784
rect 7712 36720 7728 36784
rect 7792 36720 7808 36784
rect 7872 36720 7888 36784
rect 7952 36720 7968 36784
rect 8032 36720 8048 36784
rect 8112 36720 8128 36784
rect 8192 36720 8208 36784
rect 8272 36720 8288 36784
rect 8352 36720 8368 36784
rect 8432 36720 8448 36784
rect 8512 36720 8528 36784
rect 8592 36720 8608 36784
rect 8672 36720 8688 36784
rect 8752 36720 8768 36784
rect 8832 36720 8848 36784
rect 8912 36720 8928 36784
rect 8992 36720 9000 36784
rect 5000 36704 9000 36720
rect 5000 36640 5008 36704
rect 5072 36640 5088 36704
rect 5152 36640 5168 36704
rect 5232 36640 5248 36704
rect 5312 36640 5328 36704
rect 5392 36640 5408 36704
rect 5472 36640 5488 36704
rect 5552 36640 5568 36704
rect 5632 36640 5648 36704
rect 5712 36640 5728 36704
rect 5792 36640 5808 36704
rect 5872 36640 5888 36704
rect 5952 36640 5968 36704
rect 6032 36640 6048 36704
rect 6112 36640 6128 36704
rect 6192 36640 6208 36704
rect 6272 36640 6288 36704
rect 6352 36640 6368 36704
rect 6432 36640 6448 36704
rect 6512 36640 6528 36704
rect 6592 36640 6608 36704
rect 6672 36640 6688 36704
rect 6752 36640 6768 36704
rect 6832 36640 6848 36704
rect 6912 36640 6928 36704
rect 6992 36640 7008 36704
rect 7072 36640 7088 36704
rect 7152 36640 7168 36704
rect 7232 36640 7248 36704
rect 7312 36640 7328 36704
rect 7392 36640 7408 36704
rect 7472 36640 7488 36704
rect 7552 36640 7568 36704
rect 7632 36640 7648 36704
rect 7712 36640 7728 36704
rect 7792 36640 7808 36704
rect 7872 36640 7888 36704
rect 7952 36640 7968 36704
rect 8032 36640 8048 36704
rect 8112 36640 8128 36704
rect 8192 36640 8208 36704
rect 8272 36640 8288 36704
rect 8352 36640 8368 36704
rect 8432 36640 8448 36704
rect 8512 36640 8528 36704
rect 8592 36640 8608 36704
rect 8672 36640 8688 36704
rect 8752 36640 8768 36704
rect 8832 36640 8848 36704
rect 8912 36640 8928 36704
rect 8992 36640 9000 36704
rect 5000 36624 9000 36640
rect 5000 36560 5008 36624
rect 5072 36560 5088 36624
rect 5152 36560 5168 36624
rect 5232 36560 5248 36624
rect 5312 36560 5328 36624
rect 5392 36560 5408 36624
rect 5472 36560 5488 36624
rect 5552 36560 5568 36624
rect 5632 36560 5648 36624
rect 5712 36560 5728 36624
rect 5792 36560 5808 36624
rect 5872 36560 5888 36624
rect 5952 36560 5968 36624
rect 6032 36560 6048 36624
rect 6112 36560 6128 36624
rect 6192 36560 6208 36624
rect 6272 36560 6288 36624
rect 6352 36560 6368 36624
rect 6432 36560 6448 36624
rect 6512 36560 6528 36624
rect 6592 36560 6608 36624
rect 6672 36560 6688 36624
rect 6752 36560 6768 36624
rect 6832 36560 6848 36624
rect 6912 36560 6928 36624
rect 6992 36560 7008 36624
rect 7072 36560 7088 36624
rect 7152 36560 7168 36624
rect 7232 36560 7248 36624
rect 7312 36560 7328 36624
rect 7392 36560 7408 36624
rect 7472 36560 7488 36624
rect 7552 36560 7568 36624
rect 7632 36560 7648 36624
rect 7712 36560 7728 36624
rect 7792 36560 7808 36624
rect 7872 36560 7888 36624
rect 7952 36560 7968 36624
rect 8032 36560 8048 36624
rect 8112 36560 8128 36624
rect 8192 36560 8208 36624
rect 8272 36560 8288 36624
rect 8352 36560 8368 36624
rect 8432 36560 8448 36624
rect 8512 36560 8528 36624
rect 8592 36560 8608 36624
rect 8672 36560 8688 36624
rect 8752 36560 8768 36624
rect 8832 36560 8848 36624
rect 8912 36560 8928 36624
rect 8992 36560 9000 36624
rect 5000 36544 9000 36560
rect 5000 36480 5008 36544
rect 5072 36480 5088 36544
rect 5152 36480 5168 36544
rect 5232 36480 5248 36544
rect 5312 36480 5328 36544
rect 5392 36480 5408 36544
rect 5472 36480 5488 36544
rect 5552 36480 5568 36544
rect 5632 36480 5648 36544
rect 5712 36480 5728 36544
rect 5792 36480 5808 36544
rect 5872 36480 5888 36544
rect 5952 36480 5968 36544
rect 6032 36480 6048 36544
rect 6112 36480 6128 36544
rect 6192 36480 6208 36544
rect 6272 36480 6288 36544
rect 6352 36480 6368 36544
rect 6432 36480 6448 36544
rect 6512 36480 6528 36544
rect 6592 36480 6608 36544
rect 6672 36480 6688 36544
rect 6752 36480 6768 36544
rect 6832 36480 6848 36544
rect 6912 36480 6928 36544
rect 6992 36480 7008 36544
rect 7072 36480 7088 36544
rect 7152 36480 7168 36544
rect 7232 36480 7248 36544
rect 7312 36480 7328 36544
rect 7392 36480 7408 36544
rect 7472 36480 7488 36544
rect 7552 36480 7568 36544
rect 7632 36480 7648 36544
rect 7712 36480 7728 36544
rect 7792 36480 7808 36544
rect 7872 36480 7888 36544
rect 7952 36480 7968 36544
rect 8032 36480 8048 36544
rect 8112 36480 8128 36544
rect 8192 36480 8208 36544
rect 8272 36480 8288 36544
rect 8352 36480 8368 36544
rect 8432 36480 8448 36544
rect 8512 36480 8528 36544
rect 8592 36480 8608 36544
rect 8672 36480 8688 36544
rect 8752 36480 8768 36544
rect 8832 36480 8848 36544
rect 8912 36480 8928 36544
rect 8992 36480 9000 36544
rect 5000 36464 9000 36480
rect 5000 36400 5008 36464
rect 5072 36400 5088 36464
rect 5152 36400 5168 36464
rect 5232 36400 5248 36464
rect 5312 36400 5328 36464
rect 5392 36400 5408 36464
rect 5472 36400 5488 36464
rect 5552 36400 5568 36464
rect 5632 36400 5648 36464
rect 5712 36400 5728 36464
rect 5792 36400 5808 36464
rect 5872 36400 5888 36464
rect 5952 36400 5968 36464
rect 6032 36400 6048 36464
rect 6112 36400 6128 36464
rect 6192 36400 6208 36464
rect 6272 36400 6288 36464
rect 6352 36400 6368 36464
rect 6432 36400 6448 36464
rect 6512 36400 6528 36464
rect 6592 36400 6608 36464
rect 6672 36400 6688 36464
rect 6752 36400 6768 36464
rect 6832 36400 6848 36464
rect 6912 36400 6928 36464
rect 6992 36400 7008 36464
rect 7072 36400 7088 36464
rect 7152 36400 7168 36464
rect 7232 36400 7248 36464
rect 7312 36400 7328 36464
rect 7392 36400 7408 36464
rect 7472 36400 7488 36464
rect 7552 36400 7568 36464
rect 7632 36400 7648 36464
rect 7712 36400 7728 36464
rect 7792 36400 7808 36464
rect 7872 36400 7888 36464
rect 7952 36400 7968 36464
rect 8032 36400 8048 36464
rect 8112 36400 8128 36464
rect 8192 36400 8208 36464
rect 8272 36400 8288 36464
rect 8352 36400 8368 36464
rect 8432 36400 8448 36464
rect 8512 36400 8528 36464
rect 8592 36400 8608 36464
rect 8672 36400 8688 36464
rect 8752 36400 8768 36464
rect 8832 36400 8848 36464
rect 8912 36400 8928 36464
rect 8992 36400 9000 36464
rect 5000 8992 9000 36400
rect 5000 8928 5008 8992
rect 5072 8928 5088 8992
rect 5152 8928 5168 8992
rect 5232 8928 5248 8992
rect 5312 8928 5328 8992
rect 5392 8928 5408 8992
rect 5472 8928 5488 8992
rect 5552 8928 5568 8992
rect 5632 8928 5648 8992
rect 5712 8928 5728 8992
rect 5792 8928 5808 8992
rect 5872 8928 5888 8992
rect 5952 8928 5968 8992
rect 6032 8928 6048 8992
rect 6112 8928 6128 8992
rect 6192 8928 6208 8992
rect 6272 8928 6288 8992
rect 6352 8928 6368 8992
rect 6432 8928 6448 8992
rect 6512 8928 6528 8992
rect 6592 8928 6608 8992
rect 6672 8928 6688 8992
rect 6752 8928 6768 8992
rect 6832 8928 6848 8992
rect 6912 8928 6928 8992
rect 6992 8928 7008 8992
rect 7072 8928 7088 8992
rect 7152 8928 7168 8992
rect 7232 8928 7248 8992
rect 7312 8928 7328 8992
rect 7392 8928 7408 8992
rect 7472 8928 7488 8992
rect 7552 8928 7568 8992
rect 7632 8928 7648 8992
rect 7712 8928 7728 8992
rect 7792 8928 7808 8992
rect 7872 8928 7888 8992
rect 7952 8928 7968 8992
rect 8032 8928 8048 8992
rect 8112 8928 8128 8992
rect 8192 8928 8208 8992
rect 8272 8928 8288 8992
rect 8352 8928 8368 8992
rect 8432 8928 8448 8992
rect 8512 8928 8528 8992
rect 8592 8928 8608 8992
rect 8672 8928 8688 8992
rect 8752 8928 8768 8992
rect 8832 8928 8848 8992
rect 8912 8928 8928 8992
rect 8992 8928 9000 8992
rect 5000 8912 9000 8928
rect 5000 8848 5008 8912
rect 5072 8848 5088 8912
rect 5152 8848 5168 8912
rect 5232 8848 5248 8912
rect 5312 8848 5328 8912
rect 5392 8848 5408 8912
rect 5472 8848 5488 8912
rect 5552 8848 5568 8912
rect 5632 8848 5648 8912
rect 5712 8848 5728 8912
rect 5792 8848 5808 8912
rect 5872 8848 5888 8912
rect 5952 8848 5968 8912
rect 6032 8848 6048 8912
rect 6112 8848 6128 8912
rect 6192 8848 6208 8912
rect 6272 8848 6288 8912
rect 6352 8848 6368 8912
rect 6432 8848 6448 8912
rect 6512 8848 6528 8912
rect 6592 8848 6608 8912
rect 6672 8848 6688 8912
rect 6752 8848 6768 8912
rect 6832 8848 6848 8912
rect 6912 8848 6928 8912
rect 6992 8848 7008 8912
rect 7072 8848 7088 8912
rect 7152 8848 7168 8912
rect 7232 8848 7248 8912
rect 7312 8848 7328 8912
rect 7392 8848 7408 8912
rect 7472 8848 7488 8912
rect 7552 8848 7568 8912
rect 7632 8848 7648 8912
rect 7712 8848 7728 8912
rect 7792 8848 7808 8912
rect 7872 8848 7888 8912
rect 7952 8848 7968 8912
rect 8032 8848 8048 8912
rect 8112 8848 8128 8912
rect 8192 8848 8208 8912
rect 8272 8848 8288 8912
rect 8352 8848 8368 8912
rect 8432 8848 8448 8912
rect 8512 8848 8528 8912
rect 8592 8848 8608 8912
rect 8672 8848 8688 8912
rect 8752 8848 8768 8912
rect 8832 8848 8848 8912
rect 8912 8848 8928 8912
rect 8992 8848 9000 8912
rect 5000 8832 9000 8848
rect 5000 8768 5008 8832
rect 5072 8768 5088 8832
rect 5152 8768 5168 8832
rect 5232 8768 5248 8832
rect 5312 8768 5328 8832
rect 5392 8768 5408 8832
rect 5472 8768 5488 8832
rect 5552 8768 5568 8832
rect 5632 8768 5648 8832
rect 5712 8768 5728 8832
rect 5792 8768 5808 8832
rect 5872 8768 5888 8832
rect 5952 8768 5968 8832
rect 6032 8768 6048 8832
rect 6112 8768 6128 8832
rect 6192 8768 6208 8832
rect 6272 8768 6288 8832
rect 6352 8768 6368 8832
rect 6432 8768 6448 8832
rect 6512 8768 6528 8832
rect 6592 8768 6608 8832
rect 6672 8768 6688 8832
rect 6752 8768 6768 8832
rect 6832 8768 6848 8832
rect 6912 8768 6928 8832
rect 6992 8768 7008 8832
rect 7072 8768 7088 8832
rect 7152 8768 7168 8832
rect 7232 8768 7248 8832
rect 7312 8768 7328 8832
rect 7392 8768 7408 8832
rect 7472 8768 7488 8832
rect 7552 8768 7568 8832
rect 7632 8768 7648 8832
rect 7712 8768 7728 8832
rect 7792 8768 7808 8832
rect 7872 8768 7888 8832
rect 7952 8768 7968 8832
rect 8032 8768 8048 8832
rect 8112 8768 8128 8832
rect 8192 8768 8208 8832
rect 8272 8768 8288 8832
rect 8352 8768 8368 8832
rect 8432 8768 8448 8832
rect 8512 8768 8528 8832
rect 8592 8768 8608 8832
rect 8672 8768 8688 8832
rect 8752 8768 8768 8832
rect 8832 8768 8848 8832
rect 8912 8768 8928 8832
rect 8992 8768 9000 8832
rect 5000 8752 9000 8768
rect 5000 8688 5008 8752
rect 5072 8688 5088 8752
rect 5152 8688 5168 8752
rect 5232 8688 5248 8752
rect 5312 8688 5328 8752
rect 5392 8688 5408 8752
rect 5472 8688 5488 8752
rect 5552 8688 5568 8752
rect 5632 8688 5648 8752
rect 5712 8688 5728 8752
rect 5792 8688 5808 8752
rect 5872 8688 5888 8752
rect 5952 8688 5968 8752
rect 6032 8688 6048 8752
rect 6112 8688 6128 8752
rect 6192 8688 6208 8752
rect 6272 8688 6288 8752
rect 6352 8688 6368 8752
rect 6432 8688 6448 8752
rect 6512 8688 6528 8752
rect 6592 8688 6608 8752
rect 6672 8688 6688 8752
rect 6752 8688 6768 8752
rect 6832 8688 6848 8752
rect 6912 8688 6928 8752
rect 6992 8688 7008 8752
rect 7072 8688 7088 8752
rect 7152 8688 7168 8752
rect 7232 8688 7248 8752
rect 7312 8688 7328 8752
rect 7392 8688 7408 8752
rect 7472 8688 7488 8752
rect 7552 8688 7568 8752
rect 7632 8688 7648 8752
rect 7712 8688 7728 8752
rect 7792 8688 7808 8752
rect 7872 8688 7888 8752
rect 7952 8688 7968 8752
rect 8032 8688 8048 8752
rect 8112 8688 8128 8752
rect 8192 8688 8208 8752
rect 8272 8688 8288 8752
rect 8352 8688 8368 8752
rect 8432 8688 8448 8752
rect 8512 8688 8528 8752
rect 8592 8688 8608 8752
rect 8672 8688 8688 8752
rect 8752 8688 8768 8752
rect 8832 8688 8848 8752
rect 8912 8688 8928 8752
rect 8992 8688 9000 8752
rect 5000 8672 9000 8688
rect 5000 8608 5008 8672
rect 5072 8608 5088 8672
rect 5152 8608 5168 8672
rect 5232 8608 5248 8672
rect 5312 8608 5328 8672
rect 5392 8608 5408 8672
rect 5472 8608 5488 8672
rect 5552 8608 5568 8672
rect 5632 8608 5648 8672
rect 5712 8608 5728 8672
rect 5792 8608 5808 8672
rect 5872 8608 5888 8672
rect 5952 8608 5968 8672
rect 6032 8608 6048 8672
rect 6112 8608 6128 8672
rect 6192 8608 6208 8672
rect 6272 8608 6288 8672
rect 6352 8608 6368 8672
rect 6432 8608 6448 8672
rect 6512 8608 6528 8672
rect 6592 8608 6608 8672
rect 6672 8608 6688 8672
rect 6752 8608 6768 8672
rect 6832 8608 6848 8672
rect 6912 8608 6928 8672
rect 6992 8608 7008 8672
rect 7072 8608 7088 8672
rect 7152 8608 7168 8672
rect 7232 8608 7248 8672
rect 7312 8608 7328 8672
rect 7392 8608 7408 8672
rect 7472 8608 7488 8672
rect 7552 8608 7568 8672
rect 7632 8608 7648 8672
rect 7712 8608 7728 8672
rect 7792 8608 7808 8672
rect 7872 8608 7888 8672
rect 7952 8608 7968 8672
rect 8032 8608 8048 8672
rect 8112 8608 8128 8672
rect 8192 8608 8208 8672
rect 8272 8608 8288 8672
rect 8352 8608 8368 8672
rect 8432 8608 8448 8672
rect 8512 8608 8528 8672
rect 8592 8608 8608 8672
rect 8672 8608 8688 8672
rect 8752 8608 8768 8672
rect 8832 8608 8848 8672
rect 8912 8608 8928 8672
rect 8992 8608 9000 8672
rect 5000 8592 9000 8608
rect 5000 8528 5008 8592
rect 5072 8528 5088 8592
rect 5152 8528 5168 8592
rect 5232 8528 5248 8592
rect 5312 8528 5328 8592
rect 5392 8528 5408 8592
rect 5472 8528 5488 8592
rect 5552 8528 5568 8592
rect 5632 8528 5648 8592
rect 5712 8528 5728 8592
rect 5792 8528 5808 8592
rect 5872 8528 5888 8592
rect 5952 8528 5968 8592
rect 6032 8528 6048 8592
rect 6112 8528 6128 8592
rect 6192 8528 6208 8592
rect 6272 8528 6288 8592
rect 6352 8528 6368 8592
rect 6432 8528 6448 8592
rect 6512 8528 6528 8592
rect 6592 8528 6608 8592
rect 6672 8528 6688 8592
rect 6752 8528 6768 8592
rect 6832 8528 6848 8592
rect 6912 8528 6928 8592
rect 6992 8528 7008 8592
rect 7072 8528 7088 8592
rect 7152 8528 7168 8592
rect 7232 8528 7248 8592
rect 7312 8528 7328 8592
rect 7392 8528 7408 8592
rect 7472 8528 7488 8592
rect 7552 8528 7568 8592
rect 7632 8528 7648 8592
rect 7712 8528 7728 8592
rect 7792 8528 7808 8592
rect 7872 8528 7888 8592
rect 7952 8528 7968 8592
rect 8032 8528 8048 8592
rect 8112 8528 8128 8592
rect 8192 8528 8208 8592
rect 8272 8528 8288 8592
rect 8352 8528 8368 8592
rect 8432 8528 8448 8592
rect 8512 8528 8528 8592
rect 8592 8528 8608 8592
rect 8672 8528 8688 8592
rect 8752 8528 8768 8592
rect 8832 8528 8848 8592
rect 8912 8528 8928 8592
rect 8992 8528 9000 8592
rect 5000 8512 9000 8528
rect 5000 8448 5008 8512
rect 5072 8448 5088 8512
rect 5152 8448 5168 8512
rect 5232 8448 5248 8512
rect 5312 8448 5328 8512
rect 5392 8448 5408 8512
rect 5472 8448 5488 8512
rect 5552 8448 5568 8512
rect 5632 8448 5648 8512
rect 5712 8448 5728 8512
rect 5792 8448 5808 8512
rect 5872 8448 5888 8512
rect 5952 8448 5968 8512
rect 6032 8448 6048 8512
rect 6112 8448 6128 8512
rect 6192 8448 6208 8512
rect 6272 8448 6288 8512
rect 6352 8448 6368 8512
rect 6432 8448 6448 8512
rect 6512 8448 6528 8512
rect 6592 8448 6608 8512
rect 6672 8448 6688 8512
rect 6752 8448 6768 8512
rect 6832 8448 6848 8512
rect 6912 8448 6928 8512
rect 6992 8448 7008 8512
rect 7072 8448 7088 8512
rect 7152 8448 7168 8512
rect 7232 8448 7248 8512
rect 7312 8448 7328 8512
rect 7392 8448 7408 8512
rect 7472 8448 7488 8512
rect 7552 8448 7568 8512
rect 7632 8448 7648 8512
rect 7712 8448 7728 8512
rect 7792 8448 7808 8512
rect 7872 8448 7888 8512
rect 7952 8448 7968 8512
rect 8032 8448 8048 8512
rect 8112 8448 8128 8512
rect 8192 8448 8208 8512
rect 8272 8448 8288 8512
rect 8352 8448 8368 8512
rect 8432 8448 8448 8512
rect 8512 8448 8528 8512
rect 8592 8448 8608 8512
rect 8672 8448 8688 8512
rect 8752 8448 8768 8512
rect 8832 8448 8848 8512
rect 8912 8448 8928 8512
rect 8992 8448 9000 8512
rect 5000 8432 9000 8448
rect 5000 8368 5008 8432
rect 5072 8368 5088 8432
rect 5152 8368 5168 8432
rect 5232 8368 5248 8432
rect 5312 8368 5328 8432
rect 5392 8368 5408 8432
rect 5472 8368 5488 8432
rect 5552 8368 5568 8432
rect 5632 8368 5648 8432
rect 5712 8368 5728 8432
rect 5792 8368 5808 8432
rect 5872 8368 5888 8432
rect 5952 8368 5968 8432
rect 6032 8368 6048 8432
rect 6112 8368 6128 8432
rect 6192 8368 6208 8432
rect 6272 8368 6288 8432
rect 6352 8368 6368 8432
rect 6432 8368 6448 8432
rect 6512 8368 6528 8432
rect 6592 8368 6608 8432
rect 6672 8368 6688 8432
rect 6752 8368 6768 8432
rect 6832 8368 6848 8432
rect 6912 8368 6928 8432
rect 6992 8368 7008 8432
rect 7072 8368 7088 8432
rect 7152 8368 7168 8432
rect 7232 8368 7248 8432
rect 7312 8368 7328 8432
rect 7392 8368 7408 8432
rect 7472 8368 7488 8432
rect 7552 8368 7568 8432
rect 7632 8368 7648 8432
rect 7712 8368 7728 8432
rect 7792 8368 7808 8432
rect 7872 8368 7888 8432
rect 7952 8368 7968 8432
rect 8032 8368 8048 8432
rect 8112 8368 8128 8432
rect 8192 8368 8208 8432
rect 8272 8368 8288 8432
rect 8352 8368 8368 8432
rect 8432 8368 8448 8432
rect 8512 8368 8528 8432
rect 8592 8368 8608 8432
rect 8672 8368 8688 8432
rect 8752 8368 8768 8432
rect 8832 8368 8848 8432
rect 8912 8368 8928 8432
rect 8992 8368 9000 8432
rect 5000 8352 9000 8368
rect 5000 8288 5008 8352
rect 5072 8288 5088 8352
rect 5152 8288 5168 8352
rect 5232 8288 5248 8352
rect 5312 8288 5328 8352
rect 5392 8288 5408 8352
rect 5472 8288 5488 8352
rect 5552 8288 5568 8352
rect 5632 8288 5648 8352
rect 5712 8288 5728 8352
rect 5792 8288 5808 8352
rect 5872 8288 5888 8352
rect 5952 8288 5968 8352
rect 6032 8288 6048 8352
rect 6112 8288 6128 8352
rect 6192 8288 6208 8352
rect 6272 8288 6288 8352
rect 6352 8288 6368 8352
rect 6432 8288 6448 8352
rect 6512 8288 6528 8352
rect 6592 8288 6608 8352
rect 6672 8288 6688 8352
rect 6752 8288 6768 8352
rect 6832 8288 6848 8352
rect 6912 8288 6928 8352
rect 6992 8288 7008 8352
rect 7072 8288 7088 8352
rect 7152 8288 7168 8352
rect 7232 8288 7248 8352
rect 7312 8288 7328 8352
rect 7392 8288 7408 8352
rect 7472 8288 7488 8352
rect 7552 8288 7568 8352
rect 7632 8288 7648 8352
rect 7712 8288 7728 8352
rect 7792 8288 7808 8352
rect 7872 8288 7888 8352
rect 7952 8288 7968 8352
rect 8032 8288 8048 8352
rect 8112 8288 8128 8352
rect 8192 8288 8208 8352
rect 8272 8288 8288 8352
rect 8352 8288 8368 8352
rect 8432 8288 8448 8352
rect 8512 8288 8528 8352
rect 8592 8288 8608 8352
rect 8672 8288 8688 8352
rect 8752 8288 8768 8352
rect 8832 8288 8848 8352
rect 8912 8288 8928 8352
rect 8992 8288 9000 8352
rect 5000 8272 9000 8288
rect 5000 8208 5008 8272
rect 5072 8208 5088 8272
rect 5152 8208 5168 8272
rect 5232 8208 5248 8272
rect 5312 8208 5328 8272
rect 5392 8208 5408 8272
rect 5472 8208 5488 8272
rect 5552 8208 5568 8272
rect 5632 8208 5648 8272
rect 5712 8208 5728 8272
rect 5792 8208 5808 8272
rect 5872 8208 5888 8272
rect 5952 8208 5968 8272
rect 6032 8208 6048 8272
rect 6112 8208 6128 8272
rect 6192 8208 6208 8272
rect 6272 8208 6288 8272
rect 6352 8208 6368 8272
rect 6432 8208 6448 8272
rect 6512 8208 6528 8272
rect 6592 8208 6608 8272
rect 6672 8208 6688 8272
rect 6752 8208 6768 8272
rect 6832 8208 6848 8272
rect 6912 8208 6928 8272
rect 6992 8208 7008 8272
rect 7072 8208 7088 8272
rect 7152 8208 7168 8272
rect 7232 8208 7248 8272
rect 7312 8208 7328 8272
rect 7392 8208 7408 8272
rect 7472 8208 7488 8272
rect 7552 8208 7568 8272
rect 7632 8208 7648 8272
rect 7712 8208 7728 8272
rect 7792 8208 7808 8272
rect 7872 8208 7888 8272
rect 7952 8208 7968 8272
rect 8032 8208 8048 8272
rect 8112 8208 8128 8272
rect 8192 8208 8208 8272
rect 8272 8208 8288 8272
rect 8352 8208 8368 8272
rect 8432 8208 8448 8272
rect 8512 8208 8528 8272
rect 8592 8208 8608 8272
rect 8672 8208 8688 8272
rect 8752 8208 8768 8272
rect 8832 8208 8848 8272
rect 8912 8208 8928 8272
rect 8992 8208 9000 8272
rect 5000 8192 9000 8208
rect 5000 8128 5008 8192
rect 5072 8128 5088 8192
rect 5152 8128 5168 8192
rect 5232 8128 5248 8192
rect 5312 8128 5328 8192
rect 5392 8128 5408 8192
rect 5472 8128 5488 8192
rect 5552 8128 5568 8192
rect 5632 8128 5648 8192
rect 5712 8128 5728 8192
rect 5792 8128 5808 8192
rect 5872 8128 5888 8192
rect 5952 8128 5968 8192
rect 6032 8128 6048 8192
rect 6112 8128 6128 8192
rect 6192 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6528 8192
rect 6592 8128 6608 8192
rect 6672 8128 6688 8192
rect 6752 8128 6768 8192
rect 6832 8128 6848 8192
rect 6912 8128 6928 8192
rect 6992 8128 7008 8192
rect 7072 8128 7088 8192
rect 7152 8128 7168 8192
rect 7232 8128 7248 8192
rect 7312 8128 7328 8192
rect 7392 8128 7408 8192
rect 7472 8128 7488 8192
rect 7552 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7888 8192
rect 7952 8128 7968 8192
rect 8032 8128 8048 8192
rect 8112 8128 8128 8192
rect 8192 8128 8208 8192
rect 8272 8128 8288 8192
rect 8352 8128 8368 8192
rect 8432 8128 8448 8192
rect 8512 8128 8528 8192
rect 8592 8128 8608 8192
rect 8672 8128 8688 8192
rect 8752 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9000 8192
rect 5000 8112 9000 8128
rect 5000 8048 5008 8112
rect 5072 8048 5088 8112
rect 5152 8048 5168 8112
rect 5232 8048 5248 8112
rect 5312 8048 5328 8112
rect 5392 8048 5408 8112
rect 5472 8048 5488 8112
rect 5552 8048 5568 8112
rect 5632 8048 5648 8112
rect 5712 8048 5728 8112
rect 5792 8048 5808 8112
rect 5872 8048 5888 8112
rect 5952 8048 5968 8112
rect 6032 8048 6048 8112
rect 6112 8048 6128 8112
rect 6192 8048 6208 8112
rect 6272 8048 6288 8112
rect 6352 8048 6368 8112
rect 6432 8048 6448 8112
rect 6512 8048 6528 8112
rect 6592 8048 6608 8112
rect 6672 8048 6688 8112
rect 6752 8048 6768 8112
rect 6832 8048 6848 8112
rect 6912 8048 6928 8112
rect 6992 8048 7008 8112
rect 7072 8048 7088 8112
rect 7152 8048 7168 8112
rect 7232 8048 7248 8112
rect 7312 8048 7328 8112
rect 7392 8048 7408 8112
rect 7472 8048 7488 8112
rect 7552 8048 7568 8112
rect 7632 8048 7648 8112
rect 7712 8048 7728 8112
rect 7792 8048 7808 8112
rect 7872 8048 7888 8112
rect 7952 8048 7968 8112
rect 8032 8048 8048 8112
rect 8112 8048 8128 8112
rect 8192 8048 8208 8112
rect 8272 8048 8288 8112
rect 8352 8048 8368 8112
rect 8432 8048 8448 8112
rect 8512 8048 8528 8112
rect 8592 8048 8608 8112
rect 8672 8048 8688 8112
rect 8752 8048 8768 8112
rect 8832 8048 8848 8112
rect 8912 8048 8928 8112
rect 8992 8048 9000 8112
rect 5000 8032 9000 8048
rect 5000 7968 5008 8032
rect 5072 7968 5088 8032
rect 5152 7968 5168 8032
rect 5232 7968 5248 8032
rect 5312 7968 5328 8032
rect 5392 7968 5408 8032
rect 5472 7968 5488 8032
rect 5552 7968 5568 8032
rect 5632 7968 5648 8032
rect 5712 7968 5728 8032
rect 5792 7968 5808 8032
rect 5872 7968 5888 8032
rect 5952 7968 5968 8032
rect 6032 7968 6048 8032
rect 6112 7968 6128 8032
rect 6192 7968 6208 8032
rect 6272 7968 6288 8032
rect 6352 7968 6368 8032
rect 6432 7968 6448 8032
rect 6512 7968 6528 8032
rect 6592 7968 6608 8032
rect 6672 7968 6688 8032
rect 6752 7968 6768 8032
rect 6832 7968 6848 8032
rect 6912 7968 6928 8032
rect 6992 7968 7008 8032
rect 7072 7968 7088 8032
rect 7152 7968 7168 8032
rect 7232 7968 7248 8032
rect 7312 7968 7328 8032
rect 7392 7968 7408 8032
rect 7472 7968 7488 8032
rect 7552 7968 7568 8032
rect 7632 7968 7648 8032
rect 7712 7968 7728 8032
rect 7792 7968 7808 8032
rect 7872 7968 7888 8032
rect 7952 7968 7968 8032
rect 8032 7968 8048 8032
rect 8112 7968 8128 8032
rect 8192 7968 8208 8032
rect 8272 7968 8288 8032
rect 8352 7968 8368 8032
rect 8432 7968 8448 8032
rect 8512 7968 8528 8032
rect 8592 7968 8608 8032
rect 8672 7968 8688 8032
rect 8752 7968 8768 8032
rect 8832 7968 8848 8032
rect 8912 7968 8928 8032
rect 8992 7968 9000 8032
rect 5000 7952 9000 7968
rect 5000 7888 5008 7952
rect 5072 7888 5088 7952
rect 5152 7888 5168 7952
rect 5232 7888 5248 7952
rect 5312 7888 5328 7952
rect 5392 7888 5408 7952
rect 5472 7888 5488 7952
rect 5552 7888 5568 7952
rect 5632 7888 5648 7952
rect 5712 7888 5728 7952
rect 5792 7888 5808 7952
rect 5872 7888 5888 7952
rect 5952 7888 5968 7952
rect 6032 7888 6048 7952
rect 6112 7888 6128 7952
rect 6192 7888 6208 7952
rect 6272 7888 6288 7952
rect 6352 7888 6368 7952
rect 6432 7888 6448 7952
rect 6512 7888 6528 7952
rect 6592 7888 6608 7952
rect 6672 7888 6688 7952
rect 6752 7888 6768 7952
rect 6832 7888 6848 7952
rect 6912 7888 6928 7952
rect 6992 7888 7008 7952
rect 7072 7888 7088 7952
rect 7152 7888 7168 7952
rect 7232 7888 7248 7952
rect 7312 7888 7328 7952
rect 7392 7888 7408 7952
rect 7472 7888 7488 7952
rect 7552 7888 7568 7952
rect 7632 7888 7648 7952
rect 7712 7888 7728 7952
rect 7792 7888 7808 7952
rect 7872 7888 7888 7952
rect 7952 7888 7968 7952
rect 8032 7888 8048 7952
rect 8112 7888 8128 7952
rect 8192 7888 8208 7952
rect 8272 7888 8288 7952
rect 8352 7888 8368 7952
rect 8432 7888 8448 7952
rect 8512 7888 8528 7952
rect 8592 7888 8608 7952
rect 8672 7888 8688 7952
rect 8752 7888 8768 7952
rect 8832 7888 8848 7952
rect 8912 7888 8928 7952
rect 8992 7888 9000 7952
rect 5000 7872 9000 7888
rect 5000 7808 5008 7872
rect 5072 7808 5088 7872
rect 5152 7808 5168 7872
rect 5232 7808 5248 7872
rect 5312 7808 5328 7872
rect 5392 7808 5408 7872
rect 5472 7808 5488 7872
rect 5552 7808 5568 7872
rect 5632 7808 5648 7872
rect 5712 7808 5728 7872
rect 5792 7808 5808 7872
rect 5872 7808 5888 7872
rect 5952 7808 5968 7872
rect 6032 7808 6048 7872
rect 6112 7808 6128 7872
rect 6192 7808 6208 7872
rect 6272 7808 6288 7872
rect 6352 7808 6368 7872
rect 6432 7808 6448 7872
rect 6512 7808 6528 7872
rect 6592 7808 6608 7872
rect 6672 7808 6688 7872
rect 6752 7808 6768 7872
rect 6832 7808 6848 7872
rect 6912 7808 6928 7872
rect 6992 7808 7008 7872
rect 7072 7808 7088 7872
rect 7152 7808 7168 7872
rect 7232 7808 7248 7872
rect 7312 7808 7328 7872
rect 7392 7808 7408 7872
rect 7472 7808 7488 7872
rect 7552 7808 7568 7872
rect 7632 7808 7648 7872
rect 7712 7808 7728 7872
rect 7792 7808 7808 7872
rect 7872 7808 7888 7872
rect 7952 7808 7968 7872
rect 8032 7808 8048 7872
rect 8112 7808 8128 7872
rect 8192 7808 8208 7872
rect 8272 7808 8288 7872
rect 8352 7808 8368 7872
rect 8432 7808 8448 7872
rect 8512 7808 8528 7872
rect 8592 7808 8608 7872
rect 8672 7808 8688 7872
rect 8752 7808 8768 7872
rect 8832 7808 8848 7872
rect 8912 7808 8928 7872
rect 8992 7808 9000 7872
rect 5000 7792 9000 7808
rect 5000 7728 5008 7792
rect 5072 7728 5088 7792
rect 5152 7728 5168 7792
rect 5232 7728 5248 7792
rect 5312 7728 5328 7792
rect 5392 7728 5408 7792
rect 5472 7728 5488 7792
rect 5552 7728 5568 7792
rect 5632 7728 5648 7792
rect 5712 7728 5728 7792
rect 5792 7728 5808 7792
rect 5872 7728 5888 7792
rect 5952 7728 5968 7792
rect 6032 7728 6048 7792
rect 6112 7728 6128 7792
rect 6192 7728 6208 7792
rect 6272 7728 6288 7792
rect 6352 7728 6368 7792
rect 6432 7728 6448 7792
rect 6512 7728 6528 7792
rect 6592 7728 6608 7792
rect 6672 7728 6688 7792
rect 6752 7728 6768 7792
rect 6832 7728 6848 7792
rect 6912 7728 6928 7792
rect 6992 7728 7008 7792
rect 7072 7728 7088 7792
rect 7152 7728 7168 7792
rect 7232 7728 7248 7792
rect 7312 7728 7328 7792
rect 7392 7728 7408 7792
rect 7472 7728 7488 7792
rect 7552 7728 7568 7792
rect 7632 7728 7648 7792
rect 7712 7728 7728 7792
rect 7792 7728 7808 7792
rect 7872 7728 7888 7792
rect 7952 7728 7968 7792
rect 8032 7728 8048 7792
rect 8112 7728 8128 7792
rect 8192 7728 8208 7792
rect 8272 7728 8288 7792
rect 8352 7728 8368 7792
rect 8432 7728 8448 7792
rect 8512 7728 8528 7792
rect 8592 7728 8608 7792
rect 8672 7728 8688 7792
rect 8752 7728 8768 7792
rect 8832 7728 8848 7792
rect 8912 7728 8928 7792
rect 8992 7728 9000 7792
rect 5000 7712 9000 7728
rect 5000 7648 5008 7712
rect 5072 7648 5088 7712
rect 5152 7648 5168 7712
rect 5232 7648 5248 7712
rect 5312 7648 5328 7712
rect 5392 7648 5408 7712
rect 5472 7648 5488 7712
rect 5552 7648 5568 7712
rect 5632 7648 5648 7712
rect 5712 7648 5728 7712
rect 5792 7648 5808 7712
rect 5872 7648 5888 7712
rect 5952 7648 5968 7712
rect 6032 7648 6048 7712
rect 6112 7648 6128 7712
rect 6192 7648 6208 7712
rect 6272 7648 6288 7712
rect 6352 7648 6368 7712
rect 6432 7648 6448 7712
rect 6512 7648 6528 7712
rect 6592 7648 6608 7712
rect 6672 7648 6688 7712
rect 6752 7648 6768 7712
rect 6832 7648 6848 7712
rect 6912 7648 6928 7712
rect 6992 7648 7008 7712
rect 7072 7648 7088 7712
rect 7152 7648 7168 7712
rect 7232 7648 7248 7712
rect 7312 7648 7328 7712
rect 7392 7648 7408 7712
rect 7472 7648 7488 7712
rect 7552 7648 7568 7712
rect 7632 7648 7648 7712
rect 7712 7648 7728 7712
rect 7792 7648 7808 7712
rect 7872 7648 7888 7712
rect 7952 7648 7968 7712
rect 8032 7648 8048 7712
rect 8112 7648 8128 7712
rect 8192 7648 8208 7712
rect 8272 7648 8288 7712
rect 8352 7648 8368 7712
rect 8432 7648 8448 7712
rect 8512 7648 8528 7712
rect 8592 7648 8608 7712
rect 8672 7648 8688 7712
rect 8752 7648 8768 7712
rect 8832 7648 8848 7712
rect 8912 7648 8928 7712
rect 8992 7648 9000 7712
rect 5000 7632 9000 7648
rect 5000 7568 5008 7632
rect 5072 7568 5088 7632
rect 5152 7568 5168 7632
rect 5232 7568 5248 7632
rect 5312 7568 5328 7632
rect 5392 7568 5408 7632
rect 5472 7568 5488 7632
rect 5552 7568 5568 7632
rect 5632 7568 5648 7632
rect 5712 7568 5728 7632
rect 5792 7568 5808 7632
rect 5872 7568 5888 7632
rect 5952 7568 5968 7632
rect 6032 7568 6048 7632
rect 6112 7568 6128 7632
rect 6192 7568 6208 7632
rect 6272 7568 6288 7632
rect 6352 7568 6368 7632
rect 6432 7568 6448 7632
rect 6512 7568 6528 7632
rect 6592 7568 6608 7632
rect 6672 7568 6688 7632
rect 6752 7568 6768 7632
rect 6832 7568 6848 7632
rect 6912 7568 6928 7632
rect 6992 7568 7008 7632
rect 7072 7568 7088 7632
rect 7152 7568 7168 7632
rect 7232 7568 7248 7632
rect 7312 7568 7328 7632
rect 7392 7568 7408 7632
rect 7472 7568 7488 7632
rect 7552 7568 7568 7632
rect 7632 7568 7648 7632
rect 7712 7568 7728 7632
rect 7792 7568 7808 7632
rect 7872 7568 7888 7632
rect 7952 7568 7968 7632
rect 8032 7568 8048 7632
rect 8112 7568 8128 7632
rect 8192 7568 8208 7632
rect 8272 7568 8288 7632
rect 8352 7568 8368 7632
rect 8432 7568 8448 7632
rect 8512 7568 8528 7632
rect 8592 7568 8608 7632
rect 8672 7568 8688 7632
rect 8752 7568 8768 7632
rect 8832 7568 8848 7632
rect 8912 7568 8928 7632
rect 8992 7568 9000 7632
rect 5000 7552 9000 7568
rect 5000 7488 5008 7552
rect 5072 7488 5088 7552
rect 5152 7488 5168 7552
rect 5232 7488 5248 7552
rect 5312 7488 5328 7552
rect 5392 7488 5408 7552
rect 5472 7488 5488 7552
rect 5552 7488 5568 7552
rect 5632 7488 5648 7552
rect 5712 7488 5728 7552
rect 5792 7488 5808 7552
rect 5872 7488 5888 7552
rect 5952 7488 5968 7552
rect 6032 7488 6048 7552
rect 6112 7488 6128 7552
rect 6192 7488 6208 7552
rect 6272 7488 6288 7552
rect 6352 7488 6368 7552
rect 6432 7488 6448 7552
rect 6512 7488 6528 7552
rect 6592 7488 6608 7552
rect 6672 7488 6688 7552
rect 6752 7488 6768 7552
rect 6832 7488 6848 7552
rect 6912 7488 6928 7552
rect 6992 7488 7008 7552
rect 7072 7488 7088 7552
rect 7152 7488 7168 7552
rect 7232 7488 7248 7552
rect 7312 7488 7328 7552
rect 7392 7488 7408 7552
rect 7472 7488 7488 7552
rect 7552 7488 7568 7552
rect 7632 7488 7648 7552
rect 7712 7488 7728 7552
rect 7792 7488 7808 7552
rect 7872 7488 7888 7552
rect 7952 7488 7968 7552
rect 8032 7488 8048 7552
rect 8112 7488 8128 7552
rect 8192 7488 8208 7552
rect 8272 7488 8288 7552
rect 8352 7488 8368 7552
rect 8432 7488 8448 7552
rect 8512 7488 8528 7552
rect 8592 7488 8608 7552
rect 8672 7488 8688 7552
rect 8752 7488 8768 7552
rect 8832 7488 8848 7552
rect 8912 7488 8928 7552
rect 8992 7488 9000 7552
rect 5000 7472 9000 7488
rect 5000 7408 5008 7472
rect 5072 7408 5088 7472
rect 5152 7408 5168 7472
rect 5232 7408 5248 7472
rect 5312 7408 5328 7472
rect 5392 7408 5408 7472
rect 5472 7408 5488 7472
rect 5552 7408 5568 7472
rect 5632 7408 5648 7472
rect 5712 7408 5728 7472
rect 5792 7408 5808 7472
rect 5872 7408 5888 7472
rect 5952 7408 5968 7472
rect 6032 7408 6048 7472
rect 6112 7408 6128 7472
rect 6192 7408 6208 7472
rect 6272 7408 6288 7472
rect 6352 7408 6368 7472
rect 6432 7408 6448 7472
rect 6512 7408 6528 7472
rect 6592 7408 6608 7472
rect 6672 7408 6688 7472
rect 6752 7408 6768 7472
rect 6832 7408 6848 7472
rect 6912 7408 6928 7472
rect 6992 7408 7008 7472
rect 7072 7408 7088 7472
rect 7152 7408 7168 7472
rect 7232 7408 7248 7472
rect 7312 7408 7328 7472
rect 7392 7408 7408 7472
rect 7472 7408 7488 7472
rect 7552 7408 7568 7472
rect 7632 7408 7648 7472
rect 7712 7408 7728 7472
rect 7792 7408 7808 7472
rect 7872 7408 7888 7472
rect 7952 7408 7968 7472
rect 8032 7408 8048 7472
rect 8112 7408 8128 7472
rect 8192 7408 8208 7472
rect 8272 7408 8288 7472
rect 8352 7408 8368 7472
rect 8432 7408 8448 7472
rect 8512 7408 8528 7472
rect 8592 7408 8608 7472
rect 8672 7408 8688 7472
rect 8752 7408 8768 7472
rect 8832 7408 8848 7472
rect 8912 7408 8928 7472
rect 8992 7408 9000 7472
rect 5000 7392 9000 7408
rect 5000 7328 5008 7392
rect 5072 7328 5088 7392
rect 5152 7328 5168 7392
rect 5232 7328 5248 7392
rect 5312 7328 5328 7392
rect 5392 7328 5408 7392
rect 5472 7328 5488 7392
rect 5552 7328 5568 7392
rect 5632 7328 5648 7392
rect 5712 7328 5728 7392
rect 5792 7328 5808 7392
rect 5872 7328 5888 7392
rect 5952 7328 5968 7392
rect 6032 7328 6048 7392
rect 6112 7328 6128 7392
rect 6192 7328 6208 7392
rect 6272 7328 6288 7392
rect 6352 7328 6368 7392
rect 6432 7328 6448 7392
rect 6512 7328 6528 7392
rect 6592 7328 6608 7392
rect 6672 7328 6688 7392
rect 6752 7328 6768 7392
rect 6832 7328 6848 7392
rect 6912 7328 6928 7392
rect 6992 7328 7008 7392
rect 7072 7328 7088 7392
rect 7152 7328 7168 7392
rect 7232 7328 7248 7392
rect 7312 7328 7328 7392
rect 7392 7328 7408 7392
rect 7472 7328 7488 7392
rect 7552 7328 7568 7392
rect 7632 7328 7648 7392
rect 7712 7328 7728 7392
rect 7792 7328 7808 7392
rect 7872 7328 7888 7392
rect 7952 7328 7968 7392
rect 8032 7328 8048 7392
rect 8112 7328 8128 7392
rect 8192 7328 8208 7392
rect 8272 7328 8288 7392
rect 8352 7328 8368 7392
rect 8432 7328 8448 7392
rect 8512 7328 8528 7392
rect 8592 7328 8608 7392
rect 8672 7328 8688 7392
rect 8752 7328 8768 7392
rect 8832 7328 8848 7392
rect 8912 7328 8928 7392
rect 8992 7328 9000 7392
rect 5000 7312 9000 7328
rect 5000 7248 5008 7312
rect 5072 7248 5088 7312
rect 5152 7248 5168 7312
rect 5232 7248 5248 7312
rect 5312 7248 5328 7312
rect 5392 7248 5408 7312
rect 5472 7248 5488 7312
rect 5552 7248 5568 7312
rect 5632 7248 5648 7312
rect 5712 7248 5728 7312
rect 5792 7248 5808 7312
rect 5872 7248 5888 7312
rect 5952 7248 5968 7312
rect 6032 7248 6048 7312
rect 6112 7248 6128 7312
rect 6192 7248 6208 7312
rect 6272 7248 6288 7312
rect 6352 7248 6368 7312
rect 6432 7248 6448 7312
rect 6512 7248 6528 7312
rect 6592 7248 6608 7312
rect 6672 7248 6688 7312
rect 6752 7248 6768 7312
rect 6832 7248 6848 7312
rect 6912 7248 6928 7312
rect 6992 7248 7008 7312
rect 7072 7248 7088 7312
rect 7152 7248 7168 7312
rect 7232 7248 7248 7312
rect 7312 7248 7328 7312
rect 7392 7248 7408 7312
rect 7472 7248 7488 7312
rect 7552 7248 7568 7312
rect 7632 7248 7648 7312
rect 7712 7248 7728 7312
rect 7792 7248 7808 7312
rect 7872 7248 7888 7312
rect 7952 7248 7968 7312
rect 8032 7248 8048 7312
rect 8112 7248 8128 7312
rect 8192 7248 8208 7312
rect 8272 7248 8288 7312
rect 8352 7248 8368 7312
rect 8432 7248 8448 7312
rect 8512 7248 8528 7312
rect 8592 7248 8608 7312
rect 8672 7248 8688 7312
rect 8752 7248 8768 7312
rect 8832 7248 8848 7312
rect 8912 7248 8928 7312
rect 8992 7248 9000 7312
rect 5000 7232 9000 7248
rect 5000 7168 5008 7232
rect 5072 7168 5088 7232
rect 5152 7168 5168 7232
rect 5232 7168 5248 7232
rect 5312 7168 5328 7232
rect 5392 7168 5408 7232
rect 5472 7168 5488 7232
rect 5552 7168 5568 7232
rect 5632 7168 5648 7232
rect 5712 7168 5728 7232
rect 5792 7168 5808 7232
rect 5872 7168 5888 7232
rect 5952 7168 5968 7232
rect 6032 7168 6048 7232
rect 6112 7168 6128 7232
rect 6192 7168 6208 7232
rect 6272 7168 6288 7232
rect 6352 7168 6368 7232
rect 6432 7168 6448 7232
rect 6512 7168 6528 7232
rect 6592 7168 6608 7232
rect 6672 7168 6688 7232
rect 6752 7168 6768 7232
rect 6832 7168 6848 7232
rect 6912 7168 6928 7232
rect 6992 7168 7008 7232
rect 7072 7168 7088 7232
rect 7152 7168 7168 7232
rect 7232 7168 7248 7232
rect 7312 7168 7328 7232
rect 7392 7168 7408 7232
rect 7472 7168 7488 7232
rect 7552 7168 7568 7232
rect 7632 7168 7648 7232
rect 7712 7168 7728 7232
rect 7792 7168 7808 7232
rect 7872 7168 7888 7232
rect 7952 7168 7968 7232
rect 8032 7168 8048 7232
rect 8112 7168 8128 7232
rect 8192 7168 8208 7232
rect 8272 7168 8288 7232
rect 8352 7168 8368 7232
rect 8432 7168 8448 7232
rect 8512 7168 8528 7232
rect 8592 7168 8608 7232
rect 8672 7168 8688 7232
rect 8752 7168 8768 7232
rect 8832 7168 8848 7232
rect 8912 7168 8928 7232
rect 8992 7168 9000 7232
rect 5000 7152 9000 7168
rect 5000 7088 5008 7152
rect 5072 7088 5088 7152
rect 5152 7088 5168 7152
rect 5232 7088 5248 7152
rect 5312 7088 5328 7152
rect 5392 7088 5408 7152
rect 5472 7088 5488 7152
rect 5552 7088 5568 7152
rect 5632 7088 5648 7152
rect 5712 7088 5728 7152
rect 5792 7088 5808 7152
rect 5872 7088 5888 7152
rect 5952 7088 5968 7152
rect 6032 7088 6048 7152
rect 6112 7088 6128 7152
rect 6192 7088 6208 7152
rect 6272 7088 6288 7152
rect 6352 7088 6368 7152
rect 6432 7088 6448 7152
rect 6512 7088 6528 7152
rect 6592 7088 6608 7152
rect 6672 7088 6688 7152
rect 6752 7088 6768 7152
rect 6832 7088 6848 7152
rect 6912 7088 6928 7152
rect 6992 7088 7008 7152
rect 7072 7088 7088 7152
rect 7152 7088 7168 7152
rect 7232 7088 7248 7152
rect 7312 7088 7328 7152
rect 7392 7088 7408 7152
rect 7472 7088 7488 7152
rect 7552 7088 7568 7152
rect 7632 7088 7648 7152
rect 7712 7088 7728 7152
rect 7792 7088 7808 7152
rect 7872 7088 7888 7152
rect 7952 7088 7968 7152
rect 8032 7088 8048 7152
rect 8112 7088 8128 7152
rect 8192 7088 8208 7152
rect 8272 7088 8288 7152
rect 8352 7088 8368 7152
rect 8432 7088 8448 7152
rect 8512 7088 8528 7152
rect 8592 7088 8608 7152
rect 8672 7088 8688 7152
rect 8752 7088 8768 7152
rect 8832 7088 8848 7152
rect 8912 7088 8928 7152
rect 8992 7088 9000 7152
rect 5000 7072 9000 7088
rect 5000 7008 5008 7072
rect 5072 7008 5088 7072
rect 5152 7008 5168 7072
rect 5232 7008 5248 7072
rect 5312 7008 5328 7072
rect 5392 7008 5408 7072
rect 5472 7008 5488 7072
rect 5552 7008 5568 7072
rect 5632 7008 5648 7072
rect 5712 7008 5728 7072
rect 5792 7008 5808 7072
rect 5872 7008 5888 7072
rect 5952 7008 5968 7072
rect 6032 7008 6048 7072
rect 6112 7008 6128 7072
rect 6192 7008 6208 7072
rect 6272 7008 6288 7072
rect 6352 7008 6368 7072
rect 6432 7008 6448 7072
rect 6512 7008 6528 7072
rect 6592 7008 6608 7072
rect 6672 7008 6688 7072
rect 6752 7008 6768 7072
rect 6832 7008 6848 7072
rect 6912 7008 6928 7072
rect 6992 7008 7008 7072
rect 7072 7008 7088 7072
rect 7152 7008 7168 7072
rect 7232 7008 7248 7072
rect 7312 7008 7328 7072
rect 7392 7008 7408 7072
rect 7472 7008 7488 7072
rect 7552 7008 7568 7072
rect 7632 7008 7648 7072
rect 7712 7008 7728 7072
rect 7792 7008 7808 7072
rect 7872 7008 7888 7072
rect 7952 7008 7968 7072
rect 8032 7008 8048 7072
rect 8112 7008 8128 7072
rect 8192 7008 8208 7072
rect 8272 7008 8288 7072
rect 8352 7008 8368 7072
rect 8432 7008 8448 7072
rect 8512 7008 8528 7072
rect 8592 7008 8608 7072
rect 8672 7008 8688 7072
rect 8752 7008 8768 7072
rect 8832 7008 8848 7072
rect 8912 7008 8928 7072
rect 8992 7008 9000 7072
rect 5000 6992 9000 7008
rect 5000 6928 5008 6992
rect 5072 6928 5088 6992
rect 5152 6928 5168 6992
rect 5232 6928 5248 6992
rect 5312 6928 5328 6992
rect 5392 6928 5408 6992
rect 5472 6928 5488 6992
rect 5552 6928 5568 6992
rect 5632 6928 5648 6992
rect 5712 6928 5728 6992
rect 5792 6928 5808 6992
rect 5872 6928 5888 6992
rect 5952 6928 5968 6992
rect 6032 6928 6048 6992
rect 6112 6928 6128 6992
rect 6192 6928 6208 6992
rect 6272 6928 6288 6992
rect 6352 6928 6368 6992
rect 6432 6928 6448 6992
rect 6512 6928 6528 6992
rect 6592 6928 6608 6992
rect 6672 6928 6688 6992
rect 6752 6928 6768 6992
rect 6832 6928 6848 6992
rect 6912 6928 6928 6992
rect 6992 6928 7008 6992
rect 7072 6928 7088 6992
rect 7152 6928 7168 6992
rect 7232 6928 7248 6992
rect 7312 6928 7328 6992
rect 7392 6928 7408 6992
rect 7472 6928 7488 6992
rect 7552 6928 7568 6992
rect 7632 6928 7648 6992
rect 7712 6928 7728 6992
rect 7792 6928 7808 6992
rect 7872 6928 7888 6992
rect 7952 6928 7968 6992
rect 8032 6928 8048 6992
rect 8112 6928 8128 6992
rect 8192 6928 8208 6992
rect 8272 6928 8288 6992
rect 8352 6928 8368 6992
rect 8432 6928 8448 6992
rect 8512 6928 8528 6992
rect 8592 6928 8608 6992
rect 8672 6928 8688 6992
rect 8752 6928 8768 6992
rect 8832 6928 8848 6992
rect 8912 6928 8928 6992
rect 8992 6928 9000 6992
rect 5000 6912 9000 6928
rect 5000 6848 5008 6912
rect 5072 6848 5088 6912
rect 5152 6848 5168 6912
rect 5232 6848 5248 6912
rect 5312 6848 5328 6912
rect 5392 6848 5408 6912
rect 5472 6848 5488 6912
rect 5552 6848 5568 6912
rect 5632 6848 5648 6912
rect 5712 6848 5728 6912
rect 5792 6848 5808 6912
rect 5872 6848 5888 6912
rect 5952 6848 5968 6912
rect 6032 6848 6048 6912
rect 6112 6848 6128 6912
rect 6192 6848 6208 6912
rect 6272 6848 6288 6912
rect 6352 6848 6368 6912
rect 6432 6848 6448 6912
rect 6512 6848 6528 6912
rect 6592 6848 6608 6912
rect 6672 6848 6688 6912
rect 6752 6848 6768 6912
rect 6832 6848 6848 6912
rect 6912 6848 6928 6912
rect 6992 6848 7008 6912
rect 7072 6848 7088 6912
rect 7152 6848 7168 6912
rect 7232 6848 7248 6912
rect 7312 6848 7328 6912
rect 7392 6848 7408 6912
rect 7472 6848 7488 6912
rect 7552 6848 7568 6912
rect 7632 6848 7648 6912
rect 7712 6848 7728 6912
rect 7792 6848 7808 6912
rect 7872 6848 7888 6912
rect 7952 6848 7968 6912
rect 8032 6848 8048 6912
rect 8112 6848 8128 6912
rect 8192 6848 8208 6912
rect 8272 6848 8288 6912
rect 8352 6848 8368 6912
rect 8432 6848 8448 6912
rect 8512 6848 8528 6912
rect 8592 6848 8608 6912
rect 8672 6848 8688 6912
rect 8752 6848 8768 6912
rect 8832 6848 8848 6912
rect 8912 6848 8928 6912
rect 8992 6848 9000 6912
rect 5000 6832 9000 6848
rect 5000 6768 5008 6832
rect 5072 6768 5088 6832
rect 5152 6768 5168 6832
rect 5232 6768 5248 6832
rect 5312 6768 5328 6832
rect 5392 6768 5408 6832
rect 5472 6768 5488 6832
rect 5552 6768 5568 6832
rect 5632 6768 5648 6832
rect 5712 6768 5728 6832
rect 5792 6768 5808 6832
rect 5872 6768 5888 6832
rect 5952 6768 5968 6832
rect 6032 6768 6048 6832
rect 6112 6768 6128 6832
rect 6192 6768 6208 6832
rect 6272 6768 6288 6832
rect 6352 6768 6368 6832
rect 6432 6768 6448 6832
rect 6512 6768 6528 6832
rect 6592 6768 6608 6832
rect 6672 6768 6688 6832
rect 6752 6768 6768 6832
rect 6832 6768 6848 6832
rect 6912 6768 6928 6832
rect 6992 6768 7008 6832
rect 7072 6768 7088 6832
rect 7152 6768 7168 6832
rect 7232 6768 7248 6832
rect 7312 6768 7328 6832
rect 7392 6768 7408 6832
rect 7472 6768 7488 6832
rect 7552 6768 7568 6832
rect 7632 6768 7648 6832
rect 7712 6768 7728 6832
rect 7792 6768 7808 6832
rect 7872 6768 7888 6832
rect 7952 6768 7968 6832
rect 8032 6768 8048 6832
rect 8112 6768 8128 6832
rect 8192 6768 8208 6832
rect 8272 6768 8288 6832
rect 8352 6768 8368 6832
rect 8432 6768 8448 6832
rect 8512 6768 8528 6832
rect 8592 6768 8608 6832
rect 8672 6768 8688 6832
rect 8752 6768 8768 6832
rect 8832 6768 8848 6832
rect 8912 6768 8928 6832
rect 8992 6768 9000 6832
rect 5000 6752 9000 6768
rect 5000 6688 5008 6752
rect 5072 6688 5088 6752
rect 5152 6688 5168 6752
rect 5232 6688 5248 6752
rect 5312 6688 5328 6752
rect 5392 6688 5408 6752
rect 5472 6688 5488 6752
rect 5552 6688 5568 6752
rect 5632 6688 5648 6752
rect 5712 6688 5728 6752
rect 5792 6688 5808 6752
rect 5872 6688 5888 6752
rect 5952 6688 5968 6752
rect 6032 6688 6048 6752
rect 6112 6688 6128 6752
rect 6192 6688 6208 6752
rect 6272 6688 6288 6752
rect 6352 6688 6368 6752
rect 6432 6688 6448 6752
rect 6512 6688 6528 6752
rect 6592 6688 6608 6752
rect 6672 6688 6688 6752
rect 6752 6688 6768 6752
rect 6832 6688 6848 6752
rect 6912 6688 6928 6752
rect 6992 6688 7008 6752
rect 7072 6688 7088 6752
rect 7152 6688 7168 6752
rect 7232 6688 7248 6752
rect 7312 6688 7328 6752
rect 7392 6688 7408 6752
rect 7472 6688 7488 6752
rect 7552 6688 7568 6752
rect 7632 6688 7648 6752
rect 7712 6688 7728 6752
rect 7792 6688 7808 6752
rect 7872 6688 7888 6752
rect 7952 6688 7968 6752
rect 8032 6688 8048 6752
rect 8112 6688 8128 6752
rect 8192 6688 8208 6752
rect 8272 6688 8288 6752
rect 8352 6688 8368 6752
rect 8432 6688 8448 6752
rect 8512 6688 8528 6752
rect 8592 6688 8608 6752
rect 8672 6688 8688 6752
rect 8752 6688 8768 6752
rect 8832 6688 8848 6752
rect 8912 6688 8928 6752
rect 8992 6688 9000 6752
rect 5000 6672 9000 6688
rect 5000 6608 5008 6672
rect 5072 6608 5088 6672
rect 5152 6608 5168 6672
rect 5232 6608 5248 6672
rect 5312 6608 5328 6672
rect 5392 6608 5408 6672
rect 5472 6608 5488 6672
rect 5552 6608 5568 6672
rect 5632 6608 5648 6672
rect 5712 6608 5728 6672
rect 5792 6608 5808 6672
rect 5872 6608 5888 6672
rect 5952 6608 5968 6672
rect 6032 6608 6048 6672
rect 6112 6608 6128 6672
rect 6192 6608 6208 6672
rect 6272 6608 6288 6672
rect 6352 6608 6368 6672
rect 6432 6608 6448 6672
rect 6512 6608 6528 6672
rect 6592 6608 6608 6672
rect 6672 6608 6688 6672
rect 6752 6608 6768 6672
rect 6832 6608 6848 6672
rect 6912 6608 6928 6672
rect 6992 6608 7008 6672
rect 7072 6608 7088 6672
rect 7152 6608 7168 6672
rect 7232 6608 7248 6672
rect 7312 6608 7328 6672
rect 7392 6608 7408 6672
rect 7472 6608 7488 6672
rect 7552 6608 7568 6672
rect 7632 6608 7648 6672
rect 7712 6608 7728 6672
rect 7792 6608 7808 6672
rect 7872 6608 7888 6672
rect 7952 6608 7968 6672
rect 8032 6608 8048 6672
rect 8112 6608 8128 6672
rect 8192 6608 8208 6672
rect 8272 6608 8288 6672
rect 8352 6608 8368 6672
rect 8432 6608 8448 6672
rect 8512 6608 8528 6672
rect 8592 6608 8608 6672
rect 8672 6608 8688 6672
rect 8752 6608 8768 6672
rect 8832 6608 8848 6672
rect 8912 6608 8928 6672
rect 8992 6608 9000 6672
rect 5000 6592 9000 6608
rect 5000 6528 5008 6592
rect 5072 6528 5088 6592
rect 5152 6528 5168 6592
rect 5232 6528 5248 6592
rect 5312 6528 5328 6592
rect 5392 6528 5408 6592
rect 5472 6528 5488 6592
rect 5552 6528 5568 6592
rect 5632 6528 5648 6592
rect 5712 6528 5728 6592
rect 5792 6528 5808 6592
rect 5872 6528 5888 6592
rect 5952 6528 5968 6592
rect 6032 6528 6048 6592
rect 6112 6528 6128 6592
rect 6192 6528 6208 6592
rect 6272 6528 6288 6592
rect 6352 6528 6368 6592
rect 6432 6528 6448 6592
rect 6512 6528 6528 6592
rect 6592 6528 6608 6592
rect 6672 6528 6688 6592
rect 6752 6528 6768 6592
rect 6832 6528 6848 6592
rect 6912 6528 6928 6592
rect 6992 6528 7008 6592
rect 7072 6528 7088 6592
rect 7152 6528 7168 6592
rect 7232 6528 7248 6592
rect 7312 6528 7328 6592
rect 7392 6528 7408 6592
rect 7472 6528 7488 6592
rect 7552 6528 7568 6592
rect 7632 6528 7648 6592
rect 7712 6528 7728 6592
rect 7792 6528 7808 6592
rect 7872 6528 7888 6592
rect 7952 6528 7968 6592
rect 8032 6528 8048 6592
rect 8112 6528 8128 6592
rect 8192 6528 8208 6592
rect 8272 6528 8288 6592
rect 8352 6528 8368 6592
rect 8432 6528 8448 6592
rect 8512 6528 8528 6592
rect 8592 6528 8608 6592
rect 8672 6528 8688 6592
rect 8752 6528 8768 6592
rect 8832 6528 8848 6592
rect 8912 6528 8928 6592
rect 8992 6528 9000 6592
rect 5000 6512 9000 6528
rect 5000 6448 5008 6512
rect 5072 6448 5088 6512
rect 5152 6448 5168 6512
rect 5232 6448 5248 6512
rect 5312 6448 5328 6512
rect 5392 6448 5408 6512
rect 5472 6448 5488 6512
rect 5552 6448 5568 6512
rect 5632 6448 5648 6512
rect 5712 6448 5728 6512
rect 5792 6448 5808 6512
rect 5872 6448 5888 6512
rect 5952 6448 5968 6512
rect 6032 6448 6048 6512
rect 6112 6448 6128 6512
rect 6192 6448 6208 6512
rect 6272 6448 6288 6512
rect 6352 6448 6368 6512
rect 6432 6448 6448 6512
rect 6512 6448 6528 6512
rect 6592 6448 6608 6512
rect 6672 6448 6688 6512
rect 6752 6448 6768 6512
rect 6832 6448 6848 6512
rect 6912 6448 6928 6512
rect 6992 6448 7008 6512
rect 7072 6448 7088 6512
rect 7152 6448 7168 6512
rect 7232 6448 7248 6512
rect 7312 6448 7328 6512
rect 7392 6448 7408 6512
rect 7472 6448 7488 6512
rect 7552 6448 7568 6512
rect 7632 6448 7648 6512
rect 7712 6448 7728 6512
rect 7792 6448 7808 6512
rect 7872 6448 7888 6512
rect 7952 6448 7968 6512
rect 8032 6448 8048 6512
rect 8112 6448 8128 6512
rect 8192 6448 8208 6512
rect 8272 6448 8288 6512
rect 8352 6448 8368 6512
rect 8432 6448 8448 6512
rect 8512 6448 8528 6512
rect 8592 6448 8608 6512
rect 8672 6448 8688 6512
rect 8752 6448 8768 6512
rect 8832 6448 8848 6512
rect 8912 6448 8928 6512
rect 8992 6448 9000 6512
rect 5000 6432 9000 6448
rect 5000 6368 5008 6432
rect 5072 6368 5088 6432
rect 5152 6368 5168 6432
rect 5232 6368 5248 6432
rect 5312 6368 5328 6432
rect 5392 6368 5408 6432
rect 5472 6368 5488 6432
rect 5552 6368 5568 6432
rect 5632 6368 5648 6432
rect 5712 6368 5728 6432
rect 5792 6368 5808 6432
rect 5872 6368 5888 6432
rect 5952 6368 5968 6432
rect 6032 6368 6048 6432
rect 6112 6368 6128 6432
rect 6192 6368 6208 6432
rect 6272 6368 6288 6432
rect 6352 6368 6368 6432
rect 6432 6368 6448 6432
rect 6512 6368 6528 6432
rect 6592 6368 6608 6432
rect 6672 6368 6688 6432
rect 6752 6368 6768 6432
rect 6832 6368 6848 6432
rect 6912 6368 6928 6432
rect 6992 6368 7008 6432
rect 7072 6368 7088 6432
rect 7152 6368 7168 6432
rect 7232 6368 7248 6432
rect 7312 6368 7328 6432
rect 7392 6368 7408 6432
rect 7472 6368 7488 6432
rect 7552 6368 7568 6432
rect 7632 6368 7648 6432
rect 7712 6368 7728 6432
rect 7792 6368 7808 6432
rect 7872 6368 7888 6432
rect 7952 6368 7968 6432
rect 8032 6368 8048 6432
rect 8112 6368 8128 6432
rect 8192 6368 8208 6432
rect 8272 6368 8288 6432
rect 8352 6368 8368 6432
rect 8432 6368 8448 6432
rect 8512 6368 8528 6432
rect 8592 6368 8608 6432
rect 8672 6368 8688 6432
rect 8752 6368 8768 6432
rect 8832 6368 8848 6432
rect 8912 6368 8928 6432
rect 8992 6368 9000 6432
rect 5000 6352 9000 6368
rect 5000 6288 5008 6352
rect 5072 6288 5088 6352
rect 5152 6288 5168 6352
rect 5232 6288 5248 6352
rect 5312 6288 5328 6352
rect 5392 6288 5408 6352
rect 5472 6288 5488 6352
rect 5552 6288 5568 6352
rect 5632 6288 5648 6352
rect 5712 6288 5728 6352
rect 5792 6288 5808 6352
rect 5872 6288 5888 6352
rect 5952 6288 5968 6352
rect 6032 6288 6048 6352
rect 6112 6288 6128 6352
rect 6192 6288 6208 6352
rect 6272 6288 6288 6352
rect 6352 6288 6368 6352
rect 6432 6288 6448 6352
rect 6512 6288 6528 6352
rect 6592 6288 6608 6352
rect 6672 6288 6688 6352
rect 6752 6288 6768 6352
rect 6832 6288 6848 6352
rect 6912 6288 6928 6352
rect 6992 6288 7008 6352
rect 7072 6288 7088 6352
rect 7152 6288 7168 6352
rect 7232 6288 7248 6352
rect 7312 6288 7328 6352
rect 7392 6288 7408 6352
rect 7472 6288 7488 6352
rect 7552 6288 7568 6352
rect 7632 6288 7648 6352
rect 7712 6288 7728 6352
rect 7792 6288 7808 6352
rect 7872 6288 7888 6352
rect 7952 6288 7968 6352
rect 8032 6288 8048 6352
rect 8112 6288 8128 6352
rect 8192 6288 8208 6352
rect 8272 6288 8288 6352
rect 8352 6288 8368 6352
rect 8432 6288 8448 6352
rect 8512 6288 8528 6352
rect 8592 6288 8608 6352
rect 8672 6288 8688 6352
rect 8752 6288 8768 6352
rect 8832 6288 8848 6352
rect 8912 6288 8928 6352
rect 8992 6288 9000 6352
rect 5000 6272 9000 6288
rect 5000 6208 5008 6272
rect 5072 6208 5088 6272
rect 5152 6208 5168 6272
rect 5232 6208 5248 6272
rect 5312 6208 5328 6272
rect 5392 6208 5408 6272
rect 5472 6208 5488 6272
rect 5552 6208 5568 6272
rect 5632 6208 5648 6272
rect 5712 6208 5728 6272
rect 5792 6208 5808 6272
rect 5872 6208 5888 6272
rect 5952 6208 5968 6272
rect 6032 6208 6048 6272
rect 6112 6208 6128 6272
rect 6192 6208 6208 6272
rect 6272 6208 6288 6272
rect 6352 6208 6368 6272
rect 6432 6208 6448 6272
rect 6512 6208 6528 6272
rect 6592 6208 6608 6272
rect 6672 6208 6688 6272
rect 6752 6208 6768 6272
rect 6832 6208 6848 6272
rect 6912 6208 6928 6272
rect 6992 6208 7008 6272
rect 7072 6208 7088 6272
rect 7152 6208 7168 6272
rect 7232 6208 7248 6272
rect 7312 6208 7328 6272
rect 7392 6208 7408 6272
rect 7472 6208 7488 6272
rect 7552 6208 7568 6272
rect 7632 6208 7648 6272
rect 7712 6208 7728 6272
rect 7792 6208 7808 6272
rect 7872 6208 7888 6272
rect 7952 6208 7968 6272
rect 8032 6208 8048 6272
rect 8112 6208 8128 6272
rect 8192 6208 8208 6272
rect 8272 6208 8288 6272
rect 8352 6208 8368 6272
rect 8432 6208 8448 6272
rect 8512 6208 8528 6272
rect 8592 6208 8608 6272
rect 8672 6208 8688 6272
rect 8752 6208 8768 6272
rect 8832 6208 8848 6272
rect 8912 6208 8928 6272
rect 8992 6208 9000 6272
rect 5000 6192 9000 6208
rect 5000 6128 5008 6192
rect 5072 6128 5088 6192
rect 5152 6128 5168 6192
rect 5232 6128 5248 6192
rect 5312 6128 5328 6192
rect 5392 6128 5408 6192
rect 5472 6128 5488 6192
rect 5552 6128 5568 6192
rect 5632 6128 5648 6192
rect 5712 6128 5728 6192
rect 5792 6128 5808 6192
rect 5872 6128 5888 6192
rect 5952 6128 5968 6192
rect 6032 6128 6048 6192
rect 6112 6128 6128 6192
rect 6192 6128 6208 6192
rect 6272 6128 6288 6192
rect 6352 6128 6368 6192
rect 6432 6128 6448 6192
rect 6512 6128 6528 6192
rect 6592 6128 6608 6192
rect 6672 6128 6688 6192
rect 6752 6128 6768 6192
rect 6832 6128 6848 6192
rect 6912 6128 6928 6192
rect 6992 6128 7008 6192
rect 7072 6128 7088 6192
rect 7152 6128 7168 6192
rect 7232 6128 7248 6192
rect 7312 6128 7328 6192
rect 7392 6128 7408 6192
rect 7472 6128 7488 6192
rect 7552 6128 7568 6192
rect 7632 6128 7648 6192
rect 7712 6128 7728 6192
rect 7792 6128 7808 6192
rect 7872 6128 7888 6192
rect 7952 6128 7968 6192
rect 8032 6128 8048 6192
rect 8112 6128 8128 6192
rect 8192 6128 8208 6192
rect 8272 6128 8288 6192
rect 8352 6128 8368 6192
rect 8432 6128 8448 6192
rect 8512 6128 8528 6192
rect 8592 6128 8608 6192
rect 8672 6128 8688 6192
rect 8752 6128 8768 6192
rect 8832 6128 8848 6192
rect 8912 6128 8928 6192
rect 8992 6128 9000 6192
rect 5000 6112 9000 6128
rect 5000 6048 5008 6112
rect 5072 6048 5088 6112
rect 5152 6048 5168 6112
rect 5232 6048 5248 6112
rect 5312 6048 5328 6112
rect 5392 6048 5408 6112
rect 5472 6048 5488 6112
rect 5552 6048 5568 6112
rect 5632 6048 5648 6112
rect 5712 6048 5728 6112
rect 5792 6048 5808 6112
rect 5872 6048 5888 6112
rect 5952 6048 5968 6112
rect 6032 6048 6048 6112
rect 6112 6048 6128 6112
rect 6192 6048 6208 6112
rect 6272 6048 6288 6112
rect 6352 6048 6368 6112
rect 6432 6048 6448 6112
rect 6512 6048 6528 6112
rect 6592 6048 6608 6112
rect 6672 6048 6688 6112
rect 6752 6048 6768 6112
rect 6832 6048 6848 6112
rect 6912 6048 6928 6112
rect 6992 6048 7008 6112
rect 7072 6048 7088 6112
rect 7152 6048 7168 6112
rect 7232 6048 7248 6112
rect 7312 6048 7328 6112
rect 7392 6048 7408 6112
rect 7472 6048 7488 6112
rect 7552 6048 7568 6112
rect 7632 6048 7648 6112
rect 7712 6048 7728 6112
rect 7792 6048 7808 6112
rect 7872 6048 7888 6112
rect 7952 6048 7968 6112
rect 8032 6048 8048 6112
rect 8112 6048 8128 6112
rect 8192 6048 8208 6112
rect 8272 6048 8288 6112
rect 8352 6048 8368 6112
rect 8432 6048 8448 6112
rect 8512 6048 8528 6112
rect 8592 6048 8608 6112
rect 8672 6048 8688 6112
rect 8752 6048 8768 6112
rect 8832 6048 8848 6112
rect 8912 6048 8928 6112
rect 8992 6048 9000 6112
rect 5000 6032 9000 6048
rect 5000 5968 5008 6032
rect 5072 5968 5088 6032
rect 5152 5968 5168 6032
rect 5232 5968 5248 6032
rect 5312 5968 5328 6032
rect 5392 5968 5408 6032
rect 5472 5968 5488 6032
rect 5552 5968 5568 6032
rect 5632 5968 5648 6032
rect 5712 5968 5728 6032
rect 5792 5968 5808 6032
rect 5872 5968 5888 6032
rect 5952 5968 5968 6032
rect 6032 5968 6048 6032
rect 6112 5968 6128 6032
rect 6192 5968 6208 6032
rect 6272 5968 6288 6032
rect 6352 5968 6368 6032
rect 6432 5968 6448 6032
rect 6512 5968 6528 6032
rect 6592 5968 6608 6032
rect 6672 5968 6688 6032
rect 6752 5968 6768 6032
rect 6832 5968 6848 6032
rect 6912 5968 6928 6032
rect 6992 5968 7008 6032
rect 7072 5968 7088 6032
rect 7152 5968 7168 6032
rect 7232 5968 7248 6032
rect 7312 5968 7328 6032
rect 7392 5968 7408 6032
rect 7472 5968 7488 6032
rect 7552 5968 7568 6032
rect 7632 5968 7648 6032
rect 7712 5968 7728 6032
rect 7792 5968 7808 6032
rect 7872 5968 7888 6032
rect 7952 5968 7968 6032
rect 8032 5968 8048 6032
rect 8112 5968 8128 6032
rect 8192 5968 8208 6032
rect 8272 5968 8288 6032
rect 8352 5968 8368 6032
rect 8432 5968 8448 6032
rect 8512 5968 8528 6032
rect 8592 5968 8608 6032
rect 8672 5968 8688 6032
rect 8752 5968 8768 6032
rect 8832 5968 8848 6032
rect 8912 5968 8928 6032
rect 8992 5968 9000 6032
rect 5000 5952 9000 5968
rect 5000 5888 5008 5952
rect 5072 5888 5088 5952
rect 5152 5888 5168 5952
rect 5232 5888 5248 5952
rect 5312 5888 5328 5952
rect 5392 5888 5408 5952
rect 5472 5888 5488 5952
rect 5552 5888 5568 5952
rect 5632 5888 5648 5952
rect 5712 5888 5728 5952
rect 5792 5888 5808 5952
rect 5872 5888 5888 5952
rect 5952 5888 5968 5952
rect 6032 5888 6048 5952
rect 6112 5888 6128 5952
rect 6192 5888 6208 5952
rect 6272 5888 6288 5952
rect 6352 5888 6368 5952
rect 6432 5888 6448 5952
rect 6512 5888 6528 5952
rect 6592 5888 6608 5952
rect 6672 5888 6688 5952
rect 6752 5888 6768 5952
rect 6832 5888 6848 5952
rect 6912 5888 6928 5952
rect 6992 5888 7008 5952
rect 7072 5888 7088 5952
rect 7152 5888 7168 5952
rect 7232 5888 7248 5952
rect 7312 5888 7328 5952
rect 7392 5888 7408 5952
rect 7472 5888 7488 5952
rect 7552 5888 7568 5952
rect 7632 5888 7648 5952
rect 7712 5888 7728 5952
rect 7792 5888 7808 5952
rect 7872 5888 7888 5952
rect 7952 5888 7968 5952
rect 8032 5888 8048 5952
rect 8112 5888 8128 5952
rect 8192 5888 8208 5952
rect 8272 5888 8288 5952
rect 8352 5888 8368 5952
rect 8432 5888 8448 5952
rect 8512 5888 8528 5952
rect 8592 5888 8608 5952
rect 8672 5888 8688 5952
rect 8752 5888 8768 5952
rect 8832 5888 8848 5952
rect 8912 5888 8928 5952
rect 8992 5888 9000 5952
rect 5000 5872 9000 5888
rect 5000 5808 5008 5872
rect 5072 5808 5088 5872
rect 5152 5808 5168 5872
rect 5232 5808 5248 5872
rect 5312 5808 5328 5872
rect 5392 5808 5408 5872
rect 5472 5808 5488 5872
rect 5552 5808 5568 5872
rect 5632 5808 5648 5872
rect 5712 5808 5728 5872
rect 5792 5808 5808 5872
rect 5872 5808 5888 5872
rect 5952 5808 5968 5872
rect 6032 5808 6048 5872
rect 6112 5808 6128 5872
rect 6192 5808 6208 5872
rect 6272 5808 6288 5872
rect 6352 5808 6368 5872
rect 6432 5808 6448 5872
rect 6512 5808 6528 5872
rect 6592 5808 6608 5872
rect 6672 5808 6688 5872
rect 6752 5808 6768 5872
rect 6832 5808 6848 5872
rect 6912 5808 6928 5872
rect 6992 5808 7008 5872
rect 7072 5808 7088 5872
rect 7152 5808 7168 5872
rect 7232 5808 7248 5872
rect 7312 5808 7328 5872
rect 7392 5808 7408 5872
rect 7472 5808 7488 5872
rect 7552 5808 7568 5872
rect 7632 5808 7648 5872
rect 7712 5808 7728 5872
rect 7792 5808 7808 5872
rect 7872 5808 7888 5872
rect 7952 5808 7968 5872
rect 8032 5808 8048 5872
rect 8112 5808 8128 5872
rect 8192 5808 8208 5872
rect 8272 5808 8288 5872
rect 8352 5808 8368 5872
rect 8432 5808 8448 5872
rect 8512 5808 8528 5872
rect 8592 5808 8608 5872
rect 8672 5808 8688 5872
rect 8752 5808 8768 5872
rect 8832 5808 8848 5872
rect 8912 5808 8928 5872
rect 8992 5808 9000 5872
rect 5000 5792 9000 5808
rect 5000 5728 5008 5792
rect 5072 5728 5088 5792
rect 5152 5728 5168 5792
rect 5232 5728 5248 5792
rect 5312 5728 5328 5792
rect 5392 5728 5408 5792
rect 5472 5728 5488 5792
rect 5552 5728 5568 5792
rect 5632 5728 5648 5792
rect 5712 5728 5728 5792
rect 5792 5728 5808 5792
rect 5872 5728 5888 5792
rect 5952 5728 5968 5792
rect 6032 5728 6048 5792
rect 6112 5728 6128 5792
rect 6192 5728 6208 5792
rect 6272 5728 6288 5792
rect 6352 5728 6368 5792
rect 6432 5728 6448 5792
rect 6512 5728 6528 5792
rect 6592 5728 6608 5792
rect 6672 5728 6688 5792
rect 6752 5728 6768 5792
rect 6832 5728 6848 5792
rect 6912 5728 6928 5792
rect 6992 5728 7008 5792
rect 7072 5728 7088 5792
rect 7152 5728 7168 5792
rect 7232 5728 7248 5792
rect 7312 5728 7328 5792
rect 7392 5728 7408 5792
rect 7472 5728 7488 5792
rect 7552 5728 7568 5792
rect 7632 5728 7648 5792
rect 7712 5728 7728 5792
rect 7792 5728 7808 5792
rect 7872 5728 7888 5792
rect 7952 5728 7968 5792
rect 8032 5728 8048 5792
rect 8112 5728 8128 5792
rect 8192 5728 8208 5792
rect 8272 5728 8288 5792
rect 8352 5728 8368 5792
rect 8432 5728 8448 5792
rect 8512 5728 8528 5792
rect 8592 5728 8608 5792
rect 8672 5728 8688 5792
rect 8752 5728 8768 5792
rect 8832 5728 8848 5792
rect 8912 5728 8928 5792
rect 8992 5728 9000 5792
rect 5000 5712 9000 5728
rect 5000 5648 5008 5712
rect 5072 5648 5088 5712
rect 5152 5648 5168 5712
rect 5232 5648 5248 5712
rect 5312 5648 5328 5712
rect 5392 5648 5408 5712
rect 5472 5648 5488 5712
rect 5552 5648 5568 5712
rect 5632 5648 5648 5712
rect 5712 5648 5728 5712
rect 5792 5648 5808 5712
rect 5872 5648 5888 5712
rect 5952 5648 5968 5712
rect 6032 5648 6048 5712
rect 6112 5648 6128 5712
rect 6192 5648 6208 5712
rect 6272 5648 6288 5712
rect 6352 5648 6368 5712
rect 6432 5648 6448 5712
rect 6512 5648 6528 5712
rect 6592 5648 6608 5712
rect 6672 5648 6688 5712
rect 6752 5648 6768 5712
rect 6832 5648 6848 5712
rect 6912 5648 6928 5712
rect 6992 5648 7008 5712
rect 7072 5648 7088 5712
rect 7152 5648 7168 5712
rect 7232 5648 7248 5712
rect 7312 5648 7328 5712
rect 7392 5648 7408 5712
rect 7472 5648 7488 5712
rect 7552 5648 7568 5712
rect 7632 5648 7648 5712
rect 7712 5648 7728 5712
rect 7792 5648 7808 5712
rect 7872 5648 7888 5712
rect 7952 5648 7968 5712
rect 8032 5648 8048 5712
rect 8112 5648 8128 5712
rect 8192 5648 8208 5712
rect 8272 5648 8288 5712
rect 8352 5648 8368 5712
rect 8432 5648 8448 5712
rect 8512 5648 8528 5712
rect 8592 5648 8608 5712
rect 8672 5648 8688 5712
rect 8752 5648 8768 5712
rect 8832 5648 8848 5712
rect 8912 5648 8928 5712
rect 8992 5648 9000 5712
rect 5000 5632 9000 5648
rect 5000 5568 5008 5632
rect 5072 5568 5088 5632
rect 5152 5568 5168 5632
rect 5232 5568 5248 5632
rect 5312 5568 5328 5632
rect 5392 5568 5408 5632
rect 5472 5568 5488 5632
rect 5552 5568 5568 5632
rect 5632 5568 5648 5632
rect 5712 5568 5728 5632
rect 5792 5568 5808 5632
rect 5872 5568 5888 5632
rect 5952 5568 5968 5632
rect 6032 5568 6048 5632
rect 6112 5568 6128 5632
rect 6192 5568 6208 5632
rect 6272 5568 6288 5632
rect 6352 5568 6368 5632
rect 6432 5568 6448 5632
rect 6512 5568 6528 5632
rect 6592 5568 6608 5632
rect 6672 5568 6688 5632
rect 6752 5568 6768 5632
rect 6832 5568 6848 5632
rect 6912 5568 6928 5632
rect 6992 5568 7008 5632
rect 7072 5568 7088 5632
rect 7152 5568 7168 5632
rect 7232 5568 7248 5632
rect 7312 5568 7328 5632
rect 7392 5568 7408 5632
rect 7472 5568 7488 5632
rect 7552 5568 7568 5632
rect 7632 5568 7648 5632
rect 7712 5568 7728 5632
rect 7792 5568 7808 5632
rect 7872 5568 7888 5632
rect 7952 5568 7968 5632
rect 8032 5568 8048 5632
rect 8112 5568 8128 5632
rect 8192 5568 8208 5632
rect 8272 5568 8288 5632
rect 8352 5568 8368 5632
rect 8432 5568 8448 5632
rect 8512 5568 8528 5632
rect 8592 5568 8608 5632
rect 8672 5568 8688 5632
rect 8752 5568 8768 5632
rect 8832 5568 8848 5632
rect 8912 5568 8928 5632
rect 8992 5568 9000 5632
rect 5000 5552 9000 5568
rect 5000 5488 5008 5552
rect 5072 5488 5088 5552
rect 5152 5488 5168 5552
rect 5232 5488 5248 5552
rect 5312 5488 5328 5552
rect 5392 5488 5408 5552
rect 5472 5488 5488 5552
rect 5552 5488 5568 5552
rect 5632 5488 5648 5552
rect 5712 5488 5728 5552
rect 5792 5488 5808 5552
rect 5872 5488 5888 5552
rect 5952 5488 5968 5552
rect 6032 5488 6048 5552
rect 6112 5488 6128 5552
rect 6192 5488 6208 5552
rect 6272 5488 6288 5552
rect 6352 5488 6368 5552
rect 6432 5488 6448 5552
rect 6512 5488 6528 5552
rect 6592 5488 6608 5552
rect 6672 5488 6688 5552
rect 6752 5488 6768 5552
rect 6832 5488 6848 5552
rect 6912 5488 6928 5552
rect 6992 5488 7008 5552
rect 7072 5488 7088 5552
rect 7152 5488 7168 5552
rect 7232 5488 7248 5552
rect 7312 5488 7328 5552
rect 7392 5488 7408 5552
rect 7472 5488 7488 5552
rect 7552 5488 7568 5552
rect 7632 5488 7648 5552
rect 7712 5488 7728 5552
rect 7792 5488 7808 5552
rect 7872 5488 7888 5552
rect 7952 5488 7968 5552
rect 8032 5488 8048 5552
rect 8112 5488 8128 5552
rect 8192 5488 8208 5552
rect 8272 5488 8288 5552
rect 8352 5488 8368 5552
rect 8432 5488 8448 5552
rect 8512 5488 8528 5552
rect 8592 5488 8608 5552
rect 8672 5488 8688 5552
rect 8752 5488 8768 5552
rect 8832 5488 8848 5552
rect 8912 5488 8928 5552
rect 8992 5488 9000 5552
rect 5000 5472 9000 5488
rect 5000 5408 5008 5472
rect 5072 5408 5088 5472
rect 5152 5408 5168 5472
rect 5232 5408 5248 5472
rect 5312 5408 5328 5472
rect 5392 5408 5408 5472
rect 5472 5408 5488 5472
rect 5552 5408 5568 5472
rect 5632 5408 5648 5472
rect 5712 5408 5728 5472
rect 5792 5408 5808 5472
rect 5872 5408 5888 5472
rect 5952 5408 5968 5472
rect 6032 5408 6048 5472
rect 6112 5408 6128 5472
rect 6192 5408 6208 5472
rect 6272 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6608 5472
rect 6672 5408 6688 5472
rect 6752 5408 6768 5472
rect 6832 5408 6848 5472
rect 6912 5408 6928 5472
rect 6992 5408 7008 5472
rect 7072 5408 7088 5472
rect 7152 5408 7168 5472
rect 7232 5408 7248 5472
rect 7312 5408 7328 5472
rect 7392 5408 7408 5472
rect 7472 5408 7488 5472
rect 7552 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7888 5472
rect 7952 5408 7968 5472
rect 8032 5408 8048 5472
rect 8112 5408 8128 5472
rect 8192 5408 8208 5472
rect 8272 5408 8288 5472
rect 8352 5408 8368 5472
rect 8432 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8768 5472
rect 8832 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9000 5472
rect 5000 5392 9000 5408
rect 5000 5328 5008 5392
rect 5072 5328 5088 5392
rect 5152 5328 5168 5392
rect 5232 5328 5248 5392
rect 5312 5328 5328 5392
rect 5392 5328 5408 5392
rect 5472 5328 5488 5392
rect 5552 5328 5568 5392
rect 5632 5328 5648 5392
rect 5712 5328 5728 5392
rect 5792 5328 5808 5392
rect 5872 5328 5888 5392
rect 5952 5328 5968 5392
rect 6032 5328 6048 5392
rect 6112 5328 6128 5392
rect 6192 5328 6208 5392
rect 6272 5328 6288 5392
rect 6352 5328 6368 5392
rect 6432 5328 6448 5392
rect 6512 5328 6528 5392
rect 6592 5328 6608 5392
rect 6672 5328 6688 5392
rect 6752 5328 6768 5392
rect 6832 5328 6848 5392
rect 6912 5328 6928 5392
rect 6992 5328 7008 5392
rect 7072 5328 7088 5392
rect 7152 5328 7168 5392
rect 7232 5328 7248 5392
rect 7312 5328 7328 5392
rect 7392 5328 7408 5392
rect 7472 5328 7488 5392
rect 7552 5328 7568 5392
rect 7632 5328 7648 5392
rect 7712 5328 7728 5392
rect 7792 5328 7808 5392
rect 7872 5328 7888 5392
rect 7952 5328 7968 5392
rect 8032 5328 8048 5392
rect 8112 5328 8128 5392
rect 8192 5328 8208 5392
rect 8272 5328 8288 5392
rect 8352 5328 8368 5392
rect 8432 5328 8448 5392
rect 8512 5328 8528 5392
rect 8592 5328 8608 5392
rect 8672 5328 8688 5392
rect 8752 5328 8768 5392
rect 8832 5328 8848 5392
rect 8912 5328 8928 5392
rect 8992 5328 9000 5392
rect 5000 5312 9000 5328
rect 5000 5248 5008 5312
rect 5072 5248 5088 5312
rect 5152 5248 5168 5312
rect 5232 5248 5248 5312
rect 5312 5248 5328 5312
rect 5392 5248 5408 5312
rect 5472 5248 5488 5312
rect 5552 5248 5568 5312
rect 5632 5248 5648 5312
rect 5712 5248 5728 5312
rect 5792 5248 5808 5312
rect 5872 5248 5888 5312
rect 5952 5248 5968 5312
rect 6032 5248 6048 5312
rect 6112 5248 6128 5312
rect 6192 5248 6208 5312
rect 6272 5248 6288 5312
rect 6352 5248 6368 5312
rect 6432 5248 6448 5312
rect 6512 5248 6528 5312
rect 6592 5248 6608 5312
rect 6672 5248 6688 5312
rect 6752 5248 6768 5312
rect 6832 5248 6848 5312
rect 6912 5248 6928 5312
rect 6992 5248 7008 5312
rect 7072 5248 7088 5312
rect 7152 5248 7168 5312
rect 7232 5248 7248 5312
rect 7312 5248 7328 5312
rect 7392 5248 7408 5312
rect 7472 5248 7488 5312
rect 7552 5248 7568 5312
rect 7632 5248 7648 5312
rect 7712 5248 7728 5312
rect 7792 5248 7808 5312
rect 7872 5248 7888 5312
rect 7952 5248 7968 5312
rect 8032 5248 8048 5312
rect 8112 5248 8128 5312
rect 8192 5248 8208 5312
rect 8272 5248 8288 5312
rect 8352 5248 8368 5312
rect 8432 5248 8448 5312
rect 8512 5248 8528 5312
rect 8592 5248 8608 5312
rect 8672 5248 8688 5312
rect 8752 5248 8768 5312
rect 8832 5248 8848 5312
rect 8912 5248 8928 5312
rect 8992 5248 9000 5312
rect 5000 5232 9000 5248
rect 5000 5168 5008 5232
rect 5072 5168 5088 5232
rect 5152 5168 5168 5232
rect 5232 5168 5248 5232
rect 5312 5168 5328 5232
rect 5392 5168 5408 5232
rect 5472 5168 5488 5232
rect 5552 5168 5568 5232
rect 5632 5168 5648 5232
rect 5712 5168 5728 5232
rect 5792 5168 5808 5232
rect 5872 5168 5888 5232
rect 5952 5168 5968 5232
rect 6032 5168 6048 5232
rect 6112 5168 6128 5232
rect 6192 5168 6208 5232
rect 6272 5168 6288 5232
rect 6352 5168 6368 5232
rect 6432 5168 6448 5232
rect 6512 5168 6528 5232
rect 6592 5168 6608 5232
rect 6672 5168 6688 5232
rect 6752 5168 6768 5232
rect 6832 5168 6848 5232
rect 6912 5168 6928 5232
rect 6992 5168 7008 5232
rect 7072 5168 7088 5232
rect 7152 5168 7168 5232
rect 7232 5168 7248 5232
rect 7312 5168 7328 5232
rect 7392 5168 7408 5232
rect 7472 5168 7488 5232
rect 7552 5168 7568 5232
rect 7632 5168 7648 5232
rect 7712 5168 7728 5232
rect 7792 5168 7808 5232
rect 7872 5168 7888 5232
rect 7952 5168 7968 5232
rect 8032 5168 8048 5232
rect 8112 5168 8128 5232
rect 8192 5168 8208 5232
rect 8272 5168 8288 5232
rect 8352 5168 8368 5232
rect 8432 5168 8448 5232
rect 8512 5168 8528 5232
rect 8592 5168 8608 5232
rect 8672 5168 8688 5232
rect 8752 5168 8768 5232
rect 8832 5168 8848 5232
rect 8912 5168 8928 5232
rect 8992 5168 9000 5232
rect 5000 5152 9000 5168
rect 5000 5088 5008 5152
rect 5072 5088 5088 5152
rect 5152 5088 5168 5152
rect 5232 5088 5248 5152
rect 5312 5088 5328 5152
rect 5392 5088 5408 5152
rect 5472 5088 5488 5152
rect 5552 5088 5568 5152
rect 5632 5088 5648 5152
rect 5712 5088 5728 5152
rect 5792 5088 5808 5152
rect 5872 5088 5888 5152
rect 5952 5088 5968 5152
rect 6032 5088 6048 5152
rect 6112 5088 6128 5152
rect 6192 5088 6208 5152
rect 6272 5088 6288 5152
rect 6352 5088 6368 5152
rect 6432 5088 6448 5152
rect 6512 5088 6528 5152
rect 6592 5088 6608 5152
rect 6672 5088 6688 5152
rect 6752 5088 6768 5152
rect 6832 5088 6848 5152
rect 6912 5088 6928 5152
rect 6992 5088 7008 5152
rect 7072 5088 7088 5152
rect 7152 5088 7168 5152
rect 7232 5088 7248 5152
rect 7312 5088 7328 5152
rect 7392 5088 7408 5152
rect 7472 5088 7488 5152
rect 7552 5088 7568 5152
rect 7632 5088 7648 5152
rect 7712 5088 7728 5152
rect 7792 5088 7808 5152
rect 7872 5088 7888 5152
rect 7952 5088 7968 5152
rect 8032 5088 8048 5152
rect 8112 5088 8128 5152
rect 8192 5088 8208 5152
rect 8272 5088 8288 5152
rect 8352 5088 8368 5152
rect 8432 5088 8448 5152
rect 8512 5088 8528 5152
rect 8592 5088 8608 5152
rect 8672 5088 8688 5152
rect 8752 5088 8768 5152
rect 8832 5088 8848 5152
rect 8912 5088 8928 5152
rect 8992 5088 9000 5152
rect 5000 5072 9000 5088
rect 5000 5008 5008 5072
rect 5072 5008 5088 5072
rect 5152 5008 5168 5072
rect 5232 5008 5248 5072
rect 5312 5008 5328 5072
rect 5392 5008 5408 5072
rect 5472 5008 5488 5072
rect 5552 5008 5568 5072
rect 5632 5008 5648 5072
rect 5712 5008 5728 5072
rect 5792 5008 5808 5072
rect 5872 5008 5888 5072
rect 5952 5008 5968 5072
rect 6032 5008 6048 5072
rect 6112 5008 6128 5072
rect 6192 5008 6208 5072
rect 6272 5008 6288 5072
rect 6352 5008 6368 5072
rect 6432 5008 6448 5072
rect 6512 5008 6528 5072
rect 6592 5008 6608 5072
rect 6672 5008 6688 5072
rect 6752 5008 6768 5072
rect 6832 5008 6848 5072
rect 6912 5008 6928 5072
rect 6992 5008 7008 5072
rect 7072 5008 7088 5072
rect 7152 5008 7168 5072
rect 7232 5008 7248 5072
rect 7312 5008 7328 5072
rect 7392 5008 7408 5072
rect 7472 5008 7488 5072
rect 7552 5008 7568 5072
rect 7632 5008 7648 5072
rect 7712 5008 7728 5072
rect 7792 5008 7808 5072
rect 7872 5008 7888 5072
rect 7952 5008 7968 5072
rect 8032 5008 8048 5072
rect 8112 5008 8128 5072
rect 8192 5008 8208 5072
rect 8272 5008 8288 5072
rect 8352 5008 8368 5072
rect 8432 5008 8448 5072
rect 8512 5008 8528 5072
rect 8592 5008 8608 5072
rect 8672 5008 8688 5072
rect 8752 5008 8768 5072
rect 8832 5008 8848 5072
rect 8912 5008 8928 5072
rect 8992 5008 9000 5072
rect 5000 5000 9000 5008
rect 14104 40384 14424 45392
rect 14104 40320 14112 40384
rect 14176 40320 14192 40384
rect 14256 40320 14272 40384
rect 14336 40320 14352 40384
rect 14416 40320 14424 40384
rect 14104 40304 14424 40320
rect 14104 40240 14112 40304
rect 14176 40240 14192 40304
rect 14256 40240 14272 40304
rect 14336 40240 14352 40304
rect 14416 40240 14424 40304
rect 14104 40224 14424 40240
rect 14104 40160 14112 40224
rect 14176 40160 14192 40224
rect 14256 40160 14272 40224
rect 14336 40160 14352 40224
rect 14416 40160 14424 40224
rect 14104 40144 14424 40160
rect 14104 40080 14112 40144
rect 14176 40080 14192 40144
rect 14256 40080 14272 40144
rect 14336 40080 14352 40144
rect 14416 40080 14424 40144
rect 14104 40064 14424 40080
rect 14104 40000 14112 40064
rect 14176 40000 14192 40064
rect 14256 40000 14272 40064
rect 14336 40000 14352 40064
rect 14416 40000 14424 40064
rect 14104 39984 14424 40000
rect 14104 39920 14112 39984
rect 14176 39920 14192 39984
rect 14256 39920 14272 39984
rect 14336 39920 14352 39984
rect 14416 39920 14424 39984
rect 14104 39904 14424 39920
rect 14104 39840 14112 39904
rect 14176 39840 14192 39904
rect 14256 39840 14272 39904
rect 14336 39840 14352 39904
rect 14416 39840 14424 39904
rect 14104 39824 14424 39840
rect 14104 39760 14112 39824
rect 14176 39760 14192 39824
rect 14256 39760 14272 39824
rect 14336 39760 14352 39824
rect 14416 39760 14424 39824
rect 14104 39744 14424 39760
rect 14104 39680 14112 39744
rect 14176 39680 14192 39744
rect 14256 39680 14272 39744
rect 14336 39680 14352 39744
rect 14416 39680 14424 39744
rect 14104 39664 14424 39680
rect 14104 39600 14112 39664
rect 14176 39600 14192 39664
rect 14256 39600 14272 39664
rect 14336 39600 14352 39664
rect 14416 39600 14424 39664
rect 14104 39584 14424 39600
rect 14104 39520 14112 39584
rect 14176 39520 14192 39584
rect 14256 39520 14272 39584
rect 14336 39520 14352 39584
rect 14416 39520 14424 39584
rect 14104 39504 14424 39520
rect 14104 39440 14112 39504
rect 14176 39440 14192 39504
rect 14256 39440 14272 39504
rect 14336 39440 14352 39504
rect 14416 39440 14424 39504
rect 14104 39424 14424 39440
rect 14104 39360 14112 39424
rect 14176 39360 14192 39424
rect 14256 39360 14272 39424
rect 14336 39360 14352 39424
rect 14416 39360 14424 39424
rect 14104 39344 14424 39360
rect 14104 39280 14112 39344
rect 14176 39280 14192 39344
rect 14256 39280 14272 39344
rect 14336 39280 14352 39344
rect 14416 39280 14424 39344
rect 14104 39264 14424 39280
rect 14104 39200 14112 39264
rect 14176 39200 14192 39264
rect 14256 39200 14272 39264
rect 14336 39200 14352 39264
rect 14416 39200 14424 39264
rect 14104 39184 14424 39200
rect 14104 39120 14112 39184
rect 14176 39120 14192 39184
rect 14256 39120 14272 39184
rect 14336 39120 14352 39184
rect 14416 39120 14424 39184
rect 14104 39104 14424 39120
rect 14104 39040 14112 39104
rect 14176 39040 14192 39104
rect 14256 39040 14272 39104
rect 14336 39040 14352 39104
rect 14416 39040 14424 39104
rect 14104 39024 14424 39040
rect 14104 38960 14112 39024
rect 14176 38960 14192 39024
rect 14256 38960 14272 39024
rect 14336 38960 14352 39024
rect 14416 38960 14424 39024
rect 14104 38944 14424 38960
rect 14104 38880 14112 38944
rect 14176 38880 14192 38944
rect 14256 38880 14272 38944
rect 14336 38880 14352 38944
rect 14416 38880 14424 38944
rect 14104 38864 14424 38880
rect 14104 38800 14112 38864
rect 14176 38800 14192 38864
rect 14256 38800 14272 38864
rect 14336 38800 14352 38864
rect 14416 38800 14424 38864
rect 14104 38784 14424 38800
rect 14104 38720 14112 38784
rect 14176 38720 14192 38784
rect 14256 38720 14272 38784
rect 14336 38720 14352 38784
rect 14416 38720 14424 38784
rect 14104 38704 14424 38720
rect 14104 38640 14112 38704
rect 14176 38640 14192 38704
rect 14256 38640 14272 38704
rect 14336 38640 14352 38704
rect 14416 38640 14424 38704
rect 14104 38624 14424 38640
rect 14104 38560 14112 38624
rect 14176 38560 14192 38624
rect 14256 38560 14272 38624
rect 14336 38560 14352 38624
rect 14416 38560 14424 38624
rect 14104 38544 14424 38560
rect 14104 38480 14112 38544
rect 14176 38480 14192 38544
rect 14256 38480 14272 38544
rect 14336 38480 14352 38544
rect 14416 38480 14424 38544
rect 14104 38464 14424 38480
rect 14104 38400 14112 38464
rect 14176 38400 14192 38464
rect 14256 38400 14272 38464
rect 14336 38400 14352 38464
rect 14416 38400 14424 38464
rect 14104 38384 14424 38400
rect 14104 38320 14112 38384
rect 14176 38320 14192 38384
rect 14256 38320 14272 38384
rect 14336 38320 14352 38384
rect 14416 38320 14424 38384
rect 14104 38304 14424 38320
rect 14104 38240 14112 38304
rect 14176 38240 14192 38304
rect 14256 38240 14272 38304
rect 14336 38240 14352 38304
rect 14416 38240 14424 38304
rect 14104 38224 14424 38240
rect 14104 38160 14112 38224
rect 14176 38160 14192 38224
rect 14256 38160 14272 38224
rect 14336 38160 14352 38224
rect 14416 38160 14424 38224
rect 14104 38144 14424 38160
rect 14104 38080 14112 38144
rect 14176 38080 14192 38144
rect 14256 38080 14272 38144
rect 14336 38080 14352 38144
rect 14416 38080 14424 38144
rect 14104 38064 14424 38080
rect 14104 38000 14112 38064
rect 14176 38000 14192 38064
rect 14256 38000 14272 38064
rect 14336 38000 14352 38064
rect 14416 38000 14424 38064
rect 14104 37984 14424 38000
rect 14104 37920 14112 37984
rect 14176 37920 14192 37984
rect 14256 37920 14272 37984
rect 14336 37920 14352 37984
rect 14416 37920 14424 37984
rect 14104 37904 14424 37920
rect 14104 37840 14112 37904
rect 14176 37840 14192 37904
rect 14256 37840 14272 37904
rect 14336 37840 14352 37904
rect 14416 37840 14424 37904
rect 14104 37824 14424 37840
rect 14104 37760 14112 37824
rect 14176 37760 14192 37824
rect 14256 37760 14272 37824
rect 14336 37760 14352 37824
rect 14416 37760 14424 37824
rect 14104 37744 14424 37760
rect 14104 37680 14112 37744
rect 14176 37680 14192 37744
rect 14256 37680 14272 37744
rect 14336 37680 14352 37744
rect 14416 37680 14424 37744
rect 14104 37664 14424 37680
rect 14104 37600 14112 37664
rect 14176 37600 14192 37664
rect 14256 37600 14272 37664
rect 14336 37600 14352 37664
rect 14416 37600 14424 37664
rect 14104 37584 14424 37600
rect 14104 37520 14112 37584
rect 14176 37520 14192 37584
rect 14256 37520 14272 37584
rect 14336 37520 14352 37584
rect 14416 37520 14424 37584
rect 14104 37504 14424 37520
rect 14104 37440 14112 37504
rect 14176 37440 14192 37504
rect 14256 37440 14272 37504
rect 14336 37440 14352 37504
rect 14416 37440 14424 37504
rect 14104 37424 14424 37440
rect 14104 37360 14112 37424
rect 14176 37360 14192 37424
rect 14256 37360 14272 37424
rect 14336 37360 14352 37424
rect 14416 37360 14424 37424
rect 14104 37344 14424 37360
rect 14104 37280 14112 37344
rect 14176 37280 14192 37344
rect 14256 37280 14272 37344
rect 14336 37280 14352 37344
rect 14416 37280 14424 37344
rect 14104 37264 14424 37280
rect 14104 37200 14112 37264
rect 14176 37200 14192 37264
rect 14256 37200 14272 37264
rect 14336 37200 14352 37264
rect 14416 37200 14424 37264
rect 14104 37184 14424 37200
rect 14104 37120 14112 37184
rect 14176 37120 14192 37184
rect 14256 37120 14272 37184
rect 14336 37120 14352 37184
rect 14416 37120 14424 37184
rect 14104 37104 14424 37120
rect 14104 37040 14112 37104
rect 14176 37040 14192 37104
rect 14256 37040 14272 37104
rect 14336 37040 14352 37104
rect 14416 37040 14424 37104
rect 14104 37024 14424 37040
rect 14104 36960 14112 37024
rect 14176 36960 14192 37024
rect 14256 36960 14272 37024
rect 14336 36960 14352 37024
rect 14416 36960 14424 37024
rect 14104 36944 14424 36960
rect 14104 36880 14112 36944
rect 14176 36880 14192 36944
rect 14256 36880 14272 36944
rect 14336 36880 14352 36944
rect 14416 36880 14424 36944
rect 14104 36864 14424 36880
rect 14104 36800 14112 36864
rect 14176 36800 14192 36864
rect 14256 36800 14272 36864
rect 14336 36800 14352 36864
rect 14416 36800 14424 36864
rect 14104 36784 14424 36800
rect 14104 36720 14112 36784
rect 14176 36720 14192 36784
rect 14256 36720 14272 36784
rect 14336 36720 14352 36784
rect 14416 36720 14424 36784
rect 14104 36704 14424 36720
rect 14104 36640 14112 36704
rect 14176 36640 14192 36704
rect 14256 36640 14272 36704
rect 14336 36640 14352 36704
rect 14416 36640 14424 36704
rect 14104 36624 14424 36640
rect 14104 36560 14112 36624
rect 14176 36560 14192 36624
rect 14256 36560 14272 36624
rect 14336 36560 14352 36624
rect 14416 36560 14424 36624
rect 14104 36544 14424 36560
rect 14104 36480 14112 36544
rect 14176 36480 14192 36544
rect 14256 36480 14272 36544
rect 14336 36480 14352 36544
rect 14416 36480 14424 36544
rect 14104 36464 14424 36480
rect 14104 36400 14112 36464
rect 14176 36400 14192 36464
rect 14256 36400 14272 36464
rect 14336 36400 14352 36464
rect 14416 36400 14424 36464
rect 14104 33880 14424 36400
rect 14104 33816 14112 33880
rect 14176 33816 14192 33880
rect 14256 33816 14272 33880
rect 14336 33816 14352 33880
rect 14416 33816 14424 33880
rect 14104 32792 14424 33816
rect 14104 32728 14112 32792
rect 14176 32728 14192 32792
rect 14256 32728 14272 32792
rect 14336 32728 14352 32792
rect 14416 32728 14424 32792
rect 14104 31704 14424 32728
rect 14104 31640 14112 31704
rect 14176 31640 14192 31704
rect 14256 31640 14272 31704
rect 14336 31640 14352 31704
rect 14416 31640 14424 31704
rect 14104 30616 14424 31640
rect 14104 30552 14112 30616
rect 14176 30552 14192 30616
rect 14256 30552 14272 30616
rect 14336 30552 14352 30616
rect 14416 30552 14424 30616
rect 14104 29528 14424 30552
rect 14104 29464 14112 29528
rect 14176 29464 14192 29528
rect 14256 29464 14272 29528
rect 14336 29464 14352 29528
rect 14416 29464 14424 29528
rect 14104 28440 14424 29464
rect 14104 28376 14112 28440
rect 14176 28376 14192 28440
rect 14256 28376 14272 28440
rect 14336 28376 14352 28440
rect 14416 28376 14424 28440
rect 14104 27352 14424 28376
rect 14104 27288 14112 27352
rect 14176 27288 14192 27352
rect 14256 27288 14272 27352
rect 14336 27288 14352 27352
rect 14416 27288 14424 27352
rect 14104 26264 14424 27288
rect 14104 26200 14112 26264
rect 14176 26200 14192 26264
rect 14256 26200 14272 26264
rect 14336 26200 14352 26264
rect 14416 26200 14424 26264
rect 14104 25176 14424 26200
rect 14104 25112 14112 25176
rect 14176 25112 14192 25176
rect 14256 25112 14272 25176
rect 14336 25112 14352 25176
rect 14416 25112 14424 25176
rect 14104 24088 14424 25112
rect 14104 24024 14112 24088
rect 14176 24024 14192 24088
rect 14256 24024 14272 24088
rect 14336 24024 14352 24088
rect 14416 24024 14424 24088
rect 14104 23000 14424 24024
rect 14104 22936 14112 23000
rect 14176 22936 14192 23000
rect 14256 22936 14272 23000
rect 14336 22936 14352 23000
rect 14416 22936 14424 23000
rect 14104 21912 14424 22936
rect 14104 21848 14112 21912
rect 14176 21848 14192 21912
rect 14256 21848 14272 21912
rect 14336 21848 14352 21912
rect 14416 21848 14424 21912
rect 14104 20824 14424 21848
rect 14104 20760 14112 20824
rect 14176 20760 14192 20824
rect 14256 20760 14272 20824
rect 14336 20760 14352 20824
rect 14416 20760 14424 20824
rect 14104 19736 14424 20760
rect 14104 19672 14112 19736
rect 14176 19672 14192 19736
rect 14256 19672 14272 19736
rect 14336 19672 14352 19736
rect 14416 19672 14424 19736
rect 14104 18648 14424 19672
rect 14104 18584 14112 18648
rect 14176 18584 14192 18648
rect 14256 18584 14272 18648
rect 14336 18584 14352 18648
rect 14416 18584 14424 18648
rect 14104 17560 14424 18584
rect 14104 17496 14112 17560
rect 14176 17496 14192 17560
rect 14256 17496 14272 17560
rect 14336 17496 14352 17560
rect 14416 17496 14424 17560
rect 14104 16472 14424 17496
rect 14104 16408 14112 16472
rect 14176 16408 14192 16472
rect 14256 16408 14272 16472
rect 14336 16408 14352 16472
rect 14416 16408 14424 16472
rect 14104 15384 14424 16408
rect 14104 15320 14112 15384
rect 14176 15320 14192 15384
rect 14256 15320 14272 15384
rect 14336 15320 14352 15384
rect 14416 15320 14424 15384
rect 14104 14296 14424 15320
rect 14104 14232 14112 14296
rect 14176 14232 14192 14296
rect 14256 14232 14272 14296
rect 14336 14232 14352 14296
rect 14416 14232 14424 14296
rect 14104 13208 14424 14232
rect 14104 13144 14112 13208
rect 14176 13144 14192 13208
rect 14256 13144 14272 13208
rect 14336 13144 14352 13208
rect 14416 13144 14424 13208
rect 14104 12120 14424 13144
rect 14104 12056 14112 12120
rect 14176 12056 14192 12120
rect 14256 12056 14272 12120
rect 14336 12056 14352 12120
rect 14416 12056 14424 12120
rect 14104 11032 14424 12056
rect 14104 10968 14112 11032
rect 14176 10968 14192 11032
rect 14256 10968 14272 11032
rect 14336 10968 14352 11032
rect 14416 10968 14424 11032
rect 14104 8992 14424 10968
rect 14104 8928 14112 8992
rect 14176 8928 14192 8992
rect 14256 8928 14272 8992
rect 14336 8928 14352 8992
rect 14416 8928 14424 8992
rect 14104 8912 14424 8928
rect 14104 8848 14112 8912
rect 14176 8848 14192 8912
rect 14256 8848 14272 8912
rect 14336 8848 14352 8912
rect 14416 8848 14424 8912
rect 14104 8832 14424 8848
rect 14104 8768 14112 8832
rect 14176 8768 14192 8832
rect 14256 8768 14272 8832
rect 14336 8768 14352 8832
rect 14416 8768 14424 8832
rect 14104 8752 14424 8768
rect 14104 8688 14112 8752
rect 14176 8688 14192 8752
rect 14256 8688 14272 8752
rect 14336 8688 14352 8752
rect 14416 8688 14424 8752
rect 14104 8672 14424 8688
rect 14104 8608 14112 8672
rect 14176 8608 14192 8672
rect 14256 8608 14272 8672
rect 14336 8608 14352 8672
rect 14416 8608 14424 8672
rect 14104 8592 14424 8608
rect 14104 8528 14112 8592
rect 14176 8528 14192 8592
rect 14256 8528 14272 8592
rect 14336 8528 14352 8592
rect 14416 8528 14424 8592
rect 14104 8512 14424 8528
rect 14104 8448 14112 8512
rect 14176 8448 14192 8512
rect 14256 8448 14272 8512
rect 14336 8448 14352 8512
rect 14416 8448 14424 8512
rect 14104 8432 14424 8448
rect 14104 8368 14112 8432
rect 14176 8368 14192 8432
rect 14256 8368 14272 8432
rect 14336 8368 14352 8432
rect 14416 8368 14424 8432
rect 14104 8352 14424 8368
rect 14104 8288 14112 8352
rect 14176 8288 14192 8352
rect 14256 8288 14272 8352
rect 14336 8288 14352 8352
rect 14416 8288 14424 8352
rect 14104 8272 14424 8288
rect 14104 8208 14112 8272
rect 14176 8208 14192 8272
rect 14256 8208 14272 8272
rect 14336 8208 14352 8272
rect 14416 8208 14424 8272
rect 14104 8192 14424 8208
rect 14104 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14272 8192
rect 14336 8128 14352 8192
rect 14416 8128 14424 8192
rect 14104 8112 14424 8128
rect 14104 8048 14112 8112
rect 14176 8048 14192 8112
rect 14256 8048 14272 8112
rect 14336 8048 14352 8112
rect 14416 8048 14424 8112
rect 14104 8032 14424 8048
rect 14104 7968 14112 8032
rect 14176 7968 14192 8032
rect 14256 7968 14272 8032
rect 14336 7968 14352 8032
rect 14416 7968 14424 8032
rect 14104 7952 14424 7968
rect 14104 7888 14112 7952
rect 14176 7888 14192 7952
rect 14256 7888 14272 7952
rect 14336 7888 14352 7952
rect 14416 7888 14424 7952
rect 14104 7872 14424 7888
rect 14104 7808 14112 7872
rect 14176 7808 14192 7872
rect 14256 7808 14272 7872
rect 14336 7808 14352 7872
rect 14416 7808 14424 7872
rect 14104 7792 14424 7808
rect 14104 7728 14112 7792
rect 14176 7728 14192 7792
rect 14256 7728 14272 7792
rect 14336 7728 14352 7792
rect 14416 7728 14424 7792
rect 14104 7712 14424 7728
rect 14104 7648 14112 7712
rect 14176 7648 14192 7712
rect 14256 7648 14272 7712
rect 14336 7648 14352 7712
rect 14416 7648 14424 7712
rect 14104 7632 14424 7648
rect 14104 7568 14112 7632
rect 14176 7568 14192 7632
rect 14256 7568 14272 7632
rect 14336 7568 14352 7632
rect 14416 7568 14424 7632
rect 14104 7552 14424 7568
rect 14104 7488 14112 7552
rect 14176 7488 14192 7552
rect 14256 7488 14272 7552
rect 14336 7488 14352 7552
rect 14416 7488 14424 7552
rect 14104 7472 14424 7488
rect 14104 7408 14112 7472
rect 14176 7408 14192 7472
rect 14256 7408 14272 7472
rect 14336 7408 14352 7472
rect 14416 7408 14424 7472
rect 14104 7392 14424 7408
rect 14104 7328 14112 7392
rect 14176 7328 14192 7392
rect 14256 7328 14272 7392
rect 14336 7328 14352 7392
rect 14416 7328 14424 7392
rect 14104 7312 14424 7328
rect 14104 7248 14112 7312
rect 14176 7248 14192 7312
rect 14256 7248 14272 7312
rect 14336 7248 14352 7312
rect 14416 7248 14424 7312
rect 14104 7232 14424 7248
rect 14104 7168 14112 7232
rect 14176 7168 14192 7232
rect 14256 7168 14272 7232
rect 14336 7168 14352 7232
rect 14416 7168 14424 7232
rect 14104 7152 14424 7168
rect 14104 7088 14112 7152
rect 14176 7088 14192 7152
rect 14256 7088 14272 7152
rect 14336 7088 14352 7152
rect 14416 7088 14424 7152
rect 14104 7072 14424 7088
rect 14104 7008 14112 7072
rect 14176 7008 14192 7072
rect 14256 7008 14272 7072
rect 14336 7008 14352 7072
rect 14416 7008 14424 7072
rect 14104 6992 14424 7008
rect 14104 6928 14112 6992
rect 14176 6928 14192 6992
rect 14256 6928 14272 6992
rect 14336 6928 14352 6992
rect 14416 6928 14424 6992
rect 14104 6912 14424 6928
rect 14104 6848 14112 6912
rect 14176 6848 14192 6912
rect 14256 6848 14272 6912
rect 14336 6848 14352 6912
rect 14416 6848 14424 6912
rect 14104 6832 14424 6848
rect 14104 6768 14112 6832
rect 14176 6768 14192 6832
rect 14256 6768 14272 6832
rect 14336 6768 14352 6832
rect 14416 6768 14424 6832
rect 14104 6752 14424 6768
rect 14104 6688 14112 6752
rect 14176 6688 14192 6752
rect 14256 6688 14272 6752
rect 14336 6688 14352 6752
rect 14416 6688 14424 6752
rect 14104 6672 14424 6688
rect 14104 6608 14112 6672
rect 14176 6608 14192 6672
rect 14256 6608 14272 6672
rect 14336 6608 14352 6672
rect 14416 6608 14424 6672
rect 14104 6592 14424 6608
rect 14104 6528 14112 6592
rect 14176 6528 14192 6592
rect 14256 6528 14272 6592
rect 14336 6528 14352 6592
rect 14416 6528 14424 6592
rect 14104 6512 14424 6528
rect 14104 6448 14112 6512
rect 14176 6448 14192 6512
rect 14256 6448 14272 6512
rect 14336 6448 14352 6512
rect 14416 6448 14424 6512
rect 14104 6432 14424 6448
rect 14104 6368 14112 6432
rect 14176 6368 14192 6432
rect 14256 6368 14272 6432
rect 14336 6368 14352 6432
rect 14416 6368 14424 6432
rect 14104 6352 14424 6368
rect 14104 6288 14112 6352
rect 14176 6288 14192 6352
rect 14256 6288 14272 6352
rect 14336 6288 14352 6352
rect 14416 6288 14424 6352
rect 14104 6272 14424 6288
rect 14104 6208 14112 6272
rect 14176 6208 14192 6272
rect 14256 6208 14272 6272
rect 14336 6208 14352 6272
rect 14416 6208 14424 6272
rect 14104 6192 14424 6208
rect 14104 6128 14112 6192
rect 14176 6128 14192 6192
rect 14256 6128 14272 6192
rect 14336 6128 14352 6192
rect 14416 6128 14424 6192
rect 14104 6112 14424 6128
rect 14104 6048 14112 6112
rect 14176 6048 14192 6112
rect 14256 6048 14272 6112
rect 14336 6048 14352 6112
rect 14416 6048 14424 6112
rect 14104 6032 14424 6048
rect 14104 5968 14112 6032
rect 14176 5968 14192 6032
rect 14256 5968 14272 6032
rect 14336 5968 14352 6032
rect 14416 5968 14424 6032
rect 14104 5952 14424 5968
rect 14104 5888 14112 5952
rect 14176 5888 14192 5952
rect 14256 5888 14272 5952
rect 14336 5888 14352 5952
rect 14416 5888 14424 5952
rect 14104 5872 14424 5888
rect 14104 5808 14112 5872
rect 14176 5808 14192 5872
rect 14256 5808 14272 5872
rect 14336 5808 14352 5872
rect 14416 5808 14424 5872
rect 14104 5792 14424 5808
rect 14104 5728 14112 5792
rect 14176 5728 14192 5792
rect 14256 5728 14272 5792
rect 14336 5728 14352 5792
rect 14416 5728 14424 5792
rect 14104 5712 14424 5728
rect 14104 5648 14112 5712
rect 14176 5648 14192 5712
rect 14256 5648 14272 5712
rect 14336 5648 14352 5712
rect 14416 5648 14424 5712
rect 14104 5632 14424 5648
rect 14104 5568 14112 5632
rect 14176 5568 14192 5632
rect 14256 5568 14272 5632
rect 14336 5568 14352 5632
rect 14416 5568 14424 5632
rect 14104 5552 14424 5568
rect 14104 5488 14112 5552
rect 14176 5488 14192 5552
rect 14256 5488 14272 5552
rect 14336 5488 14352 5552
rect 14416 5488 14424 5552
rect 14104 5472 14424 5488
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 5392 14424 5408
rect 14104 5328 14112 5392
rect 14176 5328 14192 5392
rect 14256 5328 14272 5392
rect 14336 5328 14352 5392
rect 14416 5328 14424 5392
rect 14104 5312 14424 5328
rect 14104 5248 14112 5312
rect 14176 5248 14192 5312
rect 14256 5248 14272 5312
rect 14336 5248 14352 5312
rect 14416 5248 14424 5312
rect 14104 5232 14424 5248
rect 14104 5168 14112 5232
rect 14176 5168 14192 5232
rect 14256 5168 14272 5232
rect 14336 5168 14352 5232
rect 14416 5168 14424 5232
rect 14104 5152 14424 5168
rect 14104 5088 14112 5152
rect 14176 5088 14192 5152
rect 14256 5088 14272 5152
rect 14336 5088 14352 5152
rect 14416 5088 14424 5152
rect 14104 5072 14424 5088
rect 14104 5008 14112 5072
rect 14176 5008 14192 5072
rect 14256 5008 14272 5072
rect 14336 5008 14352 5072
rect 14416 5008 14424 5072
rect 0 3928 8 3992
rect 72 3928 88 3992
rect 152 3928 168 3992
rect 232 3928 248 3992
rect 312 3928 328 3992
rect 392 3928 408 3992
rect 472 3928 488 3992
rect 552 3928 568 3992
rect 632 3928 648 3992
rect 712 3928 728 3992
rect 792 3928 808 3992
rect 872 3928 888 3992
rect 952 3928 968 3992
rect 1032 3928 1048 3992
rect 1112 3928 1128 3992
rect 1192 3928 1208 3992
rect 1272 3928 1288 3992
rect 1352 3928 1368 3992
rect 1432 3928 1448 3992
rect 1512 3928 1528 3992
rect 1592 3928 1608 3992
rect 1672 3928 1688 3992
rect 1752 3928 1768 3992
rect 1832 3928 1848 3992
rect 1912 3928 1928 3992
rect 1992 3928 2008 3992
rect 2072 3928 2088 3992
rect 2152 3928 2168 3992
rect 2232 3928 2248 3992
rect 2312 3928 2328 3992
rect 2392 3928 2408 3992
rect 2472 3928 2488 3992
rect 2552 3928 2568 3992
rect 2632 3928 2648 3992
rect 2712 3928 2728 3992
rect 2792 3928 2808 3992
rect 2872 3928 2888 3992
rect 2952 3928 2968 3992
rect 3032 3928 3048 3992
rect 3112 3928 3128 3992
rect 3192 3928 3208 3992
rect 3272 3928 3288 3992
rect 3352 3928 3368 3992
rect 3432 3928 3448 3992
rect 3512 3928 3528 3992
rect 3592 3928 3608 3992
rect 3672 3928 3688 3992
rect 3752 3928 3768 3992
rect 3832 3928 3848 3992
rect 3912 3928 3928 3992
rect 3992 3928 4000 3992
rect 0 3912 4000 3928
rect 0 3848 8 3912
rect 72 3848 88 3912
rect 152 3848 168 3912
rect 232 3848 248 3912
rect 312 3848 328 3912
rect 392 3848 408 3912
rect 472 3848 488 3912
rect 552 3848 568 3912
rect 632 3848 648 3912
rect 712 3848 728 3912
rect 792 3848 808 3912
rect 872 3848 888 3912
rect 952 3848 968 3912
rect 1032 3848 1048 3912
rect 1112 3848 1128 3912
rect 1192 3848 1208 3912
rect 1272 3848 1288 3912
rect 1352 3848 1368 3912
rect 1432 3848 1448 3912
rect 1512 3848 1528 3912
rect 1592 3848 1608 3912
rect 1672 3848 1688 3912
rect 1752 3848 1768 3912
rect 1832 3848 1848 3912
rect 1912 3848 1928 3912
rect 1992 3848 2008 3912
rect 2072 3848 2088 3912
rect 2152 3848 2168 3912
rect 2232 3848 2248 3912
rect 2312 3848 2328 3912
rect 2392 3848 2408 3912
rect 2472 3848 2488 3912
rect 2552 3848 2568 3912
rect 2632 3848 2648 3912
rect 2712 3848 2728 3912
rect 2792 3848 2808 3912
rect 2872 3848 2888 3912
rect 2952 3848 2968 3912
rect 3032 3848 3048 3912
rect 3112 3848 3128 3912
rect 3192 3848 3208 3912
rect 3272 3848 3288 3912
rect 3352 3848 3368 3912
rect 3432 3848 3448 3912
rect 3512 3848 3528 3912
rect 3592 3848 3608 3912
rect 3672 3848 3688 3912
rect 3752 3848 3768 3912
rect 3832 3848 3848 3912
rect 3912 3848 3928 3912
rect 3992 3848 4000 3912
rect 0 3832 4000 3848
rect 0 3768 8 3832
rect 72 3768 88 3832
rect 152 3768 168 3832
rect 232 3768 248 3832
rect 312 3768 328 3832
rect 392 3768 408 3832
rect 472 3768 488 3832
rect 552 3768 568 3832
rect 632 3768 648 3832
rect 712 3768 728 3832
rect 792 3768 808 3832
rect 872 3768 888 3832
rect 952 3768 968 3832
rect 1032 3768 1048 3832
rect 1112 3768 1128 3832
rect 1192 3768 1208 3832
rect 1272 3768 1288 3832
rect 1352 3768 1368 3832
rect 1432 3768 1448 3832
rect 1512 3768 1528 3832
rect 1592 3768 1608 3832
rect 1672 3768 1688 3832
rect 1752 3768 1768 3832
rect 1832 3768 1848 3832
rect 1912 3768 1928 3832
rect 1992 3768 2008 3832
rect 2072 3768 2088 3832
rect 2152 3768 2168 3832
rect 2232 3768 2248 3832
rect 2312 3768 2328 3832
rect 2392 3768 2408 3832
rect 2472 3768 2488 3832
rect 2552 3768 2568 3832
rect 2632 3768 2648 3832
rect 2712 3768 2728 3832
rect 2792 3768 2808 3832
rect 2872 3768 2888 3832
rect 2952 3768 2968 3832
rect 3032 3768 3048 3832
rect 3112 3768 3128 3832
rect 3192 3768 3208 3832
rect 3272 3768 3288 3832
rect 3352 3768 3368 3832
rect 3432 3768 3448 3832
rect 3512 3768 3528 3832
rect 3592 3768 3608 3832
rect 3672 3768 3688 3832
rect 3752 3768 3768 3832
rect 3832 3768 3848 3832
rect 3912 3768 3928 3832
rect 3992 3768 4000 3832
rect 0 3752 4000 3768
rect 0 3688 8 3752
rect 72 3688 88 3752
rect 152 3688 168 3752
rect 232 3688 248 3752
rect 312 3688 328 3752
rect 392 3688 408 3752
rect 472 3688 488 3752
rect 552 3688 568 3752
rect 632 3688 648 3752
rect 712 3688 728 3752
rect 792 3688 808 3752
rect 872 3688 888 3752
rect 952 3688 968 3752
rect 1032 3688 1048 3752
rect 1112 3688 1128 3752
rect 1192 3688 1208 3752
rect 1272 3688 1288 3752
rect 1352 3688 1368 3752
rect 1432 3688 1448 3752
rect 1512 3688 1528 3752
rect 1592 3688 1608 3752
rect 1672 3688 1688 3752
rect 1752 3688 1768 3752
rect 1832 3688 1848 3752
rect 1912 3688 1928 3752
rect 1992 3688 2008 3752
rect 2072 3688 2088 3752
rect 2152 3688 2168 3752
rect 2232 3688 2248 3752
rect 2312 3688 2328 3752
rect 2392 3688 2408 3752
rect 2472 3688 2488 3752
rect 2552 3688 2568 3752
rect 2632 3688 2648 3752
rect 2712 3688 2728 3752
rect 2792 3688 2808 3752
rect 2872 3688 2888 3752
rect 2952 3688 2968 3752
rect 3032 3688 3048 3752
rect 3112 3688 3128 3752
rect 3192 3688 3208 3752
rect 3272 3688 3288 3752
rect 3352 3688 3368 3752
rect 3432 3688 3448 3752
rect 3512 3688 3528 3752
rect 3592 3688 3608 3752
rect 3672 3688 3688 3752
rect 3752 3688 3768 3752
rect 3832 3688 3848 3752
rect 3912 3688 3928 3752
rect 3992 3688 4000 3752
rect 0 3672 4000 3688
rect 0 3608 8 3672
rect 72 3608 88 3672
rect 152 3608 168 3672
rect 232 3608 248 3672
rect 312 3608 328 3672
rect 392 3608 408 3672
rect 472 3608 488 3672
rect 552 3608 568 3672
rect 632 3608 648 3672
rect 712 3608 728 3672
rect 792 3608 808 3672
rect 872 3608 888 3672
rect 952 3608 968 3672
rect 1032 3608 1048 3672
rect 1112 3608 1128 3672
rect 1192 3608 1208 3672
rect 1272 3608 1288 3672
rect 1352 3608 1368 3672
rect 1432 3608 1448 3672
rect 1512 3608 1528 3672
rect 1592 3608 1608 3672
rect 1672 3608 1688 3672
rect 1752 3608 1768 3672
rect 1832 3608 1848 3672
rect 1912 3608 1928 3672
rect 1992 3608 2008 3672
rect 2072 3608 2088 3672
rect 2152 3608 2168 3672
rect 2232 3608 2248 3672
rect 2312 3608 2328 3672
rect 2392 3608 2408 3672
rect 2472 3608 2488 3672
rect 2552 3608 2568 3672
rect 2632 3608 2648 3672
rect 2712 3608 2728 3672
rect 2792 3608 2808 3672
rect 2872 3608 2888 3672
rect 2952 3608 2968 3672
rect 3032 3608 3048 3672
rect 3112 3608 3128 3672
rect 3192 3608 3208 3672
rect 3272 3608 3288 3672
rect 3352 3608 3368 3672
rect 3432 3608 3448 3672
rect 3512 3608 3528 3672
rect 3592 3608 3608 3672
rect 3672 3608 3688 3672
rect 3752 3608 3768 3672
rect 3832 3608 3848 3672
rect 3912 3608 3928 3672
rect 3992 3608 4000 3672
rect 0 3592 4000 3608
rect 0 3528 8 3592
rect 72 3528 88 3592
rect 152 3528 168 3592
rect 232 3528 248 3592
rect 312 3528 328 3592
rect 392 3528 408 3592
rect 472 3528 488 3592
rect 552 3528 568 3592
rect 632 3528 648 3592
rect 712 3528 728 3592
rect 792 3528 808 3592
rect 872 3528 888 3592
rect 952 3528 968 3592
rect 1032 3528 1048 3592
rect 1112 3528 1128 3592
rect 1192 3528 1208 3592
rect 1272 3528 1288 3592
rect 1352 3528 1368 3592
rect 1432 3528 1448 3592
rect 1512 3528 1528 3592
rect 1592 3528 1608 3592
rect 1672 3528 1688 3592
rect 1752 3528 1768 3592
rect 1832 3528 1848 3592
rect 1912 3528 1928 3592
rect 1992 3528 2008 3592
rect 2072 3528 2088 3592
rect 2152 3528 2168 3592
rect 2232 3528 2248 3592
rect 2312 3528 2328 3592
rect 2392 3528 2408 3592
rect 2472 3528 2488 3592
rect 2552 3528 2568 3592
rect 2632 3528 2648 3592
rect 2712 3528 2728 3592
rect 2792 3528 2808 3592
rect 2872 3528 2888 3592
rect 2952 3528 2968 3592
rect 3032 3528 3048 3592
rect 3112 3528 3128 3592
rect 3192 3528 3208 3592
rect 3272 3528 3288 3592
rect 3352 3528 3368 3592
rect 3432 3528 3448 3592
rect 3512 3528 3528 3592
rect 3592 3528 3608 3592
rect 3672 3528 3688 3592
rect 3752 3528 3768 3592
rect 3832 3528 3848 3592
rect 3912 3528 3928 3592
rect 3992 3528 4000 3592
rect 0 3512 4000 3528
rect 0 3448 8 3512
rect 72 3448 88 3512
rect 152 3448 168 3512
rect 232 3448 248 3512
rect 312 3448 328 3512
rect 392 3448 408 3512
rect 472 3448 488 3512
rect 552 3448 568 3512
rect 632 3448 648 3512
rect 712 3448 728 3512
rect 792 3448 808 3512
rect 872 3448 888 3512
rect 952 3448 968 3512
rect 1032 3448 1048 3512
rect 1112 3448 1128 3512
rect 1192 3448 1208 3512
rect 1272 3448 1288 3512
rect 1352 3448 1368 3512
rect 1432 3448 1448 3512
rect 1512 3448 1528 3512
rect 1592 3448 1608 3512
rect 1672 3448 1688 3512
rect 1752 3448 1768 3512
rect 1832 3448 1848 3512
rect 1912 3448 1928 3512
rect 1992 3448 2008 3512
rect 2072 3448 2088 3512
rect 2152 3448 2168 3512
rect 2232 3448 2248 3512
rect 2312 3448 2328 3512
rect 2392 3448 2408 3512
rect 2472 3448 2488 3512
rect 2552 3448 2568 3512
rect 2632 3448 2648 3512
rect 2712 3448 2728 3512
rect 2792 3448 2808 3512
rect 2872 3448 2888 3512
rect 2952 3448 2968 3512
rect 3032 3448 3048 3512
rect 3112 3448 3128 3512
rect 3192 3448 3208 3512
rect 3272 3448 3288 3512
rect 3352 3448 3368 3512
rect 3432 3448 3448 3512
rect 3512 3448 3528 3512
rect 3592 3448 3608 3512
rect 3672 3448 3688 3512
rect 3752 3448 3768 3512
rect 3832 3448 3848 3512
rect 3912 3448 3928 3512
rect 3992 3448 4000 3512
rect 0 3432 4000 3448
rect 0 3368 8 3432
rect 72 3368 88 3432
rect 152 3368 168 3432
rect 232 3368 248 3432
rect 312 3368 328 3432
rect 392 3368 408 3432
rect 472 3368 488 3432
rect 552 3368 568 3432
rect 632 3368 648 3432
rect 712 3368 728 3432
rect 792 3368 808 3432
rect 872 3368 888 3432
rect 952 3368 968 3432
rect 1032 3368 1048 3432
rect 1112 3368 1128 3432
rect 1192 3368 1208 3432
rect 1272 3368 1288 3432
rect 1352 3368 1368 3432
rect 1432 3368 1448 3432
rect 1512 3368 1528 3432
rect 1592 3368 1608 3432
rect 1672 3368 1688 3432
rect 1752 3368 1768 3432
rect 1832 3368 1848 3432
rect 1912 3368 1928 3432
rect 1992 3368 2008 3432
rect 2072 3368 2088 3432
rect 2152 3368 2168 3432
rect 2232 3368 2248 3432
rect 2312 3368 2328 3432
rect 2392 3368 2408 3432
rect 2472 3368 2488 3432
rect 2552 3368 2568 3432
rect 2632 3368 2648 3432
rect 2712 3368 2728 3432
rect 2792 3368 2808 3432
rect 2872 3368 2888 3432
rect 2952 3368 2968 3432
rect 3032 3368 3048 3432
rect 3112 3368 3128 3432
rect 3192 3368 3208 3432
rect 3272 3368 3288 3432
rect 3352 3368 3368 3432
rect 3432 3368 3448 3432
rect 3512 3368 3528 3432
rect 3592 3368 3608 3432
rect 3672 3368 3688 3432
rect 3752 3368 3768 3432
rect 3832 3368 3848 3432
rect 3912 3368 3928 3432
rect 3992 3368 4000 3432
rect 0 3352 4000 3368
rect 0 3288 8 3352
rect 72 3288 88 3352
rect 152 3288 168 3352
rect 232 3288 248 3352
rect 312 3288 328 3352
rect 392 3288 408 3352
rect 472 3288 488 3352
rect 552 3288 568 3352
rect 632 3288 648 3352
rect 712 3288 728 3352
rect 792 3288 808 3352
rect 872 3288 888 3352
rect 952 3288 968 3352
rect 1032 3288 1048 3352
rect 1112 3288 1128 3352
rect 1192 3288 1208 3352
rect 1272 3288 1288 3352
rect 1352 3288 1368 3352
rect 1432 3288 1448 3352
rect 1512 3288 1528 3352
rect 1592 3288 1608 3352
rect 1672 3288 1688 3352
rect 1752 3288 1768 3352
rect 1832 3288 1848 3352
rect 1912 3288 1928 3352
rect 1992 3288 2008 3352
rect 2072 3288 2088 3352
rect 2152 3288 2168 3352
rect 2232 3288 2248 3352
rect 2312 3288 2328 3352
rect 2392 3288 2408 3352
rect 2472 3288 2488 3352
rect 2552 3288 2568 3352
rect 2632 3288 2648 3352
rect 2712 3288 2728 3352
rect 2792 3288 2808 3352
rect 2872 3288 2888 3352
rect 2952 3288 2968 3352
rect 3032 3288 3048 3352
rect 3112 3288 3128 3352
rect 3192 3288 3208 3352
rect 3272 3288 3288 3352
rect 3352 3288 3368 3352
rect 3432 3288 3448 3352
rect 3512 3288 3528 3352
rect 3592 3288 3608 3352
rect 3672 3288 3688 3352
rect 3752 3288 3768 3352
rect 3832 3288 3848 3352
rect 3912 3288 3928 3352
rect 3992 3288 4000 3352
rect 0 3272 4000 3288
rect 0 3208 8 3272
rect 72 3208 88 3272
rect 152 3208 168 3272
rect 232 3208 248 3272
rect 312 3208 328 3272
rect 392 3208 408 3272
rect 472 3208 488 3272
rect 552 3208 568 3272
rect 632 3208 648 3272
rect 712 3208 728 3272
rect 792 3208 808 3272
rect 872 3208 888 3272
rect 952 3208 968 3272
rect 1032 3208 1048 3272
rect 1112 3208 1128 3272
rect 1192 3208 1208 3272
rect 1272 3208 1288 3272
rect 1352 3208 1368 3272
rect 1432 3208 1448 3272
rect 1512 3208 1528 3272
rect 1592 3208 1608 3272
rect 1672 3208 1688 3272
rect 1752 3208 1768 3272
rect 1832 3208 1848 3272
rect 1912 3208 1928 3272
rect 1992 3208 2008 3272
rect 2072 3208 2088 3272
rect 2152 3208 2168 3272
rect 2232 3208 2248 3272
rect 2312 3208 2328 3272
rect 2392 3208 2408 3272
rect 2472 3208 2488 3272
rect 2552 3208 2568 3272
rect 2632 3208 2648 3272
rect 2712 3208 2728 3272
rect 2792 3208 2808 3272
rect 2872 3208 2888 3272
rect 2952 3208 2968 3272
rect 3032 3208 3048 3272
rect 3112 3208 3128 3272
rect 3192 3208 3208 3272
rect 3272 3208 3288 3272
rect 3352 3208 3368 3272
rect 3432 3208 3448 3272
rect 3512 3208 3528 3272
rect 3592 3208 3608 3272
rect 3672 3208 3688 3272
rect 3752 3208 3768 3272
rect 3832 3208 3848 3272
rect 3912 3208 3928 3272
rect 3992 3208 4000 3272
rect 0 3192 4000 3208
rect 0 3128 8 3192
rect 72 3128 88 3192
rect 152 3128 168 3192
rect 232 3128 248 3192
rect 312 3128 328 3192
rect 392 3128 408 3192
rect 472 3128 488 3192
rect 552 3128 568 3192
rect 632 3128 648 3192
rect 712 3128 728 3192
rect 792 3128 808 3192
rect 872 3128 888 3192
rect 952 3128 968 3192
rect 1032 3128 1048 3192
rect 1112 3128 1128 3192
rect 1192 3128 1208 3192
rect 1272 3128 1288 3192
rect 1352 3128 1368 3192
rect 1432 3128 1448 3192
rect 1512 3128 1528 3192
rect 1592 3128 1608 3192
rect 1672 3128 1688 3192
rect 1752 3128 1768 3192
rect 1832 3128 1848 3192
rect 1912 3128 1928 3192
rect 1992 3128 2008 3192
rect 2072 3128 2088 3192
rect 2152 3128 2168 3192
rect 2232 3128 2248 3192
rect 2312 3128 2328 3192
rect 2392 3128 2408 3192
rect 2472 3128 2488 3192
rect 2552 3128 2568 3192
rect 2632 3128 2648 3192
rect 2712 3128 2728 3192
rect 2792 3128 2808 3192
rect 2872 3128 2888 3192
rect 2952 3128 2968 3192
rect 3032 3128 3048 3192
rect 3112 3128 3128 3192
rect 3192 3128 3208 3192
rect 3272 3128 3288 3192
rect 3352 3128 3368 3192
rect 3432 3128 3448 3192
rect 3512 3128 3528 3192
rect 3592 3128 3608 3192
rect 3672 3128 3688 3192
rect 3752 3128 3768 3192
rect 3832 3128 3848 3192
rect 3912 3128 3928 3192
rect 3992 3128 4000 3192
rect 0 3112 4000 3128
rect 0 3048 8 3112
rect 72 3048 88 3112
rect 152 3048 168 3112
rect 232 3048 248 3112
rect 312 3048 328 3112
rect 392 3048 408 3112
rect 472 3048 488 3112
rect 552 3048 568 3112
rect 632 3048 648 3112
rect 712 3048 728 3112
rect 792 3048 808 3112
rect 872 3048 888 3112
rect 952 3048 968 3112
rect 1032 3048 1048 3112
rect 1112 3048 1128 3112
rect 1192 3048 1208 3112
rect 1272 3048 1288 3112
rect 1352 3048 1368 3112
rect 1432 3048 1448 3112
rect 1512 3048 1528 3112
rect 1592 3048 1608 3112
rect 1672 3048 1688 3112
rect 1752 3048 1768 3112
rect 1832 3048 1848 3112
rect 1912 3048 1928 3112
rect 1992 3048 2008 3112
rect 2072 3048 2088 3112
rect 2152 3048 2168 3112
rect 2232 3048 2248 3112
rect 2312 3048 2328 3112
rect 2392 3048 2408 3112
rect 2472 3048 2488 3112
rect 2552 3048 2568 3112
rect 2632 3048 2648 3112
rect 2712 3048 2728 3112
rect 2792 3048 2808 3112
rect 2872 3048 2888 3112
rect 2952 3048 2968 3112
rect 3032 3048 3048 3112
rect 3112 3048 3128 3112
rect 3192 3048 3208 3112
rect 3272 3048 3288 3112
rect 3352 3048 3368 3112
rect 3432 3048 3448 3112
rect 3512 3048 3528 3112
rect 3592 3048 3608 3112
rect 3672 3048 3688 3112
rect 3752 3048 3768 3112
rect 3832 3048 3848 3112
rect 3912 3048 3928 3112
rect 3992 3048 4000 3112
rect 0 3032 4000 3048
rect 0 2968 8 3032
rect 72 2968 88 3032
rect 152 2968 168 3032
rect 232 2968 248 3032
rect 312 2968 328 3032
rect 392 2968 408 3032
rect 472 2968 488 3032
rect 552 2968 568 3032
rect 632 2968 648 3032
rect 712 2968 728 3032
rect 792 2968 808 3032
rect 872 2968 888 3032
rect 952 2968 968 3032
rect 1032 2968 1048 3032
rect 1112 2968 1128 3032
rect 1192 2968 1208 3032
rect 1272 2968 1288 3032
rect 1352 2968 1368 3032
rect 1432 2968 1448 3032
rect 1512 2968 1528 3032
rect 1592 2968 1608 3032
rect 1672 2968 1688 3032
rect 1752 2968 1768 3032
rect 1832 2968 1848 3032
rect 1912 2968 1928 3032
rect 1992 2968 2008 3032
rect 2072 2968 2088 3032
rect 2152 2968 2168 3032
rect 2232 2968 2248 3032
rect 2312 2968 2328 3032
rect 2392 2968 2408 3032
rect 2472 2968 2488 3032
rect 2552 2968 2568 3032
rect 2632 2968 2648 3032
rect 2712 2968 2728 3032
rect 2792 2968 2808 3032
rect 2872 2968 2888 3032
rect 2952 2968 2968 3032
rect 3032 2968 3048 3032
rect 3112 2968 3128 3032
rect 3192 2968 3208 3032
rect 3272 2968 3288 3032
rect 3352 2968 3368 3032
rect 3432 2968 3448 3032
rect 3512 2968 3528 3032
rect 3592 2968 3608 3032
rect 3672 2968 3688 3032
rect 3752 2968 3768 3032
rect 3832 2968 3848 3032
rect 3912 2968 3928 3032
rect 3992 2968 4000 3032
rect 0 2952 4000 2968
rect 0 2888 8 2952
rect 72 2888 88 2952
rect 152 2888 168 2952
rect 232 2888 248 2952
rect 312 2888 328 2952
rect 392 2888 408 2952
rect 472 2888 488 2952
rect 552 2888 568 2952
rect 632 2888 648 2952
rect 712 2888 728 2952
rect 792 2888 808 2952
rect 872 2888 888 2952
rect 952 2888 968 2952
rect 1032 2888 1048 2952
rect 1112 2888 1128 2952
rect 1192 2888 1208 2952
rect 1272 2888 1288 2952
rect 1352 2888 1368 2952
rect 1432 2888 1448 2952
rect 1512 2888 1528 2952
rect 1592 2888 1608 2952
rect 1672 2888 1688 2952
rect 1752 2888 1768 2952
rect 1832 2888 1848 2952
rect 1912 2888 1928 2952
rect 1992 2888 2008 2952
rect 2072 2888 2088 2952
rect 2152 2888 2168 2952
rect 2232 2888 2248 2952
rect 2312 2888 2328 2952
rect 2392 2888 2408 2952
rect 2472 2888 2488 2952
rect 2552 2888 2568 2952
rect 2632 2888 2648 2952
rect 2712 2888 2728 2952
rect 2792 2888 2808 2952
rect 2872 2888 2888 2952
rect 2952 2888 2968 2952
rect 3032 2888 3048 2952
rect 3112 2888 3128 2952
rect 3192 2888 3208 2952
rect 3272 2888 3288 2952
rect 3352 2888 3368 2952
rect 3432 2888 3448 2952
rect 3512 2888 3528 2952
rect 3592 2888 3608 2952
rect 3672 2888 3688 2952
rect 3752 2888 3768 2952
rect 3832 2888 3848 2952
rect 3912 2888 3928 2952
rect 3992 2888 4000 2952
rect 0 2872 4000 2888
rect 0 2808 8 2872
rect 72 2808 88 2872
rect 152 2808 168 2872
rect 232 2808 248 2872
rect 312 2808 328 2872
rect 392 2808 408 2872
rect 472 2808 488 2872
rect 552 2808 568 2872
rect 632 2808 648 2872
rect 712 2808 728 2872
rect 792 2808 808 2872
rect 872 2808 888 2872
rect 952 2808 968 2872
rect 1032 2808 1048 2872
rect 1112 2808 1128 2872
rect 1192 2808 1208 2872
rect 1272 2808 1288 2872
rect 1352 2808 1368 2872
rect 1432 2808 1448 2872
rect 1512 2808 1528 2872
rect 1592 2808 1608 2872
rect 1672 2808 1688 2872
rect 1752 2808 1768 2872
rect 1832 2808 1848 2872
rect 1912 2808 1928 2872
rect 1992 2808 2008 2872
rect 2072 2808 2088 2872
rect 2152 2808 2168 2872
rect 2232 2808 2248 2872
rect 2312 2808 2328 2872
rect 2392 2808 2408 2872
rect 2472 2808 2488 2872
rect 2552 2808 2568 2872
rect 2632 2808 2648 2872
rect 2712 2808 2728 2872
rect 2792 2808 2808 2872
rect 2872 2808 2888 2872
rect 2952 2808 2968 2872
rect 3032 2808 3048 2872
rect 3112 2808 3128 2872
rect 3192 2808 3208 2872
rect 3272 2808 3288 2872
rect 3352 2808 3368 2872
rect 3432 2808 3448 2872
rect 3512 2808 3528 2872
rect 3592 2808 3608 2872
rect 3672 2808 3688 2872
rect 3752 2808 3768 2872
rect 3832 2808 3848 2872
rect 3912 2808 3928 2872
rect 3992 2808 4000 2872
rect 0 2792 4000 2808
rect 0 2728 8 2792
rect 72 2728 88 2792
rect 152 2728 168 2792
rect 232 2728 248 2792
rect 312 2728 328 2792
rect 392 2728 408 2792
rect 472 2728 488 2792
rect 552 2728 568 2792
rect 632 2728 648 2792
rect 712 2728 728 2792
rect 792 2728 808 2792
rect 872 2728 888 2792
rect 952 2728 968 2792
rect 1032 2728 1048 2792
rect 1112 2728 1128 2792
rect 1192 2728 1208 2792
rect 1272 2728 1288 2792
rect 1352 2728 1368 2792
rect 1432 2728 1448 2792
rect 1512 2728 1528 2792
rect 1592 2728 1608 2792
rect 1672 2728 1688 2792
rect 1752 2728 1768 2792
rect 1832 2728 1848 2792
rect 1912 2728 1928 2792
rect 1992 2728 2008 2792
rect 2072 2728 2088 2792
rect 2152 2728 2168 2792
rect 2232 2728 2248 2792
rect 2312 2728 2328 2792
rect 2392 2728 2408 2792
rect 2472 2728 2488 2792
rect 2552 2728 2568 2792
rect 2632 2728 2648 2792
rect 2712 2728 2728 2792
rect 2792 2728 2808 2792
rect 2872 2728 2888 2792
rect 2952 2728 2968 2792
rect 3032 2728 3048 2792
rect 3112 2728 3128 2792
rect 3192 2728 3208 2792
rect 3272 2728 3288 2792
rect 3352 2728 3368 2792
rect 3432 2728 3448 2792
rect 3512 2728 3528 2792
rect 3592 2728 3608 2792
rect 3672 2728 3688 2792
rect 3752 2728 3768 2792
rect 3832 2728 3848 2792
rect 3912 2728 3928 2792
rect 3992 2728 4000 2792
rect 0 2712 4000 2728
rect 0 2648 8 2712
rect 72 2648 88 2712
rect 152 2648 168 2712
rect 232 2648 248 2712
rect 312 2648 328 2712
rect 392 2648 408 2712
rect 472 2648 488 2712
rect 552 2648 568 2712
rect 632 2648 648 2712
rect 712 2648 728 2712
rect 792 2648 808 2712
rect 872 2648 888 2712
rect 952 2648 968 2712
rect 1032 2648 1048 2712
rect 1112 2648 1128 2712
rect 1192 2648 1208 2712
rect 1272 2648 1288 2712
rect 1352 2648 1368 2712
rect 1432 2648 1448 2712
rect 1512 2648 1528 2712
rect 1592 2648 1608 2712
rect 1672 2648 1688 2712
rect 1752 2648 1768 2712
rect 1832 2648 1848 2712
rect 1912 2648 1928 2712
rect 1992 2648 2008 2712
rect 2072 2648 2088 2712
rect 2152 2648 2168 2712
rect 2232 2648 2248 2712
rect 2312 2648 2328 2712
rect 2392 2648 2408 2712
rect 2472 2648 2488 2712
rect 2552 2648 2568 2712
rect 2632 2648 2648 2712
rect 2712 2648 2728 2712
rect 2792 2648 2808 2712
rect 2872 2648 2888 2712
rect 2952 2648 2968 2712
rect 3032 2648 3048 2712
rect 3112 2648 3128 2712
rect 3192 2648 3208 2712
rect 3272 2648 3288 2712
rect 3352 2648 3368 2712
rect 3432 2648 3448 2712
rect 3512 2648 3528 2712
rect 3592 2648 3608 2712
rect 3672 2648 3688 2712
rect 3752 2648 3768 2712
rect 3832 2648 3848 2712
rect 3912 2648 3928 2712
rect 3992 2648 4000 2712
rect 0 2632 4000 2648
rect 0 2568 8 2632
rect 72 2568 88 2632
rect 152 2568 168 2632
rect 232 2568 248 2632
rect 312 2568 328 2632
rect 392 2568 408 2632
rect 472 2568 488 2632
rect 552 2568 568 2632
rect 632 2568 648 2632
rect 712 2568 728 2632
rect 792 2568 808 2632
rect 872 2568 888 2632
rect 952 2568 968 2632
rect 1032 2568 1048 2632
rect 1112 2568 1128 2632
rect 1192 2568 1208 2632
rect 1272 2568 1288 2632
rect 1352 2568 1368 2632
rect 1432 2568 1448 2632
rect 1512 2568 1528 2632
rect 1592 2568 1608 2632
rect 1672 2568 1688 2632
rect 1752 2568 1768 2632
rect 1832 2568 1848 2632
rect 1912 2568 1928 2632
rect 1992 2568 2008 2632
rect 2072 2568 2088 2632
rect 2152 2568 2168 2632
rect 2232 2568 2248 2632
rect 2312 2568 2328 2632
rect 2392 2568 2408 2632
rect 2472 2568 2488 2632
rect 2552 2568 2568 2632
rect 2632 2568 2648 2632
rect 2712 2568 2728 2632
rect 2792 2568 2808 2632
rect 2872 2568 2888 2632
rect 2952 2568 2968 2632
rect 3032 2568 3048 2632
rect 3112 2568 3128 2632
rect 3192 2568 3208 2632
rect 3272 2568 3288 2632
rect 3352 2568 3368 2632
rect 3432 2568 3448 2632
rect 3512 2568 3528 2632
rect 3592 2568 3608 2632
rect 3672 2568 3688 2632
rect 3752 2568 3768 2632
rect 3832 2568 3848 2632
rect 3912 2568 3928 2632
rect 3992 2568 4000 2632
rect 0 2552 4000 2568
rect 0 2488 8 2552
rect 72 2488 88 2552
rect 152 2488 168 2552
rect 232 2488 248 2552
rect 312 2488 328 2552
rect 392 2488 408 2552
rect 472 2488 488 2552
rect 552 2488 568 2552
rect 632 2488 648 2552
rect 712 2488 728 2552
rect 792 2488 808 2552
rect 872 2488 888 2552
rect 952 2488 968 2552
rect 1032 2488 1048 2552
rect 1112 2488 1128 2552
rect 1192 2488 1208 2552
rect 1272 2488 1288 2552
rect 1352 2488 1368 2552
rect 1432 2488 1448 2552
rect 1512 2488 1528 2552
rect 1592 2488 1608 2552
rect 1672 2488 1688 2552
rect 1752 2488 1768 2552
rect 1832 2488 1848 2552
rect 1912 2488 1928 2552
rect 1992 2488 2008 2552
rect 2072 2488 2088 2552
rect 2152 2488 2168 2552
rect 2232 2488 2248 2552
rect 2312 2488 2328 2552
rect 2392 2488 2408 2552
rect 2472 2488 2488 2552
rect 2552 2488 2568 2552
rect 2632 2488 2648 2552
rect 2712 2488 2728 2552
rect 2792 2488 2808 2552
rect 2872 2488 2888 2552
rect 2952 2488 2968 2552
rect 3032 2488 3048 2552
rect 3112 2488 3128 2552
rect 3192 2488 3208 2552
rect 3272 2488 3288 2552
rect 3352 2488 3368 2552
rect 3432 2488 3448 2552
rect 3512 2488 3528 2552
rect 3592 2488 3608 2552
rect 3672 2488 3688 2552
rect 3752 2488 3768 2552
rect 3832 2488 3848 2552
rect 3912 2488 3928 2552
rect 3992 2488 4000 2552
rect 0 2472 4000 2488
rect 0 2408 8 2472
rect 72 2408 88 2472
rect 152 2408 168 2472
rect 232 2408 248 2472
rect 312 2408 328 2472
rect 392 2408 408 2472
rect 472 2408 488 2472
rect 552 2408 568 2472
rect 632 2408 648 2472
rect 712 2408 728 2472
rect 792 2408 808 2472
rect 872 2408 888 2472
rect 952 2408 968 2472
rect 1032 2408 1048 2472
rect 1112 2408 1128 2472
rect 1192 2408 1208 2472
rect 1272 2408 1288 2472
rect 1352 2408 1368 2472
rect 1432 2408 1448 2472
rect 1512 2408 1528 2472
rect 1592 2408 1608 2472
rect 1672 2408 1688 2472
rect 1752 2408 1768 2472
rect 1832 2408 1848 2472
rect 1912 2408 1928 2472
rect 1992 2408 2008 2472
rect 2072 2408 2088 2472
rect 2152 2408 2168 2472
rect 2232 2408 2248 2472
rect 2312 2408 2328 2472
rect 2392 2408 2408 2472
rect 2472 2408 2488 2472
rect 2552 2408 2568 2472
rect 2632 2408 2648 2472
rect 2712 2408 2728 2472
rect 2792 2408 2808 2472
rect 2872 2408 2888 2472
rect 2952 2408 2968 2472
rect 3032 2408 3048 2472
rect 3112 2408 3128 2472
rect 3192 2408 3208 2472
rect 3272 2408 3288 2472
rect 3352 2408 3368 2472
rect 3432 2408 3448 2472
rect 3512 2408 3528 2472
rect 3592 2408 3608 2472
rect 3672 2408 3688 2472
rect 3752 2408 3768 2472
rect 3832 2408 3848 2472
rect 3912 2408 3928 2472
rect 3992 2408 4000 2472
rect 0 2392 4000 2408
rect 0 2328 8 2392
rect 72 2328 88 2392
rect 152 2328 168 2392
rect 232 2328 248 2392
rect 312 2328 328 2392
rect 392 2328 408 2392
rect 472 2328 488 2392
rect 552 2328 568 2392
rect 632 2328 648 2392
rect 712 2328 728 2392
rect 792 2328 808 2392
rect 872 2328 888 2392
rect 952 2328 968 2392
rect 1032 2328 1048 2392
rect 1112 2328 1128 2392
rect 1192 2328 1208 2392
rect 1272 2328 1288 2392
rect 1352 2328 1368 2392
rect 1432 2328 1448 2392
rect 1512 2328 1528 2392
rect 1592 2328 1608 2392
rect 1672 2328 1688 2392
rect 1752 2328 1768 2392
rect 1832 2328 1848 2392
rect 1912 2328 1928 2392
rect 1992 2328 2008 2392
rect 2072 2328 2088 2392
rect 2152 2328 2168 2392
rect 2232 2328 2248 2392
rect 2312 2328 2328 2392
rect 2392 2328 2408 2392
rect 2472 2328 2488 2392
rect 2552 2328 2568 2392
rect 2632 2328 2648 2392
rect 2712 2328 2728 2392
rect 2792 2328 2808 2392
rect 2872 2328 2888 2392
rect 2952 2328 2968 2392
rect 3032 2328 3048 2392
rect 3112 2328 3128 2392
rect 3192 2328 3208 2392
rect 3272 2328 3288 2392
rect 3352 2328 3368 2392
rect 3432 2328 3448 2392
rect 3512 2328 3528 2392
rect 3592 2328 3608 2392
rect 3672 2328 3688 2392
rect 3752 2328 3768 2392
rect 3832 2328 3848 2392
rect 3912 2328 3928 2392
rect 3992 2328 4000 2392
rect 0 2312 4000 2328
rect 0 2248 8 2312
rect 72 2248 88 2312
rect 152 2248 168 2312
rect 232 2248 248 2312
rect 312 2248 328 2312
rect 392 2248 408 2312
rect 472 2248 488 2312
rect 552 2248 568 2312
rect 632 2248 648 2312
rect 712 2248 728 2312
rect 792 2248 808 2312
rect 872 2248 888 2312
rect 952 2248 968 2312
rect 1032 2248 1048 2312
rect 1112 2248 1128 2312
rect 1192 2248 1208 2312
rect 1272 2248 1288 2312
rect 1352 2248 1368 2312
rect 1432 2248 1448 2312
rect 1512 2248 1528 2312
rect 1592 2248 1608 2312
rect 1672 2248 1688 2312
rect 1752 2248 1768 2312
rect 1832 2248 1848 2312
rect 1912 2248 1928 2312
rect 1992 2248 2008 2312
rect 2072 2248 2088 2312
rect 2152 2248 2168 2312
rect 2232 2248 2248 2312
rect 2312 2248 2328 2312
rect 2392 2248 2408 2312
rect 2472 2248 2488 2312
rect 2552 2248 2568 2312
rect 2632 2248 2648 2312
rect 2712 2248 2728 2312
rect 2792 2248 2808 2312
rect 2872 2248 2888 2312
rect 2952 2248 2968 2312
rect 3032 2248 3048 2312
rect 3112 2248 3128 2312
rect 3192 2248 3208 2312
rect 3272 2248 3288 2312
rect 3352 2248 3368 2312
rect 3432 2248 3448 2312
rect 3512 2248 3528 2312
rect 3592 2248 3608 2312
rect 3672 2248 3688 2312
rect 3752 2248 3768 2312
rect 3832 2248 3848 2312
rect 3912 2248 3928 2312
rect 3992 2248 4000 2312
rect 0 2232 4000 2248
rect 0 2168 8 2232
rect 72 2168 88 2232
rect 152 2168 168 2232
rect 232 2168 248 2232
rect 312 2168 328 2232
rect 392 2168 408 2232
rect 472 2168 488 2232
rect 552 2168 568 2232
rect 632 2168 648 2232
rect 712 2168 728 2232
rect 792 2168 808 2232
rect 872 2168 888 2232
rect 952 2168 968 2232
rect 1032 2168 1048 2232
rect 1112 2168 1128 2232
rect 1192 2168 1208 2232
rect 1272 2168 1288 2232
rect 1352 2168 1368 2232
rect 1432 2168 1448 2232
rect 1512 2168 1528 2232
rect 1592 2168 1608 2232
rect 1672 2168 1688 2232
rect 1752 2168 1768 2232
rect 1832 2168 1848 2232
rect 1912 2168 1928 2232
rect 1992 2168 2008 2232
rect 2072 2168 2088 2232
rect 2152 2168 2168 2232
rect 2232 2168 2248 2232
rect 2312 2168 2328 2232
rect 2392 2168 2408 2232
rect 2472 2168 2488 2232
rect 2552 2168 2568 2232
rect 2632 2168 2648 2232
rect 2712 2168 2728 2232
rect 2792 2168 2808 2232
rect 2872 2168 2888 2232
rect 2952 2168 2968 2232
rect 3032 2168 3048 2232
rect 3112 2168 3128 2232
rect 3192 2168 3208 2232
rect 3272 2168 3288 2232
rect 3352 2168 3368 2232
rect 3432 2168 3448 2232
rect 3512 2168 3528 2232
rect 3592 2168 3608 2232
rect 3672 2168 3688 2232
rect 3752 2168 3768 2232
rect 3832 2168 3848 2232
rect 3912 2168 3928 2232
rect 3992 2168 4000 2232
rect 0 2152 4000 2168
rect 0 2088 8 2152
rect 72 2088 88 2152
rect 152 2088 168 2152
rect 232 2088 248 2152
rect 312 2088 328 2152
rect 392 2088 408 2152
rect 472 2088 488 2152
rect 552 2088 568 2152
rect 632 2088 648 2152
rect 712 2088 728 2152
rect 792 2088 808 2152
rect 872 2088 888 2152
rect 952 2088 968 2152
rect 1032 2088 1048 2152
rect 1112 2088 1128 2152
rect 1192 2088 1208 2152
rect 1272 2088 1288 2152
rect 1352 2088 1368 2152
rect 1432 2088 1448 2152
rect 1512 2088 1528 2152
rect 1592 2088 1608 2152
rect 1672 2088 1688 2152
rect 1752 2088 1768 2152
rect 1832 2088 1848 2152
rect 1912 2088 1928 2152
rect 1992 2088 2008 2152
rect 2072 2088 2088 2152
rect 2152 2088 2168 2152
rect 2232 2088 2248 2152
rect 2312 2088 2328 2152
rect 2392 2088 2408 2152
rect 2472 2088 2488 2152
rect 2552 2088 2568 2152
rect 2632 2088 2648 2152
rect 2712 2088 2728 2152
rect 2792 2088 2808 2152
rect 2872 2088 2888 2152
rect 2952 2088 2968 2152
rect 3032 2088 3048 2152
rect 3112 2088 3128 2152
rect 3192 2088 3208 2152
rect 3272 2088 3288 2152
rect 3352 2088 3368 2152
rect 3432 2088 3448 2152
rect 3512 2088 3528 2152
rect 3592 2088 3608 2152
rect 3672 2088 3688 2152
rect 3752 2088 3768 2152
rect 3832 2088 3848 2152
rect 3912 2088 3928 2152
rect 3992 2088 4000 2152
rect 0 2072 4000 2088
rect 0 2008 8 2072
rect 72 2008 88 2072
rect 152 2008 168 2072
rect 232 2008 248 2072
rect 312 2008 328 2072
rect 392 2008 408 2072
rect 472 2008 488 2072
rect 552 2008 568 2072
rect 632 2008 648 2072
rect 712 2008 728 2072
rect 792 2008 808 2072
rect 872 2008 888 2072
rect 952 2008 968 2072
rect 1032 2008 1048 2072
rect 1112 2008 1128 2072
rect 1192 2008 1208 2072
rect 1272 2008 1288 2072
rect 1352 2008 1368 2072
rect 1432 2008 1448 2072
rect 1512 2008 1528 2072
rect 1592 2008 1608 2072
rect 1672 2008 1688 2072
rect 1752 2008 1768 2072
rect 1832 2008 1848 2072
rect 1912 2008 1928 2072
rect 1992 2008 2008 2072
rect 2072 2008 2088 2072
rect 2152 2008 2168 2072
rect 2232 2008 2248 2072
rect 2312 2008 2328 2072
rect 2392 2008 2408 2072
rect 2472 2008 2488 2072
rect 2552 2008 2568 2072
rect 2632 2008 2648 2072
rect 2712 2008 2728 2072
rect 2792 2008 2808 2072
rect 2872 2008 2888 2072
rect 2952 2008 2968 2072
rect 3032 2008 3048 2072
rect 3112 2008 3128 2072
rect 3192 2008 3208 2072
rect 3272 2008 3288 2072
rect 3352 2008 3368 2072
rect 3432 2008 3448 2072
rect 3512 2008 3528 2072
rect 3592 2008 3608 2072
rect 3672 2008 3688 2072
rect 3752 2008 3768 2072
rect 3832 2008 3848 2072
rect 3912 2008 3928 2072
rect 3992 2008 4000 2072
rect 0 1992 4000 2008
rect 0 1928 8 1992
rect 72 1928 88 1992
rect 152 1928 168 1992
rect 232 1928 248 1992
rect 312 1928 328 1992
rect 392 1928 408 1992
rect 472 1928 488 1992
rect 552 1928 568 1992
rect 632 1928 648 1992
rect 712 1928 728 1992
rect 792 1928 808 1992
rect 872 1928 888 1992
rect 952 1928 968 1992
rect 1032 1928 1048 1992
rect 1112 1928 1128 1992
rect 1192 1928 1208 1992
rect 1272 1928 1288 1992
rect 1352 1928 1368 1992
rect 1432 1928 1448 1992
rect 1512 1928 1528 1992
rect 1592 1928 1608 1992
rect 1672 1928 1688 1992
rect 1752 1928 1768 1992
rect 1832 1928 1848 1992
rect 1912 1928 1928 1992
rect 1992 1928 2008 1992
rect 2072 1928 2088 1992
rect 2152 1928 2168 1992
rect 2232 1928 2248 1992
rect 2312 1928 2328 1992
rect 2392 1928 2408 1992
rect 2472 1928 2488 1992
rect 2552 1928 2568 1992
rect 2632 1928 2648 1992
rect 2712 1928 2728 1992
rect 2792 1928 2808 1992
rect 2872 1928 2888 1992
rect 2952 1928 2968 1992
rect 3032 1928 3048 1992
rect 3112 1928 3128 1992
rect 3192 1928 3208 1992
rect 3272 1928 3288 1992
rect 3352 1928 3368 1992
rect 3432 1928 3448 1992
rect 3512 1928 3528 1992
rect 3592 1928 3608 1992
rect 3672 1928 3688 1992
rect 3752 1928 3768 1992
rect 3832 1928 3848 1992
rect 3912 1928 3928 1992
rect 3992 1928 4000 1992
rect 0 1912 4000 1928
rect 0 1848 8 1912
rect 72 1848 88 1912
rect 152 1848 168 1912
rect 232 1848 248 1912
rect 312 1848 328 1912
rect 392 1848 408 1912
rect 472 1848 488 1912
rect 552 1848 568 1912
rect 632 1848 648 1912
rect 712 1848 728 1912
rect 792 1848 808 1912
rect 872 1848 888 1912
rect 952 1848 968 1912
rect 1032 1848 1048 1912
rect 1112 1848 1128 1912
rect 1192 1848 1208 1912
rect 1272 1848 1288 1912
rect 1352 1848 1368 1912
rect 1432 1848 1448 1912
rect 1512 1848 1528 1912
rect 1592 1848 1608 1912
rect 1672 1848 1688 1912
rect 1752 1848 1768 1912
rect 1832 1848 1848 1912
rect 1912 1848 1928 1912
rect 1992 1848 2008 1912
rect 2072 1848 2088 1912
rect 2152 1848 2168 1912
rect 2232 1848 2248 1912
rect 2312 1848 2328 1912
rect 2392 1848 2408 1912
rect 2472 1848 2488 1912
rect 2552 1848 2568 1912
rect 2632 1848 2648 1912
rect 2712 1848 2728 1912
rect 2792 1848 2808 1912
rect 2872 1848 2888 1912
rect 2952 1848 2968 1912
rect 3032 1848 3048 1912
rect 3112 1848 3128 1912
rect 3192 1848 3208 1912
rect 3272 1848 3288 1912
rect 3352 1848 3368 1912
rect 3432 1848 3448 1912
rect 3512 1848 3528 1912
rect 3592 1848 3608 1912
rect 3672 1848 3688 1912
rect 3752 1848 3768 1912
rect 3832 1848 3848 1912
rect 3912 1848 3928 1912
rect 3992 1848 4000 1912
rect 0 1832 4000 1848
rect 0 1768 8 1832
rect 72 1768 88 1832
rect 152 1768 168 1832
rect 232 1768 248 1832
rect 312 1768 328 1832
rect 392 1768 408 1832
rect 472 1768 488 1832
rect 552 1768 568 1832
rect 632 1768 648 1832
rect 712 1768 728 1832
rect 792 1768 808 1832
rect 872 1768 888 1832
rect 952 1768 968 1832
rect 1032 1768 1048 1832
rect 1112 1768 1128 1832
rect 1192 1768 1208 1832
rect 1272 1768 1288 1832
rect 1352 1768 1368 1832
rect 1432 1768 1448 1832
rect 1512 1768 1528 1832
rect 1592 1768 1608 1832
rect 1672 1768 1688 1832
rect 1752 1768 1768 1832
rect 1832 1768 1848 1832
rect 1912 1768 1928 1832
rect 1992 1768 2008 1832
rect 2072 1768 2088 1832
rect 2152 1768 2168 1832
rect 2232 1768 2248 1832
rect 2312 1768 2328 1832
rect 2392 1768 2408 1832
rect 2472 1768 2488 1832
rect 2552 1768 2568 1832
rect 2632 1768 2648 1832
rect 2712 1768 2728 1832
rect 2792 1768 2808 1832
rect 2872 1768 2888 1832
rect 2952 1768 2968 1832
rect 3032 1768 3048 1832
rect 3112 1768 3128 1832
rect 3192 1768 3208 1832
rect 3272 1768 3288 1832
rect 3352 1768 3368 1832
rect 3432 1768 3448 1832
rect 3512 1768 3528 1832
rect 3592 1768 3608 1832
rect 3672 1768 3688 1832
rect 3752 1768 3768 1832
rect 3832 1768 3848 1832
rect 3912 1768 3928 1832
rect 3992 1768 4000 1832
rect 0 1752 4000 1768
rect 0 1688 8 1752
rect 72 1688 88 1752
rect 152 1688 168 1752
rect 232 1688 248 1752
rect 312 1688 328 1752
rect 392 1688 408 1752
rect 472 1688 488 1752
rect 552 1688 568 1752
rect 632 1688 648 1752
rect 712 1688 728 1752
rect 792 1688 808 1752
rect 872 1688 888 1752
rect 952 1688 968 1752
rect 1032 1688 1048 1752
rect 1112 1688 1128 1752
rect 1192 1688 1208 1752
rect 1272 1688 1288 1752
rect 1352 1688 1368 1752
rect 1432 1688 1448 1752
rect 1512 1688 1528 1752
rect 1592 1688 1608 1752
rect 1672 1688 1688 1752
rect 1752 1688 1768 1752
rect 1832 1688 1848 1752
rect 1912 1688 1928 1752
rect 1992 1688 2008 1752
rect 2072 1688 2088 1752
rect 2152 1688 2168 1752
rect 2232 1688 2248 1752
rect 2312 1688 2328 1752
rect 2392 1688 2408 1752
rect 2472 1688 2488 1752
rect 2552 1688 2568 1752
rect 2632 1688 2648 1752
rect 2712 1688 2728 1752
rect 2792 1688 2808 1752
rect 2872 1688 2888 1752
rect 2952 1688 2968 1752
rect 3032 1688 3048 1752
rect 3112 1688 3128 1752
rect 3192 1688 3208 1752
rect 3272 1688 3288 1752
rect 3352 1688 3368 1752
rect 3432 1688 3448 1752
rect 3512 1688 3528 1752
rect 3592 1688 3608 1752
rect 3672 1688 3688 1752
rect 3752 1688 3768 1752
rect 3832 1688 3848 1752
rect 3912 1688 3928 1752
rect 3992 1688 4000 1752
rect 0 1672 4000 1688
rect 0 1608 8 1672
rect 72 1608 88 1672
rect 152 1608 168 1672
rect 232 1608 248 1672
rect 312 1608 328 1672
rect 392 1608 408 1672
rect 472 1608 488 1672
rect 552 1608 568 1672
rect 632 1608 648 1672
rect 712 1608 728 1672
rect 792 1608 808 1672
rect 872 1608 888 1672
rect 952 1608 968 1672
rect 1032 1608 1048 1672
rect 1112 1608 1128 1672
rect 1192 1608 1208 1672
rect 1272 1608 1288 1672
rect 1352 1608 1368 1672
rect 1432 1608 1448 1672
rect 1512 1608 1528 1672
rect 1592 1608 1608 1672
rect 1672 1608 1688 1672
rect 1752 1608 1768 1672
rect 1832 1608 1848 1672
rect 1912 1608 1928 1672
rect 1992 1608 2008 1672
rect 2072 1608 2088 1672
rect 2152 1608 2168 1672
rect 2232 1608 2248 1672
rect 2312 1608 2328 1672
rect 2392 1608 2408 1672
rect 2472 1608 2488 1672
rect 2552 1608 2568 1672
rect 2632 1608 2648 1672
rect 2712 1608 2728 1672
rect 2792 1608 2808 1672
rect 2872 1608 2888 1672
rect 2952 1608 2968 1672
rect 3032 1608 3048 1672
rect 3112 1608 3128 1672
rect 3192 1608 3208 1672
rect 3272 1608 3288 1672
rect 3352 1608 3368 1672
rect 3432 1608 3448 1672
rect 3512 1608 3528 1672
rect 3592 1608 3608 1672
rect 3672 1608 3688 1672
rect 3752 1608 3768 1672
rect 3832 1608 3848 1672
rect 3912 1608 3928 1672
rect 3992 1608 4000 1672
rect 0 1592 4000 1608
rect 0 1528 8 1592
rect 72 1528 88 1592
rect 152 1528 168 1592
rect 232 1528 248 1592
rect 312 1528 328 1592
rect 392 1528 408 1592
rect 472 1528 488 1592
rect 552 1528 568 1592
rect 632 1528 648 1592
rect 712 1528 728 1592
rect 792 1528 808 1592
rect 872 1528 888 1592
rect 952 1528 968 1592
rect 1032 1528 1048 1592
rect 1112 1528 1128 1592
rect 1192 1528 1208 1592
rect 1272 1528 1288 1592
rect 1352 1528 1368 1592
rect 1432 1528 1448 1592
rect 1512 1528 1528 1592
rect 1592 1528 1608 1592
rect 1672 1528 1688 1592
rect 1752 1528 1768 1592
rect 1832 1528 1848 1592
rect 1912 1528 1928 1592
rect 1992 1528 2008 1592
rect 2072 1528 2088 1592
rect 2152 1528 2168 1592
rect 2232 1528 2248 1592
rect 2312 1528 2328 1592
rect 2392 1528 2408 1592
rect 2472 1528 2488 1592
rect 2552 1528 2568 1592
rect 2632 1528 2648 1592
rect 2712 1528 2728 1592
rect 2792 1528 2808 1592
rect 2872 1528 2888 1592
rect 2952 1528 2968 1592
rect 3032 1528 3048 1592
rect 3112 1528 3128 1592
rect 3192 1528 3208 1592
rect 3272 1528 3288 1592
rect 3352 1528 3368 1592
rect 3432 1528 3448 1592
rect 3512 1528 3528 1592
rect 3592 1528 3608 1592
rect 3672 1528 3688 1592
rect 3752 1528 3768 1592
rect 3832 1528 3848 1592
rect 3912 1528 3928 1592
rect 3992 1528 4000 1592
rect 0 1512 4000 1528
rect 0 1448 8 1512
rect 72 1448 88 1512
rect 152 1448 168 1512
rect 232 1448 248 1512
rect 312 1448 328 1512
rect 392 1448 408 1512
rect 472 1448 488 1512
rect 552 1448 568 1512
rect 632 1448 648 1512
rect 712 1448 728 1512
rect 792 1448 808 1512
rect 872 1448 888 1512
rect 952 1448 968 1512
rect 1032 1448 1048 1512
rect 1112 1448 1128 1512
rect 1192 1448 1208 1512
rect 1272 1448 1288 1512
rect 1352 1448 1368 1512
rect 1432 1448 1448 1512
rect 1512 1448 1528 1512
rect 1592 1448 1608 1512
rect 1672 1448 1688 1512
rect 1752 1448 1768 1512
rect 1832 1448 1848 1512
rect 1912 1448 1928 1512
rect 1992 1448 2008 1512
rect 2072 1448 2088 1512
rect 2152 1448 2168 1512
rect 2232 1448 2248 1512
rect 2312 1448 2328 1512
rect 2392 1448 2408 1512
rect 2472 1448 2488 1512
rect 2552 1448 2568 1512
rect 2632 1448 2648 1512
rect 2712 1448 2728 1512
rect 2792 1448 2808 1512
rect 2872 1448 2888 1512
rect 2952 1448 2968 1512
rect 3032 1448 3048 1512
rect 3112 1448 3128 1512
rect 3192 1448 3208 1512
rect 3272 1448 3288 1512
rect 3352 1448 3368 1512
rect 3432 1448 3448 1512
rect 3512 1448 3528 1512
rect 3592 1448 3608 1512
rect 3672 1448 3688 1512
rect 3752 1448 3768 1512
rect 3832 1448 3848 1512
rect 3912 1448 3928 1512
rect 3992 1448 4000 1512
rect 0 1432 4000 1448
rect 0 1368 8 1432
rect 72 1368 88 1432
rect 152 1368 168 1432
rect 232 1368 248 1432
rect 312 1368 328 1432
rect 392 1368 408 1432
rect 472 1368 488 1432
rect 552 1368 568 1432
rect 632 1368 648 1432
rect 712 1368 728 1432
rect 792 1368 808 1432
rect 872 1368 888 1432
rect 952 1368 968 1432
rect 1032 1368 1048 1432
rect 1112 1368 1128 1432
rect 1192 1368 1208 1432
rect 1272 1368 1288 1432
rect 1352 1368 1368 1432
rect 1432 1368 1448 1432
rect 1512 1368 1528 1432
rect 1592 1368 1608 1432
rect 1672 1368 1688 1432
rect 1752 1368 1768 1432
rect 1832 1368 1848 1432
rect 1912 1368 1928 1432
rect 1992 1368 2008 1432
rect 2072 1368 2088 1432
rect 2152 1368 2168 1432
rect 2232 1368 2248 1432
rect 2312 1368 2328 1432
rect 2392 1368 2408 1432
rect 2472 1368 2488 1432
rect 2552 1368 2568 1432
rect 2632 1368 2648 1432
rect 2712 1368 2728 1432
rect 2792 1368 2808 1432
rect 2872 1368 2888 1432
rect 2952 1368 2968 1432
rect 3032 1368 3048 1432
rect 3112 1368 3128 1432
rect 3192 1368 3208 1432
rect 3272 1368 3288 1432
rect 3352 1368 3368 1432
rect 3432 1368 3448 1432
rect 3512 1368 3528 1432
rect 3592 1368 3608 1432
rect 3672 1368 3688 1432
rect 3752 1368 3768 1432
rect 3832 1368 3848 1432
rect 3912 1368 3928 1432
rect 3992 1368 4000 1432
rect 0 1352 4000 1368
rect 0 1288 8 1352
rect 72 1288 88 1352
rect 152 1288 168 1352
rect 232 1288 248 1352
rect 312 1288 328 1352
rect 392 1288 408 1352
rect 472 1288 488 1352
rect 552 1288 568 1352
rect 632 1288 648 1352
rect 712 1288 728 1352
rect 792 1288 808 1352
rect 872 1288 888 1352
rect 952 1288 968 1352
rect 1032 1288 1048 1352
rect 1112 1288 1128 1352
rect 1192 1288 1208 1352
rect 1272 1288 1288 1352
rect 1352 1288 1368 1352
rect 1432 1288 1448 1352
rect 1512 1288 1528 1352
rect 1592 1288 1608 1352
rect 1672 1288 1688 1352
rect 1752 1288 1768 1352
rect 1832 1288 1848 1352
rect 1912 1288 1928 1352
rect 1992 1288 2008 1352
rect 2072 1288 2088 1352
rect 2152 1288 2168 1352
rect 2232 1288 2248 1352
rect 2312 1288 2328 1352
rect 2392 1288 2408 1352
rect 2472 1288 2488 1352
rect 2552 1288 2568 1352
rect 2632 1288 2648 1352
rect 2712 1288 2728 1352
rect 2792 1288 2808 1352
rect 2872 1288 2888 1352
rect 2952 1288 2968 1352
rect 3032 1288 3048 1352
rect 3112 1288 3128 1352
rect 3192 1288 3208 1352
rect 3272 1288 3288 1352
rect 3352 1288 3368 1352
rect 3432 1288 3448 1352
rect 3512 1288 3528 1352
rect 3592 1288 3608 1352
rect 3672 1288 3688 1352
rect 3752 1288 3768 1352
rect 3832 1288 3848 1352
rect 3912 1288 3928 1352
rect 3992 1288 4000 1352
rect 0 1272 4000 1288
rect 0 1208 8 1272
rect 72 1208 88 1272
rect 152 1208 168 1272
rect 232 1208 248 1272
rect 312 1208 328 1272
rect 392 1208 408 1272
rect 472 1208 488 1272
rect 552 1208 568 1272
rect 632 1208 648 1272
rect 712 1208 728 1272
rect 792 1208 808 1272
rect 872 1208 888 1272
rect 952 1208 968 1272
rect 1032 1208 1048 1272
rect 1112 1208 1128 1272
rect 1192 1208 1208 1272
rect 1272 1208 1288 1272
rect 1352 1208 1368 1272
rect 1432 1208 1448 1272
rect 1512 1208 1528 1272
rect 1592 1208 1608 1272
rect 1672 1208 1688 1272
rect 1752 1208 1768 1272
rect 1832 1208 1848 1272
rect 1912 1208 1928 1272
rect 1992 1208 2008 1272
rect 2072 1208 2088 1272
rect 2152 1208 2168 1272
rect 2232 1208 2248 1272
rect 2312 1208 2328 1272
rect 2392 1208 2408 1272
rect 2472 1208 2488 1272
rect 2552 1208 2568 1272
rect 2632 1208 2648 1272
rect 2712 1208 2728 1272
rect 2792 1208 2808 1272
rect 2872 1208 2888 1272
rect 2952 1208 2968 1272
rect 3032 1208 3048 1272
rect 3112 1208 3128 1272
rect 3192 1208 3208 1272
rect 3272 1208 3288 1272
rect 3352 1208 3368 1272
rect 3432 1208 3448 1272
rect 3512 1208 3528 1272
rect 3592 1208 3608 1272
rect 3672 1208 3688 1272
rect 3752 1208 3768 1272
rect 3832 1208 3848 1272
rect 3912 1208 3928 1272
rect 3992 1208 4000 1272
rect 0 1192 4000 1208
rect 0 1128 8 1192
rect 72 1128 88 1192
rect 152 1128 168 1192
rect 232 1128 248 1192
rect 312 1128 328 1192
rect 392 1128 408 1192
rect 472 1128 488 1192
rect 552 1128 568 1192
rect 632 1128 648 1192
rect 712 1128 728 1192
rect 792 1128 808 1192
rect 872 1128 888 1192
rect 952 1128 968 1192
rect 1032 1128 1048 1192
rect 1112 1128 1128 1192
rect 1192 1128 1208 1192
rect 1272 1128 1288 1192
rect 1352 1128 1368 1192
rect 1432 1128 1448 1192
rect 1512 1128 1528 1192
rect 1592 1128 1608 1192
rect 1672 1128 1688 1192
rect 1752 1128 1768 1192
rect 1832 1128 1848 1192
rect 1912 1128 1928 1192
rect 1992 1128 2008 1192
rect 2072 1128 2088 1192
rect 2152 1128 2168 1192
rect 2232 1128 2248 1192
rect 2312 1128 2328 1192
rect 2392 1128 2408 1192
rect 2472 1128 2488 1192
rect 2552 1128 2568 1192
rect 2632 1128 2648 1192
rect 2712 1128 2728 1192
rect 2792 1128 2808 1192
rect 2872 1128 2888 1192
rect 2952 1128 2968 1192
rect 3032 1128 3048 1192
rect 3112 1128 3128 1192
rect 3192 1128 3208 1192
rect 3272 1128 3288 1192
rect 3352 1128 3368 1192
rect 3432 1128 3448 1192
rect 3512 1128 3528 1192
rect 3592 1128 3608 1192
rect 3672 1128 3688 1192
rect 3752 1128 3768 1192
rect 3832 1128 3848 1192
rect 3912 1128 3928 1192
rect 3992 1128 4000 1192
rect 0 1112 4000 1128
rect 0 1048 8 1112
rect 72 1048 88 1112
rect 152 1048 168 1112
rect 232 1048 248 1112
rect 312 1048 328 1112
rect 392 1048 408 1112
rect 472 1048 488 1112
rect 552 1048 568 1112
rect 632 1048 648 1112
rect 712 1048 728 1112
rect 792 1048 808 1112
rect 872 1048 888 1112
rect 952 1048 968 1112
rect 1032 1048 1048 1112
rect 1112 1048 1128 1112
rect 1192 1048 1208 1112
rect 1272 1048 1288 1112
rect 1352 1048 1368 1112
rect 1432 1048 1448 1112
rect 1512 1048 1528 1112
rect 1592 1048 1608 1112
rect 1672 1048 1688 1112
rect 1752 1048 1768 1112
rect 1832 1048 1848 1112
rect 1912 1048 1928 1112
rect 1992 1048 2008 1112
rect 2072 1048 2088 1112
rect 2152 1048 2168 1112
rect 2232 1048 2248 1112
rect 2312 1048 2328 1112
rect 2392 1048 2408 1112
rect 2472 1048 2488 1112
rect 2552 1048 2568 1112
rect 2632 1048 2648 1112
rect 2712 1048 2728 1112
rect 2792 1048 2808 1112
rect 2872 1048 2888 1112
rect 2952 1048 2968 1112
rect 3032 1048 3048 1112
rect 3112 1048 3128 1112
rect 3192 1048 3208 1112
rect 3272 1048 3288 1112
rect 3352 1048 3368 1112
rect 3432 1048 3448 1112
rect 3512 1048 3528 1112
rect 3592 1048 3608 1112
rect 3672 1048 3688 1112
rect 3752 1048 3768 1112
rect 3832 1048 3848 1112
rect 3912 1048 3928 1112
rect 3992 1048 4000 1112
rect 0 1032 4000 1048
rect 0 968 8 1032
rect 72 968 88 1032
rect 152 968 168 1032
rect 232 968 248 1032
rect 312 968 328 1032
rect 392 968 408 1032
rect 472 968 488 1032
rect 552 968 568 1032
rect 632 968 648 1032
rect 712 968 728 1032
rect 792 968 808 1032
rect 872 968 888 1032
rect 952 968 968 1032
rect 1032 968 1048 1032
rect 1112 968 1128 1032
rect 1192 968 1208 1032
rect 1272 968 1288 1032
rect 1352 968 1368 1032
rect 1432 968 1448 1032
rect 1512 968 1528 1032
rect 1592 968 1608 1032
rect 1672 968 1688 1032
rect 1752 968 1768 1032
rect 1832 968 1848 1032
rect 1912 968 1928 1032
rect 1992 968 2008 1032
rect 2072 968 2088 1032
rect 2152 968 2168 1032
rect 2232 968 2248 1032
rect 2312 968 2328 1032
rect 2392 968 2408 1032
rect 2472 968 2488 1032
rect 2552 968 2568 1032
rect 2632 968 2648 1032
rect 2712 968 2728 1032
rect 2792 968 2808 1032
rect 2872 968 2888 1032
rect 2952 968 2968 1032
rect 3032 968 3048 1032
rect 3112 968 3128 1032
rect 3192 968 3208 1032
rect 3272 968 3288 1032
rect 3352 968 3368 1032
rect 3432 968 3448 1032
rect 3512 968 3528 1032
rect 3592 968 3608 1032
rect 3672 968 3688 1032
rect 3752 968 3768 1032
rect 3832 968 3848 1032
rect 3912 968 3928 1032
rect 3992 968 4000 1032
rect 0 952 4000 968
rect 0 888 8 952
rect 72 888 88 952
rect 152 888 168 952
rect 232 888 248 952
rect 312 888 328 952
rect 392 888 408 952
rect 472 888 488 952
rect 552 888 568 952
rect 632 888 648 952
rect 712 888 728 952
rect 792 888 808 952
rect 872 888 888 952
rect 952 888 968 952
rect 1032 888 1048 952
rect 1112 888 1128 952
rect 1192 888 1208 952
rect 1272 888 1288 952
rect 1352 888 1368 952
rect 1432 888 1448 952
rect 1512 888 1528 952
rect 1592 888 1608 952
rect 1672 888 1688 952
rect 1752 888 1768 952
rect 1832 888 1848 952
rect 1912 888 1928 952
rect 1992 888 2008 952
rect 2072 888 2088 952
rect 2152 888 2168 952
rect 2232 888 2248 952
rect 2312 888 2328 952
rect 2392 888 2408 952
rect 2472 888 2488 952
rect 2552 888 2568 952
rect 2632 888 2648 952
rect 2712 888 2728 952
rect 2792 888 2808 952
rect 2872 888 2888 952
rect 2952 888 2968 952
rect 3032 888 3048 952
rect 3112 888 3128 952
rect 3192 888 3208 952
rect 3272 888 3288 952
rect 3352 888 3368 952
rect 3432 888 3448 952
rect 3512 888 3528 952
rect 3592 888 3608 952
rect 3672 888 3688 952
rect 3752 888 3768 952
rect 3832 888 3848 952
rect 3912 888 3928 952
rect 3992 888 4000 952
rect 0 872 4000 888
rect 0 808 8 872
rect 72 808 88 872
rect 152 808 168 872
rect 232 808 248 872
rect 312 808 328 872
rect 392 808 408 872
rect 472 808 488 872
rect 552 808 568 872
rect 632 808 648 872
rect 712 808 728 872
rect 792 808 808 872
rect 872 808 888 872
rect 952 808 968 872
rect 1032 808 1048 872
rect 1112 808 1128 872
rect 1192 808 1208 872
rect 1272 808 1288 872
rect 1352 808 1368 872
rect 1432 808 1448 872
rect 1512 808 1528 872
rect 1592 808 1608 872
rect 1672 808 1688 872
rect 1752 808 1768 872
rect 1832 808 1848 872
rect 1912 808 1928 872
rect 1992 808 2008 872
rect 2072 808 2088 872
rect 2152 808 2168 872
rect 2232 808 2248 872
rect 2312 808 2328 872
rect 2392 808 2408 872
rect 2472 808 2488 872
rect 2552 808 2568 872
rect 2632 808 2648 872
rect 2712 808 2728 872
rect 2792 808 2808 872
rect 2872 808 2888 872
rect 2952 808 2968 872
rect 3032 808 3048 872
rect 3112 808 3128 872
rect 3192 808 3208 872
rect 3272 808 3288 872
rect 3352 808 3368 872
rect 3432 808 3448 872
rect 3512 808 3528 872
rect 3592 808 3608 872
rect 3672 808 3688 872
rect 3752 808 3768 872
rect 3832 808 3848 872
rect 3912 808 3928 872
rect 3992 808 4000 872
rect 0 792 4000 808
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 808 792
rect 872 728 888 792
rect 952 728 968 792
rect 1032 728 1048 792
rect 1112 728 1128 792
rect 1192 728 1208 792
rect 1272 728 1288 792
rect 1352 728 1368 792
rect 1432 728 1448 792
rect 1512 728 1528 792
rect 1592 728 1608 792
rect 1672 728 1688 792
rect 1752 728 1768 792
rect 1832 728 1848 792
rect 1912 728 1928 792
rect 1992 728 2008 792
rect 2072 728 2088 792
rect 2152 728 2168 792
rect 2232 728 2248 792
rect 2312 728 2328 792
rect 2392 728 2408 792
rect 2472 728 2488 792
rect 2552 728 2568 792
rect 2632 728 2648 792
rect 2712 728 2728 792
rect 2792 728 2808 792
rect 2872 728 2888 792
rect 2952 728 2968 792
rect 3032 728 3048 792
rect 3112 728 3128 792
rect 3192 728 3208 792
rect 3272 728 3288 792
rect 3352 728 3368 792
rect 3432 728 3448 792
rect 3512 728 3528 792
rect 3592 728 3608 792
rect 3672 728 3688 792
rect 3752 728 3768 792
rect 3832 728 3848 792
rect 3912 728 3928 792
rect 3992 728 4000 792
rect 0 712 4000 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 808 712
rect 872 648 888 712
rect 952 648 968 712
rect 1032 648 1048 712
rect 1112 648 1128 712
rect 1192 648 1208 712
rect 1272 648 1288 712
rect 1352 648 1368 712
rect 1432 648 1448 712
rect 1512 648 1528 712
rect 1592 648 1608 712
rect 1672 648 1688 712
rect 1752 648 1768 712
rect 1832 648 1848 712
rect 1912 648 1928 712
rect 1992 648 2008 712
rect 2072 648 2088 712
rect 2152 648 2168 712
rect 2232 648 2248 712
rect 2312 648 2328 712
rect 2392 648 2408 712
rect 2472 648 2488 712
rect 2552 648 2568 712
rect 2632 648 2648 712
rect 2712 648 2728 712
rect 2792 648 2808 712
rect 2872 648 2888 712
rect 2952 648 2968 712
rect 3032 648 3048 712
rect 3112 648 3128 712
rect 3192 648 3208 712
rect 3272 648 3288 712
rect 3352 648 3368 712
rect 3432 648 3448 712
rect 3512 648 3528 712
rect 3592 648 3608 712
rect 3672 648 3688 712
rect 3752 648 3768 712
rect 3832 648 3848 712
rect 3912 648 3928 712
rect 3992 648 4000 712
rect 0 632 4000 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 808 632
rect 872 568 888 632
rect 952 568 968 632
rect 1032 568 1048 632
rect 1112 568 1128 632
rect 1192 568 1208 632
rect 1272 568 1288 632
rect 1352 568 1368 632
rect 1432 568 1448 632
rect 1512 568 1528 632
rect 1592 568 1608 632
rect 1672 568 1688 632
rect 1752 568 1768 632
rect 1832 568 1848 632
rect 1912 568 1928 632
rect 1992 568 2008 632
rect 2072 568 2088 632
rect 2152 568 2168 632
rect 2232 568 2248 632
rect 2312 568 2328 632
rect 2392 568 2408 632
rect 2472 568 2488 632
rect 2552 568 2568 632
rect 2632 568 2648 632
rect 2712 568 2728 632
rect 2792 568 2808 632
rect 2872 568 2888 632
rect 2952 568 2968 632
rect 3032 568 3048 632
rect 3112 568 3128 632
rect 3192 568 3208 632
rect 3272 568 3288 632
rect 3352 568 3368 632
rect 3432 568 3448 632
rect 3512 568 3528 632
rect 3592 568 3608 632
rect 3672 568 3688 632
rect 3752 568 3768 632
rect 3832 568 3848 632
rect 3912 568 3928 632
rect 3992 568 4000 632
rect 0 552 4000 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 808 552
rect 872 488 888 552
rect 952 488 968 552
rect 1032 488 1048 552
rect 1112 488 1128 552
rect 1192 488 1208 552
rect 1272 488 1288 552
rect 1352 488 1368 552
rect 1432 488 1448 552
rect 1512 488 1528 552
rect 1592 488 1608 552
rect 1672 488 1688 552
rect 1752 488 1768 552
rect 1832 488 1848 552
rect 1912 488 1928 552
rect 1992 488 2008 552
rect 2072 488 2088 552
rect 2152 488 2168 552
rect 2232 488 2248 552
rect 2312 488 2328 552
rect 2392 488 2408 552
rect 2472 488 2488 552
rect 2552 488 2568 552
rect 2632 488 2648 552
rect 2712 488 2728 552
rect 2792 488 2808 552
rect 2872 488 2888 552
rect 2952 488 2968 552
rect 3032 488 3048 552
rect 3112 488 3128 552
rect 3192 488 3208 552
rect 3272 488 3288 552
rect 3352 488 3368 552
rect 3432 488 3448 552
rect 3512 488 3528 552
rect 3592 488 3608 552
rect 3672 488 3688 552
rect 3752 488 3768 552
rect 3832 488 3848 552
rect 3912 488 3928 552
rect 3992 488 4000 552
rect 0 472 4000 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 808 472
rect 872 408 888 472
rect 952 408 968 472
rect 1032 408 1048 472
rect 1112 408 1128 472
rect 1192 408 1208 472
rect 1272 408 1288 472
rect 1352 408 1368 472
rect 1432 408 1448 472
rect 1512 408 1528 472
rect 1592 408 1608 472
rect 1672 408 1688 472
rect 1752 408 1768 472
rect 1832 408 1848 472
rect 1912 408 1928 472
rect 1992 408 2008 472
rect 2072 408 2088 472
rect 2152 408 2168 472
rect 2232 408 2248 472
rect 2312 408 2328 472
rect 2392 408 2408 472
rect 2472 408 2488 472
rect 2552 408 2568 472
rect 2632 408 2648 472
rect 2712 408 2728 472
rect 2792 408 2808 472
rect 2872 408 2888 472
rect 2952 408 2968 472
rect 3032 408 3048 472
rect 3112 408 3128 472
rect 3192 408 3208 472
rect 3272 408 3288 472
rect 3352 408 3368 472
rect 3432 408 3448 472
rect 3512 408 3528 472
rect 3592 408 3608 472
rect 3672 408 3688 472
rect 3752 408 3768 472
rect 3832 408 3848 472
rect 3912 408 3928 472
rect 3992 408 4000 472
rect 0 392 4000 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 808 392
rect 872 328 888 392
rect 952 328 968 392
rect 1032 328 1048 392
rect 1112 328 1128 392
rect 1192 328 1208 392
rect 1272 328 1288 392
rect 1352 328 1368 392
rect 1432 328 1448 392
rect 1512 328 1528 392
rect 1592 328 1608 392
rect 1672 328 1688 392
rect 1752 328 1768 392
rect 1832 328 1848 392
rect 1912 328 1928 392
rect 1992 328 2008 392
rect 2072 328 2088 392
rect 2152 328 2168 392
rect 2232 328 2248 392
rect 2312 328 2328 392
rect 2392 328 2408 392
rect 2472 328 2488 392
rect 2552 328 2568 392
rect 2632 328 2648 392
rect 2712 328 2728 392
rect 2792 328 2808 392
rect 2872 328 2888 392
rect 2952 328 2968 392
rect 3032 328 3048 392
rect 3112 328 3128 392
rect 3192 328 3208 392
rect 3272 328 3288 392
rect 3352 328 3368 392
rect 3432 328 3448 392
rect 3512 328 3528 392
rect 3592 328 3608 392
rect 3672 328 3688 392
rect 3752 328 3768 392
rect 3832 328 3848 392
rect 3912 328 3928 392
rect 3992 328 4000 392
rect 0 312 4000 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 808 312
rect 872 248 888 312
rect 952 248 968 312
rect 1032 248 1048 312
rect 1112 248 1128 312
rect 1192 248 1208 312
rect 1272 248 1288 312
rect 1352 248 1368 312
rect 1432 248 1448 312
rect 1512 248 1528 312
rect 1592 248 1608 312
rect 1672 248 1688 312
rect 1752 248 1768 312
rect 1832 248 1848 312
rect 1912 248 1928 312
rect 1992 248 2008 312
rect 2072 248 2088 312
rect 2152 248 2168 312
rect 2232 248 2248 312
rect 2312 248 2328 312
rect 2392 248 2408 312
rect 2472 248 2488 312
rect 2552 248 2568 312
rect 2632 248 2648 312
rect 2712 248 2728 312
rect 2792 248 2808 312
rect 2872 248 2888 312
rect 2952 248 2968 312
rect 3032 248 3048 312
rect 3112 248 3128 312
rect 3192 248 3208 312
rect 3272 248 3288 312
rect 3352 248 3368 312
rect 3432 248 3448 312
rect 3512 248 3528 312
rect 3592 248 3608 312
rect 3672 248 3688 312
rect 3752 248 3768 312
rect 3832 248 3848 312
rect 3912 248 3928 312
rect 3992 248 4000 312
rect 0 232 4000 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 808 232
rect 872 168 888 232
rect 952 168 968 232
rect 1032 168 1048 232
rect 1112 168 1128 232
rect 1192 168 1208 232
rect 1272 168 1288 232
rect 1352 168 1368 232
rect 1432 168 1448 232
rect 1512 168 1528 232
rect 1592 168 1608 232
rect 1672 168 1688 232
rect 1752 168 1768 232
rect 1832 168 1848 232
rect 1912 168 1928 232
rect 1992 168 2008 232
rect 2072 168 2088 232
rect 2152 168 2168 232
rect 2232 168 2248 232
rect 2312 168 2328 232
rect 2392 168 2408 232
rect 2472 168 2488 232
rect 2552 168 2568 232
rect 2632 168 2648 232
rect 2712 168 2728 232
rect 2792 168 2808 232
rect 2872 168 2888 232
rect 2952 168 2968 232
rect 3032 168 3048 232
rect 3112 168 3128 232
rect 3192 168 3208 232
rect 3272 168 3288 232
rect 3352 168 3368 232
rect 3432 168 3448 232
rect 3512 168 3528 232
rect 3592 168 3608 232
rect 3672 168 3688 232
rect 3752 168 3768 232
rect 3832 168 3848 232
rect 3912 168 3928 232
rect 3992 168 4000 232
rect 0 152 4000 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 808 152
rect 872 88 888 152
rect 952 88 968 152
rect 1032 88 1048 152
rect 1112 88 1128 152
rect 1192 88 1208 152
rect 1272 88 1288 152
rect 1352 88 1368 152
rect 1432 88 1448 152
rect 1512 88 1528 152
rect 1592 88 1608 152
rect 1672 88 1688 152
rect 1752 88 1768 152
rect 1832 88 1848 152
rect 1912 88 1928 152
rect 1992 88 2008 152
rect 2072 88 2088 152
rect 2152 88 2168 152
rect 2232 88 2248 152
rect 2312 88 2328 152
rect 2392 88 2408 152
rect 2472 88 2488 152
rect 2552 88 2568 152
rect 2632 88 2648 152
rect 2712 88 2728 152
rect 2792 88 2808 152
rect 2872 88 2888 152
rect 2952 88 2968 152
rect 3032 88 3048 152
rect 3112 88 3128 152
rect 3192 88 3208 152
rect 3272 88 3288 152
rect 3352 88 3368 152
rect 3432 88 3448 152
rect 3512 88 3528 152
rect 3592 88 3608 152
rect 3672 88 3688 152
rect 3752 88 3768 152
rect 3832 88 3848 152
rect 3912 88 3928 152
rect 3992 88 4000 152
rect 0 72 4000 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 808 72
rect 872 8 888 72
rect 952 8 968 72
rect 1032 8 1048 72
rect 1112 8 1128 72
rect 1192 8 1208 72
rect 1272 8 1288 72
rect 1352 8 1368 72
rect 1432 8 1448 72
rect 1512 8 1528 72
rect 1592 8 1608 72
rect 1672 8 1688 72
rect 1752 8 1768 72
rect 1832 8 1848 72
rect 1912 8 1928 72
rect 1992 8 2008 72
rect 2072 8 2088 72
rect 2152 8 2168 72
rect 2232 8 2248 72
rect 2312 8 2328 72
rect 2392 8 2408 72
rect 2472 8 2488 72
rect 2552 8 2568 72
rect 2632 8 2648 72
rect 2712 8 2728 72
rect 2792 8 2808 72
rect 2872 8 2888 72
rect 2952 8 2968 72
rect 3032 8 3048 72
rect 3112 8 3128 72
rect 3192 8 3208 72
rect 3272 8 3288 72
rect 3352 8 3368 72
rect 3432 8 3448 72
rect 3512 8 3528 72
rect 3592 8 3608 72
rect 3672 8 3688 72
rect 3752 8 3768 72
rect 3832 8 3848 72
rect 3912 8 3928 72
rect 3992 8 4000 72
rect 0 0 4000 8
rect 14104 0 14424 5008
rect 19104 45384 19424 45392
rect 19104 45320 19112 45384
rect 19176 45320 19192 45384
rect 19256 45320 19272 45384
rect 19336 45320 19352 45384
rect 19416 45320 19424 45384
rect 19104 45304 19424 45320
rect 19104 45240 19112 45304
rect 19176 45240 19192 45304
rect 19256 45240 19272 45304
rect 19336 45240 19352 45304
rect 19416 45240 19424 45304
rect 19104 45224 19424 45240
rect 19104 45160 19112 45224
rect 19176 45160 19192 45224
rect 19256 45160 19272 45224
rect 19336 45160 19352 45224
rect 19416 45160 19424 45224
rect 19104 45144 19424 45160
rect 19104 45080 19112 45144
rect 19176 45080 19192 45144
rect 19256 45080 19272 45144
rect 19336 45080 19352 45144
rect 19416 45080 19424 45144
rect 19104 45064 19424 45080
rect 19104 45000 19112 45064
rect 19176 45000 19192 45064
rect 19256 45000 19272 45064
rect 19336 45000 19352 45064
rect 19416 45000 19424 45064
rect 19104 44984 19424 45000
rect 19104 44920 19112 44984
rect 19176 44920 19192 44984
rect 19256 44920 19272 44984
rect 19336 44920 19352 44984
rect 19416 44920 19424 44984
rect 19104 44904 19424 44920
rect 19104 44840 19112 44904
rect 19176 44840 19192 44904
rect 19256 44840 19272 44904
rect 19336 44840 19352 44904
rect 19416 44840 19424 44904
rect 19104 44824 19424 44840
rect 19104 44760 19112 44824
rect 19176 44760 19192 44824
rect 19256 44760 19272 44824
rect 19336 44760 19352 44824
rect 19416 44760 19424 44824
rect 19104 44744 19424 44760
rect 19104 44680 19112 44744
rect 19176 44680 19192 44744
rect 19256 44680 19272 44744
rect 19336 44680 19352 44744
rect 19416 44680 19424 44744
rect 19104 44664 19424 44680
rect 19104 44600 19112 44664
rect 19176 44600 19192 44664
rect 19256 44600 19272 44664
rect 19336 44600 19352 44664
rect 19416 44600 19424 44664
rect 19104 44584 19424 44600
rect 19104 44520 19112 44584
rect 19176 44520 19192 44584
rect 19256 44520 19272 44584
rect 19336 44520 19352 44584
rect 19416 44520 19424 44584
rect 19104 44504 19424 44520
rect 19104 44440 19112 44504
rect 19176 44440 19192 44504
rect 19256 44440 19272 44504
rect 19336 44440 19352 44504
rect 19416 44440 19424 44504
rect 19104 44424 19424 44440
rect 19104 44360 19112 44424
rect 19176 44360 19192 44424
rect 19256 44360 19272 44424
rect 19336 44360 19352 44424
rect 19416 44360 19424 44424
rect 19104 44344 19424 44360
rect 19104 44280 19112 44344
rect 19176 44280 19192 44344
rect 19256 44280 19272 44344
rect 19336 44280 19352 44344
rect 19416 44280 19424 44344
rect 19104 44264 19424 44280
rect 19104 44200 19112 44264
rect 19176 44200 19192 44264
rect 19256 44200 19272 44264
rect 19336 44200 19352 44264
rect 19416 44200 19424 44264
rect 19104 44184 19424 44200
rect 19104 44120 19112 44184
rect 19176 44120 19192 44184
rect 19256 44120 19272 44184
rect 19336 44120 19352 44184
rect 19416 44120 19424 44184
rect 19104 44104 19424 44120
rect 19104 44040 19112 44104
rect 19176 44040 19192 44104
rect 19256 44040 19272 44104
rect 19336 44040 19352 44104
rect 19416 44040 19424 44104
rect 19104 44024 19424 44040
rect 19104 43960 19112 44024
rect 19176 43960 19192 44024
rect 19256 43960 19272 44024
rect 19336 43960 19352 44024
rect 19416 43960 19424 44024
rect 19104 43944 19424 43960
rect 19104 43880 19112 43944
rect 19176 43880 19192 43944
rect 19256 43880 19272 43944
rect 19336 43880 19352 43944
rect 19416 43880 19424 43944
rect 19104 43864 19424 43880
rect 19104 43800 19112 43864
rect 19176 43800 19192 43864
rect 19256 43800 19272 43864
rect 19336 43800 19352 43864
rect 19416 43800 19424 43864
rect 19104 43784 19424 43800
rect 19104 43720 19112 43784
rect 19176 43720 19192 43784
rect 19256 43720 19272 43784
rect 19336 43720 19352 43784
rect 19416 43720 19424 43784
rect 19104 43704 19424 43720
rect 19104 43640 19112 43704
rect 19176 43640 19192 43704
rect 19256 43640 19272 43704
rect 19336 43640 19352 43704
rect 19416 43640 19424 43704
rect 19104 43624 19424 43640
rect 19104 43560 19112 43624
rect 19176 43560 19192 43624
rect 19256 43560 19272 43624
rect 19336 43560 19352 43624
rect 19416 43560 19424 43624
rect 19104 43544 19424 43560
rect 19104 43480 19112 43544
rect 19176 43480 19192 43544
rect 19256 43480 19272 43544
rect 19336 43480 19352 43544
rect 19416 43480 19424 43544
rect 19104 43464 19424 43480
rect 19104 43400 19112 43464
rect 19176 43400 19192 43464
rect 19256 43400 19272 43464
rect 19336 43400 19352 43464
rect 19416 43400 19424 43464
rect 19104 43384 19424 43400
rect 19104 43320 19112 43384
rect 19176 43320 19192 43384
rect 19256 43320 19272 43384
rect 19336 43320 19352 43384
rect 19416 43320 19424 43384
rect 19104 43304 19424 43320
rect 19104 43240 19112 43304
rect 19176 43240 19192 43304
rect 19256 43240 19272 43304
rect 19336 43240 19352 43304
rect 19416 43240 19424 43304
rect 19104 43224 19424 43240
rect 19104 43160 19112 43224
rect 19176 43160 19192 43224
rect 19256 43160 19272 43224
rect 19336 43160 19352 43224
rect 19416 43160 19424 43224
rect 19104 43144 19424 43160
rect 19104 43080 19112 43144
rect 19176 43080 19192 43144
rect 19256 43080 19272 43144
rect 19336 43080 19352 43144
rect 19416 43080 19424 43144
rect 19104 43064 19424 43080
rect 19104 43000 19112 43064
rect 19176 43000 19192 43064
rect 19256 43000 19272 43064
rect 19336 43000 19352 43064
rect 19416 43000 19424 43064
rect 19104 42984 19424 43000
rect 19104 42920 19112 42984
rect 19176 42920 19192 42984
rect 19256 42920 19272 42984
rect 19336 42920 19352 42984
rect 19416 42920 19424 42984
rect 19104 42904 19424 42920
rect 19104 42840 19112 42904
rect 19176 42840 19192 42904
rect 19256 42840 19272 42904
rect 19336 42840 19352 42904
rect 19416 42840 19424 42904
rect 19104 42824 19424 42840
rect 19104 42760 19112 42824
rect 19176 42760 19192 42824
rect 19256 42760 19272 42824
rect 19336 42760 19352 42824
rect 19416 42760 19424 42824
rect 19104 42744 19424 42760
rect 19104 42680 19112 42744
rect 19176 42680 19192 42744
rect 19256 42680 19272 42744
rect 19336 42680 19352 42744
rect 19416 42680 19424 42744
rect 19104 42664 19424 42680
rect 19104 42600 19112 42664
rect 19176 42600 19192 42664
rect 19256 42600 19272 42664
rect 19336 42600 19352 42664
rect 19416 42600 19424 42664
rect 19104 42584 19424 42600
rect 19104 42520 19112 42584
rect 19176 42520 19192 42584
rect 19256 42520 19272 42584
rect 19336 42520 19352 42584
rect 19416 42520 19424 42584
rect 19104 42504 19424 42520
rect 19104 42440 19112 42504
rect 19176 42440 19192 42504
rect 19256 42440 19272 42504
rect 19336 42440 19352 42504
rect 19416 42440 19424 42504
rect 19104 42424 19424 42440
rect 19104 42360 19112 42424
rect 19176 42360 19192 42424
rect 19256 42360 19272 42424
rect 19336 42360 19352 42424
rect 19416 42360 19424 42424
rect 19104 42344 19424 42360
rect 19104 42280 19112 42344
rect 19176 42280 19192 42344
rect 19256 42280 19272 42344
rect 19336 42280 19352 42344
rect 19416 42280 19424 42344
rect 19104 42264 19424 42280
rect 19104 42200 19112 42264
rect 19176 42200 19192 42264
rect 19256 42200 19272 42264
rect 19336 42200 19352 42264
rect 19416 42200 19424 42264
rect 19104 42184 19424 42200
rect 19104 42120 19112 42184
rect 19176 42120 19192 42184
rect 19256 42120 19272 42184
rect 19336 42120 19352 42184
rect 19416 42120 19424 42184
rect 19104 42104 19424 42120
rect 19104 42040 19112 42104
rect 19176 42040 19192 42104
rect 19256 42040 19272 42104
rect 19336 42040 19352 42104
rect 19416 42040 19424 42104
rect 19104 42024 19424 42040
rect 19104 41960 19112 42024
rect 19176 41960 19192 42024
rect 19256 41960 19272 42024
rect 19336 41960 19352 42024
rect 19416 41960 19424 42024
rect 19104 41944 19424 41960
rect 19104 41880 19112 41944
rect 19176 41880 19192 41944
rect 19256 41880 19272 41944
rect 19336 41880 19352 41944
rect 19416 41880 19424 41944
rect 19104 41864 19424 41880
rect 19104 41800 19112 41864
rect 19176 41800 19192 41864
rect 19256 41800 19272 41864
rect 19336 41800 19352 41864
rect 19416 41800 19424 41864
rect 19104 41784 19424 41800
rect 19104 41720 19112 41784
rect 19176 41720 19192 41784
rect 19256 41720 19272 41784
rect 19336 41720 19352 41784
rect 19416 41720 19424 41784
rect 19104 41704 19424 41720
rect 19104 41640 19112 41704
rect 19176 41640 19192 41704
rect 19256 41640 19272 41704
rect 19336 41640 19352 41704
rect 19416 41640 19424 41704
rect 19104 41624 19424 41640
rect 19104 41560 19112 41624
rect 19176 41560 19192 41624
rect 19256 41560 19272 41624
rect 19336 41560 19352 41624
rect 19416 41560 19424 41624
rect 19104 41544 19424 41560
rect 19104 41480 19112 41544
rect 19176 41480 19192 41544
rect 19256 41480 19272 41544
rect 19336 41480 19352 41544
rect 19416 41480 19424 41544
rect 19104 41464 19424 41480
rect 19104 41400 19112 41464
rect 19176 41400 19192 41464
rect 19256 41400 19272 41464
rect 19336 41400 19352 41464
rect 19416 41400 19424 41464
rect 19104 34424 19424 41400
rect 19104 34360 19112 34424
rect 19176 34360 19192 34424
rect 19256 34360 19272 34424
rect 19336 34360 19352 34424
rect 19416 34360 19424 34424
rect 19104 33336 19424 34360
rect 19104 33272 19112 33336
rect 19176 33272 19192 33336
rect 19256 33272 19272 33336
rect 19336 33272 19352 33336
rect 19416 33272 19424 33336
rect 19104 32248 19424 33272
rect 19104 32184 19112 32248
rect 19176 32184 19192 32248
rect 19256 32184 19272 32248
rect 19336 32184 19352 32248
rect 19416 32184 19424 32248
rect 19104 31160 19424 32184
rect 19104 31096 19112 31160
rect 19176 31096 19192 31160
rect 19256 31096 19272 31160
rect 19336 31096 19352 31160
rect 19416 31096 19424 31160
rect 19104 30072 19424 31096
rect 19104 30008 19112 30072
rect 19176 30008 19192 30072
rect 19256 30008 19272 30072
rect 19336 30008 19352 30072
rect 19416 30008 19424 30072
rect 19104 28984 19424 30008
rect 19104 28920 19112 28984
rect 19176 28920 19192 28984
rect 19256 28920 19272 28984
rect 19336 28920 19352 28984
rect 19416 28920 19424 28984
rect 19104 27896 19424 28920
rect 19104 27832 19112 27896
rect 19176 27832 19192 27896
rect 19256 27832 19272 27896
rect 19336 27832 19352 27896
rect 19416 27832 19424 27896
rect 19104 26808 19424 27832
rect 19104 26744 19112 26808
rect 19176 26744 19192 26808
rect 19256 26744 19272 26808
rect 19336 26744 19352 26808
rect 19416 26744 19424 26808
rect 19104 25720 19424 26744
rect 19104 25656 19112 25720
rect 19176 25656 19192 25720
rect 19256 25656 19272 25720
rect 19336 25656 19352 25720
rect 19416 25656 19424 25720
rect 19104 24632 19424 25656
rect 19104 24568 19112 24632
rect 19176 24568 19192 24632
rect 19256 24568 19272 24632
rect 19336 24568 19352 24632
rect 19416 24568 19424 24632
rect 19104 23544 19424 24568
rect 19104 23480 19112 23544
rect 19176 23480 19192 23544
rect 19256 23480 19272 23544
rect 19336 23480 19352 23544
rect 19416 23480 19424 23544
rect 19104 22456 19424 23480
rect 19104 22392 19112 22456
rect 19176 22392 19192 22456
rect 19256 22392 19272 22456
rect 19336 22392 19352 22456
rect 19416 22392 19424 22456
rect 19104 21368 19424 22392
rect 19104 21304 19112 21368
rect 19176 21304 19192 21368
rect 19256 21304 19272 21368
rect 19336 21304 19352 21368
rect 19416 21304 19424 21368
rect 19104 20280 19424 21304
rect 19104 20216 19112 20280
rect 19176 20216 19192 20280
rect 19256 20216 19272 20280
rect 19336 20216 19352 20280
rect 19416 20216 19424 20280
rect 19104 19192 19424 20216
rect 19104 19128 19112 19192
rect 19176 19128 19192 19192
rect 19256 19128 19272 19192
rect 19336 19128 19352 19192
rect 19416 19128 19424 19192
rect 19104 18104 19424 19128
rect 19104 18040 19112 18104
rect 19176 18040 19192 18104
rect 19256 18040 19272 18104
rect 19336 18040 19352 18104
rect 19416 18040 19424 18104
rect 19104 17016 19424 18040
rect 19104 16952 19112 17016
rect 19176 16952 19192 17016
rect 19256 16952 19272 17016
rect 19336 16952 19352 17016
rect 19416 16952 19424 17016
rect 19104 15928 19424 16952
rect 19104 15864 19112 15928
rect 19176 15864 19192 15928
rect 19256 15864 19272 15928
rect 19336 15864 19352 15928
rect 19416 15864 19424 15928
rect 19104 14840 19424 15864
rect 19104 14776 19112 14840
rect 19176 14776 19192 14840
rect 19256 14776 19272 14840
rect 19336 14776 19352 14840
rect 19416 14776 19424 14840
rect 19104 13752 19424 14776
rect 19104 13688 19112 13752
rect 19176 13688 19192 13752
rect 19256 13688 19272 13752
rect 19336 13688 19352 13752
rect 19416 13688 19424 13752
rect 19104 12664 19424 13688
rect 19104 12600 19112 12664
rect 19176 12600 19192 12664
rect 19256 12600 19272 12664
rect 19336 12600 19352 12664
rect 19416 12600 19424 12664
rect 19104 11576 19424 12600
rect 19104 11512 19112 11576
rect 19176 11512 19192 11576
rect 19256 11512 19272 11576
rect 19336 11512 19352 11576
rect 19416 11512 19424 11576
rect 19104 3992 19424 11512
rect 19104 3928 19112 3992
rect 19176 3928 19192 3992
rect 19256 3928 19272 3992
rect 19336 3928 19352 3992
rect 19416 3928 19424 3992
rect 19104 3912 19424 3928
rect 19104 3848 19112 3912
rect 19176 3848 19192 3912
rect 19256 3848 19272 3912
rect 19336 3848 19352 3912
rect 19416 3848 19424 3912
rect 19104 3832 19424 3848
rect 19104 3768 19112 3832
rect 19176 3768 19192 3832
rect 19256 3768 19272 3832
rect 19336 3768 19352 3832
rect 19416 3768 19424 3832
rect 19104 3752 19424 3768
rect 19104 3688 19112 3752
rect 19176 3688 19192 3752
rect 19256 3688 19272 3752
rect 19336 3688 19352 3752
rect 19416 3688 19424 3752
rect 19104 3672 19424 3688
rect 19104 3608 19112 3672
rect 19176 3608 19192 3672
rect 19256 3608 19272 3672
rect 19336 3608 19352 3672
rect 19416 3608 19424 3672
rect 19104 3592 19424 3608
rect 19104 3528 19112 3592
rect 19176 3528 19192 3592
rect 19256 3528 19272 3592
rect 19336 3528 19352 3592
rect 19416 3528 19424 3592
rect 19104 3512 19424 3528
rect 19104 3448 19112 3512
rect 19176 3448 19192 3512
rect 19256 3448 19272 3512
rect 19336 3448 19352 3512
rect 19416 3448 19424 3512
rect 19104 3432 19424 3448
rect 19104 3368 19112 3432
rect 19176 3368 19192 3432
rect 19256 3368 19272 3432
rect 19336 3368 19352 3432
rect 19416 3368 19424 3432
rect 19104 3352 19424 3368
rect 19104 3288 19112 3352
rect 19176 3288 19192 3352
rect 19256 3288 19272 3352
rect 19336 3288 19352 3352
rect 19416 3288 19424 3352
rect 19104 3272 19424 3288
rect 19104 3208 19112 3272
rect 19176 3208 19192 3272
rect 19256 3208 19272 3272
rect 19336 3208 19352 3272
rect 19416 3208 19424 3272
rect 19104 3192 19424 3208
rect 19104 3128 19112 3192
rect 19176 3128 19192 3192
rect 19256 3128 19272 3192
rect 19336 3128 19352 3192
rect 19416 3128 19424 3192
rect 19104 3112 19424 3128
rect 19104 3048 19112 3112
rect 19176 3048 19192 3112
rect 19256 3048 19272 3112
rect 19336 3048 19352 3112
rect 19416 3048 19424 3112
rect 19104 3032 19424 3048
rect 19104 2968 19112 3032
rect 19176 2968 19192 3032
rect 19256 2968 19272 3032
rect 19336 2968 19352 3032
rect 19416 2968 19424 3032
rect 19104 2952 19424 2968
rect 19104 2888 19112 2952
rect 19176 2888 19192 2952
rect 19256 2888 19272 2952
rect 19336 2888 19352 2952
rect 19416 2888 19424 2952
rect 19104 2872 19424 2888
rect 19104 2808 19112 2872
rect 19176 2808 19192 2872
rect 19256 2808 19272 2872
rect 19336 2808 19352 2872
rect 19416 2808 19424 2872
rect 19104 2792 19424 2808
rect 19104 2728 19112 2792
rect 19176 2728 19192 2792
rect 19256 2728 19272 2792
rect 19336 2728 19352 2792
rect 19416 2728 19424 2792
rect 19104 2712 19424 2728
rect 19104 2648 19112 2712
rect 19176 2648 19192 2712
rect 19256 2648 19272 2712
rect 19336 2648 19352 2712
rect 19416 2648 19424 2712
rect 19104 2632 19424 2648
rect 19104 2568 19112 2632
rect 19176 2568 19192 2632
rect 19256 2568 19272 2632
rect 19336 2568 19352 2632
rect 19416 2568 19424 2632
rect 19104 2552 19424 2568
rect 19104 2488 19112 2552
rect 19176 2488 19192 2552
rect 19256 2488 19272 2552
rect 19336 2488 19352 2552
rect 19416 2488 19424 2552
rect 19104 2472 19424 2488
rect 19104 2408 19112 2472
rect 19176 2408 19192 2472
rect 19256 2408 19272 2472
rect 19336 2408 19352 2472
rect 19416 2408 19424 2472
rect 19104 2392 19424 2408
rect 19104 2328 19112 2392
rect 19176 2328 19192 2392
rect 19256 2328 19272 2392
rect 19336 2328 19352 2392
rect 19416 2328 19424 2392
rect 19104 2312 19424 2328
rect 19104 2248 19112 2312
rect 19176 2248 19192 2312
rect 19256 2248 19272 2312
rect 19336 2248 19352 2312
rect 19416 2248 19424 2312
rect 19104 2232 19424 2248
rect 19104 2168 19112 2232
rect 19176 2168 19192 2232
rect 19256 2168 19272 2232
rect 19336 2168 19352 2232
rect 19416 2168 19424 2232
rect 19104 2152 19424 2168
rect 19104 2088 19112 2152
rect 19176 2088 19192 2152
rect 19256 2088 19272 2152
rect 19336 2088 19352 2152
rect 19416 2088 19424 2152
rect 19104 2072 19424 2088
rect 19104 2008 19112 2072
rect 19176 2008 19192 2072
rect 19256 2008 19272 2072
rect 19336 2008 19352 2072
rect 19416 2008 19424 2072
rect 19104 1992 19424 2008
rect 19104 1928 19112 1992
rect 19176 1928 19192 1992
rect 19256 1928 19272 1992
rect 19336 1928 19352 1992
rect 19416 1928 19424 1992
rect 19104 1912 19424 1928
rect 19104 1848 19112 1912
rect 19176 1848 19192 1912
rect 19256 1848 19272 1912
rect 19336 1848 19352 1912
rect 19416 1848 19424 1912
rect 19104 1832 19424 1848
rect 19104 1768 19112 1832
rect 19176 1768 19192 1832
rect 19256 1768 19272 1832
rect 19336 1768 19352 1832
rect 19416 1768 19424 1832
rect 19104 1752 19424 1768
rect 19104 1688 19112 1752
rect 19176 1688 19192 1752
rect 19256 1688 19272 1752
rect 19336 1688 19352 1752
rect 19416 1688 19424 1752
rect 19104 1672 19424 1688
rect 19104 1608 19112 1672
rect 19176 1608 19192 1672
rect 19256 1608 19272 1672
rect 19336 1608 19352 1672
rect 19416 1608 19424 1672
rect 19104 1592 19424 1608
rect 19104 1528 19112 1592
rect 19176 1528 19192 1592
rect 19256 1528 19272 1592
rect 19336 1528 19352 1592
rect 19416 1528 19424 1592
rect 19104 1512 19424 1528
rect 19104 1448 19112 1512
rect 19176 1448 19192 1512
rect 19256 1448 19272 1512
rect 19336 1448 19352 1512
rect 19416 1448 19424 1512
rect 19104 1432 19424 1448
rect 19104 1368 19112 1432
rect 19176 1368 19192 1432
rect 19256 1368 19272 1432
rect 19336 1368 19352 1432
rect 19416 1368 19424 1432
rect 19104 1352 19424 1368
rect 19104 1288 19112 1352
rect 19176 1288 19192 1352
rect 19256 1288 19272 1352
rect 19336 1288 19352 1352
rect 19416 1288 19424 1352
rect 19104 1272 19424 1288
rect 19104 1208 19112 1272
rect 19176 1208 19192 1272
rect 19256 1208 19272 1272
rect 19336 1208 19352 1272
rect 19416 1208 19424 1272
rect 19104 1192 19424 1208
rect 19104 1128 19112 1192
rect 19176 1128 19192 1192
rect 19256 1128 19272 1192
rect 19336 1128 19352 1192
rect 19416 1128 19424 1192
rect 19104 1112 19424 1128
rect 19104 1048 19112 1112
rect 19176 1048 19192 1112
rect 19256 1048 19272 1112
rect 19336 1048 19352 1112
rect 19416 1048 19424 1112
rect 19104 1032 19424 1048
rect 19104 968 19112 1032
rect 19176 968 19192 1032
rect 19256 968 19272 1032
rect 19336 968 19352 1032
rect 19416 968 19424 1032
rect 19104 952 19424 968
rect 19104 888 19112 952
rect 19176 888 19192 952
rect 19256 888 19272 952
rect 19336 888 19352 952
rect 19416 888 19424 952
rect 19104 872 19424 888
rect 19104 808 19112 872
rect 19176 808 19192 872
rect 19256 808 19272 872
rect 19336 808 19352 872
rect 19416 808 19424 872
rect 19104 792 19424 808
rect 19104 728 19112 792
rect 19176 728 19192 792
rect 19256 728 19272 792
rect 19336 728 19352 792
rect 19416 728 19424 792
rect 19104 712 19424 728
rect 19104 648 19112 712
rect 19176 648 19192 712
rect 19256 648 19272 712
rect 19336 648 19352 712
rect 19416 648 19424 712
rect 19104 632 19424 648
rect 19104 568 19112 632
rect 19176 568 19192 632
rect 19256 568 19272 632
rect 19336 568 19352 632
rect 19416 568 19424 632
rect 19104 552 19424 568
rect 19104 488 19112 552
rect 19176 488 19192 552
rect 19256 488 19272 552
rect 19336 488 19352 552
rect 19416 488 19424 552
rect 19104 472 19424 488
rect 19104 408 19112 472
rect 19176 408 19192 472
rect 19256 408 19272 472
rect 19336 408 19352 472
rect 19416 408 19424 472
rect 19104 392 19424 408
rect 19104 328 19112 392
rect 19176 328 19192 392
rect 19256 328 19272 392
rect 19336 328 19352 392
rect 19416 328 19424 392
rect 19104 312 19424 328
rect 19104 248 19112 312
rect 19176 248 19192 312
rect 19256 248 19272 312
rect 19336 248 19352 312
rect 19416 248 19424 312
rect 19104 232 19424 248
rect 19104 168 19112 232
rect 19176 168 19192 232
rect 19256 168 19272 232
rect 19336 168 19352 232
rect 19416 168 19424 232
rect 19104 152 19424 168
rect 19104 88 19112 152
rect 19176 88 19192 152
rect 19256 88 19272 152
rect 19336 88 19352 152
rect 19416 88 19424 152
rect 19104 72 19424 88
rect 19104 8 19112 72
rect 19176 8 19192 72
rect 19256 8 19272 72
rect 19336 8 19352 72
rect 19416 8 19424 72
rect 19104 0 19424 8
rect 24104 40384 24424 45392
rect 24104 40320 24112 40384
rect 24176 40320 24192 40384
rect 24256 40320 24272 40384
rect 24336 40320 24352 40384
rect 24416 40320 24424 40384
rect 24104 40304 24424 40320
rect 24104 40240 24112 40304
rect 24176 40240 24192 40304
rect 24256 40240 24272 40304
rect 24336 40240 24352 40304
rect 24416 40240 24424 40304
rect 24104 40224 24424 40240
rect 24104 40160 24112 40224
rect 24176 40160 24192 40224
rect 24256 40160 24272 40224
rect 24336 40160 24352 40224
rect 24416 40160 24424 40224
rect 24104 40144 24424 40160
rect 24104 40080 24112 40144
rect 24176 40080 24192 40144
rect 24256 40080 24272 40144
rect 24336 40080 24352 40144
rect 24416 40080 24424 40144
rect 24104 40064 24424 40080
rect 24104 40000 24112 40064
rect 24176 40000 24192 40064
rect 24256 40000 24272 40064
rect 24336 40000 24352 40064
rect 24416 40000 24424 40064
rect 24104 39984 24424 40000
rect 24104 39920 24112 39984
rect 24176 39920 24192 39984
rect 24256 39920 24272 39984
rect 24336 39920 24352 39984
rect 24416 39920 24424 39984
rect 24104 39904 24424 39920
rect 24104 39840 24112 39904
rect 24176 39840 24192 39904
rect 24256 39840 24272 39904
rect 24336 39840 24352 39904
rect 24416 39840 24424 39904
rect 24104 39824 24424 39840
rect 24104 39760 24112 39824
rect 24176 39760 24192 39824
rect 24256 39760 24272 39824
rect 24336 39760 24352 39824
rect 24416 39760 24424 39824
rect 24104 39744 24424 39760
rect 24104 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 24424 39744
rect 24104 39664 24424 39680
rect 24104 39600 24112 39664
rect 24176 39600 24192 39664
rect 24256 39600 24272 39664
rect 24336 39600 24352 39664
rect 24416 39600 24424 39664
rect 24104 39584 24424 39600
rect 24104 39520 24112 39584
rect 24176 39520 24192 39584
rect 24256 39520 24272 39584
rect 24336 39520 24352 39584
rect 24416 39520 24424 39584
rect 24104 39504 24424 39520
rect 24104 39440 24112 39504
rect 24176 39440 24192 39504
rect 24256 39440 24272 39504
rect 24336 39440 24352 39504
rect 24416 39440 24424 39504
rect 24104 39424 24424 39440
rect 24104 39360 24112 39424
rect 24176 39360 24192 39424
rect 24256 39360 24272 39424
rect 24336 39360 24352 39424
rect 24416 39360 24424 39424
rect 24104 39344 24424 39360
rect 24104 39280 24112 39344
rect 24176 39280 24192 39344
rect 24256 39280 24272 39344
rect 24336 39280 24352 39344
rect 24416 39280 24424 39344
rect 24104 39264 24424 39280
rect 24104 39200 24112 39264
rect 24176 39200 24192 39264
rect 24256 39200 24272 39264
rect 24336 39200 24352 39264
rect 24416 39200 24424 39264
rect 24104 39184 24424 39200
rect 24104 39120 24112 39184
rect 24176 39120 24192 39184
rect 24256 39120 24272 39184
rect 24336 39120 24352 39184
rect 24416 39120 24424 39184
rect 24104 39104 24424 39120
rect 24104 39040 24112 39104
rect 24176 39040 24192 39104
rect 24256 39040 24272 39104
rect 24336 39040 24352 39104
rect 24416 39040 24424 39104
rect 24104 39024 24424 39040
rect 24104 38960 24112 39024
rect 24176 38960 24192 39024
rect 24256 38960 24272 39024
rect 24336 38960 24352 39024
rect 24416 38960 24424 39024
rect 24104 38944 24424 38960
rect 24104 38880 24112 38944
rect 24176 38880 24192 38944
rect 24256 38880 24272 38944
rect 24336 38880 24352 38944
rect 24416 38880 24424 38944
rect 24104 38864 24424 38880
rect 24104 38800 24112 38864
rect 24176 38800 24192 38864
rect 24256 38800 24272 38864
rect 24336 38800 24352 38864
rect 24416 38800 24424 38864
rect 24104 38784 24424 38800
rect 24104 38720 24112 38784
rect 24176 38720 24192 38784
rect 24256 38720 24272 38784
rect 24336 38720 24352 38784
rect 24416 38720 24424 38784
rect 24104 38704 24424 38720
rect 24104 38640 24112 38704
rect 24176 38640 24192 38704
rect 24256 38640 24272 38704
rect 24336 38640 24352 38704
rect 24416 38640 24424 38704
rect 24104 38624 24424 38640
rect 24104 38560 24112 38624
rect 24176 38560 24192 38624
rect 24256 38560 24272 38624
rect 24336 38560 24352 38624
rect 24416 38560 24424 38624
rect 24104 38544 24424 38560
rect 24104 38480 24112 38544
rect 24176 38480 24192 38544
rect 24256 38480 24272 38544
rect 24336 38480 24352 38544
rect 24416 38480 24424 38544
rect 24104 38464 24424 38480
rect 24104 38400 24112 38464
rect 24176 38400 24192 38464
rect 24256 38400 24272 38464
rect 24336 38400 24352 38464
rect 24416 38400 24424 38464
rect 24104 38384 24424 38400
rect 24104 38320 24112 38384
rect 24176 38320 24192 38384
rect 24256 38320 24272 38384
rect 24336 38320 24352 38384
rect 24416 38320 24424 38384
rect 24104 38304 24424 38320
rect 24104 38240 24112 38304
rect 24176 38240 24192 38304
rect 24256 38240 24272 38304
rect 24336 38240 24352 38304
rect 24416 38240 24424 38304
rect 24104 38224 24424 38240
rect 24104 38160 24112 38224
rect 24176 38160 24192 38224
rect 24256 38160 24272 38224
rect 24336 38160 24352 38224
rect 24416 38160 24424 38224
rect 24104 38144 24424 38160
rect 24104 38080 24112 38144
rect 24176 38080 24192 38144
rect 24256 38080 24272 38144
rect 24336 38080 24352 38144
rect 24416 38080 24424 38144
rect 24104 38064 24424 38080
rect 24104 38000 24112 38064
rect 24176 38000 24192 38064
rect 24256 38000 24272 38064
rect 24336 38000 24352 38064
rect 24416 38000 24424 38064
rect 24104 37984 24424 38000
rect 24104 37920 24112 37984
rect 24176 37920 24192 37984
rect 24256 37920 24272 37984
rect 24336 37920 24352 37984
rect 24416 37920 24424 37984
rect 24104 37904 24424 37920
rect 24104 37840 24112 37904
rect 24176 37840 24192 37904
rect 24256 37840 24272 37904
rect 24336 37840 24352 37904
rect 24416 37840 24424 37904
rect 24104 37824 24424 37840
rect 24104 37760 24112 37824
rect 24176 37760 24192 37824
rect 24256 37760 24272 37824
rect 24336 37760 24352 37824
rect 24416 37760 24424 37824
rect 24104 37744 24424 37760
rect 24104 37680 24112 37744
rect 24176 37680 24192 37744
rect 24256 37680 24272 37744
rect 24336 37680 24352 37744
rect 24416 37680 24424 37744
rect 24104 37664 24424 37680
rect 24104 37600 24112 37664
rect 24176 37600 24192 37664
rect 24256 37600 24272 37664
rect 24336 37600 24352 37664
rect 24416 37600 24424 37664
rect 24104 37584 24424 37600
rect 24104 37520 24112 37584
rect 24176 37520 24192 37584
rect 24256 37520 24272 37584
rect 24336 37520 24352 37584
rect 24416 37520 24424 37584
rect 24104 37504 24424 37520
rect 24104 37440 24112 37504
rect 24176 37440 24192 37504
rect 24256 37440 24272 37504
rect 24336 37440 24352 37504
rect 24416 37440 24424 37504
rect 24104 37424 24424 37440
rect 24104 37360 24112 37424
rect 24176 37360 24192 37424
rect 24256 37360 24272 37424
rect 24336 37360 24352 37424
rect 24416 37360 24424 37424
rect 24104 37344 24424 37360
rect 24104 37280 24112 37344
rect 24176 37280 24192 37344
rect 24256 37280 24272 37344
rect 24336 37280 24352 37344
rect 24416 37280 24424 37344
rect 24104 37264 24424 37280
rect 24104 37200 24112 37264
rect 24176 37200 24192 37264
rect 24256 37200 24272 37264
rect 24336 37200 24352 37264
rect 24416 37200 24424 37264
rect 24104 37184 24424 37200
rect 24104 37120 24112 37184
rect 24176 37120 24192 37184
rect 24256 37120 24272 37184
rect 24336 37120 24352 37184
rect 24416 37120 24424 37184
rect 24104 37104 24424 37120
rect 24104 37040 24112 37104
rect 24176 37040 24192 37104
rect 24256 37040 24272 37104
rect 24336 37040 24352 37104
rect 24416 37040 24424 37104
rect 24104 37024 24424 37040
rect 24104 36960 24112 37024
rect 24176 36960 24192 37024
rect 24256 36960 24272 37024
rect 24336 36960 24352 37024
rect 24416 36960 24424 37024
rect 24104 36944 24424 36960
rect 24104 36880 24112 36944
rect 24176 36880 24192 36944
rect 24256 36880 24272 36944
rect 24336 36880 24352 36944
rect 24416 36880 24424 36944
rect 24104 36864 24424 36880
rect 24104 36800 24112 36864
rect 24176 36800 24192 36864
rect 24256 36800 24272 36864
rect 24336 36800 24352 36864
rect 24416 36800 24424 36864
rect 24104 36784 24424 36800
rect 24104 36720 24112 36784
rect 24176 36720 24192 36784
rect 24256 36720 24272 36784
rect 24336 36720 24352 36784
rect 24416 36720 24424 36784
rect 24104 36704 24424 36720
rect 24104 36640 24112 36704
rect 24176 36640 24192 36704
rect 24256 36640 24272 36704
rect 24336 36640 24352 36704
rect 24416 36640 24424 36704
rect 24104 36624 24424 36640
rect 24104 36560 24112 36624
rect 24176 36560 24192 36624
rect 24256 36560 24272 36624
rect 24336 36560 24352 36624
rect 24416 36560 24424 36624
rect 24104 36544 24424 36560
rect 24104 36480 24112 36544
rect 24176 36480 24192 36544
rect 24256 36480 24272 36544
rect 24336 36480 24352 36544
rect 24416 36480 24424 36544
rect 24104 36464 24424 36480
rect 24104 36400 24112 36464
rect 24176 36400 24192 36464
rect 24256 36400 24272 36464
rect 24336 36400 24352 36464
rect 24416 36400 24424 36464
rect 24104 33880 24424 36400
rect 24104 33816 24112 33880
rect 24176 33816 24192 33880
rect 24256 33816 24272 33880
rect 24336 33816 24352 33880
rect 24416 33816 24424 33880
rect 24104 32792 24424 33816
rect 24104 32728 24112 32792
rect 24176 32728 24192 32792
rect 24256 32728 24272 32792
rect 24336 32728 24352 32792
rect 24416 32728 24424 32792
rect 24104 31704 24424 32728
rect 24104 31640 24112 31704
rect 24176 31640 24192 31704
rect 24256 31640 24272 31704
rect 24336 31640 24352 31704
rect 24416 31640 24424 31704
rect 24104 30616 24424 31640
rect 24104 30552 24112 30616
rect 24176 30552 24192 30616
rect 24256 30552 24272 30616
rect 24336 30552 24352 30616
rect 24416 30552 24424 30616
rect 24104 29528 24424 30552
rect 24104 29464 24112 29528
rect 24176 29464 24192 29528
rect 24256 29464 24272 29528
rect 24336 29464 24352 29528
rect 24416 29464 24424 29528
rect 24104 28440 24424 29464
rect 24104 28376 24112 28440
rect 24176 28376 24192 28440
rect 24256 28376 24272 28440
rect 24336 28376 24352 28440
rect 24416 28376 24424 28440
rect 24104 27352 24424 28376
rect 24104 27288 24112 27352
rect 24176 27288 24192 27352
rect 24256 27288 24272 27352
rect 24336 27288 24352 27352
rect 24416 27288 24424 27352
rect 24104 26264 24424 27288
rect 24104 26200 24112 26264
rect 24176 26200 24192 26264
rect 24256 26200 24272 26264
rect 24336 26200 24352 26264
rect 24416 26200 24424 26264
rect 24104 25176 24424 26200
rect 24104 25112 24112 25176
rect 24176 25112 24192 25176
rect 24256 25112 24272 25176
rect 24336 25112 24352 25176
rect 24416 25112 24424 25176
rect 24104 24088 24424 25112
rect 24104 24024 24112 24088
rect 24176 24024 24192 24088
rect 24256 24024 24272 24088
rect 24336 24024 24352 24088
rect 24416 24024 24424 24088
rect 24104 23000 24424 24024
rect 24104 22936 24112 23000
rect 24176 22936 24192 23000
rect 24256 22936 24272 23000
rect 24336 22936 24352 23000
rect 24416 22936 24424 23000
rect 24104 21912 24424 22936
rect 24104 21848 24112 21912
rect 24176 21848 24192 21912
rect 24256 21848 24272 21912
rect 24336 21848 24352 21912
rect 24416 21848 24424 21912
rect 24104 20824 24424 21848
rect 24104 20760 24112 20824
rect 24176 20760 24192 20824
rect 24256 20760 24272 20824
rect 24336 20760 24352 20824
rect 24416 20760 24424 20824
rect 24104 19736 24424 20760
rect 24104 19672 24112 19736
rect 24176 19672 24192 19736
rect 24256 19672 24272 19736
rect 24336 19672 24352 19736
rect 24416 19672 24424 19736
rect 24104 18648 24424 19672
rect 24104 18584 24112 18648
rect 24176 18584 24192 18648
rect 24256 18584 24272 18648
rect 24336 18584 24352 18648
rect 24416 18584 24424 18648
rect 24104 17560 24424 18584
rect 24104 17496 24112 17560
rect 24176 17496 24192 17560
rect 24256 17496 24272 17560
rect 24336 17496 24352 17560
rect 24416 17496 24424 17560
rect 24104 16472 24424 17496
rect 24104 16408 24112 16472
rect 24176 16408 24192 16472
rect 24256 16408 24272 16472
rect 24336 16408 24352 16472
rect 24416 16408 24424 16472
rect 24104 15384 24424 16408
rect 24104 15320 24112 15384
rect 24176 15320 24192 15384
rect 24256 15320 24272 15384
rect 24336 15320 24352 15384
rect 24416 15320 24424 15384
rect 24104 14296 24424 15320
rect 24104 14232 24112 14296
rect 24176 14232 24192 14296
rect 24256 14232 24272 14296
rect 24336 14232 24352 14296
rect 24416 14232 24424 14296
rect 24104 13208 24424 14232
rect 24104 13144 24112 13208
rect 24176 13144 24192 13208
rect 24256 13144 24272 13208
rect 24336 13144 24352 13208
rect 24416 13144 24424 13208
rect 24104 12120 24424 13144
rect 24104 12056 24112 12120
rect 24176 12056 24192 12120
rect 24256 12056 24272 12120
rect 24336 12056 24352 12120
rect 24416 12056 24424 12120
rect 24104 11032 24424 12056
rect 24104 10968 24112 11032
rect 24176 10968 24192 11032
rect 24256 10968 24272 11032
rect 24336 10968 24352 11032
rect 24416 10968 24424 11032
rect 24104 8992 24424 10968
rect 24104 8928 24112 8992
rect 24176 8928 24192 8992
rect 24256 8928 24272 8992
rect 24336 8928 24352 8992
rect 24416 8928 24424 8992
rect 24104 8912 24424 8928
rect 24104 8848 24112 8912
rect 24176 8848 24192 8912
rect 24256 8848 24272 8912
rect 24336 8848 24352 8912
rect 24416 8848 24424 8912
rect 24104 8832 24424 8848
rect 24104 8768 24112 8832
rect 24176 8768 24192 8832
rect 24256 8768 24272 8832
rect 24336 8768 24352 8832
rect 24416 8768 24424 8832
rect 24104 8752 24424 8768
rect 24104 8688 24112 8752
rect 24176 8688 24192 8752
rect 24256 8688 24272 8752
rect 24336 8688 24352 8752
rect 24416 8688 24424 8752
rect 24104 8672 24424 8688
rect 24104 8608 24112 8672
rect 24176 8608 24192 8672
rect 24256 8608 24272 8672
rect 24336 8608 24352 8672
rect 24416 8608 24424 8672
rect 24104 8592 24424 8608
rect 24104 8528 24112 8592
rect 24176 8528 24192 8592
rect 24256 8528 24272 8592
rect 24336 8528 24352 8592
rect 24416 8528 24424 8592
rect 24104 8512 24424 8528
rect 24104 8448 24112 8512
rect 24176 8448 24192 8512
rect 24256 8448 24272 8512
rect 24336 8448 24352 8512
rect 24416 8448 24424 8512
rect 24104 8432 24424 8448
rect 24104 8368 24112 8432
rect 24176 8368 24192 8432
rect 24256 8368 24272 8432
rect 24336 8368 24352 8432
rect 24416 8368 24424 8432
rect 24104 8352 24424 8368
rect 24104 8288 24112 8352
rect 24176 8288 24192 8352
rect 24256 8288 24272 8352
rect 24336 8288 24352 8352
rect 24416 8288 24424 8352
rect 24104 8272 24424 8288
rect 24104 8208 24112 8272
rect 24176 8208 24192 8272
rect 24256 8208 24272 8272
rect 24336 8208 24352 8272
rect 24416 8208 24424 8272
rect 24104 8192 24424 8208
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 8112 24424 8128
rect 24104 8048 24112 8112
rect 24176 8048 24192 8112
rect 24256 8048 24272 8112
rect 24336 8048 24352 8112
rect 24416 8048 24424 8112
rect 24104 8032 24424 8048
rect 24104 7968 24112 8032
rect 24176 7968 24192 8032
rect 24256 7968 24272 8032
rect 24336 7968 24352 8032
rect 24416 7968 24424 8032
rect 24104 7952 24424 7968
rect 24104 7888 24112 7952
rect 24176 7888 24192 7952
rect 24256 7888 24272 7952
rect 24336 7888 24352 7952
rect 24416 7888 24424 7952
rect 24104 7872 24424 7888
rect 24104 7808 24112 7872
rect 24176 7808 24192 7872
rect 24256 7808 24272 7872
rect 24336 7808 24352 7872
rect 24416 7808 24424 7872
rect 24104 7792 24424 7808
rect 24104 7728 24112 7792
rect 24176 7728 24192 7792
rect 24256 7728 24272 7792
rect 24336 7728 24352 7792
rect 24416 7728 24424 7792
rect 24104 7712 24424 7728
rect 24104 7648 24112 7712
rect 24176 7648 24192 7712
rect 24256 7648 24272 7712
rect 24336 7648 24352 7712
rect 24416 7648 24424 7712
rect 24104 7632 24424 7648
rect 24104 7568 24112 7632
rect 24176 7568 24192 7632
rect 24256 7568 24272 7632
rect 24336 7568 24352 7632
rect 24416 7568 24424 7632
rect 24104 7552 24424 7568
rect 24104 7488 24112 7552
rect 24176 7488 24192 7552
rect 24256 7488 24272 7552
rect 24336 7488 24352 7552
rect 24416 7488 24424 7552
rect 24104 7472 24424 7488
rect 24104 7408 24112 7472
rect 24176 7408 24192 7472
rect 24256 7408 24272 7472
rect 24336 7408 24352 7472
rect 24416 7408 24424 7472
rect 24104 7392 24424 7408
rect 24104 7328 24112 7392
rect 24176 7328 24192 7392
rect 24256 7328 24272 7392
rect 24336 7328 24352 7392
rect 24416 7328 24424 7392
rect 24104 7312 24424 7328
rect 24104 7248 24112 7312
rect 24176 7248 24192 7312
rect 24256 7248 24272 7312
rect 24336 7248 24352 7312
rect 24416 7248 24424 7312
rect 24104 7232 24424 7248
rect 24104 7168 24112 7232
rect 24176 7168 24192 7232
rect 24256 7168 24272 7232
rect 24336 7168 24352 7232
rect 24416 7168 24424 7232
rect 24104 7152 24424 7168
rect 24104 7088 24112 7152
rect 24176 7088 24192 7152
rect 24256 7088 24272 7152
rect 24336 7088 24352 7152
rect 24416 7088 24424 7152
rect 24104 7072 24424 7088
rect 24104 7008 24112 7072
rect 24176 7008 24192 7072
rect 24256 7008 24272 7072
rect 24336 7008 24352 7072
rect 24416 7008 24424 7072
rect 24104 6992 24424 7008
rect 24104 6928 24112 6992
rect 24176 6928 24192 6992
rect 24256 6928 24272 6992
rect 24336 6928 24352 6992
rect 24416 6928 24424 6992
rect 24104 6912 24424 6928
rect 24104 6848 24112 6912
rect 24176 6848 24192 6912
rect 24256 6848 24272 6912
rect 24336 6848 24352 6912
rect 24416 6848 24424 6912
rect 24104 6832 24424 6848
rect 24104 6768 24112 6832
rect 24176 6768 24192 6832
rect 24256 6768 24272 6832
rect 24336 6768 24352 6832
rect 24416 6768 24424 6832
rect 24104 6752 24424 6768
rect 24104 6688 24112 6752
rect 24176 6688 24192 6752
rect 24256 6688 24272 6752
rect 24336 6688 24352 6752
rect 24416 6688 24424 6752
rect 24104 6672 24424 6688
rect 24104 6608 24112 6672
rect 24176 6608 24192 6672
rect 24256 6608 24272 6672
rect 24336 6608 24352 6672
rect 24416 6608 24424 6672
rect 24104 6592 24424 6608
rect 24104 6528 24112 6592
rect 24176 6528 24192 6592
rect 24256 6528 24272 6592
rect 24336 6528 24352 6592
rect 24416 6528 24424 6592
rect 24104 6512 24424 6528
rect 24104 6448 24112 6512
rect 24176 6448 24192 6512
rect 24256 6448 24272 6512
rect 24336 6448 24352 6512
rect 24416 6448 24424 6512
rect 24104 6432 24424 6448
rect 24104 6368 24112 6432
rect 24176 6368 24192 6432
rect 24256 6368 24272 6432
rect 24336 6368 24352 6432
rect 24416 6368 24424 6432
rect 24104 6352 24424 6368
rect 24104 6288 24112 6352
rect 24176 6288 24192 6352
rect 24256 6288 24272 6352
rect 24336 6288 24352 6352
rect 24416 6288 24424 6352
rect 24104 6272 24424 6288
rect 24104 6208 24112 6272
rect 24176 6208 24192 6272
rect 24256 6208 24272 6272
rect 24336 6208 24352 6272
rect 24416 6208 24424 6272
rect 24104 6192 24424 6208
rect 24104 6128 24112 6192
rect 24176 6128 24192 6192
rect 24256 6128 24272 6192
rect 24336 6128 24352 6192
rect 24416 6128 24424 6192
rect 24104 6112 24424 6128
rect 24104 6048 24112 6112
rect 24176 6048 24192 6112
rect 24256 6048 24272 6112
rect 24336 6048 24352 6112
rect 24416 6048 24424 6112
rect 24104 6032 24424 6048
rect 24104 5968 24112 6032
rect 24176 5968 24192 6032
rect 24256 5968 24272 6032
rect 24336 5968 24352 6032
rect 24416 5968 24424 6032
rect 24104 5952 24424 5968
rect 24104 5888 24112 5952
rect 24176 5888 24192 5952
rect 24256 5888 24272 5952
rect 24336 5888 24352 5952
rect 24416 5888 24424 5952
rect 24104 5872 24424 5888
rect 24104 5808 24112 5872
rect 24176 5808 24192 5872
rect 24256 5808 24272 5872
rect 24336 5808 24352 5872
rect 24416 5808 24424 5872
rect 24104 5792 24424 5808
rect 24104 5728 24112 5792
rect 24176 5728 24192 5792
rect 24256 5728 24272 5792
rect 24336 5728 24352 5792
rect 24416 5728 24424 5792
rect 24104 5712 24424 5728
rect 24104 5648 24112 5712
rect 24176 5648 24192 5712
rect 24256 5648 24272 5712
rect 24336 5648 24352 5712
rect 24416 5648 24424 5712
rect 24104 5632 24424 5648
rect 24104 5568 24112 5632
rect 24176 5568 24192 5632
rect 24256 5568 24272 5632
rect 24336 5568 24352 5632
rect 24416 5568 24424 5632
rect 24104 5552 24424 5568
rect 24104 5488 24112 5552
rect 24176 5488 24192 5552
rect 24256 5488 24272 5552
rect 24336 5488 24352 5552
rect 24416 5488 24424 5552
rect 24104 5472 24424 5488
rect 24104 5408 24112 5472
rect 24176 5408 24192 5472
rect 24256 5408 24272 5472
rect 24336 5408 24352 5472
rect 24416 5408 24424 5472
rect 24104 5392 24424 5408
rect 24104 5328 24112 5392
rect 24176 5328 24192 5392
rect 24256 5328 24272 5392
rect 24336 5328 24352 5392
rect 24416 5328 24424 5392
rect 24104 5312 24424 5328
rect 24104 5248 24112 5312
rect 24176 5248 24192 5312
rect 24256 5248 24272 5312
rect 24336 5248 24352 5312
rect 24416 5248 24424 5312
rect 24104 5232 24424 5248
rect 24104 5168 24112 5232
rect 24176 5168 24192 5232
rect 24256 5168 24272 5232
rect 24336 5168 24352 5232
rect 24416 5168 24424 5232
rect 24104 5152 24424 5168
rect 24104 5088 24112 5152
rect 24176 5088 24192 5152
rect 24256 5088 24272 5152
rect 24336 5088 24352 5152
rect 24416 5088 24424 5152
rect 24104 5072 24424 5088
rect 24104 5008 24112 5072
rect 24176 5008 24192 5072
rect 24256 5008 24272 5072
rect 24336 5008 24352 5072
rect 24416 5008 24424 5072
rect 24104 0 24424 5008
rect 29104 45384 29424 45392
rect 29104 45320 29112 45384
rect 29176 45320 29192 45384
rect 29256 45320 29272 45384
rect 29336 45320 29352 45384
rect 29416 45320 29424 45384
rect 29104 45304 29424 45320
rect 29104 45240 29112 45304
rect 29176 45240 29192 45304
rect 29256 45240 29272 45304
rect 29336 45240 29352 45304
rect 29416 45240 29424 45304
rect 29104 45224 29424 45240
rect 29104 45160 29112 45224
rect 29176 45160 29192 45224
rect 29256 45160 29272 45224
rect 29336 45160 29352 45224
rect 29416 45160 29424 45224
rect 29104 45144 29424 45160
rect 29104 45080 29112 45144
rect 29176 45080 29192 45144
rect 29256 45080 29272 45144
rect 29336 45080 29352 45144
rect 29416 45080 29424 45144
rect 29104 45064 29424 45080
rect 29104 45000 29112 45064
rect 29176 45000 29192 45064
rect 29256 45000 29272 45064
rect 29336 45000 29352 45064
rect 29416 45000 29424 45064
rect 29104 44984 29424 45000
rect 29104 44920 29112 44984
rect 29176 44920 29192 44984
rect 29256 44920 29272 44984
rect 29336 44920 29352 44984
rect 29416 44920 29424 44984
rect 29104 44904 29424 44920
rect 29104 44840 29112 44904
rect 29176 44840 29192 44904
rect 29256 44840 29272 44904
rect 29336 44840 29352 44904
rect 29416 44840 29424 44904
rect 29104 44824 29424 44840
rect 29104 44760 29112 44824
rect 29176 44760 29192 44824
rect 29256 44760 29272 44824
rect 29336 44760 29352 44824
rect 29416 44760 29424 44824
rect 29104 44744 29424 44760
rect 29104 44680 29112 44744
rect 29176 44680 29192 44744
rect 29256 44680 29272 44744
rect 29336 44680 29352 44744
rect 29416 44680 29424 44744
rect 29104 44664 29424 44680
rect 29104 44600 29112 44664
rect 29176 44600 29192 44664
rect 29256 44600 29272 44664
rect 29336 44600 29352 44664
rect 29416 44600 29424 44664
rect 29104 44584 29424 44600
rect 29104 44520 29112 44584
rect 29176 44520 29192 44584
rect 29256 44520 29272 44584
rect 29336 44520 29352 44584
rect 29416 44520 29424 44584
rect 29104 44504 29424 44520
rect 29104 44440 29112 44504
rect 29176 44440 29192 44504
rect 29256 44440 29272 44504
rect 29336 44440 29352 44504
rect 29416 44440 29424 44504
rect 29104 44424 29424 44440
rect 29104 44360 29112 44424
rect 29176 44360 29192 44424
rect 29256 44360 29272 44424
rect 29336 44360 29352 44424
rect 29416 44360 29424 44424
rect 29104 44344 29424 44360
rect 29104 44280 29112 44344
rect 29176 44280 29192 44344
rect 29256 44280 29272 44344
rect 29336 44280 29352 44344
rect 29416 44280 29424 44344
rect 29104 44264 29424 44280
rect 29104 44200 29112 44264
rect 29176 44200 29192 44264
rect 29256 44200 29272 44264
rect 29336 44200 29352 44264
rect 29416 44200 29424 44264
rect 29104 44184 29424 44200
rect 29104 44120 29112 44184
rect 29176 44120 29192 44184
rect 29256 44120 29272 44184
rect 29336 44120 29352 44184
rect 29416 44120 29424 44184
rect 29104 44104 29424 44120
rect 29104 44040 29112 44104
rect 29176 44040 29192 44104
rect 29256 44040 29272 44104
rect 29336 44040 29352 44104
rect 29416 44040 29424 44104
rect 29104 44024 29424 44040
rect 29104 43960 29112 44024
rect 29176 43960 29192 44024
rect 29256 43960 29272 44024
rect 29336 43960 29352 44024
rect 29416 43960 29424 44024
rect 29104 43944 29424 43960
rect 29104 43880 29112 43944
rect 29176 43880 29192 43944
rect 29256 43880 29272 43944
rect 29336 43880 29352 43944
rect 29416 43880 29424 43944
rect 29104 43864 29424 43880
rect 29104 43800 29112 43864
rect 29176 43800 29192 43864
rect 29256 43800 29272 43864
rect 29336 43800 29352 43864
rect 29416 43800 29424 43864
rect 29104 43784 29424 43800
rect 29104 43720 29112 43784
rect 29176 43720 29192 43784
rect 29256 43720 29272 43784
rect 29336 43720 29352 43784
rect 29416 43720 29424 43784
rect 29104 43704 29424 43720
rect 29104 43640 29112 43704
rect 29176 43640 29192 43704
rect 29256 43640 29272 43704
rect 29336 43640 29352 43704
rect 29416 43640 29424 43704
rect 29104 43624 29424 43640
rect 29104 43560 29112 43624
rect 29176 43560 29192 43624
rect 29256 43560 29272 43624
rect 29336 43560 29352 43624
rect 29416 43560 29424 43624
rect 29104 43544 29424 43560
rect 29104 43480 29112 43544
rect 29176 43480 29192 43544
rect 29256 43480 29272 43544
rect 29336 43480 29352 43544
rect 29416 43480 29424 43544
rect 29104 43464 29424 43480
rect 29104 43400 29112 43464
rect 29176 43400 29192 43464
rect 29256 43400 29272 43464
rect 29336 43400 29352 43464
rect 29416 43400 29424 43464
rect 29104 43384 29424 43400
rect 29104 43320 29112 43384
rect 29176 43320 29192 43384
rect 29256 43320 29272 43384
rect 29336 43320 29352 43384
rect 29416 43320 29424 43384
rect 29104 43304 29424 43320
rect 29104 43240 29112 43304
rect 29176 43240 29192 43304
rect 29256 43240 29272 43304
rect 29336 43240 29352 43304
rect 29416 43240 29424 43304
rect 29104 43224 29424 43240
rect 29104 43160 29112 43224
rect 29176 43160 29192 43224
rect 29256 43160 29272 43224
rect 29336 43160 29352 43224
rect 29416 43160 29424 43224
rect 29104 43144 29424 43160
rect 29104 43080 29112 43144
rect 29176 43080 29192 43144
rect 29256 43080 29272 43144
rect 29336 43080 29352 43144
rect 29416 43080 29424 43144
rect 29104 43064 29424 43080
rect 29104 43000 29112 43064
rect 29176 43000 29192 43064
rect 29256 43000 29272 43064
rect 29336 43000 29352 43064
rect 29416 43000 29424 43064
rect 29104 42984 29424 43000
rect 29104 42920 29112 42984
rect 29176 42920 29192 42984
rect 29256 42920 29272 42984
rect 29336 42920 29352 42984
rect 29416 42920 29424 42984
rect 29104 42904 29424 42920
rect 29104 42840 29112 42904
rect 29176 42840 29192 42904
rect 29256 42840 29272 42904
rect 29336 42840 29352 42904
rect 29416 42840 29424 42904
rect 29104 42824 29424 42840
rect 29104 42760 29112 42824
rect 29176 42760 29192 42824
rect 29256 42760 29272 42824
rect 29336 42760 29352 42824
rect 29416 42760 29424 42824
rect 29104 42744 29424 42760
rect 29104 42680 29112 42744
rect 29176 42680 29192 42744
rect 29256 42680 29272 42744
rect 29336 42680 29352 42744
rect 29416 42680 29424 42744
rect 29104 42664 29424 42680
rect 29104 42600 29112 42664
rect 29176 42600 29192 42664
rect 29256 42600 29272 42664
rect 29336 42600 29352 42664
rect 29416 42600 29424 42664
rect 29104 42584 29424 42600
rect 29104 42520 29112 42584
rect 29176 42520 29192 42584
rect 29256 42520 29272 42584
rect 29336 42520 29352 42584
rect 29416 42520 29424 42584
rect 29104 42504 29424 42520
rect 29104 42440 29112 42504
rect 29176 42440 29192 42504
rect 29256 42440 29272 42504
rect 29336 42440 29352 42504
rect 29416 42440 29424 42504
rect 29104 42424 29424 42440
rect 29104 42360 29112 42424
rect 29176 42360 29192 42424
rect 29256 42360 29272 42424
rect 29336 42360 29352 42424
rect 29416 42360 29424 42424
rect 29104 42344 29424 42360
rect 29104 42280 29112 42344
rect 29176 42280 29192 42344
rect 29256 42280 29272 42344
rect 29336 42280 29352 42344
rect 29416 42280 29424 42344
rect 29104 42264 29424 42280
rect 29104 42200 29112 42264
rect 29176 42200 29192 42264
rect 29256 42200 29272 42264
rect 29336 42200 29352 42264
rect 29416 42200 29424 42264
rect 29104 42184 29424 42200
rect 29104 42120 29112 42184
rect 29176 42120 29192 42184
rect 29256 42120 29272 42184
rect 29336 42120 29352 42184
rect 29416 42120 29424 42184
rect 29104 42104 29424 42120
rect 29104 42040 29112 42104
rect 29176 42040 29192 42104
rect 29256 42040 29272 42104
rect 29336 42040 29352 42104
rect 29416 42040 29424 42104
rect 29104 42024 29424 42040
rect 29104 41960 29112 42024
rect 29176 41960 29192 42024
rect 29256 41960 29272 42024
rect 29336 41960 29352 42024
rect 29416 41960 29424 42024
rect 29104 41944 29424 41960
rect 29104 41880 29112 41944
rect 29176 41880 29192 41944
rect 29256 41880 29272 41944
rect 29336 41880 29352 41944
rect 29416 41880 29424 41944
rect 29104 41864 29424 41880
rect 29104 41800 29112 41864
rect 29176 41800 29192 41864
rect 29256 41800 29272 41864
rect 29336 41800 29352 41864
rect 29416 41800 29424 41864
rect 29104 41784 29424 41800
rect 29104 41720 29112 41784
rect 29176 41720 29192 41784
rect 29256 41720 29272 41784
rect 29336 41720 29352 41784
rect 29416 41720 29424 41784
rect 29104 41704 29424 41720
rect 29104 41640 29112 41704
rect 29176 41640 29192 41704
rect 29256 41640 29272 41704
rect 29336 41640 29352 41704
rect 29416 41640 29424 41704
rect 29104 41624 29424 41640
rect 29104 41560 29112 41624
rect 29176 41560 29192 41624
rect 29256 41560 29272 41624
rect 29336 41560 29352 41624
rect 29416 41560 29424 41624
rect 29104 41544 29424 41560
rect 29104 41480 29112 41544
rect 29176 41480 29192 41544
rect 29256 41480 29272 41544
rect 29336 41480 29352 41544
rect 29416 41480 29424 41544
rect 29104 41464 29424 41480
rect 29104 41400 29112 41464
rect 29176 41400 29192 41464
rect 29256 41400 29272 41464
rect 29336 41400 29352 41464
rect 29416 41400 29424 41464
rect 29104 34424 29424 41400
rect 41368 45384 45368 45392
rect 41368 45320 41376 45384
rect 41440 45320 41456 45384
rect 41520 45320 41536 45384
rect 41600 45320 41616 45384
rect 41680 45320 41696 45384
rect 41760 45320 41776 45384
rect 41840 45320 41856 45384
rect 41920 45320 41936 45384
rect 42000 45320 42016 45384
rect 42080 45320 42096 45384
rect 42160 45320 42176 45384
rect 42240 45320 42256 45384
rect 42320 45320 42336 45384
rect 42400 45320 42416 45384
rect 42480 45320 42496 45384
rect 42560 45320 42576 45384
rect 42640 45320 42656 45384
rect 42720 45320 42736 45384
rect 42800 45320 42816 45384
rect 42880 45320 42896 45384
rect 42960 45320 42976 45384
rect 43040 45320 43056 45384
rect 43120 45320 43136 45384
rect 43200 45320 43216 45384
rect 43280 45320 43296 45384
rect 43360 45320 43376 45384
rect 43440 45320 43456 45384
rect 43520 45320 43536 45384
rect 43600 45320 43616 45384
rect 43680 45320 43696 45384
rect 43760 45320 43776 45384
rect 43840 45320 43856 45384
rect 43920 45320 43936 45384
rect 44000 45320 44016 45384
rect 44080 45320 44096 45384
rect 44160 45320 44176 45384
rect 44240 45320 44256 45384
rect 44320 45320 44336 45384
rect 44400 45320 44416 45384
rect 44480 45320 44496 45384
rect 44560 45320 44576 45384
rect 44640 45320 44656 45384
rect 44720 45320 44736 45384
rect 44800 45320 44816 45384
rect 44880 45320 44896 45384
rect 44960 45320 44976 45384
rect 45040 45320 45056 45384
rect 45120 45320 45136 45384
rect 45200 45320 45216 45384
rect 45280 45320 45296 45384
rect 45360 45320 45368 45384
rect 41368 45304 45368 45320
rect 41368 45240 41376 45304
rect 41440 45240 41456 45304
rect 41520 45240 41536 45304
rect 41600 45240 41616 45304
rect 41680 45240 41696 45304
rect 41760 45240 41776 45304
rect 41840 45240 41856 45304
rect 41920 45240 41936 45304
rect 42000 45240 42016 45304
rect 42080 45240 42096 45304
rect 42160 45240 42176 45304
rect 42240 45240 42256 45304
rect 42320 45240 42336 45304
rect 42400 45240 42416 45304
rect 42480 45240 42496 45304
rect 42560 45240 42576 45304
rect 42640 45240 42656 45304
rect 42720 45240 42736 45304
rect 42800 45240 42816 45304
rect 42880 45240 42896 45304
rect 42960 45240 42976 45304
rect 43040 45240 43056 45304
rect 43120 45240 43136 45304
rect 43200 45240 43216 45304
rect 43280 45240 43296 45304
rect 43360 45240 43376 45304
rect 43440 45240 43456 45304
rect 43520 45240 43536 45304
rect 43600 45240 43616 45304
rect 43680 45240 43696 45304
rect 43760 45240 43776 45304
rect 43840 45240 43856 45304
rect 43920 45240 43936 45304
rect 44000 45240 44016 45304
rect 44080 45240 44096 45304
rect 44160 45240 44176 45304
rect 44240 45240 44256 45304
rect 44320 45240 44336 45304
rect 44400 45240 44416 45304
rect 44480 45240 44496 45304
rect 44560 45240 44576 45304
rect 44640 45240 44656 45304
rect 44720 45240 44736 45304
rect 44800 45240 44816 45304
rect 44880 45240 44896 45304
rect 44960 45240 44976 45304
rect 45040 45240 45056 45304
rect 45120 45240 45136 45304
rect 45200 45240 45216 45304
rect 45280 45240 45296 45304
rect 45360 45240 45368 45304
rect 41368 45224 45368 45240
rect 41368 45160 41376 45224
rect 41440 45160 41456 45224
rect 41520 45160 41536 45224
rect 41600 45160 41616 45224
rect 41680 45160 41696 45224
rect 41760 45160 41776 45224
rect 41840 45160 41856 45224
rect 41920 45160 41936 45224
rect 42000 45160 42016 45224
rect 42080 45160 42096 45224
rect 42160 45160 42176 45224
rect 42240 45160 42256 45224
rect 42320 45160 42336 45224
rect 42400 45160 42416 45224
rect 42480 45160 42496 45224
rect 42560 45160 42576 45224
rect 42640 45160 42656 45224
rect 42720 45160 42736 45224
rect 42800 45160 42816 45224
rect 42880 45160 42896 45224
rect 42960 45160 42976 45224
rect 43040 45160 43056 45224
rect 43120 45160 43136 45224
rect 43200 45160 43216 45224
rect 43280 45160 43296 45224
rect 43360 45160 43376 45224
rect 43440 45160 43456 45224
rect 43520 45160 43536 45224
rect 43600 45160 43616 45224
rect 43680 45160 43696 45224
rect 43760 45160 43776 45224
rect 43840 45160 43856 45224
rect 43920 45160 43936 45224
rect 44000 45160 44016 45224
rect 44080 45160 44096 45224
rect 44160 45160 44176 45224
rect 44240 45160 44256 45224
rect 44320 45160 44336 45224
rect 44400 45160 44416 45224
rect 44480 45160 44496 45224
rect 44560 45160 44576 45224
rect 44640 45160 44656 45224
rect 44720 45160 44736 45224
rect 44800 45160 44816 45224
rect 44880 45160 44896 45224
rect 44960 45160 44976 45224
rect 45040 45160 45056 45224
rect 45120 45160 45136 45224
rect 45200 45160 45216 45224
rect 45280 45160 45296 45224
rect 45360 45160 45368 45224
rect 41368 45144 45368 45160
rect 41368 45080 41376 45144
rect 41440 45080 41456 45144
rect 41520 45080 41536 45144
rect 41600 45080 41616 45144
rect 41680 45080 41696 45144
rect 41760 45080 41776 45144
rect 41840 45080 41856 45144
rect 41920 45080 41936 45144
rect 42000 45080 42016 45144
rect 42080 45080 42096 45144
rect 42160 45080 42176 45144
rect 42240 45080 42256 45144
rect 42320 45080 42336 45144
rect 42400 45080 42416 45144
rect 42480 45080 42496 45144
rect 42560 45080 42576 45144
rect 42640 45080 42656 45144
rect 42720 45080 42736 45144
rect 42800 45080 42816 45144
rect 42880 45080 42896 45144
rect 42960 45080 42976 45144
rect 43040 45080 43056 45144
rect 43120 45080 43136 45144
rect 43200 45080 43216 45144
rect 43280 45080 43296 45144
rect 43360 45080 43376 45144
rect 43440 45080 43456 45144
rect 43520 45080 43536 45144
rect 43600 45080 43616 45144
rect 43680 45080 43696 45144
rect 43760 45080 43776 45144
rect 43840 45080 43856 45144
rect 43920 45080 43936 45144
rect 44000 45080 44016 45144
rect 44080 45080 44096 45144
rect 44160 45080 44176 45144
rect 44240 45080 44256 45144
rect 44320 45080 44336 45144
rect 44400 45080 44416 45144
rect 44480 45080 44496 45144
rect 44560 45080 44576 45144
rect 44640 45080 44656 45144
rect 44720 45080 44736 45144
rect 44800 45080 44816 45144
rect 44880 45080 44896 45144
rect 44960 45080 44976 45144
rect 45040 45080 45056 45144
rect 45120 45080 45136 45144
rect 45200 45080 45216 45144
rect 45280 45080 45296 45144
rect 45360 45080 45368 45144
rect 41368 45064 45368 45080
rect 41368 45000 41376 45064
rect 41440 45000 41456 45064
rect 41520 45000 41536 45064
rect 41600 45000 41616 45064
rect 41680 45000 41696 45064
rect 41760 45000 41776 45064
rect 41840 45000 41856 45064
rect 41920 45000 41936 45064
rect 42000 45000 42016 45064
rect 42080 45000 42096 45064
rect 42160 45000 42176 45064
rect 42240 45000 42256 45064
rect 42320 45000 42336 45064
rect 42400 45000 42416 45064
rect 42480 45000 42496 45064
rect 42560 45000 42576 45064
rect 42640 45000 42656 45064
rect 42720 45000 42736 45064
rect 42800 45000 42816 45064
rect 42880 45000 42896 45064
rect 42960 45000 42976 45064
rect 43040 45000 43056 45064
rect 43120 45000 43136 45064
rect 43200 45000 43216 45064
rect 43280 45000 43296 45064
rect 43360 45000 43376 45064
rect 43440 45000 43456 45064
rect 43520 45000 43536 45064
rect 43600 45000 43616 45064
rect 43680 45000 43696 45064
rect 43760 45000 43776 45064
rect 43840 45000 43856 45064
rect 43920 45000 43936 45064
rect 44000 45000 44016 45064
rect 44080 45000 44096 45064
rect 44160 45000 44176 45064
rect 44240 45000 44256 45064
rect 44320 45000 44336 45064
rect 44400 45000 44416 45064
rect 44480 45000 44496 45064
rect 44560 45000 44576 45064
rect 44640 45000 44656 45064
rect 44720 45000 44736 45064
rect 44800 45000 44816 45064
rect 44880 45000 44896 45064
rect 44960 45000 44976 45064
rect 45040 45000 45056 45064
rect 45120 45000 45136 45064
rect 45200 45000 45216 45064
rect 45280 45000 45296 45064
rect 45360 45000 45368 45064
rect 41368 44984 45368 45000
rect 41368 44920 41376 44984
rect 41440 44920 41456 44984
rect 41520 44920 41536 44984
rect 41600 44920 41616 44984
rect 41680 44920 41696 44984
rect 41760 44920 41776 44984
rect 41840 44920 41856 44984
rect 41920 44920 41936 44984
rect 42000 44920 42016 44984
rect 42080 44920 42096 44984
rect 42160 44920 42176 44984
rect 42240 44920 42256 44984
rect 42320 44920 42336 44984
rect 42400 44920 42416 44984
rect 42480 44920 42496 44984
rect 42560 44920 42576 44984
rect 42640 44920 42656 44984
rect 42720 44920 42736 44984
rect 42800 44920 42816 44984
rect 42880 44920 42896 44984
rect 42960 44920 42976 44984
rect 43040 44920 43056 44984
rect 43120 44920 43136 44984
rect 43200 44920 43216 44984
rect 43280 44920 43296 44984
rect 43360 44920 43376 44984
rect 43440 44920 43456 44984
rect 43520 44920 43536 44984
rect 43600 44920 43616 44984
rect 43680 44920 43696 44984
rect 43760 44920 43776 44984
rect 43840 44920 43856 44984
rect 43920 44920 43936 44984
rect 44000 44920 44016 44984
rect 44080 44920 44096 44984
rect 44160 44920 44176 44984
rect 44240 44920 44256 44984
rect 44320 44920 44336 44984
rect 44400 44920 44416 44984
rect 44480 44920 44496 44984
rect 44560 44920 44576 44984
rect 44640 44920 44656 44984
rect 44720 44920 44736 44984
rect 44800 44920 44816 44984
rect 44880 44920 44896 44984
rect 44960 44920 44976 44984
rect 45040 44920 45056 44984
rect 45120 44920 45136 44984
rect 45200 44920 45216 44984
rect 45280 44920 45296 44984
rect 45360 44920 45368 44984
rect 41368 44904 45368 44920
rect 41368 44840 41376 44904
rect 41440 44840 41456 44904
rect 41520 44840 41536 44904
rect 41600 44840 41616 44904
rect 41680 44840 41696 44904
rect 41760 44840 41776 44904
rect 41840 44840 41856 44904
rect 41920 44840 41936 44904
rect 42000 44840 42016 44904
rect 42080 44840 42096 44904
rect 42160 44840 42176 44904
rect 42240 44840 42256 44904
rect 42320 44840 42336 44904
rect 42400 44840 42416 44904
rect 42480 44840 42496 44904
rect 42560 44840 42576 44904
rect 42640 44840 42656 44904
rect 42720 44840 42736 44904
rect 42800 44840 42816 44904
rect 42880 44840 42896 44904
rect 42960 44840 42976 44904
rect 43040 44840 43056 44904
rect 43120 44840 43136 44904
rect 43200 44840 43216 44904
rect 43280 44840 43296 44904
rect 43360 44840 43376 44904
rect 43440 44840 43456 44904
rect 43520 44840 43536 44904
rect 43600 44840 43616 44904
rect 43680 44840 43696 44904
rect 43760 44840 43776 44904
rect 43840 44840 43856 44904
rect 43920 44840 43936 44904
rect 44000 44840 44016 44904
rect 44080 44840 44096 44904
rect 44160 44840 44176 44904
rect 44240 44840 44256 44904
rect 44320 44840 44336 44904
rect 44400 44840 44416 44904
rect 44480 44840 44496 44904
rect 44560 44840 44576 44904
rect 44640 44840 44656 44904
rect 44720 44840 44736 44904
rect 44800 44840 44816 44904
rect 44880 44840 44896 44904
rect 44960 44840 44976 44904
rect 45040 44840 45056 44904
rect 45120 44840 45136 44904
rect 45200 44840 45216 44904
rect 45280 44840 45296 44904
rect 45360 44840 45368 44904
rect 41368 44824 45368 44840
rect 41368 44760 41376 44824
rect 41440 44760 41456 44824
rect 41520 44760 41536 44824
rect 41600 44760 41616 44824
rect 41680 44760 41696 44824
rect 41760 44760 41776 44824
rect 41840 44760 41856 44824
rect 41920 44760 41936 44824
rect 42000 44760 42016 44824
rect 42080 44760 42096 44824
rect 42160 44760 42176 44824
rect 42240 44760 42256 44824
rect 42320 44760 42336 44824
rect 42400 44760 42416 44824
rect 42480 44760 42496 44824
rect 42560 44760 42576 44824
rect 42640 44760 42656 44824
rect 42720 44760 42736 44824
rect 42800 44760 42816 44824
rect 42880 44760 42896 44824
rect 42960 44760 42976 44824
rect 43040 44760 43056 44824
rect 43120 44760 43136 44824
rect 43200 44760 43216 44824
rect 43280 44760 43296 44824
rect 43360 44760 43376 44824
rect 43440 44760 43456 44824
rect 43520 44760 43536 44824
rect 43600 44760 43616 44824
rect 43680 44760 43696 44824
rect 43760 44760 43776 44824
rect 43840 44760 43856 44824
rect 43920 44760 43936 44824
rect 44000 44760 44016 44824
rect 44080 44760 44096 44824
rect 44160 44760 44176 44824
rect 44240 44760 44256 44824
rect 44320 44760 44336 44824
rect 44400 44760 44416 44824
rect 44480 44760 44496 44824
rect 44560 44760 44576 44824
rect 44640 44760 44656 44824
rect 44720 44760 44736 44824
rect 44800 44760 44816 44824
rect 44880 44760 44896 44824
rect 44960 44760 44976 44824
rect 45040 44760 45056 44824
rect 45120 44760 45136 44824
rect 45200 44760 45216 44824
rect 45280 44760 45296 44824
rect 45360 44760 45368 44824
rect 41368 44744 45368 44760
rect 41368 44680 41376 44744
rect 41440 44680 41456 44744
rect 41520 44680 41536 44744
rect 41600 44680 41616 44744
rect 41680 44680 41696 44744
rect 41760 44680 41776 44744
rect 41840 44680 41856 44744
rect 41920 44680 41936 44744
rect 42000 44680 42016 44744
rect 42080 44680 42096 44744
rect 42160 44680 42176 44744
rect 42240 44680 42256 44744
rect 42320 44680 42336 44744
rect 42400 44680 42416 44744
rect 42480 44680 42496 44744
rect 42560 44680 42576 44744
rect 42640 44680 42656 44744
rect 42720 44680 42736 44744
rect 42800 44680 42816 44744
rect 42880 44680 42896 44744
rect 42960 44680 42976 44744
rect 43040 44680 43056 44744
rect 43120 44680 43136 44744
rect 43200 44680 43216 44744
rect 43280 44680 43296 44744
rect 43360 44680 43376 44744
rect 43440 44680 43456 44744
rect 43520 44680 43536 44744
rect 43600 44680 43616 44744
rect 43680 44680 43696 44744
rect 43760 44680 43776 44744
rect 43840 44680 43856 44744
rect 43920 44680 43936 44744
rect 44000 44680 44016 44744
rect 44080 44680 44096 44744
rect 44160 44680 44176 44744
rect 44240 44680 44256 44744
rect 44320 44680 44336 44744
rect 44400 44680 44416 44744
rect 44480 44680 44496 44744
rect 44560 44680 44576 44744
rect 44640 44680 44656 44744
rect 44720 44680 44736 44744
rect 44800 44680 44816 44744
rect 44880 44680 44896 44744
rect 44960 44680 44976 44744
rect 45040 44680 45056 44744
rect 45120 44680 45136 44744
rect 45200 44680 45216 44744
rect 45280 44680 45296 44744
rect 45360 44680 45368 44744
rect 41368 44664 45368 44680
rect 41368 44600 41376 44664
rect 41440 44600 41456 44664
rect 41520 44600 41536 44664
rect 41600 44600 41616 44664
rect 41680 44600 41696 44664
rect 41760 44600 41776 44664
rect 41840 44600 41856 44664
rect 41920 44600 41936 44664
rect 42000 44600 42016 44664
rect 42080 44600 42096 44664
rect 42160 44600 42176 44664
rect 42240 44600 42256 44664
rect 42320 44600 42336 44664
rect 42400 44600 42416 44664
rect 42480 44600 42496 44664
rect 42560 44600 42576 44664
rect 42640 44600 42656 44664
rect 42720 44600 42736 44664
rect 42800 44600 42816 44664
rect 42880 44600 42896 44664
rect 42960 44600 42976 44664
rect 43040 44600 43056 44664
rect 43120 44600 43136 44664
rect 43200 44600 43216 44664
rect 43280 44600 43296 44664
rect 43360 44600 43376 44664
rect 43440 44600 43456 44664
rect 43520 44600 43536 44664
rect 43600 44600 43616 44664
rect 43680 44600 43696 44664
rect 43760 44600 43776 44664
rect 43840 44600 43856 44664
rect 43920 44600 43936 44664
rect 44000 44600 44016 44664
rect 44080 44600 44096 44664
rect 44160 44600 44176 44664
rect 44240 44600 44256 44664
rect 44320 44600 44336 44664
rect 44400 44600 44416 44664
rect 44480 44600 44496 44664
rect 44560 44600 44576 44664
rect 44640 44600 44656 44664
rect 44720 44600 44736 44664
rect 44800 44600 44816 44664
rect 44880 44600 44896 44664
rect 44960 44600 44976 44664
rect 45040 44600 45056 44664
rect 45120 44600 45136 44664
rect 45200 44600 45216 44664
rect 45280 44600 45296 44664
rect 45360 44600 45368 44664
rect 41368 44584 45368 44600
rect 41368 44520 41376 44584
rect 41440 44520 41456 44584
rect 41520 44520 41536 44584
rect 41600 44520 41616 44584
rect 41680 44520 41696 44584
rect 41760 44520 41776 44584
rect 41840 44520 41856 44584
rect 41920 44520 41936 44584
rect 42000 44520 42016 44584
rect 42080 44520 42096 44584
rect 42160 44520 42176 44584
rect 42240 44520 42256 44584
rect 42320 44520 42336 44584
rect 42400 44520 42416 44584
rect 42480 44520 42496 44584
rect 42560 44520 42576 44584
rect 42640 44520 42656 44584
rect 42720 44520 42736 44584
rect 42800 44520 42816 44584
rect 42880 44520 42896 44584
rect 42960 44520 42976 44584
rect 43040 44520 43056 44584
rect 43120 44520 43136 44584
rect 43200 44520 43216 44584
rect 43280 44520 43296 44584
rect 43360 44520 43376 44584
rect 43440 44520 43456 44584
rect 43520 44520 43536 44584
rect 43600 44520 43616 44584
rect 43680 44520 43696 44584
rect 43760 44520 43776 44584
rect 43840 44520 43856 44584
rect 43920 44520 43936 44584
rect 44000 44520 44016 44584
rect 44080 44520 44096 44584
rect 44160 44520 44176 44584
rect 44240 44520 44256 44584
rect 44320 44520 44336 44584
rect 44400 44520 44416 44584
rect 44480 44520 44496 44584
rect 44560 44520 44576 44584
rect 44640 44520 44656 44584
rect 44720 44520 44736 44584
rect 44800 44520 44816 44584
rect 44880 44520 44896 44584
rect 44960 44520 44976 44584
rect 45040 44520 45056 44584
rect 45120 44520 45136 44584
rect 45200 44520 45216 44584
rect 45280 44520 45296 44584
rect 45360 44520 45368 44584
rect 41368 44504 45368 44520
rect 41368 44440 41376 44504
rect 41440 44440 41456 44504
rect 41520 44440 41536 44504
rect 41600 44440 41616 44504
rect 41680 44440 41696 44504
rect 41760 44440 41776 44504
rect 41840 44440 41856 44504
rect 41920 44440 41936 44504
rect 42000 44440 42016 44504
rect 42080 44440 42096 44504
rect 42160 44440 42176 44504
rect 42240 44440 42256 44504
rect 42320 44440 42336 44504
rect 42400 44440 42416 44504
rect 42480 44440 42496 44504
rect 42560 44440 42576 44504
rect 42640 44440 42656 44504
rect 42720 44440 42736 44504
rect 42800 44440 42816 44504
rect 42880 44440 42896 44504
rect 42960 44440 42976 44504
rect 43040 44440 43056 44504
rect 43120 44440 43136 44504
rect 43200 44440 43216 44504
rect 43280 44440 43296 44504
rect 43360 44440 43376 44504
rect 43440 44440 43456 44504
rect 43520 44440 43536 44504
rect 43600 44440 43616 44504
rect 43680 44440 43696 44504
rect 43760 44440 43776 44504
rect 43840 44440 43856 44504
rect 43920 44440 43936 44504
rect 44000 44440 44016 44504
rect 44080 44440 44096 44504
rect 44160 44440 44176 44504
rect 44240 44440 44256 44504
rect 44320 44440 44336 44504
rect 44400 44440 44416 44504
rect 44480 44440 44496 44504
rect 44560 44440 44576 44504
rect 44640 44440 44656 44504
rect 44720 44440 44736 44504
rect 44800 44440 44816 44504
rect 44880 44440 44896 44504
rect 44960 44440 44976 44504
rect 45040 44440 45056 44504
rect 45120 44440 45136 44504
rect 45200 44440 45216 44504
rect 45280 44440 45296 44504
rect 45360 44440 45368 44504
rect 41368 44424 45368 44440
rect 41368 44360 41376 44424
rect 41440 44360 41456 44424
rect 41520 44360 41536 44424
rect 41600 44360 41616 44424
rect 41680 44360 41696 44424
rect 41760 44360 41776 44424
rect 41840 44360 41856 44424
rect 41920 44360 41936 44424
rect 42000 44360 42016 44424
rect 42080 44360 42096 44424
rect 42160 44360 42176 44424
rect 42240 44360 42256 44424
rect 42320 44360 42336 44424
rect 42400 44360 42416 44424
rect 42480 44360 42496 44424
rect 42560 44360 42576 44424
rect 42640 44360 42656 44424
rect 42720 44360 42736 44424
rect 42800 44360 42816 44424
rect 42880 44360 42896 44424
rect 42960 44360 42976 44424
rect 43040 44360 43056 44424
rect 43120 44360 43136 44424
rect 43200 44360 43216 44424
rect 43280 44360 43296 44424
rect 43360 44360 43376 44424
rect 43440 44360 43456 44424
rect 43520 44360 43536 44424
rect 43600 44360 43616 44424
rect 43680 44360 43696 44424
rect 43760 44360 43776 44424
rect 43840 44360 43856 44424
rect 43920 44360 43936 44424
rect 44000 44360 44016 44424
rect 44080 44360 44096 44424
rect 44160 44360 44176 44424
rect 44240 44360 44256 44424
rect 44320 44360 44336 44424
rect 44400 44360 44416 44424
rect 44480 44360 44496 44424
rect 44560 44360 44576 44424
rect 44640 44360 44656 44424
rect 44720 44360 44736 44424
rect 44800 44360 44816 44424
rect 44880 44360 44896 44424
rect 44960 44360 44976 44424
rect 45040 44360 45056 44424
rect 45120 44360 45136 44424
rect 45200 44360 45216 44424
rect 45280 44360 45296 44424
rect 45360 44360 45368 44424
rect 41368 44344 45368 44360
rect 41368 44280 41376 44344
rect 41440 44280 41456 44344
rect 41520 44280 41536 44344
rect 41600 44280 41616 44344
rect 41680 44280 41696 44344
rect 41760 44280 41776 44344
rect 41840 44280 41856 44344
rect 41920 44280 41936 44344
rect 42000 44280 42016 44344
rect 42080 44280 42096 44344
rect 42160 44280 42176 44344
rect 42240 44280 42256 44344
rect 42320 44280 42336 44344
rect 42400 44280 42416 44344
rect 42480 44280 42496 44344
rect 42560 44280 42576 44344
rect 42640 44280 42656 44344
rect 42720 44280 42736 44344
rect 42800 44280 42816 44344
rect 42880 44280 42896 44344
rect 42960 44280 42976 44344
rect 43040 44280 43056 44344
rect 43120 44280 43136 44344
rect 43200 44280 43216 44344
rect 43280 44280 43296 44344
rect 43360 44280 43376 44344
rect 43440 44280 43456 44344
rect 43520 44280 43536 44344
rect 43600 44280 43616 44344
rect 43680 44280 43696 44344
rect 43760 44280 43776 44344
rect 43840 44280 43856 44344
rect 43920 44280 43936 44344
rect 44000 44280 44016 44344
rect 44080 44280 44096 44344
rect 44160 44280 44176 44344
rect 44240 44280 44256 44344
rect 44320 44280 44336 44344
rect 44400 44280 44416 44344
rect 44480 44280 44496 44344
rect 44560 44280 44576 44344
rect 44640 44280 44656 44344
rect 44720 44280 44736 44344
rect 44800 44280 44816 44344
rect 44880 44280 44896 44344
rect 44960 44280 44976 44344
rect 45040 44280 45056 44344
rect 45120 44280 45136 44344
rect 45200 44280 45216 44344
rect 45280 44280 45296 44344
rect 45360 44280 45368 44344
rect 41368 44264 45368 44280
rect 41368 44200 41376 44264
rect 41440 44200 41456 44264
rect 41520 44200 41536 44264
rect 41600 44200 41616 44264
rect 41680 44200 41696 44264
rect 41760 44200 41776 44264
rect 41840 44200 41856 44264
rect 41920 44200 41936 44264
rect 42000 44200 42016 44264
rect 42080 44200 42096 44264
rect 42160 44200 42176 44264
rect 42240 44200 42256 44264
rect 42320 44200 42336 44264
rect 42400 44200 42416 44264
rect 42480 44200 42496 44264
rect 42560 44200 42576 44264
rect 42640 44200 42656 44264
rect 42720 44200 42736 44264
rect 42800 44200 42816 44264
rect 42880 44200 42896 44264
rect 42960 44200 42976 44264
rect 43040 44200 43056 44264
rect 43120 44200 43136 44264
rect 43200 44200 43216 44264
rect 43280 44200 43296 44264
rect 43360 44200 43376 44264
rect 43440 44200 43456 44264
rect 43520 44200 43536 44264
rect 43600 44200 43616 44264
rect 43680 44200 43696 44264
rect 43760 44200 43776 44264
rect 43840 44200 43856 44264
rect 43920 44200 43936 44264
rect 44000 44200 44016 44264
rect 44080 44200 44096 44264
rect 44160 44200 44176 44264
rect 44240 44200 44256 44264
rect 44320 44200 44336 44264
rect 44400 44200 44416 44264
rect 44480 44200 44496 44264
rect 44560 44200 44576 44264
rect 44640 44200 44656 44264
rect 44720 44200 44736 44264
rect 44800 44200 44816 44264
rect 44880 44200 44896 44264
rect 44960 44200 44976 44264
rect 45040 44200 45056 44264
rect 45120 44200 45136 44264
rect 45200 44200 45216 44264
rect 45280 44200 45296 44264
rect 45360 44200 45368 44264
rect 41368 44184 45368 44200
rect 41368 44120 41376 44184
rect 41440 44120 41456 44184
rect 41520 44120 41536 44184
rect 41600 44120 41616 44184
rect 41680 44120 41696 44184
rect 41760 44120 41776 44184
rect 41840 44120 41856 44184
rect 41920 44120 41936 44184
rect 42000 44120 42016 44184
rect 42080 44120 42096 44184
rect 42160 44120 42176 44184
rect 42240 44120 42256 44184
rect 42320 44120 42336 44184
rect 42400 44120 42416 44184
rect 42480 44120 42496 44184
rect 42560 44120 42576 44184
rect 42640 44120 42656 44184
rect 42720 44120 42736 44184
rect 42800 44120 42816 44184
rect 42880 44120 42896 44184
rect 42960 44120 42976 44184
rect 43040 44120 43056 44184
rect 43120 44120 43136 44184
rect 43200 44120 43216 44184
rect 43280 44120 43296 44184
rect 43360 44120 43376 44184
rect 43440 44120 43456 44184
rect 43520 44120 43536 44184
rect 43600 44120 43616 44184
rect 43680 44120 43696 44184
rect 43760 44120 43776 44184
rect 43840 44120 43856 44184
rect 43920 44120 43936 44184
rect 44000 44120 44016 44184
rect 44080 44120 44096 44184
rect 44160 44120 44176 44184
rect 44240 44120 44256 44184
rect 44320 44120 44336 44184
rect 44400 44120 44416 44184
rect 44480 44120 44496 44184
rect 44560 44120 44576 44184
rect 44640 44120 44656 44184
rect 44720 44120 44736 44184
rect 44800 44120 44816 44184
rect 44880 44120 44896 44184
rect 44960 44120 44976 44184
rect 45040 44120 45056 44184
rect 45120 44120 45136 44184
rect 45200 44120 45216 44184
rect 45280 44120 45296 44184
rect 45360 44120 45368 44184
rect 41368 44104 45368 44120
rect 41368 44040 41376 44104
rect 41440 44040 41456 44104
rect 41520 44040 41536 44104
rect 41600 44040 41616 44104
rect 41680 44040 41696 44104
rect 41760 44040 41776 44104
rect 41840 44040 41856 44104
rect 41920 44040 41936 44104
rect 42000 44040 42016 44104
rect 42080 44040 42096 44104
rect 42160 44040 42176 44104
rect 42240 44040 42256 44104
rect 42320 44040 42336 44104
rect 42400 44040 42416 44104
rect 42480 44040 42496 44104
rect 42560 44040 42576 44104
rect 42640 44040 42656 44104
rect 42720 44040 42736 44104
rect 42800 44040 42816 44104
rect 42880 44040 42896 44104
rect 42960 44040 42976 44104
rect 43040 44040 43056 44104
rect 43120 44040 43136 44104
rect 43200 44040 43216 44104
rect 43280 44040 43296 44104
rect 43360 44040 43376 44104
rect 43440 44040 43456 44104
rect 43520 44040 43536 44104
rect 43600 44040 43616 44104
rect 43680 44040 43696 44104
rect 43760 44040 43776 44104
rect 43840 44040 43856 44104
rect 43920 44040 43936 44104
rect 44000 44040 44016 44104
rect 44080 44040 44096 44104
rect 44160 44040 44176 44104
rect 44240 44040 44256 44104
rect 44320 44040 44336 44104
rect 44400 44040 44416 44104
rect 44480 44040 44496 44104
rect 44560 44040 44576 44104
rect 44640 44040 44656 44104
rect 44720 44040 44736 44104
rect 44800 44040 44816 44104
rect 44880 44040 44896 44104
rect 44960 44040 44976 44104
rect 45040 44040 45056 44104
rect 45120 44040 45136 44104
rect 45200 44040 45216 44104
rect 45280 44040 45296 44104
rect 45360 44040 45368 44104
rect 41368 44024 45368 44040
rect 41368 43960 41376 44024
rect 41440 43960 41456 44024
rect 41520 43960 41536 44024
rect 41600 43960 41616 44024
rect 41680 43960 41696 44024
rect 41760 43960 41776 44024
rect 41840 43960 41856 44024
rect 41920 43960 41936 44024
rect 42000 43960 42016 44024
rect 42080 43960 42096 44024
rect 42160 43960 42176 44024
rect 42240 43960 42256 44024
rect 42320 43960 42336 44024
rect 42400 43960 42416 44024
rect 42480 43960 42496 44024
rect 42560 43960 42576 44024
rect 42640 43960 42656 44024
rect 42720 43960 42736 44024
rect 42800 43960 42816 44024
rect 42880 43960 42896 44024
rect 42960 43960 42976 44024
rect 43040 43960 43056 44024
rect 43120 43960 43136 44024
rect 43200 43960 43216 44024
rect 43280 43960 43296 44024
rect 43360 43960 43376 44024
rect 43440 43960 43456 44024
rect 43520 43960 43536 44024
rect 43600 43960 43616 44024
rect 43680 43960 43696 44024
rect 43760 43960 43776 44024
rect 43840 43960 43856 44024
rect 43920 43960 43936 44024
rect 44000 43960 44016 44024
rect 44080 43960 44096 44024
rect 44160 43960 44176 44024
rect 44240 43960 44256 44024
rect 44320 43960 44336 44024
rect 44400 43960 44416 44024
rect 44480 43960 44496 44024
rect 44560 43960 44576 44024
rect 44640 43960 44656 44024
rect 44720 43960 44736 44024
rect 44800 43960 44816 44024
rect 44880 43960 44896 44024
rect 44960 43960 44976 44024
rect 45040 43960 45056 44024
rect 45120 43960 45136 44024
rect 45200 43960 45216 44024
rect 45280 43960 45296 44024
rect 45360 43960 45368 44024
rect 41368 43944 45368 43960
rect 41368 43880 41376 43944
rect 41440 43880 41456 43944
rect 41520 43880 41536 43944
rect 41600 43880 41616 43944
rect 41680 43880 41696 43944
rect 41760 43880 41776 43944
rect 41840 43880 41856 43944
rect 41920 43880 41936 43944
rect 42000 43880 42016 43944
rect 42080 43880 42096 43944
rect 42160 43880 42176 43944
rect 42240 43880 42256 43944
rect 42320 43880 42336 43944
rect 42400 43880 42416 43944
rect 42480 43880 42496 43944
rect 42560 43880 42576 43944
rect 42640 43880 42656 43944
rect 42720 43880 42736 43944
rect 42800 43880 42816 43944
rect 42880 43880 42896 43944
rect 42960 43880 42976 43944
rect 43040 43880 43056 43944
rect 43120 43880 43136 43944
rect 43200 43880 43216 43944
rect 43280 43880 43296 43944
rect 43360 43880 43376 43944
rect 43440 43880 43456 43944
rect 43520 43880 43536 43944
rect 43600 43880 43616 43944
rect 43680 43880 43696 43944
rect 43760 43880 43776 43944
rect 43840 43880 43856 43944
rect 43920 43880 43936 43944
rect 44000 43880 44016 43944
rect 44080 43880 44096 43944
rect 44160 43880 44176 43944
rect 44240 43880 44256 43944
rect 44320 43880 44336 43944
rect 44400 43880 44416 43944
rect 44480 43880 44496 43944
rect 44560 43880 44576 43944
rect 44640 43880 44656 43944
rect 44720 43880 44736 43944
rect 44800 43880 44816 43944
rect 44880 43880 44896 43944
rect 44960 43880 44976 43944
rect 45040 43880 45056 43944
rect 45120 43880 45136 43944
rect 45200 43880 45216 43944
rect 45280 43880 45296 43944
rect 45360 43880 45368 43944
rect 41368 43864 45368 43880
rect 41368 43800 41376 43864
rect 41440 43800 41456 43864
rect 41520 43800 41536 43864
rect 41600 43800 41616 43864
rect 41680 43800 41696 43864
rect 41760 43800 41776 43864
rect 41840 43800 41856 43864
rect 41920 43800 41936 43864
rect 42000 43800 42016 43864
rect 42080 43800 42096 43864
rect 42160 43800 42176 43864
rect 42240 43800 42256 43864
rect 42320 43800 42336 43864
rect 42400 43800 42416 43864
rect 42480 43800 42496 43864
rect 42560 43800 42576 43864
rect 42640 43800 42656 43864
rect 42720 43800 42736 43864
rect 42800 43800 42816 43864
rect 42880 43800 42896 43864
rect 42960 43800 42976 43864
rect 43040 43800 43056 43864
rect 43120 43800 43136 43864
rect 43200 43800 43216 43864
rect 43280 43800 43296 43864
rect 43360 43800 43376 43864
rect 43440 43800 43456 43864
rect 43520 43800 43536 43864
rect 43600 43800 43616 43864
rect 43680 43800 43696 43864
rect 43760 43800 43776 43864
rect 43840 43800 43856 43864
rect 43920 43800 43936 43864
rect 44000 43800 44016 43864
rect 44080 43800 44096 43864
rect 44160 43800 44176 43864
rect 44240 43800 44256 43864
rect 44320 43800 44336 43864
rect 44400 43800 44416 43864
rect 44480 43800 44496 43864
rect 44560 43800 44576 43864
rect 44640 43800 44656 43864
rect 44720 43800 44736 43864
rect 44800 43800 44816 43864
rect 44880 43800 44896 43864
rect 44960 43800 44976 43864
rect 45040 43800 45056 43864
rect 45120 43800 45136 43864
rect 45200 43800 45216 43864
rect 45280 43800 45296 43864
rect 45360 43800 45368 43864
rect 41368 43784 45368 43800
rect 41368 43720 41376 43784
rect 41440 43720 41456 43784
rect 41520 43720 41536 43784
rect 41600 43720 41616 43784
rect 41680 43720 41696 43784
rect 41760 43720 41776 43784
rect 41840 43720 41856 43784
rect 41920 43720 41936 43784
rect 42000 43720 42016 43784
rect 42080 43720 42096 43784
rect 42160 43720 42176 43784
rect 42240 43720 42256 43784
rect 42320 43720 42336 43784
rect 42400 43720 42416 43784
rect 42480 43720 42496 43784
rect 42560 43720 42576 43784
rect 42640 43720 42656 43784
rect 42720 43720 42736 43784
rect 42800 43720 42816 43784
rect 42880 43720 42896 43784
rect 42960 43720 42976 43784
rect 43040 43720 43056 43784
rect 43120 43720 43136 43784
rect 43200 43720 43216 43784
rect 43280 43720 43296 43784
rect 43360 43720 43376 43784
rect 43440 43720 43456 43784
rect 43520 43720 43536 43784
rect 43600 43720 43616 43784
rect 43680 43720 43696 43784
rect 43760 43720 43776 43784
rect 43840 43720 43856 43784
rect 43920 43720 43936 43784
rect 44000 43720 44016 43784
rect 44080 43720 44096 43784
rect 44160 43720 44176 43784
rect 44240 43720 44256 43784
rect 44320 43720 44336 43784
rect 44400 43720 44416 43784
rect 44480 43720 44496 43784
rect 44560 43720 44576 43784
rect 44640 43720 44656 43784
rect 44720 43720 44736 43784
rect 44800 43720 44816 43784
rect 44880 43720 44896 43784
rect 44960 43720 44976 43784
rect 45040 43720 45056 43784
rect 45120 43720 45136 43784
rect 45200 43720 45216 43784
rect 45280 43720 45296 43784
rect 45360 43720 45368 43784
rect 41368 43704 45368 43720
rect 41368 43640 41376 43704
rect 41440 43640 41456 43704
rect 41520 43640 41536 43704
rect 41600 43640 41616 43704
rect 41680 43640 41696 43704
rect 41760 43640 41776 43704
rect 41840 43640 41856 43704
rect 41920 43640 41936 43704
rect 42000 43640 42016 43704
rect 42080 43640 42096 43704
rect 42160 43640 42176 43704
rect 42240 43640 42256 43704
rect 42320 43640 42336 43704
rect 42400 43640 42416 43704
rect 42480 43640 42496 43704
rect 42560 43640 42576 43704
rect 42640 43640 42656 43704
rect 42720 43640 42736 43704
rect 42800 43640 42816 43704
rect 42880 43640 42896 43704
rect 42960 43640 42976 43704
rect 43040 43640 43056 43704
rect 43120 43640 43136 43704
rect 43200 43640 43216 43704
rect 43280 43640 43296 43704
rect 43360 43640 43376 43704
rect 43440 43640 43456 43704
rect 43520 43640 43536 43704
rect 43600 43640 43616 43704
rect 43680 43640 43696 43704
rect 43760 43640 43776 43704
rect 43840 43640 43856 43704
rect 43920 43640 43936 43704
rect 44000 43640 44016 43704
rect 44080 43640 44096 43704
rect 44160 43640 44176 43704
rect 44240 43640 44256 43704
rect 44320 43640 44336 43704
rect 44400 43640 44416 43704
rect 44480 43640 44496 43704
rect 44560 43640 44576 43704
rect 44640 43640 44656 43704
rect 44720 43640 44736 43704
rect 44800 43640 44816 43704
rect 44880 43640 44896 43704
rect 44960 43640 44976 43704
rect 45040 43640 45056 43704
rect 45120 43640 45136 43704
rect 45200 43640 45216 43704
rect 45280 43640 45296 43704
rect 45360 43640 45368 43704
rect 41368 43624 45368 43640
rect 41368 43560 41376 43624
rect 41440 43560 41456 43624
rect 41520 43560 41536 43624
rect 41600 43560 41616 43624
rect 41680 43560 41696 43624
rect 41760 43560 41776 43624
rect 41840 43560 41856 43624
rect 41920 43560 41936 43624
rect 42000 43560 42016 43624
rect 42080 43560 42096 43624
rect 42160 43560 42176 43624
rect 42240 43560 42256 43624
rect 42320 43560 42336 43624
rect 42400 43560 42416 43624
rect 42480 43560 42496 43624
rect 42560 43560 42576 43624
rect 42640 43560 42656 43624
rect 42720 43560 42736 43624
rect 42800 43560 42816 43624
rect 42880 43560 42896 43624
rect 42960 43560 42976 43624
rect 43040 43560 43056 43624
rect 43120 43560 43136 43624
rect 43200 43560 43216 43624
rect 43280 43560 43296 43624
rect 43360 43560 43376 43624
rect 43440 43560 43456 43624
rect 43520 43560 43536 43624
rect 43600 43560 43616 43624
rect 43680 43560 43696 43624
rect 43760 43560 43776 43624
rect 43840 43560 43856 43624
rect 43920 43560 43936 43624
rect 44000 43560 44016 43624
rect 44080 43560 44096 43624
rect 44160 43560 44176 43624
rect 44240 43560 44256 43624
rect 44320 43560 44336 43624
rect 44400 43560 44416 43624
rect 44480 43560 44496 43624
rect 44560 43560 44576 43624
rect 44640 43560 44656 43624
rect 44720 43560 44736 43624
rect 44800 43560 44816 43624
rect 44880 43560 44896 43624
rect 44960 43560 44976 43624
rect 45040 43560 45056 43624
rect 45120 43560 45136 43624
rect 45200 43560 45216 43624
rect 45280 43560 45296 43624
rect 45360 43560 45368 43624
rect 41368 43544 45368 43560
rect 41368 43480 41376 43544
rect 41440 43480 41456 43544
rect 41520 43480 41536 43544
rect 41600 43480 41616 43544
rect 41680 43480 41696 43544
rect 41760 43480 41776 43544
rect 41840 43480 41856 43544
rect 41920 43480 41936 43544
rect 42000 43480 42016 43544
rect 42080 43480 42096 43544
rect 42160 43480 42176 43544
rect 42240 43480 42256 43544
rect 42320 43480 42336 43544
rect 42400 43480 42416 43544
rect 42480 43480 42496 43544
rect 42560 43480 42576 43544
rect 42640 43480 42656 43544
rect 42720 43480 42736 43544
rect 42800 43480 42816 43544
rect 42880 43480 42896 43544
rect 42960 43480 42976 43544
rect 43040 43480 43056 43544
rect 43120 43480 43136 43544
rect 43200 43480 43216 43544
rect 43280 43480 43296 43544
rect 43360 43480 43376 43544
rect 43440 43480 43456 43544
rect 43520 43480 43536 43544
rect 43600 43480 43616 43544
rect 43680 43480 43696 43544
rect 43760 43480 43776 43544
rect 43840 43480 43856 43544
rect 43920 43480 43936 43544
rect 44000 43480 44016 43544
rect 44080 43480 44096 43544
rect 44160 43480 44176 43544
rect 44240 43480 44256 43544
rect 44320 43480 44336 43544
rect 44400 43480 44416 43544
rect 44480 43480 44496 43544
rect 44560 43480 44576 43544
rect 44640 43480 44656 43544
rect 44720 43480 44736 43544
rect 44800 43480 44816 43544
rect 44880 43480 44896 43544
rect 44960 43480 44976 43544
rect 45040 43480 45056 43544
rect 45120 43480 45136 43544
rect 45200 43480 45216 43544
rect 45280 43480 45296 43544
rect 45360 43480 45368 43544
rect 41368 43464 45368 43480
rect 41368 43400 41376 43464
rect 41440 43400 41456 43464
rect 41520 43400 41536 43464
rect 41600 43400 41616 43464
rect 41680 43400 41696 43464
rect 41760 43400 41776 43464
rect 41840 43400 41856 43464
rect 41920 43400 41936 43464
rect 42000 43400 42016 43464
rect 42080 43400 42096 43464
rect 42160 43400 42176 43464
rect 42240 43400 42256 43464
rect 42320 43400 42336 43464
rect 42400 43400 42416 43464
rect 42480 43400 42496 43464
rect 42560 43400 42576 43464
rect 42640 43400 42656 43464
rect 42720 43400 42736 43464
rect 42800 43400 42816 43464
rect 42880 43400 42896 43464
rect 42960 43400 42976 43464
rect 43040 43400 43056 43464
rect 43120 43400 43136 43464
rect 43200 43400 43216 43464
rect 43280 43400 43296 43464
rect 43360 43400 43376 43464
rect 43440 43400 43456 43464
rect 43520 43400 43536 43464
rect 43600 43400 43616 43464
rect 43680 43400 43696 43464
rect 43760 43400 43776 43464
rect 43840 43400 43856 43464
rect 43920 43400 43936 43464
rect 44000 43400 44016 43464
rect 44080 43400 44096 43464
rect 44160 43400 44176 43464
rect 44240 43400 44256 43464
rect 44320 43400 44336 43464
rect 44400 43400 44416 43464
rect 44480 43400 44496 43464
rect 44560 43400 44576 43464
rect 44640 43400 44656 43464
rect 44720 43400 44736 43464
rect 44800 43400 44816 43464
rect 44880 43400 44896 43464
rect 44960 43400 44976 43464
rect 45040 43400 45056 43464
rect 45120 43400 45136 43464
rect 45200 43400 45216 43464
rect 45280 43400 45296 43464
rect 45360 43400 45368 43464
rect 41368 43384 45368 43400
rect 41368 43320 41376 43384
rect 41440 43320 41456 43384
rect 41520 43320 41536 43384
rect 41600 43320 41616 43384
rect 41680 43320 41696 43384
rect 41760 43320 41776 43384
rect 41840 43320 41856 43384
rect 41920 43320 41936 43384
rect 42000 43320 42016 43384
rect 42080 43320 42096 43384
rect 42160 43320 42176 43384
rect 42240 43320 42256 43384
rect 42320 43320 42336 43384
rect 42400 43320 42416 43384
rect 42480 43320 42496 43384
rect 42560 43320 42576 43384
rect 42640 43320 42656 43384
rect 42720 43320 42736 43384
rect 42800 43320 42816 43384
rect 42880 43320 42896 43384
rect 42960 43320 42976 43384
rect 43040 43320 43056 43384
rect 43120 43320 43136 43384
rect 43200 43320 43216 43384
rect 43280 43320 43296 43384
rect 43360 43320 43376 43384
rect 43440 43320 43456 43384
rect 43520 43320 43536 43384
rect 43600 43320 43616 43384
rect 43680 43320 43696 43384
rect 43760 43320 43776 43384
rect 43840 43320 43856 43384
rect 43920 43320 43936 43384
rect 44000 43320 44016 43384
rect 44080 43320 44096 43384
rect 44160 43320 44176 43384
rect 44240 43320 44256 43384
rect 44320 43320 44336 43384
rect 44400 43320 44416 43384
rect 44480 43320 44496 43384
rect 44560 43320 44576 43384
rect 44640 43320 44656 43384
rect 44720 43320 44736 43384
rect 44800 43320 44816 43384
rect 44880 43320 44896 43384
rect 44960 43320 44976 43384
rect 45040 43320 45056 43384
rect 45120 43320 45136 43384
rect 45200 43320 45216 43384
rect 45280 43320 45296 43384
rect 45360 43320 45368 43384
rect 41368 43304 45368 43320
rect 41368 43240 41376 43304
rect 41440 43240 41456 43304
rect 41520 43240 41536 43304
rect 41600 43240 41616 43304
rect 41680 43240 41696 43304
rect 41760 43240 41776 43304
rect 41840 43240 41856 43304
rect 41920 43240 41936 43304
rect 42000 43240 42016 43304
rect 42080 43240 42096 43304
rect 42160 43240 42176 43304
rect 42240 43240 42256 43304
rect 42320 43240 42336 43304
rect 42400 43240 42416 43304
rect 42480 43240 42496 43304
rect 42560 43240 42576 43304
rect 42640 43240 42656 43304
rect 42720 43240 42736 43304
rect 42800 43240 42816 43304
rect 42880 43240 42896 43304
rect 42960 43240 42976 43304
rect 43040 43240 43056 43304
rect 43120 43240 43136 43304
rect 43200 43240 43216 43304
rect 43280 43240 43296 43304
rect 43360 43240 43376 43304
rect 43440 43240 43456 43304
rect 43520 43240 43536 43304
rect 43600 43240 43616 43304
rect 43680 43240 43696 43304
rect 43760 43240 43776 43304
rect 43840 43240 43856 43304
rect 43920 43240 43936 43304
rect 44000 43240 44016 43304
rect 44080 43240 44096 43304
rect 44160 43240 44176 43304
rect 44240 43240 44256 43304
rect 44320 43240 44336 43304
rect 44400 43240 44416 43304
rect 44480 43240 44496 43304
rect 44560 43240 44576 43304
rect 44640 43240 44656 43304
rect 44720 43240 44736 43304
rect 44800 43240 44816 43304
rect 44880 43240 44896 43304
rect 44960 43240 44976 43304
rect 45040 43240 45056 43304
rect 45120 43240 45136 43304
rect 45200 43240 45216 43304
rect 45280 43240 45296 43304
rect 45360 43240 45368 43304
rect 41368 43224 45368 43240
rect 41368 43160 41376 43224
rect 41440 43160 41456 43224
rect 41520 43160 41536 43224
rect 41600 43160 41616 43224
rect 41680 43160 41696 43224
rect 41760 43160 41776 43224
rect 41840 43160 41856 43224
rect 41920 43160 41936 43224
rect 42000 43160 42016 43224
rect 42080 43160 42096 43224
rect 42160 43160 42176 43224
rect 42240 43160 42256 43224
rect 42320 43160 42336 43224
rect 42400 43160 42416 43224
rect 42480 43160 42496 43224
rect 42560 43160 42576 43224
rect 42640 43160 42656 43224
rect 42720 43160 42736 43224
rect 42800 43160 42816 43224
rect 42880 43160 42896 43224
rect 42960 43160 42976 43224
rect 43040 43160 43056 43224
rect 43120 43160 43136 43224
rect 43200 43160 43216 43224
rect 43280 43160 43296 43224
rect 43360 43160 43376 43224
rect 43440 43160 43456 43224
rect 43520 43160 43536 43224
rect 43600 43160 43616 43224
rect 43680 43160 43696 43224
rect 43760 43160 43776 43224
rect 43840 43160 43856 43224
rect 43920 43160 43936 43224
rect 44000 43160 44016 43224
rect 44080 43160 44096 43224
rect 44160 43160 44176 43224
rect 44240 43160 44256 43224
rect 44320 43160 44336 43224
rect 44400 43160 44416 43224
rect 44480 43160 44496 43224
rect 44560 43160 44576 43224
rect 44640 43160 44656 43224
rect 44720 43160 44736 43224
rect 44800 43160 44816 43224
rect 44880 43160 44896 43224
rect 44960 43160 44976 43224
rect 45040 43160 45056 43224
rect 45120 43160 45136 43224
rect 45200 43160 45216 43224
rect 45280 43160 45296 43224
rect 45360 43160 45368 43224
rect 41368 43144 45368 43160
rect 41368 43080 41376 43144
rect 41440 43080 41456 43144
rect 41520 43080 41536 43144
rect 41600 43080 41616 43144
rect 41680 43080 41696 43144
rect 41760 43080 41776 43144
rect 41840 43080 41856 43144
rect 41920 43080 41936 43144
rect 42000 43080 42016 43144
rect 42080 43080 42096 43144
rect 42160 43080 42176 43144
rect 42240 43080 42256 43144
rect 42320 43080 42336 43144
rect 42400 43080 42416 43144
rect 42480 43080 42496 43144
rect 42560 43080 42576 43144
rect 42640 43080 42656 43144
rect 42720 43080 42736 43144
rect 42800 43080 42816 43144
rect 42880 43080 42896 43144
rect 42960 43080 42976 43144
rect 43040 43080 43056 43144
rect 43120 43080 43136 43144
rect 43200 43080 43216 43144
rect 43280 43080 43296 43144
rect 43360 43080 43376 43144
rect 43440 43080 43456 43144
rect 43520 43080 43536 43144
rect 43600 43080 43616 43144
rect 43680 43080 43696 43144
rect 43760 43080 43776 43144
rect 43840 43080 43856 43144
rect 43920 43080 43936 43144
rect 44000 43080 44016 43144
rect 44080 43080 44096 43144
rect 44160 43080 44176 43144
rect 44240 43080 44256 43144
rect 44320 43080 44336 43144
rect 44400 43080 44416 43144
rect 44480 43080 44496 43144
rect 44560 43080 44576 43144
rect 44640 43080 44656 43144
rect 44720 43080 44736 43144
rect 44800 43080 44816 43144
rect 44880 43080 44896 43144
rect 44960 43080 44976 43144
rect 45040 43080 45056 43144
rect 45120 43080 45136 43144
rect 45200 43080 45216 43144
rect 45280 43080 45296 43144
rect 45360 43080 45368 43144
rect 41368 43064 45368 43080
rect 41368 43000 41376 43064
rect 41440 43000 41456 43064
rect 41520 43000 41536 43064
rect 41600 43000 41616 43064
rect 41680 43000 41696 43064
rect 41760 43000 41776 43064
rect 41840 43000 41856 43064
rect 41920 43000 41936 43064
rect 42000 43000 42016 43064
rect 42080 43000 42096 43064
rect 42160 43000 42176 43064
rect 42240 43000 42256 43064
rect 42320 43000 42336 43064
rect 42400 43000 42416 43064
rect 42480 43000 42496 43064
rect 42560 43000 42576 43064
rect 42640 43000 42656 43064
rect 42720 43000 42736 43064
rect 42800 43000 42816 43064
rect 42880 43000 42896 43064
rect 42960 43000 42976 43064
rect 43040 43000 43056 43064
rect 43120 43000 43136 43064
rect 43200 43000 43216 43064
rect 43280 43000 43296 43064
rect 43360 43000 43376 43064
rect 43440 43000 43456 43064
rect 43520 43000 43536 43064
rect 43600 43000 43616 43064
rect 43680 43000 43696 43064
rect 43760 43000 43776 43064
rect 43840 43000 43856 43064
rect 43920 43000 43936 43064
rect 44000 43000 44016 43064
rect 44080 43000 44096 43064
rect 44160 43000 44176 43064
rect 44240 43000 44256 43064
rect 44320 43000 44336 43064
rect 44400 43000 44416 43064
rect 44480 43000 44496 43064
rect 44560 43000 44576 43064
rect 44640 43000 44656 43064
rect 44720 43000 44736 43064
rect 44800 43000 44816 43064
rect 44880 43000 44896 43064
rect 44960 43000 44976 43064
rect 45040 43000 45056 43064
rect 45120 43000 45136 43064
rect 45200 43000 45216 43064
rect 45280 43000 45296 43064
rect 45360 43000 45368 43064
rect 41368 42984 45368 43000
rect 41368 42920 41376 42984
rect 41440 42920 41456 42984
rect 41520 42920 41536 42984
rect 41600 42920 41616 42984
rect 41680 42920 41696 42984
rect 41760 42920 41776 42984
rect 41840 42920 41856 42984
rect 41920 42920 41936 42984
rect 42000 42920 42016 42984
rect 42080 42920 42096 42984
rect 42160 42920 42176 42984
rect 42240 42920 42256 42984
rect 42320 42920 42336 42984
rect 42400 42920 42416 42984
rect 42480 42920 42496 42984
rect 42560 42920 42576 42984
rect 42640 42920 42656 42984
rect 42720 42920 42736 42984
rect 42800 42920 42816 42984
rect 42880 42920 42896 42984
rect 42960 42920 42976 42984
rect 43040 42920 43056 42984
rect 43120 42920 43136 42984
rect 43200 42920 43216 42984
rect 43280 42920 43296 42984
rect 43360 42920 43376 42984
rect 43440 42920 43456 42984
rect 43520 42920 43536 42984
rect 43600 42920 43616 42984
rect 43680 42920 43696 42984
rect 43760 42920 43776 42984
rect 43840 42920 43856 42984
rect 43920 42920 43936 42984
rect 44000 42920 44016 42984
rect 44080 42920 44096 42984
rect 44160 42920 44176 42984
rect 44240 42920 44256 42984
rect 44320 42920 44336 42984
rect 44400 42920 44416 42984
rect 44480 42920 44496 42984
rect 44560 42920 44576 42984
rect 44640 42920 44656 42984
rect 44720 42920 44736 42984
rect 44800 42920 44816 42984
rect 44880 42920 44896 42984
rect 44960 42920 44976 42984
rect 45040 42920 45056 42984
rect 45120 42920 45136 42984
rect 45200 42920 45216 42984
rect 45280 42920 45296 42984
rect 45360 42920 45368 42984
rect 41368 42904 45368 42920
rect 41368 42840 41376 42904
rect 41440 42840 41456 42904
rect 41520 42840 41536 42904
rect 41600 42840 41616 42904
rect 41680 42840 41696 42904
rect 41760 42840 41776 42904
rect 41840 42840 41856 42904
rect 41920 42840 41936 42904
rect 42000 42840 42016 42904
rect 42080 42840 42096 42904
rect 42160 42840 42176 42904
rect 42240 42840 42256 42904
rect 42320 42840 42336 42904
rect 42400 42840 42416 42904
rect 42480 42840 42496 42904
rect 42560 42840 42576 42904
rect 42640 42840 42656 42904
rect 42720 42840 42736 42904
rect 42800 42840 42816 42904
rect 42880 42840 42896 42904
rect 42960 42840 42976 42904
rect 43040 42840 43056 42904
rect 43120 42840 43136 42904
rect 43200 42840 43216 42904
rect 43280 42840 43296 42904
rect 43360 42840 43376 42904
rect 43440 42840 43456 42904
rect 43520 42840 43536 42904
rect 43600 42840 43616 42904
rect 43680 42840 43696 42904
rect 43760 42840 43776 42904
rect 43840 42840 43856 42904
rect 43920 42840 43936 42904
rect 44000 42840 44016 42904
rect 44080 42840 44096 42904
rect 44160 42840 44176 42904
rect 44240 42840 44256 42904
rect 44320 42840 44336 42904
rect 44400 42840 44416 42904
rect 44480 42840 44496 42904
rect 44560 42840 44576 42904
rect 44640 42840 44656 42904
rect 44720 42840 44736 42904
rect 44800 42840 44816 42904
rect 44880 42840 44896 42904
rect 44960 42840 44976 42904
rect 45040 42840 45056 42904
rect 45120 42840 45136 42904
rect 45200 42840 45216 42904
rect 45280 42840 45296 42904
rect 45360 42840 45368 42904
rect 41368 42824 45368 42840
rect 41368 42760 41376 42824
rect 41440 42760 41456 42824
rect 41520 42760 41536 42824
rect 41600 42760 41616 42824
rect 41680 42760 41696 42824
rect 41760 42760 41776 42824
rect 41840 42760 41856 42824
rect 41920 42760 41936 42824
rect 42000 42760 42016 42824
rect 42080 42760 42096 42824
rect 42160 42760 42176 42824
rect 42240 42760 42256 42824
rect 42320 42760 42336 42824
rect 42400 42760 42416 42824
rect 42480 42760 42496 42824
rect 42560 42760 42576 42824
rect 42640 42760 42656 42824
rect 42720 42760 42736 42824
rect 42800 42760 42816 42824
rect 42880 42760 42896 42824
rect 42960 42760 42976 42824
rect 43040 42760 43056 42824
rect 43120 42760 43136 42824
rect 43200 42760 43216 42824
rect 43280 42760 43296 42824
rect 43360 42760 43376 42824
rect 43440 42760 43456 42824
rect 43520 42760 43536 42824
rect 43600 42760 43616 42824
rect 43680 42760 43696 42824
rect 43760 42760 43776 42824
rect 43840 42760 43856 42824
rect 43920 42760 43936 42824
rect 44000 42760 44016 42824
rect 44080 42760 44096 42824
rect 44160 42760 44176 42824
rect 44240 42760 44256 42824
rect 44320 42760 44336 42824
rect 44400 42760 44416 42824
rect 44480 42760 44496 42824
rect 44560 42760 44576 42824
rect 44640 42760 44656 42824
rect 44720 42760 44736 42824
rect 44800 42760 44816 42824
rect 44880 42760 44896 42824
rect 44960 42760 44976 42824
rect 45040 42760 45056 42824
rect 45120 42760 45136 42824
rect 45200 42760 45216 42824
rect 45280 42760 45296 42824
rect 45360 42760 45368 42824
rect 41368 42744 45368 42760
rect 41368 42680 41376 42744
rect 41440 42680 41456 42744
rect 41520 42680 41536 42744
rect 41600 42680 41616 42744
rect 41680 42680 41696 42744
rect 41760 42680 41776 42744
rect 41840 42680 41856 42744
rect 41920 42680 41936 42744
rect 42000 42680 42016 42744
rect 42080 42680 42096 42744
rect 42160 42680 42176 42744
rect 42240 42680 42256 42744
rect 42320 42680 42336 42744
rect 42400 42680 42416 42744
rect 42480 42680 42496 42744
rect 42560 42680 42576 42744
rect 42640 42680 42656 42744
rect 42720 42680 42736 42744
rect 42800 42680 42816 42744
rect 42880 42680 42896 42744
rect 42960 42680 42976 42744
rect 43040 42680 43056 42744
rect 43120 42680 43136 42744
rect 43200 42680 43216 42744
rect 43280 42680 43296 42744
rect 43360 42680 43376 42744
rect 43440 42680 43456 42744
rect 43520 42680 43536 42744
rect 43600 42680 43616 42744
rect 43680 42680 43696 42744
rect 43760 42680 43776 42744
rect 43840 42680 43856 42744
rect 43920 42680 43936 42744
rect 44000 42680 44016 42744
rect 44080 42680 44096 42744
rect 44160 42680 44176 42744
rect 44240 42680 44256 42744
rect 44320 42680 44336 42744
rect 44400 42680 44416 42744
rect 44480 42680 44496 42744
rect 44560 42680 44576 42744
rect 44640 42680 44656 42744
rect 44720 42680 44736 42744
rect 44800 42680 44816 42744
rect 44880 42680 44896 42744
rect 44960 42680 44976 42744
rect 45040 42680 45056 42744
rect 45120 42680 45136 42744
rect 45200 42680 45216 42744
rect 45280 42680 45296 42744
rect 45360 42680 45368 42744
rect 41368 42664 45368 42680
rect 41368 42600 41376 42664
rect 41440 42600 41456 42664
rect 41520 42600 41536 42664
rect 41600 42600 41616 42664
rect 41680 42600 41696 42664
rect 41760 42600 41776 42664
rect 41840 42600 41856 42664
rect 41920 42600 41936 42664
rect 42000 42600 42016 42664
rect 42080 42600 42096 42664
rect 42160 42600 42176 42664
rect 42240 42600 42256 42664
rect 42320 42600 42336 42664
rect 42400 42600 42416 42664
rect 42480 42600 42496 42664
rect 42560 42600 42576 42664
rect 42640 42600 42656 42664
rect 42720 42600 42736 42664
rect 42800 42600 42816 42664
rect 42880 42600 42896 42664
rect 42960 42600 42976 42664
rect 43040 42600 43056 42664
rect 43120 42600 43136 42664
rect 43200 42600 43216 42664
rect 43280 42600 43296 42664
rect 43360 42600 43376 42664
rect 43440 42600 43456 42664
rect 43520 42600 43536 42664
rect 43600 42600 43616 42664
rect 43680 42600 43696 42664
rect 43760 42600 43776 42664
rect 43840 42600 43856 42664
rect 43920 42600 43936 42664
rect 44000 42600 44016 42664
rect 44080 42600 44096 42664
rect 44160 42600 44176 42664
rect 44240 42600 44256 42664
rect 44320 42600 44336 42664
rect 44400 42600 44416 42664
rect 44480 42600 44496 42664
rect 44560 42600 44576 42664
rect 44640 42600 44656 42664
rect 44720 42600 44736 42664
rect 44800 42600 44816 42664
rect 44880 42600 44896 42664
rect 44960 42600 44976 42664
rect 45040 42600 45056 42664
rect 45120 42600 45136 42664
rect 45200 42600 45216 42664
rect 45280 42600 45296 42664
rect 45360 42600 45368 42664
rect 41368 42584 45368 42600
rect 41368 42520 41376 42584
rect 41440 42520 41456 42584
rect 41520 42520 41536 42584
rect 41600 42520 41616 42584
rect 41680 42520 41696 42584
rect 41760 42520 41776 42584
rect 41840 42520 41856 42584
rect 41920 42520 41936 42584
rect 42000 42520 42016 42584
rect 42080 42520 42096 42584
rect 42160 42520 42176 42584
rect 42240 42520 42256 42584
rect 42320 42520 42336 42584
rect 42400 42520 42416 42584
rect 42480 42520 42496 42584
rect 42560 42520 42576 42584
rect 42640 42520 42656 42584
rect 42720 42520 42736 42584
rect 42800 42520 42816 42584
rect 42880 42520 42896 42584
rect 42960 42520 42976 42584
rect 43040 42520 43056 42584
rect 43120 42520 43136 42584
rect 43200 42520 43216 42584
rect 43280 42520 43296 42584
rect 43360 42520 43376 42584
rect 43440 42520 43456 42584
rect 43520 42520 43536 42584
rect 43600 42520 43616 42584
rect 43680 42520 43696 42584
rect 43760 42520 43776 42584
rect 43840 42520 43856 42584
rect 43920 42520 43936 42584
rect 44000 42520 44016 42584
rect 44080 42520 44096 42584
rect 44160 42520 44176 42584
rect 44240 42520 44256 42584
rect 44320 42520 44336 42584
rect 44400 42520 44416 42584
rect 44480 42520 44496 42584
rect 44560 42520 44576 42584
rect 44640 42520 44656 42584
rect 44720 42520 44736 42584
rect 44800 42520 44816 42584
rect 44880 42520 44896 42584
rect 44960 42520 44976 42584
rect 45040 42520 45056 42584
rect 45120 42520 45136 42584
rect 45200 42520 45216 42584
rect 45280 42520 45296 42584
rect 45360 42520 45368 42584
rect 41368 42504 45368 42520
rect 41368 42440 41376 42504
rect 41440 42440 41456 42504
rect 41520 42440 41536 42504
rect 41600 42440 41616 42504
rect 41680 42440 41696 42504
rect 41760 42440 41776 42504
rect 41840 42440 41856 42504
rect 41920 42440 41936 42504
rect 42000 42440 42016 42504
rect 42080 42440 42096 42504
rect 42160 42440 42176 42504
rect 42240 42440 42256 42504
rect 42320 42440 42336 42504
rect 42400 42440 42416 42504
rect 42480 42440 42496 42504
rect 42560 42440 42576 42504
rect 42640 42440 42656 42504
rect 42720 42440 42736 42504
rect 42800 42440 42816 42504
rect 42880 42440 42896 42504
rect 42960 42440 42976 42504
rect 43040 42440 43056 42504
rect 43120 42440 43136 42504
rect 43200 42440 43216 42504
rect 43280 42440 43296 42504
rect 43360 42440 43376 42504
rect 43440 42440 43456 42504
rect 43520 42440 43536 42504
rect 43600 42440 43616 42504
rect 43680 42440 43696 42504
rect 43760 42440 43776 42504
rect 43840 42440 43856 42504
rect 43920 42440 43936 42504
rect 44000 42440 44016 42504
rect 44080 42440 44096 42504
rect 44160 42440 44176 42504
rect 44240 42440 44256 42504
rect 44320 42440 44336 42504
rect 44400 42440 44416 42504
rect 44480 42440 44496 42504
rect 44560 42440 44576 42504
rect 44640 42440 44656 42504
rect 44720 42440 44736 42504
rect 44800 42440 44816 42504
rect 44880 42440 44896 42504
rect 44960 42440 44976 42504
rect 45040 42440 45056 42504
rect 45120 42440 45136 42504
rect 45200 42440 45216 42504
rect 45280 42440 45296 42504
rect 45360 42440 45368 42504
rect 41368 42424 45368 42440
rect 41368 42360 41376 42424
rect 41440 42360 41456 42424
rect 41520 42360 41536 42424
rect 41600 42360 41616 42424
rect 41680 42360 41696 42424
rect 41760 42360 41776 42424
rect 41840 42360 41856 42424
rect 41920 42360 41936 42424
rect 42000 42360 42016 42424
rect 42080 42360 42096 42424
rect 42160 42360 42176 42424
rect 42240 42360 42256 42424
rect 42320 42360 42336 42424
rect 42400 42360 42416 42424
rect 42480 42360 42496 42424
rect 42560 42360 42576 42424
rect 42640 42360 42656 42424
rect 42720 42360 42736 42424
rect 42800 42360 42816 42424
rect 42880 42360 42896 42424
rect 42960 42360 42976 42424
rect 43040 42360 43056 42424
rect 43120 42360 43136 42424
rect 43200 42360 43216 42424
rect 43280 42360 43296 42424
rect 43360 42360 43376 42424
rect 43440 42360 43456 42424
rect 43520 42360 43536 42424
rect 43600 42360 43616 42424
rect 43680 42360 43696 42424
rect 43760 42360 43776 42424
rect 43840 42360 43856 42424
rect 43920 42360 43936 42424
rect 44000 42360 44016 42424
rect 44080 42360 44096 42424
rect 44160 42360 44176 42424
rect 44240 42360 44256 42424
rect 44320 42360 44336 42424
rect 44400 42360 44416 42424
rect 44480 42360 44496 42424
rect 44560 42360 44576 42424
rect 44640 42360 44656 42424
rect 44720 42360 44736 42424
rect 44800 42360 44816 42424
rect 44880 42360 44896 42424
rect 44960 42360 44976 42424
rect 45040 42360 45056 42424
rect 45120 42360 45136 42424
rect 45200 42360 45216 42424
rect 45280 42360 45296 42424
rect 45360 42360 45368 42424
rect 41368 42344 45368 42360
rect 41368 42280 41376 42344
rect 41440 42280 41456 42344
rect 41520 42280 41536 42344
rect 41600 42280 41616 42344
rect 41680 42280 41696 42344
rect 41760 42280 41776 42344
rect 41840 42280 41856 42344
rect 41920 42280 41936 42344
rect 42000 42280 42016 42344
rect 42080 42280 42096 42344
rect 42160 42280 42176 42344
rect 42240 42280 42256 42344
rect 42320 42280 42336 42344
rect 42400 42280 42416 42344
rect 42480 42280 42496 42344
rect 42560 42280 42576 42344
rect 42640 42280 42656 42344
rect 42720 42280 42736 42344
rect 42800 42280 42816 42344
rect 42880 42280 42896 42344
rect 42960 42280 42976 42344
rect 43040 42280 43056 42344
rect 43120 42280 43136 42344
rect 43200 42280 43216 42344
rect 43280 42280 43296 42344
rect 43360 42280 43376 42344
rect 43440 42280 43456 42344
rect 43520 42280 43536 42344
rect 43600 42280 43616 42344
rect 43680 42280 43696 42344
rect 43760 42280 43776 42344
rect 43840 42280 43856 42344
rect 43920 42280 43936 42344
rect 44000 42280 44016 42344
rect 44080 42280 44096 42344
rect 44160 42280 44176 42344
rect 44240 42280 44256 42344
rect 44320 42280 44336 42344
rect 44400 42280 44416 42344
rect 44480 42280 44496 42344
rect 44560 42280 44576 42344
rect 44640 42280 44656 42344
rect 44720 42280 44736 42344
rect 44800 42280 44816 42344
rect 44880 42280 44896 42344
rect 44960 42280 44976 42344
rect 45040 42280 45056 42344
rect 45120 42280 45136 42344
rect 45200 42280 45216 42344
rect 45280 42280 45296 42344
rect 45360 42280 45368 42344
rect 41368 42264 45368 42280
rect 41368 42200 41376 42264
rect 41440 42200 41456 42264
rect 41520 42200 41536 42264
rect 41600 42200 41616 42264
rect 41680 42200 41696 42264
rect 41760 42200 41776 42264
rect 41840 42200 41856 42264
rect 41920 42200 41936 42264
rect 42000 42200 42016 42264
rect 42080 42200 42096 42264
rect 42160 42200 42176 42264
rect 42240 42200 42256 42264
rect 42320 42200 42336 42264
rect 42400 42200 42416 42264
rect 42480 42200 42496 42264
rect 42560 42200 42576 42264
rect 42640 42200 42656 42264
rect 42720 42200 42736 42264
rect 42800 42200 42816 42264
rect 42880 42200 42896 42264
rect 42960 42200 42976 42264
rect 43040 42200 43056 42264
rect 43120 42200 43136 42264
rect 43200 42200 43216 42264
rect 43280 42200 43296 42264
rect 43360 42200 43376 42264
rect 43440 42200 43456 42264
rect 43520 42200 43536 42264
rect 43600 42200 43616 42264
rect 43680 42200 43696 42264
rect 43760 42200 43776 42264
rect 43840 42200 43856 42264
rect 43920 42200 43936 42264
rect 44000 42200 44016 42264
rect 44080 42200 44096 42264
rect 44160 42200 44176 42264
rect 44240 42200 44256 42264
rect 44320 42200 44336 42264
rect 44400 42200 44416 42264
rect 44480 42200 44496 42264
rect 44560 42200 44576 42264
rect 44640 42200 44656 42264
rect 44720 42200 44736 42264
rect 44800 42200 44816 42264
rect 44880 42200 44896 42264
rect 44960 42200 44976 42264
rect 45040 42200 45056 42264
rect 45120 42200 45136 42264
rect 45200 42200 45216 42264
rect 45280 42200 45296 42264
rect 45360 42200 45368 42264
rect 41368 42184 45368 42200
rect 41368 42120 41376 42184
rect 41440 42120 41456 42184
rect 41520 42120 41536 42184
rect 41600 42120 41616 42184
rect 41680 42120 41696 42184
rect 41760 42120 41776 42184
rect 41840 42120 41856 42184
rect 41920 42120 41936 42184
rect 42000 42120 42016 42184
rect 42080 42120 42096 42184
rect 42160 42120 42176 42184
rect 42240 42120 42256 42184
rect 42320 42120 42336 42184
rect 42400 42120 42416 42184
rect 42480 42120 42496 42184
rect 42560 42120 42576 42184
rect 42640 42120 42656 42184
rect 42720 42120 42736 42184
rect 42800 42120 42816 42184
rect 42880 42120 42896 42184
rect 42960 42120 42976 42184
rect 43040 42120 43056 42184
rect 43120 42120 43136 42184
rect 43200 42120 43216 42184
rect 43280 42120 43296 42184
rect 43360 42120 43376 42184
rect 43440 42120 43456 42184
rect 43520 42120 43536 42184
rect 43600 42120 43616 42184
rect 43680 42120 43696 42184
rect 43760 42120 43776 42184
rect 43840 42120 43856 42184
rect 43920 42120 43936 42184
rect 44000 42120 44016 42184
rect 44080 42120 44096 42184
rect 44160 42120 44176 42184
rect 44240 42120 44256 42184
rect 44320 42120 44336 42184
rect 44400 42120 44416 42184
rect 44480 42120 44496 42184
rect 44560 42120 44576 42184
rect 44640 42120 44656 42184
rect 44720 42120 44736 42184
rect 44800 42120 44816 42184
rect 44880 42120 44896 42184
rect 44960 42120 44976 42184
rect 45040 42120 45056 42184
rect 45120 42120 45136 42184
rect 45200 42120 45216 42184
rect 45280 42120 45296 42184
rect 45360 42120 45368 42184
rect 41368 42104 45368 42120
rect 41368 42040 41376 42104
rect 41440 42040 41456 42104
rect 41520 42040 41536 42104
rect 41600 42040 41616 42104
rect 41680 42040 41696 42104
rect 41760 42040 41776 42104
rect 41840 42040 41856 42104
rect 41920 42040 41936 42104
rect 42000 42040 42016 42104
rect 42080 42040 42096 42104
rect 42160 42040 42176 42104
rect 42240 42040 42256 42104
rect 42320 42040 42336 42104
rect 42400 42040 42416 42104
rect 42480 42040 42496 42104
rect 42560 42040 42576 42104
rect 42640 42040 42656 42104
rect 42720 42040 42736 42104
rect 42800 42040 42816 42104
rect 42880 42040 42896 42104
rect 42960 42040 42976 42104
rect 43040 42040 43056 42104
rect 43120 42040 43136 42104
rect 43200 42040 43216 42104
rect 43280 42040 43296 42104
rect 43360 42040 43376 42104
rect 43440 42040 43456 42104
rect 43520 42040 43536 42104
rect 43600 42040 43616 42104
rect 43680 42040 43696 42104
rect 43760 42040 43776 42104
rect 43840 42040 43856 42104
rect 43920 42040 43936 42104
rect 44000 42040 44016 42104
rect 44080 42040 44096 42104
rect 44160 42040 44176 42104
rect 44240 42040 44256 42104
rect 44320 42040 44336 42104
rect 44400 42040 44416 42104
rect 44480 42040 44496 42104
rect 44560 42040 44576 42104
rect 44640 42040 44656 42104
rect 44720 42040 44736 42104
rect 44800 42040 44816 42104
rect 44880 42040 44896 42104
rect 44960 42040 44976 42104
rect 45040 42040 45056 42104
rect 45120 42040 45136 42104
rect 45200 42040 45216 42104
rect 45280 42040 45296 42104
rect 45360 42040 45368 42104
rect 41368 42024 45368 42040
rect 41368 41960 41376 42024
rect 41440 41960 41456 42024
rect 41520 41960 41536 42024
rect 41600 41960 41616 42024
rect 41680 41960 41696 42024
rect 41760 41960 41776 42024
rect 41840 41960 41856 42024
rect 41920 41960 41936 42024
rect 42000 41960 42016 42024
rect 42080 41960 42096 42024
rect 42160 41960 42176 42024
rect 42240 41960 42256 42024
rect 42320 41960 42336 42024
rect 42400 41960 42416 42024
rect 42480 41960 42496 42024
rect 42560 41960 42576 42024
rect 42640 41960 42656 42024
rect 42720 41960 42736 42024
rect 42800 41960 42816 42024
rect 42880 41960 42896 42024
rect 42960 41960 42976 42024
rect 43040 41960 43056 42024
rect 43120 41960 43136 42024
rect 43200 41960 43216 42024
rect 43280 41960 43296 42024
rect 43360 41960 43376 42024
rect 43440 41960 43456 42024
rect 43520 41960 43536 42024
rect 43600 41960 43616 42024
rect 43680 41960 43696 42024
rect 43760 41960 43776 42024
rect 43840 41960 43856 42024
rect 43920 41960 43936 42024
rect 44000 41960 44016 42024
rect 44080 41960 44096 42024
rect 44160 41960 44176 42024
rect 44240 41960 44256 42024
rect 44320 41960 44336 42024
rect 44400 41960 44416 42024
rect 44480 41960 44496 42024
rect 44560 41960 44576 42024
rect 44640 41960 44656 42024
rect 44720 41960 44736 42024
rect 44800 41960 44816 42024
rect 44880 41960 44896 42024
rect 44960 41960 44976 42024
rect 45040 41960 45056 42024
rect 45120 41960 45136 42024
rect 45200 41960 45216 42024
rect 45280 41960 45296 42024
rect 45360 41960 45368 42024
rect 41368 41944 45368 41960
rect 41368 41880 41376 41944
rect 41440 41880 41456 41944
rect 41520 41880 41536 41944
rect 41600 41880 41616 41944
rect 41680 41880 41696 41944
rect 41760 41880 41776 41944
rect 41840 41880 41856 41944
rect 41920 41880 41936 41944
rect 42000 41880 42016 41944
rect 42080 41880 42096 41944
rect 42160 41880 42176 41944
rect 42240 41880 42256 41944
rect 42320 41880 42336 41944
rect 42400 41880 42416 41944
rect 42480 41880 42496 41944
rect 42560 41880 42576 41944
rect 42640 41880 42656 41944
rect 42720 41880 42736 41944
rect 42800 41880 42816 41944
rect 42880 41880 42896 41944
rect 42960 41880 42976 41944
rect 43040 41880 43056 41944
rect 43120 41880 43136 41944
rect 43200 41880 43216 41944
rect 43280 41880 43296 41944
rect 43360 41880 43376 41944
rect 43440 41880 43456 41944
rect 43520 41880 43536 41944
rect 43600 41880 43616 41944
rect 43680 41880 43696 41944
rect 43760 41880 43776 41944
rect 43840 41880 43856 41944
rect 43920 41880 43936 41944
rect 44000 41880 44016 41944
rect 44080 41880 44096 41944
rect 44160 41880 44176 41944
rect 44240 41880 44256 41944
rect 44320 41880 44336 41944
rect 44400 41880 44416 41944
rect 44480 41880 44496 41944
rect 44560 41880 44576 41944
rect 44640 41880 44656 41944
rect 44720 41880 44736 41944
rect 44800 41880 44816 41944
rect 44880 41880 44896 41944
rect 44960 41880 44976 41944
rect 45040 41880 45056 41944
rect 45120 41880 45136 41944
rect 45200 41880 45216 41944
rect 45280 41880 45296 41944
rect 45360 41880 45368 41944
rect 41368 41864 45368 41880
rect 41368 41800 41376 41864
rect 41440 41800 41456 41864
rect 41520 41800 41536 41864
rect 41600 41800 41616 41864
rect 41680 41800 41696 41864
rect 41760 41800 41776 41864
rect 41840 41800 41856 41864
rect 41920 41800 41936 41864
rect 42000 41800 42016 41864
rect 42080 41800 42096 41864
rect 42160 41800 42176 41864
rect 42240 41800 42256 41864
rect 42320 41800 42336 41864
rect 42400 41800 42416 41864
rect 42480 41800 42496 41864
rect 42560 41800 42576 41864
rect 42640 41800 42656 41864
rect 42720 41800 42736 41864
rect 42800 41800 42816 41864
rect 42880 41800 42896 41864
rect 42960 41800 42976 41864
rect 43040 41800 43056 41864
rect 43120 41800 43136 41864
rect 43200 41800 43216 41864
rect 43280 41800 43296 41864
rect 43360 41800 43376 41864
rect 43440 41800 43456 41864
rect 43520 41800 43536 41864
rect 43600 41800 43616 41864
rect 43680 41800 43696 41864
rect 43760 41800 43776 41864
rect 43840 41800 43856 41864
rect 43920 41800 43936 41864
rect 44000 41800 44016 41864
rect 44080 41800 44096 41864
rect 44160 41800 44176 41864
rect 44240 41800 44256 41864
rect 44320 41800 44336 41864
rect 44400 41800 44416 41864
rect 44480 41800 44496 41864
rect 44560 41800 44576 41864
rect 44640 41800 44656 41864
rect 44720 41800 44736 41864
rect 44800 41800 44816 41864
rect 44880 41800 44896 41864
rect 44960 41800 44976 41864
rect 45040 41800 45056 41864
rect 45120 41800 45136 41864
rect 45200 41800 45216 41864
rect 45280 41800 45296 41864
rect 45360 41800 45368 41864
rect 41368 41784 45368 41800
rect 41368 41720 41376 41784
rect 41440 41720 41456 41784
rect 41520 41720 41536 41784
rect 41600 41720 41616 41784
rect 41680 41720 41696 41784
rect 41760 41720 41776 41784
rect 41840 41720 41856 41784
rect 41920 41720 41936 41784
rect 42000 41720 42016 41784
rect 42080 41720 42096 41784
rect 42160 41720 42176 41784
rect 42240 41720 42256 41784
rect 42320 41720 42336 41784
rect 42400 41720 42416 41784
rect 42480 41720 42496 41784
rect 42560 41720 42576 41784
rect 42640 41720 42656 41784
rect 42720 41720 42736 41784
rect 42800 41720 42816 41784
rect 42880 41720 42896 41784
rect 42960 41720 42976 41784
rect 43040 41720 43056 41784
rect 43120 41720 43136 41784
rect 43200 41720 43216 41784
rect 43280 41720 43296 41784
rect 43360 41720 43376 41784
rect 43440 41720 43456 41784
rect 43520 41720 43536 41784
rect 43600 41720 43616 41784
rect 43680 41720 43696 41784
rect 43760 41720 43776 41784
rect 43840 41720 43856 41784
rect 43920 41720 43936 41784
rect 44000 41720 44016 41784
rect 44080 41720 44096 41784
rect 44160 41720 44176 41784
rect 44240 41720 44256 41784
rect 44320 41720 44336 41784
rect 44400 41720 44416 41784
rect 44480 41720 44496 41784
rect 44560 41720 44576 41784
rect 44640 41720 44656 41784
rect 44720 41720 44736 41784
rect 44800 41720 44816 41784
rect 44880 41720 44896 41784
rect 44960 41720 44976 41784
rect 45040 41720 45056 41784
rect 45120 41720 45136 41784
rect 45200 41720 45216 41784
rect 45280 41720 45296 41784
rect 45360 41720 45368 41784
rect 41368 41704 45368 41720
rect 41368 41640 41376 41704
rect 41440 41640 41456 41704
rect 41520 41640 41536 41704
rect 41600 41640 41616 41704
rect 41680 41640 41696 41704
rect 41760 41640 41776 41704
rect 41840 41640 41856 41704
rect 41920 41640 41936 41704
rect 42000 41640 42016 41704
rect 42080 41640 42096 41704
rect 42160 41640 42176 41704
rect 42240 41640 42256 41704
rect 42320 41640 42336 41704
rect 42400 41640 42416 41704
rect 42480 41640 42496 41704
rect 42560 41640 42576 41704
rect 42640 41640 42656 41704
rect 42720 41640 42736 41704
rect 42800 41640 42816 41704
rect 42880 41640 42896 41704
rect 42960 41640 42976 41704
rect 43040 41640 43056 41704
rect 43120 41640 43136 41704
rect 43200 41640 43216 41704
rect 43280 41640 43296 41704
rect 43360 41640 43376 41704
rect 43440 41640 43456 41704
rect 43520 41640 43536 41704
rect 43600 41640 43616 41704
rect 43680 41640 43696 41704
rect 43760 41640 43776 41704
rect 43840 41640 43856 41704
rect 43920 41640 43936 41704
rect 44000 41640 44016 41704
rect 44080 41640 44096 41704
rect 44160 41640 44176 41704
rect 44240 41640 44256 41704
rect 44320 41640 44336 41704
rect 44400 41640 44416 41704
rect 44480 41640 44496 41704
rect 44560 41640 44576 41704
rect 44640 41640 44656 41704
rect 44720 41640 44736 41704
rect 44800 41640 44816 41704
rect 44880 41640 44896 41704
rect 44960 41640 44976 41704
rect 45040 41640 45056 41704
rect 45120 41640 45136 41704
rect 45200 41640 45216 41704
rect 45280 41640 45296 41704
rect 45360 41640 45368 41704
rect 41368 41624 45368 41640
rect 41368 41560 41376 41624
rect 41440 41560 41456 41624
rect 41520 41560 41536 41624
rect 41600 41560 41616 41624
rect 41680 41560 41696 41624
rect 41760 41560 41776 41624
rect 41840 41560 41856 41624
rect 41920 41560 41936 41624
rect 42000 41560 42016 41624
rect 42080 41560 42096 41624
rect 42160 41560 42176 41624
rect 42240 41560 42256 41624
rect 42320 41560 42336 41624
rect 42400 41560 42416 41624
rect 42480 41560 42496 41624
rect 42560 41560 42576 41624
rect 42640 41560 42656 41624
rect 42720 41560 42736 41624
rect 42800 41560 42816 41624
rect 42880 41560 42896 41624
rect 42960 41560 42976 41624
rect 43040 41560 43056 41624
rect 43120 41560 43136 41624
rect 43200 41560 43216 41624
rect 43280 41560 43296 41624
rect 43360 41560 43376 41624
rect 43440 41560 43456 41624
rect 43520 41560 43536 41624
rect 43600 41560 43616 41624
rect 43680 41560 43696 41624
rect 43760 41560 43776 41624
rect 43840 41560 43856 41624
rect 43920 41560 43936 41624
rect 44000 41560 44016 41624
rect 44080 41560 44096 41624
rect 44160 41560 44176 41624
rect 44240 41560 44256 41624
rect 44320 41560 44336 41624
rect 44400 41560 44416 41624
rect 44480 41560 44496 41624
rect 44560 41560 44576 41624
rect 44640 41560 44656 41624
rect 44720 41560 44736 41624
rect 44800 41560 44816 41624
rect 44880 41560 44896 41624
rect 44960 41560 44976 41624
rect 45040 41560 45056 41624
rect 45120 41560 45136 41624
rect 45200 41560 45216 41624
rect 45280 41560 45296 41624
rect 45360 41560 45368 41624
rect 41368 41544 45368 41560
rect 41368 41480 41376 41544
rect 41440 41480 41456 41544
rect 41520 41480 41536 41544
rect 41600 41480 41616 41544
rect 41680 41480 41696 41544
rect 41760 41480 41776 41544
rect 41840 41480 41856 41544
rect 41920 41480 41936 41544
rect 42000 41480 42016 41544
rect 42080 41480 42096 41544
rect 42160 41480 42176 41544
rect 42240 41480 42256 41544
rect 42320 41480 42336 41544
rect 42400 41480 42416 41544
rect 42480 41480 42496 41544
rect 42560 41480 42576 41544
rect 42640 41480 42656 41544
rect 42720 41480 42736 41544
rect 42800 41480 42816 41544
rect 42880 41480 42896 41544
rect 42960 41480 42976 41544
rect 43040 41480 43056 41544
rect 43120 41480 43136 41544
rect 43200 41480 43216 41544
rect 43280 41480 43296 41544
rect 43360 41480 43376 41544
rect 43440 41480 43456 41544
rect 43520 41480 43536 41544
rect 43600 41480 43616 41544
rect 43680 41480 43696 41544
rect 43760 41480 43776 41544
rect 43840 41480 43856 41544
rect 43920 41480 43936 41544
rect 44000 41480 44016 41544
rect 44080 41480 44096 41544
rect 44160 41480 44176 41544
rect 44240 41480 44256 41544
rect 44320 41480 44336 41544
rect 44400 41480 44416 41544
rect 44480 41480 44496 41544
rect 44560 41480 44576 41544
rect 44640 41480 44656 41544
rect 44720 41480 44736 41544
rect 44800 41480 44816 41544
rect 44880 41480 44896 41544
rect 44960 41480 44976 41544
rect 45040 41480 45056 41544
rect 45120 41480 45136 41544
rect 45200 41480 45216 41544
rect 45280 41480 45296 41544
rect 45360 41480 45368 41544
rect 41368 41464 45368 41480
rect 41368 41400 41376 41464
rect 41440 41400 41456 41464
rect 41520 41400 41536 41464
rect 41600 41400 41616 41464
rect 41680 41400 41696 41464
rect 41760 41400 41776 41464
rect 41840 41400 41856 41464
rect 41920 41400 41936 41464
rect 42000 41400 42016 41464
rect 42080 41400 42096 41464
rect 42160 41400 42176 41464
rect 42240 41400 42256 41464
rect 42320 41400 42336 41464
rect 42400 41400 42416 41464
rect 42480 41400 42496 41464
rect 42560 41400 42576 41464
rect 42640 41400 42656 41464
rect 42720 41400 42736 41464
rect 42800 41400 42816 41464
rect 42880 41400 42896 41464
rect 42960 41400 42976 41464
rect 43040 41400 43056 41464
rect 43120 41400 43136 41464
rect 43200 41400 43216 41464
rect 43280 41400 43296 41464
rect 43360 41400 43376 41464
rect 43440 41400 43456 41464
rect 43520 41400 43536 41464
rect 43600 41400 43616 41464
rect 43680 41400 43696 41464
rect 43760 41400 43776 41464
rect 43840 41400 43856 41464
rect 43920 41400 43936 41464
rect 44000 41400 44016 41464
rect 44080 41400 44096 41464
rect 44160 41400 44176 41464
rect 44240 41400 44256 41464
rect 44320 41400 44336 41464
rect 44400 41400 44416 41464
rect 44480 41400 44496 41464
rect 44560 41400 44576 41464
rect 44640 41400 44656 41464
rect 44720 41400 44736 41464
rect 44800 41400 44816 41464
rect 44880 41400 44896 41464
rect 44960 41400 44976 41464
rect 45040 41400 45056 41464
rect 45120 41400 45136 41464
rect 45200 41400 45216 41464
rect 45280 41400 45296 41464
rect 45360 41400 45368 41464
rect 29104 34360 29112 34424
rect 29176 34360 29192 34424
rect 29256 34360 29272 34424
rect 29336 34360 29352 34424
rect 29416 34360 29424 34424
rect 29104 33336 29424 34360
rect 29104 33272 29112 33336
rect 29176 33272 29192 33336
rect 29256 33272 29272 33336
rect 29336 33272 29352 33336
rect 29416 33272 29424 33336
rect 29104 32248 29424 33272
rect 29104 32184 29112 32248
rect 29176 32184 29192 32248
rect 29256 32184 29272 32248
rect 29336 32184 29352 32248
rect 29416 32184 29424 32248
rect 29104 31160 29424 32184
rect 29104 31096 29112 31160
rect 29176 31096 29192 31160
rect 29256 31096 29272 31160
rect 29336 31096 29352 31160
rect 29416 31096 29424 31160
rect 29104 30072 29424 31096
rect 29104 30008 29112 30072
rect 29176 30008 29192 30072
rect 29256 30008 29272 30072
rect 29336 30008 29352 30072
rect 29416 30008 29424 30072
rect 29104 28984 29424 30008
rect 29104 28920 29112 28984
rect 29176 28920 29192 28984
rect 29256 28920 29272 28984
rect 29336 28920 29352 28984
rect 29416 28920 29424 28984
rect 29104 27896 29424 28920
rect 29104 27832 29112 27896
rect 29176 27832 29192 27896
rect 29256 27832 29272 27896
rect 29336 27832 29352 27896
rect 29416 27832 29424 27896
rect 29104 26808 29424 27832
rect 29104 26744 29112 26808
rect 29176 26744 29192 26808
rect 29256 26744 29272 26808
rect 29336 26744 29352 26808
rect 29416 26744 29424 26808
rect 29104 25720 29424 26744
rect 29104 25656 29112 25720
rect 29176 25656 29192 25720
rect 29256 25656 29272 25720
rect 29336 25656 29352 25720
rect 29416 25656 29424 25720
rect 29104 24632 29424 25656
rect 29104 24568 29112 24632
rect 29176 24568 29192 24632
rect 29256 24568 29272 24632
rect 29336 24568 29352 24632
rect 29416 24568 29424 24632
rect 29104 23544 29424 24568
rect 29104 23480 29112 23544
rect 29176 23480 29192 23544
rect 29256 23480 29272 23544
rect 29336 23480 29352 23544
rect 29416 23480 29424 23544
rect 29104 22456 29424 23480
rect 29104 22392 29112 22456
rect 29176 22392 29192 22456
rect 29256 22392 29272 22456
rect 29336 22392 29352 22456
rect 29416 22392 29424 22456
rect 29104 21368 29424 22392
rect 29104 21304 29112 21368
rect 29176 21304 29192 21368
rect 29256 21304 29272 21368
rect 29336 21304 29352 21368
rect 29416 21304 29424 21368
rect 29104 20280 29424 21304
rect 29104 20216 29112 20280
rect 29176 20216 29192 20280
rect 29256 20216 29272 20280
rect 29336 20216 29352 20280
rect 29416 20216 29424 20280
rect 29104 19192 29424 20216
rect 29104 19128 29112 19192
rect 29176 19128 29192 19192
rect 29256 19128 29272 19192
rect 29336 19128 29352 19192
rect 29416 19128 29424 19192
rect 29104 18104 29424 19128
rect 29104 18040 29112 18104
rect 29176 18040 29192 18104
rect 29256 18040 29272 18104
rect 29336 18040 29352 18104
rect 29416 18040 29424 18104
rect 29104 17016 29424 18040
rect 29104 16952 29112 17016
rect 29176 16952 29192 17016
rect 29256 16952 29272 17016
rect 29336 16952 29352 17016
rect 29416 16952 29424 17016
rect 29104 15928 29424 16952
rect 29104 15864 29112 15928
rect 29176 15864 29192 15928
rect 29256 15864 29272 15928
rect 29336 15864 29352 15928
rect 29416 15864 29424 15928
rect 29104 14840 29424 15864
rect 29104 14776 29112 14840
rect 29176 14776 29192 14840
rect 29256 14776 29272 14840
rect 29336 14776 29352 14840
rect 29416 14776 29424 14840
rect 29104 13752 29424 14776
rect 29104 13688 29112 13752
rect 29176 13688 29192 13752
rect 29256 13688 29272 13752
rect 29336 13688 29352 13752
rect 29416 13688 29424 13752
rect 29104 12664 29424 13688
rect 29104 12600 29112 12664
rect 29176 12600 29192 12664
rect 29256 12600 29272 12664
rect 29336 12600 29352 12664
rect 29416 12600 29424 12664
rect 29104 11576 29424 12600
rect 29104 11512 29112 11576
rect 29176 11512 29192 11576
rect 29256 11512 29272 11576
rect 29336 11512 29352 11576
rect 29416 11512 29424 11576
rect 29104 3992 29424 11512
rect 36368 40384 40368 40392
rect 36368 40320 36376 40384
rect 36440 40320 36456 40384
rect 36520 40320 36536 40384
rect 36600 40320 36616 40384
rect 36680 40320 36696 40384
rect 36760 40320 36776 40384
rect 36840 40320 36856 40384
rect 36920 40320 36936 40384
rect 37000 40320 37016 40384
rect 37080 40320 37096 40384
rect 37160 40320 37176 40384
rect 37240 40320 37256 40384
rect 37320 40320 37336 40384
rect 37400 40320 37416 40384
rect 37480 40320 37496 40384
rect 37560 40320 37576 40384
rect 37640 40320 37656 40384
rect 37720 40320 37736 40384
rect 37800 40320 37816 40384
rect 37880 40320 37896 40384
rect 37960 40320 37976 40384
rect 38040 40320 38056 40384
rect 38120 40320 38136 40384
rect 38200 40320 38216 40384
rect 38280 40320 38296 40384
rect 38360 40320 38376 40384
rect 38440 40320 38456 40384
rect 38520 40320 38536 40384
rect 38600 40320 38616 40384
rect 38680 40320 38696 40384
rect 38760 40320 38776 40384
rect 38840 40320 38856 40384
rect 38920 40320 38936 40384
rect 39000 40320 39016 40384
rect 39080 40320 39096 40384
rect 39160 40320 39176 40384
rect 39240 40320 39256 40384
rect 39320 40320 39336 40384
rect 39400 40320 39416 40384
rect 39480 40320 39496 40384
rect 39560 40320 39576 40384
rect 39640 40320 39656 40384
rect 39720 40320 39736 40384
rect 39800 40320 39816 40384
rect 39880 40320 39896 40384
rect 39960 40320 39976 40384
rect 40040 40320 40056 40384
rect 40120 40320 40136 40384
rect 40200 40320 40216 40384
rect 40280 40320 40296 40384
rect 40360 40320 40368 40384
rect 36368 40304 40368 40320
rect 36368 40240 36376 40304
rect 36440 40240 36456 40304
rect 36520 40240 36536 40304
rect 36600 40240 36616 40304
rect 36680 40240 36696 40304
rect 36760 40240 36776 40304
rect 36840 40240 36856 40304
rect 36920 40240 36936 40304
rect 37000 40240 37016 40304
rect 37080 40240 37096 40304
rect 37160 40240 37176 40304
rect 37240 40240 37256 40304
rect 37320 40240 37336 40304
rect 37400 40240 37416 40304
rect 37480 40240 37496 40304
rect 37560 40240 37576 40304
rect 37640 40240 37656 40304
rect 37720 40240 37736 40304
rect 37800 40240 37816 40304
rect 37880 40240 37896 40304
rect 37960 40240 37976 40304
rect 38040 40240 38056 40304
rect 38120 40240 38136 40304
rect 38200 40240 38216 40304
rect 38280 40240 38296 40304
rect 38360 40240 38376 40304
rect 38440 40240 38456 40304
rect 38520 40240 38536 40304
rect 38600 40240 38616 40304
rect 38680 40240 38696 40304
rect 38760 40240 38776 40304
rect 38840 40240 38856 40304
rect 38920 40240 38936 40304
rect 39000 40240 39016 40304
rect 39080 40240 39096 40304
rect 39160 40240 39176 40304
rect 39240 40240 39256 40304
rect 39320 40240 39336 40304
rect 39400 40240 39416 40304
rect 39480 40240 39496 40304
rect 39560 40240 39576 40304
rect 39640 40240 39656 40304
rect 39720 40240 39736 40304
rect 39800 40240 39816 40304
rect 39880 40240 39896 40304
rect 39960 40240 39976 40304
rect 40040 40240 40056 40304
rect 40120 40240 40136 40304
rect 40200 40240 40216 40304
rect 40280 40240 40296 40304
rect 40360 40240 40368 40304
rect 36368 40224 40368 40240
rect 36368 40160 36376 40224
rect 36440 40160 36456 40224
rect 36520 40160 36536 40224
rect 36600 40160 36616 40224
rect 36680 40160 36696 40224
rect 36760 40160 36776 40224
rect 36840 40160 36856 40224
rect 36920 40160 36936 40224
rect 37000 40160 37016 40224
rect 37080 40160 37096 40224
rect 37160 40160 37176 40224
rect 37240 40160 37256 40224
rect 37320 40160 37336 40224
rect 37400 40160 37416 40224
rect 37480 40160 37496 40224
rect 37560 40160 37576 40224
rect 37640 40160 37656 40224
rect 37720 40160 37736 40224
rect 37800 40160 37816 40224
rect 37880 40160 37896 40224
rect 37960 40160 37976 40224
rect 38040 40160 38056 40224
rect 38120 40160 38136 40224
rect 38200 40160 38216 40224
rect 38280 40160 38296 40224
rect 38360 40160 38376 40224
rect 38440 40160 38456 40224
rect 38520 40160 38536 40224
rect 38600 40160 38616 40224
rect 38680 40160 38696 40224
rect 38760 40160 38776 40224
rect 38840 40160 38856 40224
rect 38920 40160 38936 40224
rect 39000 40160 39016 40224
rect 39080 40160 39096 40224
rect 39160 40160 39176 40224
rect 39240 40160 39256 40224
rect 39320 40160 39336 40224
rect 39400 40160 39416 40224
rect 39480 40160 39496 40224
rect 39560 40160 39576 40224
rect 39640 40160 39656 40224
rect 39720 40160 39736 40224
rect 39800 40160 39816 40224
rect 39880 40160 39896 40224
rect 39960 40160 39976 40224
rect 40040 40160 40056 40224
rect 40120 40160 40136 40224
rect 40200 40160 40216 40224
rect 40280 40160 40296 40224
rect 40360 40160 40368 40224
rect 36368 40144 40368 40160
rect 36368 40080 36376 40144
rect 36440 40080 36456 40144
rect 36520 40080 36536 40144
rect 36600 40080 36616 40144
rect 36680 40080 36696 40144
rect 36760 40080 36776 40144
rect 36840 40080 36856 40144
rect 36920 40080 36936 40144
rect 37000 40080 37016 40144
rect 37080 40080 37096 40144
rect 37160 40080 37176 40144
rect 37240 40080 37256 40144
rect 37320 40080 37336 40144
rect 37400 40080 37416 40144
rect 37480 40080 37496 40144
rect 37560 40080 37576 40144
rect 37640 40080 37656 40144
rect 37720 40080 37736 40144
rect 37800 40080 37816 40144
rect 37880 40080 37896 40144
rect 37960 40080 37976 40144
rect 38040 40080 38056 40144
rect 38120 40080 38136 40144
rect 38200 40080 38216 40144
rect 38280 40080 38296 40144
rect 38360 40080 38376 40144
rect 38440 40080 38456 40144
rect 38520 40080 38536 40144
rect 38600 40080 38616 40144
rect 38680 40080 38696 40144
rect 38760 40080 38776 40144
rect 38840 40080 38856 40144
rect 38920 40080 38936 40144
rect 39000 40080 39016 40144
rect 39080 40080 39096 40144
rect 39160 40080 39176 40144
rect 39240 40080 39256 40144
rect 39320 40080 39336 40144
rect 39400 40080 39416 40144
rect 39480 40080 39496 40144
rect 39560 40080 39576 40144
rect 39640 40080 39656 40144
rect 39720 40080 39736 40144
rect 39800 40080 39816 40144
rect 39880 40080 39896 40144
rect 39960 40080 39976 40144
rect 40040 40080 40056 40144
rect 40120 40080 40136 40144
rect 40200 40080 40216 40144
rect 40280 40080 40296 40144
rect 40360 40080 40368 40144
rect 36368 40064 40368 40080
rect 36368 40000 36376 40064
rect 36440 40000 36456 40064
rect 36520 40000 36536 40064
rect 36600 40000 36616 40064
rect 36680 40000 36696 40064
rect 36760 40000 36776 40064
rect 36840 40000 36856 40064
rect 36920 40000 36936 40064
rect 37000 40000 37016 40064
rect 37080 40000 37096 40064
rect 37160 40000 37176 40064
rect 37240 40000 37256 40064
rect 37320 40000 37336 40064
rect 37400 40000 37416 40064
rect 37480 40000 37496 40064
rect 37560 40000 37576 40064
rect 37640 40000 37656 40064
rect 37720 40000 37736 40064
rect 37800 40000 37816 40064
rect 37880 40000 37896 40064
rect 37960 40000 37976 40064
rect 38040 40000 38056 40064
rect 38120 40000 38136 40064
rect 38200 40000 38216 40064
rect 38280 40000 38296 40064
rect 38360 40000 38376 40064
rect 38440 40000 38456 40064
rect 38520 40000 38536 40064
rect 38600 40000 38616 40064
rect 38680 40000 38696 40064
rect 38760 40000 38776 40064
rect 38840 40000 38856 40064
rect 38920 40000 38936 40064
rect 39000 40000 39016 40064
rect 39080 40000 39096 40064
rect 39160 40000 39176 40064
rect 39240 40000 39256 40064
rect 39320 40000 39336 40064
rect 39400 40000 39416 40064
rect 39480 40000 39496 40064
rect 39560 40000 39576 40064
rect 39640 40000 39656 40064
rect 39720 40000 39736 40064
rect 39800 40000 39816 40064
rect 39880 40000 39896 40064
rect 39960 40000 39976 40064
rect 40040 40000 40056 40064
rect 40120 40000 40136 40064
rect 40200 40000 40216 40064
rect 40280 40000 40296 40064
rect 40360 40000 40368 40064
rect 36368 39984 40368 40000
rect 36368 39920 36376 39984
rect 36440 39920 36456 39984
rect 36520 39920 36536 39984
rect 36600 39920 36616 39984
rect 36680 39920 36696 39984
rect 36760 39920 36776 39984
rect 36840 39920 36856 39984
rect 36920 39920 36936 39984
rect 37000 39920 37016 39984
rect 37080 39920 37096 39984
rect 37160 39920 37176 39984
rect 37240 39920 37256 39984
rect 37320 39920 37336 39984
rect 37400 39920 37416 39984
rect 37480 39920 37496 39984
rect 37560 39920 37576 39984
rect 37640 39920 37656 39984
rect 37720 39920 37736 39984
rect 37800 39920 37816 39984
rect 37880 39920 37896 39984
rect 37960 39920 37976 39984
rect 38040 39920 38056 39984
rect 38120 39920 38136 39984
rect 38200 39920 38216 39984
rect 38280 39920 38296 39984
rect 38360 39920 38376 39984
rect 38440 39920 38456 39984
rect 38520 39920 38536 39984
rect 38600 39920 38616 39984
rect 38680 39920 38696 39984
rect 38760 39920 38776 39984
rect 38840 39920 38856 39984
rect 38920 39920 38936 39984
rect 39000 39920 39016 39984
rect 39080 39920 39096 39984
rect 39160 39920 39176 39984
rect 39240 39920 39256 39984
rect 39320 39920 39336 39984
rect 39400 39920 39416 39984
rect 39480 39920 39496 39984
rect 39560 39920 39576 39984
rect 39640 39920 39656 39984
rect 39720 39920 39736 39984
rect 39800 39920 39816 39984
rect 39880 39920 39896 39984
rect 39960 39920 39976 39984
rect 40040 39920 40056 39984
rect 40120 39920 40136 39984
rect 40200 39920 40216 39984
rect 40280 39920 40296 39984
rect 40360 39920 40368 39984
rect 36368 39904 40368 39920
rect 36368 39840 36376 39904
rect 36440 39840 36456 39904
rect 36520 39840 36536 39904
rect 36600 39840 36616 39904
rect 36680 39840 36696 39904
rect 36760 39840 36776 39904
rect 36840 39840 36856 39904
rect 36920 39840 36936 39904
rect 37000 39840 37016 39904
rect 37080 39840 37096 39904
rect 37160 39840 37176 39904
rect 37240 39840 37256 39904
rect 37320 39840 37336 39904
rect 37400 39840 37416 39904
rect 37480 39840 37496 39904
rect 37560 39840 37576 39904
rect 37640 39840 37656 39904
rect 37720 39840 37736 39904
rect 37800 39840 37816 39904
rect 37880 39840 37896 39904
rect 37960 39840 37976 39904
rect 38040 39840 38056 39904
rect 38120 39840 38136 39904
rect 38200 39840 38216 39904
rect 38280 39840 38296 39904
rect 38360 39840 38376 39904
rect 38440 39840 38456 39904
rect 38520 39840 38536 39904
rect 38600 39840 38616 39904
rect 38680 39840 38696 39904
rect 38760 39840 38776 39904
rect 38840 39840 38856 39904
rect 38920 39840 38936 39904
rect 39000 39840 39016 39904
rect 39080 39840 39096 39904
rect 39160 39840 39176 39904
rect 39240 39840 39256 39904
rect 39320 39840 39336 39904
rect 39400 39840 39416 39904
rect 39480 39840 39496 39904
rect 39560 39840 39576 39904
rect 39640 39840 39656 39904
rect 39720 39840 39736 39904
rect 39800 39840 39816 39904
rect 39880 39840 39896 39904
rect 39960 39840 39976 39904
rect 40040 39840 40056 39904
rect 40120 39840 40136 39904
rect 40200 39840 40216 39904
rect 40280 39840 40296 39904
rect 40360 39840 40368 39904
rect 36368 39824 40368 39840
rect 36368 39760 36376 39824
rect 36440 39760 36456 39824
rect 36520 39760 36536 39824
rect 36600 39760 36616 39824
rect 36680 39760 36696 39824
rect 36760 39760 36776 39824
rect 36840 39760 36856 39824
rect 36920 39760 36936 39824
rect 37000 39760 37016 39824
rect 37080 39760 37096 39824
rect 37160 39760 37176 39824
rect 37240 39760 37256 39824
rect 37320 39760 37336 39824
rect 37400 39760 37416 39824
rect 37480 39760 37496 39824
rect 37560 39760 37576 39824
rect 37640 39760 37656 39824
rect 37720 39760 37736 39824
rect 37800 39760 37816 39824
rect 37880 39760 37896 39824
rect 37960 39760 37976 39824
rect 38040 39760 38056 39824
rect 38120 39760 38136 39824
rect 38200 39760 38216 39824
rect 38280 39760 38296 39824
rect 38360 39760 38376 39824
rect 38440 39760 38456 39824
rect 38520 39760 38536 39824
rect 38600 39760 38616 39824
rect 38680 39760 38696 39824
rect 38760 39760 38776 39824
rect 38840 39760 38856 39824
rect 38920 39760 38936 39824
rect 39000 39760 39016 39824
rect 39080 39760 39096 39824
rect 39160 39760 39176 39824
rect 39240 39760 39256 39824
rect 39320 39760 39336 39824
rect 39400 39760 39416 39824
rect 39480 39760 39496 39824
rect 39560 39760 39576 39824
rect 39640 39760 39656 39824
rect 39720 39760 39736 39824
rect 39800 39760 39816 39824
rect 39880 39760 39896 39824
rect 39960 39760 39976 39824
rect 40040 39760 40056 39824
rect 40120 39760 40136 39824
rect 40200 39760 40216 39824
rect 40280 39760 40296 39824
rect 40360 39760 40368 39824
rect 36368 39744 40368 39760
rect 36368 39680 36376 39744
rect 36440 39680 36456 39744
rect 36520 39680 36536 39744
rect 36600 39680 36616 39744
rect 36680 39680 36696 39744
rect 36760 39680 36776 39744
rect 36840 39680 36856 39744
rect 36920 39680 36936 39744
rect 37000 39680 37016 39744
rect 37080 39680 37096 39744
rect 37160 39680 37176 39744
rect 37240 39680 37256 39744
rect 37320 39680 37336 39744
rect 37400 39680 37416 39744
rect 37480 39680 37496 39744
rect 37560 39680 37576 39744
rect 37640 39680 37656 39744
rect 37720 39680 37736 39744
rect 37800 39680 37816 39744
rect 37880 39680 37896 39744
rect 37960 39680 37976 39744
rect 38040 39680 38056 39744
rect 38120 39680 38136 39744
rect 38200 39680 38216 39744
rect 38280 39680 38296 39744
rect 38360 39680 38376 39744
rect 38440 39680 38456 39744
rect 38520 39680 38536 39744
rect 38600 39680 38616 39744
rect 38680 39680 38696 39744
rect 38760 39680 38776 39744
rect 38840 39680 38856 39744
rect 38920 39680 38936 39744
rect 39000 39680 39016 39744
rect 39080 39680 39096 39744
rect 39160 39680 39176 39744
rect 39240 39680 39256 39744
rect 39320 39680 39336 39744
rect 39400 39680 39416 39744
rect 39480 39680 39496 39744
rect 39560 39680 39576 39744
rect 39640 39680 39656 39744
rect 39720 39680 39736 39744
rect 39800 39680 39816 39744
rect 39880 39680 39896 39744
rect 39960 39680 39976 39744
rect 40040 39680 40056 39744
rect 40120 39680 40136 39744
rect 40200 39680 40216 39744
rect 40280 39680 40296 39744
rect 40360 39680 40368 39744
rect 36368 39664 40368 39680
rect 36368 39600 36376 39664
rect 36440 39600 36456 39664
rect 36520 39600 36536 39664
rect 36600 39600 36616 39664
rect 36680 39600 36696 39664
rect 36760 39600 36776 39664
rect 36840 39600 36856 39664
rect 36920 39600 36936 39664
rect 37000 39600 37016 39664
rect 37080 39600 37096 39664
rect 37160 39600 37176 39664
rect 37240 39600 37256 39664
rect 37320 39600 37336 39664
rect 37400 39600 37416 39664
rect 37480 39600 37496 39664
rect 37560 39600 37576 39664
rect 37640 39600 37656 39664
rect 37720 39600 37736 39664
rect 37800 39600 37816 39664
rect 37880 39600 37896 39664
rect 37960 39600 37976 39664
rect 38040 39600 38056 39664
rect 38120 39600 38136 39664
rect 38200 39600 38216 39664
rect 38280 39600 38296 39664
rect 38360 39600 38376 39664
rect 38440 39600 38456 39664
rect 38520 39600 38536 39664
rect 38600 39600 38616 39664
rect 38680 39600 38696 39664
rect 38760 39600 38776 39664
rect 38840 39600 38856 39664
rect 38920 39600 38936 39664
rect 39000 39600 39016 39664
rect 39080 39600 39096 39664
rect 39160 39600 39176 39664
rect 39240 39600 39256 39664
rect 39320 39600 39336 39664
rect 39400 39600 39416 39664
rect 39480 39600 39496 39664
rect 39560 39600 39576 39664
rect 39640 39600 39656 39664
rect 39720 39600 39736 39664
rect 39800 39600 39816 39664
rect 39880 39600 39896 39664
rect 39960 39600 39976 39664
rect 40040 39600 40056 39664
rect 40120 39600 40136 39664
rect 40200 39600 40216 39664
rect 40280 39600 40296 39664
rect 40360 39600 40368 39664
rect 36368 39584 40368 39600
rect 36368 39520 36376 39584
rect 36440 39520 36456 39584
rect 36520 39520 36536 39584
rect 36600 39520 36616 39584
rect 36680 39520 36696 39584
rect 36760 39520 36776 39584
rect 36840 39520 36856 39584
rect 36920 39520 36936 39584
rect 37000 39520 37016 39584
rect 37080 39520 37096 39584
rect 37160 39520 37176 39584
rect 37240 39520 37256 39584
rect 37320 39520 37336 39584
rect 37400 39520 37416 39584
rect 37480 39520 37496 39584
rect 37560 39520 37576 39584
rect 37640 39520 37656 39584
rect 37720 39520 37736 39584
rect 37800 39520 37816 39584
rect 37880 39520 37896 39584
rect 37960 39520 37976 39584
rect 38040 39520 38056 39584
rect 38120 39520 38136 39584
rect 38200 39520 38216 39584
rect 38280 39520 38296 39584
rect 38360 39520 38376 39584
rect 38440 39520 38456 39584
rect 38520 39520 38536 39584
rect 38600 39520 38616 39584
rect 38680 39520 38696 39584
rect 38760 39520 38776 39584
rect 38840 39520 38856 39584
rect 38920 39520 38936 39584
rect 39000 39520 39016 39584
rect 39080 39520 39096 39584
rect 39160 39520 39176 39584
rect 39240 39520 39256 39584
rect 39320 39520 39336 39584
rect 39400 39520 39416 39584
rect 39480 39520 39496 39584
rect 39560 39520 39576 39584
rect 39640 39520 39656 39584
rect 39720 39520 39736 39584
rect 39800 39520 39816 39584
rect 39880 39520 39896 39584
rect 39960 39520 39976 39584
rect 40040 39520 40056 39584
rect 40120 39520 40136 39584
rect 40200 39520 40216 39584
rect 40280 39520 40296 39584
rect 40360 39520 40368 39584
rect 36368 39504 40368 39520
rect 36368 39440 36376 39504
rect 36440 39440 36456 39504
rect 36520 39440 36536 39504
rect 36600 39440 36616 39504
rect 36680 39440 36696 39504
rect 36760 39440 36776 39504
rect 36840 39440 36856 39504
rect 36920 39440 36936 39504
rect 37000 39440 37016 39504
rect 37080 39440 37096 39504
rect 37160 39440 37176 39504
rect 37240 39440 37256 39504
rect 37320 39440 37336 39504
rect 37400 39440 37416 39504
rect 37480 39440 37496 39504
rect 37560 39440 37576 39504
rect 37640 39440 37656 39504
rect 37720 39440 37736 39504
rect 37800 39440 37816 39504
rect 37880 39440 37896 39504
rect 37960 39440 37976 39504
rect 38040 39440 38056 39504
rect 38120 39440 38136 39504
rect 38200 39440 38216 39504
rect 38280 39440 38296 39504
rect 38360 39440 38376 39504
rect 38440 39440 38456 39504
rect 38520 39440 38536 39504
rect 38600 39440 38616 39504
rect 38680 39440 38696 39504
rect 38760 39440 38776 39504
rect 38840 39440 38856 39504
rect 38920 39440 38936 39504
rect 39000 39440 39016 39504
rect 39080 39440 39096 39504
rect 39160 39440 39176 39504
rect 39240 39440 39256 39504
rect 39320 39440 39336 39504
rect 39400 39440 39416 39504
rect 39480 39440 39496 39504
rect 39560 39440 39576 39504
rect 39640 39440 39656 39504
rect 39720 39440 39736 39504
rect 39800 39440 39816 39504
rect 39880 39440 39896 39504
rect 39960 39440 39976 39504
rect 40040 39440 40056 39504
rect 40120 39440 40136 39504
rect 40200 39440 40216 39504
rect 40280 39440 40296 39504
rect 40360 39440 40368 39504
rect 36368 39424 40368 39440
rect 36368 39360 36376 39424
rect 36440 39360 36456 39424
rect 36520 39360 36536 39424
rect 36600 39360 36616 39424
rect 36680 39360 36696 39424
rect 36760 39360 36776 39424
rect 36840 39360 36856 39424
rect 36920 39360 36936 39424
rect 37000 39360 37016 39424
rect 37080 39360 37096 39424
rect 37160 39360 37176 39424
rect 37240 39360 37256 39424
rect 37320 39360 37336 39424
rect 37400 39360 37416 39424
rect 37480 39360 37496 39424
rect 37560 39360 37576 39424
rect 37640 39360 37656 39424
rect 37720 39360 37736 39424
rect 37800 39360 37816 39424
rect 37880 39360 37896 39424
rect 37960 39360 37976 39424
rect 38040 39360 38056 39424
rect 38120 39360 38136 39424
rect 38200 39360 38216 39424
rect 38280 39360 38296 39424
rect 38360 39360 38376 39424
rect 38440 39360 38456 39424
rect 38520 39360 38536 39424
rect 38600 39360 38616 39424
rect 38680 39360 38696 39424
rect 38760 39360 38776 39424
rect 38840 39360 38856 39424
rect 38920 39360 38936 39424
rect 39000 39360 39016 39424
rect 39080 39360 39096 39424
rect 39160 39360 39176 39424
rect 39240 39360 39256 39424
rect 39320 39360 39336 39424
rect 39400 39360 39416 39424
rect 39480 39360 39496 39424
rect 39560 39360 39576 39424
rect 39640 39360 39656 39424
rect 39720 39360 39736 39424
rect 39800 39360 39816 39424
rect 39880 39360 39896 39424
rect 39960 39360 39976 39424
rect 40040 39360 40056 39424
rect 40120 39360 40136 39424
rect 40200 39360 40216 39424
rect 40280 39360 40296 39424
rect 40360 39360 40368 39424
rect 36368 39344 40368 39360
rect 36368 39280 36376 39344
rect 36440 39280 36456 39344
rect 36520 39280 36536 39344
rect 36600 39280 36616 39344
rect 36680 39280 36696 39344
rect 36760 39280 36776 39344
rect 36840 39280 36856 39344
rect 36920 39280 36936 39344
rect 37000 39280 37016 39344
rect 37080 39280 37096 39344
rect 37160 39280 37176 39344
rect 37240 39280 37256 39344
rect 37320 39280 37336 39344
rect 37400 39280 37416 39344
rect 37480 39280 37496 39344
rect 37560 39280 37576 39344
rect 37640 39280 37656 39344
rect 37720 39280 37736 39344
rect 37800 39280 37816 39344
rect 37880 39280 37896 39344
rect 37960 39280 37976 39344
rect 38040 39280 38056 39344
rect 38120 39280 38136 39344
rect 38200 39280 38216 39344
rect 38280 39280 38296 39344
rect 38360 39280 38376 39344
rect 38440 39280 38456 39344
rect 38520 39280 38536 39344
rect 38600 39280 38616 39344
rect 38680 39280 38696 39344
rect 38760 39280 38776 39344
rect 38840 39280 38856 39344
rect 38920 39280 38936 39344
rect 39000 39280 39016 39344
rect 39080 39280 39096 39344
rect 39160 39280 39176 39344
rect 39240 39280 39256 39344
rect 39320 39280 39336 39344
rect 39400 39280 39416 39344
rect 39480 39280 39496 39344
rect 39560 39280 39576 39344
rect 39640 39280 39656 39344
rect 39720 39280 39736 39344
rect 39800 39280 39816 39344
rect 39880 39280 39896 39344
rect 39960 39280 39976 39344
rect 40040 39280 40056 39344
rect 40120 39280 40136 39344
rect 40200 39280 40216 39344
rect 40280 39280 40296 39344
rect 40360 39280 40368 39344
rect 36368 39264 40368 39280
rect 36368 39200 36376 39264
rect 36440 39200 36456 39264
rect 36520 39200 36536 39264
rect 36600 39200 36616 39264
rect 36680 39200 36696 39264
rect 36760 39200 36776 39264
rect 36840 39200 36856 39264
rect 36920 39200 36936 39264
rect 37000 39200 37016 39264
rect 37080 39200 37096 39264
rect 37160 39200 37176 39264
rect 37240 39200 37256 39264
rect 37320 39200 37336 39264
rect 37400 39200 37416 39264
rect 37480 39200 37496 39264
rect 37560 39200 37576 39264
rect 37640 39200 37656 39264
rect 37720 39200 37736 39264
rect 37800 39200 37816 39264
rect 37880 39200 37896 39264
rect 37960 39200 37976 39264
rect 38040 39200 38056 39264
rect 38120 39200 38136 39264
rect 38200 39200 38216 39264
rect 38280 39200 38296 39264
rect 38360 39200 38376 39264
rect 38440 39200 38456 39264
rect 38520 39200 38536 39264
rect 38600 39200 38616 39264
rect 38680 39200 38696 39264
rect 38760 39200 38776 39264
rect 38840 39200 38856 39264
rect 38920 39200 38936 39264
rect 39000 39200 39016 39264
rect 39080 39200 39096 39264
rect 39160 39200 39176 39264
rect 39240 39200 39256 39264
rect 39320 39200 39336 39264
rect 39400 39200 39416 39264
rect 39480 39200 39496 39264
rect 39560 39200 39576 39264
rect 39640 39200 39656 39264
rect 39720 39200 39736 39264
rect 39800 39200 39816 39264
rect 39880 39200 39896 39264
rect 39960 39200 39976 39264
rect 40040 39200 40056 39264
rect 40120 39200 40136 39264
rect 40200 39200 40216 39264
rect 40280 39200 40296 39264
rect 40360 39200 40368 39264
rect 36368 39184 40368 39200
rect 36368 39120 36376 39184
rect 36440 39120 36456 39184
rect 36520 39120 36536 39184
rect 36600 39120 36616 39184
rect 36680 39120 36696 39184
rect 36760 39120 36776 39184
rect 36840 39120 36856 39184
rect 36920 39120 36936 39184
rect 37000 39120 37016 39184
rect 37080 39120 37096 39184
rect 37160 39120 37176 39184
rect 37240 39120 37256 39184
rect 37320 39120 37336 39184
rect 37400 39120 37416 39184
rect 37480 39120 37496 39184
rect 37560 39120 37576 39184
rect 37640 39120 37656 39184
rect 37720 39120 37736 39184
rect 37800 39120 37816 39184
rect 37880 39120 37896 39184
rect 37960 39120 37976 39184
rect 38040 39120 38056 39184
rect 38120 39120 38136 39184
rect 38200 39120 38216 39184
rect 38280 39120 38296 39184
rect 38360 39120 38376 39184
rect 38440 39120 38456 39184
rect 38520 39120 38536 39184
rect 38600 39120 38616 39184
rect 38680 39120 38696 39184
rect 38760 39120 38776 39184
rect 38840 39120 38856 39184
rect 38920 39120 38936 39184
rect 39000 39120 39016 39184
rect 39080 39120 39096 39184
rect 39160 39120 39176 39184
rect 39240 39120 39256 39184
rect 39320 39120 39336 39184
rect 39400 39120 39416 39184
rect 39480 39120 39496 39184
rect 39560 39120 39576 39184
rect 39640 39120 39656 39184
rect 39720 39120 39736 39184
rect 39800 39120 39816 39184
rect 39880 39120 39896 39184
rect 39960 39120 39976 39184
rect 40040 39120 40056 39184
rect 40120 39120 40136 39184
rect 40200 39120 40216 39184
rect 40280 39120 40296 39184
rect 40360 39120 40368 39184
rect 36368 39104 40368 39120
rect 36368 39040 36376 39104
rect 36440 39040 36456 39104
rect 36520 39040 36536 39104
rect 36600 39040 36616 39104
rect 36680 39040 36696 39104
rect 36760 39040 36776 39104
rect 36840 39040 36856 39104
rect 36920 39040 36936 39104
rect 37000 39040 37016 39104
rect 37080 39040 37096 39104
rect 37160 39040 37176 39104
rect 37240 39040 37256 39104
rect 37320 39040 37336 39104
rect 37400 39040 37416 39104
rect 37480 39040 37496 39104
rect 37560 39040 37576 39104
rect 37640 39040 37656 39104
rect 37720 39040 37736 39104
rect 37800 39040 37816 39104
rect 37880 39040 37896 39104
rect 37960 39040 37976 39104
rect 38040 39040 38056 39104
rect 38120 39040 38136 39104
rect 38200 39040 38216 39104
rect 38280 39040 38296 39104
rect 38360 39040 38376 39104
rect 38440 39040 38456 39104
rect 38520 39040 38536 39104
rect 38600 39040 38616 39104
rect 38680 39040 38696 39104
rect 38760 39040 38776 39104
rect 38840 39040 38856 39104
rect 38920 39040 38936 39104
rect 39000 39040 39016 39104
rect 39080 39040 39096 39104
rect 39160 39040 39176 39104
rect 39240 39040 39256 39104
rect 39320 39040 39336 39104
rect 39400 39040 39416 39104
rect 39480 39040 39496 39104
rect 39560 39040 39576 39104
rect 39640 39040 39656 39104
rect 39720 39040 39736 39104
rect 39800 39040 39816 39104
rect 39880 39040 39896 39104
rect 39960 39040 39976 39104
rect 40040 39040 40056 39104
rect 40120 39040 40136 39104
rect 40200 39040 40216 39104
rect 40280 39040 40296 39104
rect 40360 39040 40368 39104
rect 36368 39024 40368 39040
rect 36368 38960 36376 39024
rect 36440 38960 36456 39024
rect 36520 38960 36536 39024
rect 36600 38960 36616 39024
rect 36680 38960 36696 39024
rect 36760 38960 36776 39024
rect 36840 38960 36856 39024
rect 36920 38960 36936 39024
rect 37000 38960 37016 39024
rect 37080 38960 37096 39024
rect 37160 38960 37176 39024
rect 37240 38960 37256 39024
rect 37320 38960 37336 39024
rect 37400 38960 37416 39024
rect 37480 38960 37496 39024
rect 37560 38960 37576 39024
rect 37640 38960 37656 39024
rect 37720 38960 37736 39024
rect 37800 38960 37816 39024
rect 37880 38960 37896 39024
rect 37960 38960 37976 39024
rect 38040 38960 38056 39024
rect 38120 38960 38136 39024
rect 38200 38960 38216 39024
rect 38280 38960 38296 39024
rect 38360 38960 38376 39024
rect 38440 38960 38456 39024
rect 38520 38960 38536 39024
rect 38600 38960 38616 39024
rect 38680 38960 38696 39024
rect 38760 38960 38776 39024
rect 38840 38960 38856 39024
rect 38920 38960 38936 39024
rect 39000 38960 39016 39024
rect 39080 38960 39096 39024
rect 39160 38960 39176 39024
rect 39240 38960 39256 39024
rect 39320 38960 39336 39024
rect 39400 38960 39416 39024
rect 39480 38960 39496 39024
rect 39560 38960 39576 39024
rect 39640 38960 39656 39024
rect 39720 38960 39736 39024
rect 39800 38960 39816 39024
rect 39880 38960 39896 39024
rect 39960 38960 39976 39024
rect 40040 38960 40056 39024
rect 40120 38960 40136 39024
rect 40200 38960 40216 39024
rect 40280 38960 40296 39024
rect 40360 38960 40368 39024
rect 36368 38944 40368 38960
rect 36368 38880 36376 38944
rect 36440 38880 36456 38944
rect 36520 38880 36536 38944
rect 36600 38880 36616 38944
rect 36680 38880 36696 38944
rect 36760 38880 36776 38944
rect 36840 38880 36856 38944
rect 36920 38880 36936 38944
rect 37000 38880 37016 38944
rect 37080 38880 37096 38944
rect 37160 38880 37176 38944
rect 37240 38880 37256 38944
rect 37320 38880 37336 38944
rect 37400 38880 37416 38944
rect 37480 38880 37496 38944
rect 37560 38880 37576 38944
rect 37640 38880 37656 38944
rect 37720 38880 37736 38944
rect 37800 38880 37816 38944
rect 37880 38880 37896 38944
rect 37960 38880 37976 38944
rect 38040 38880 38056 38944
rect 38120 38880 38136 38944
rect 38200 38880 38216 38944
rect 38280 38880 38296 38944
rect 38360 38880 38376 38944
rect 38440 38880 38456 38944
rect 38520 38880 38536 38944
rect 38600 38880 38616 38944
rect 38680 38880 38696 38944
rect 38760 38880 38776 38944
rect 38840 38880 38856 38944
rect 38920 38880 38936 38944
rect 39000 38880 39016 38944
rect 39080 38880 39096 38944
rect 39160 38880 39176 38944
rect 39240 38880 39256 38944
rect 39320 38880 39336 38944
rect 39400 38880 39416 38944
rect 39480 38880 39496 38944
rect 39560 38880 39576 38944
rect 39640 38880 39656 38944
rect 39720 38880 39736 38944
rect 39800 38880 39816 38944
rect 39880 38880 39896 38944
rect 39960 38880 39976 38944
rect 40040 38880 40056 38944
rect 40120 38880 40136 38944
rect 40200 38880 40216 38944
rect 40280 38880 40296 38944
rect 40360 38880 40368 38944
rect 36368 38864 40368 38880
rect 36368 38800 36376 38864
rect 36440 38800 36456 38864
rect 36520 38800 36536 38864
rect 36600 38800 36616 38864
rect 36680 38800 36696 38864
rect 36760 38800 36776 38864
rect 36840 38800 36856 38864
rect 36920 38800 36936 38864
rect 37000 38800 37016 38864
rect 37080 38800 37096 38864
rect 37160 38800 37176 38864
rect 37240 38800 37256 38864
rect 37320 38800 37336 38864
rect 37400 38800 37416 38864
rect 37480 38800 37496 38864
rect 37560 38800 37576 38864
rect 37640 38800 37656 38864
rect 37720 38800 37736 38864
rect 37800 38800 37816 38864
rect 37880 38800 37896 38864
rect 37960 38800 37976 38864
rect 38040 38800 38056 38864
rect 38120 38800 38136 38864
rect 38200 38800 38216 38864
rect 38280 38800 38296 38864
rect 38360 38800 38376 38864
rect 38440 38800 38456 38864
rect 38520 38800 38536 38864
rect 38600 38800 38616 38864
rect 38680 38800 38696 38864
rect 38760 38800 38776 38864
rect 38840 38800 38856 38864
rect 38920 38800 38936 38864
rect 39000 38800 39016 38864
rect 39080 38800 39096 38864
rect 39160 38800 39176 38864
rect 39240 38800 39256 38864
rect 39320 38800 39336 38864
rect 39400 38800 39416 38864
rect 39480 38800 39496 38864
rect 39560 38800 39576 38864
rect 39640 38800 39656 38864
rect 39720 38800 39736 38864
rect 39800 38800 39816 38864
rect 39880 38800 39896 38864
rect 39960 38800 39976 38864
rect 40040 38800 40056 38864
rect 40120 38800 40136 38864
rect 40200 38800 40216 38864
rect 40280 38800 40296 38864
rect 40360 38800 40368 38864
rect 36368 38784 40368 38800
rect 36368 38720 36376 38784
rect 36440 38720 36456 38784
rect 36520 38720 36536 38784
rect 36600 38720 36616 38784
rect 36680 38720 36696 38784
rect 36760 38720 36776 38784
rect 36840 38720 36856 38784
rect 36920 38720 36936 38784
rect 37000 38720 37016 38784
rect 37080 38720 37096 38784
rect 37160 38720 37176 38784
rect 37240 38720 37256 38784
rect 37320 38720 37336 38784
rect 37400 38720 37416 38784
rect 37480 38720 37496 38784
rect 37560 38720 37576 38784
rect 37640 38720 37656 38784
rect 37720 38720 37736 38784
rect 37800 38720 37816 38784
rect 37880 38720 37896 38784
rect 37960 38720 37976 38784
rect 38040 38720 38056 38784
rect 38120 38720 38136 38784
rect 38200 38720 38216 38784
rect 38280 38720 38296 38784
rect 38360 38720 38376 38784
rect 38440 38720 38456 38784
rect 38520 38720 38536 38784
rect 38600 38720 38616 38784
rect 38680 38720 38696 38784
rect 38760 38720 38776 38784
rect 38840 38720 38856 38784
rect 38920 38720 38936 38784
rect 39000 38720 39016 38784
rect 39080 38720 39096 38784
rect 39160 38720 39176 38784
rect 39240 38720 39256 38784
rect 39320 38720 39336 38784
rect 39400 38720 39416 38784
rect 39480 38720 39496 38784
rect 39560 38720 39576 38784
rect 39640 38720 39656 38784
rect 39720 38720 39736 38784
rect 39800 38720 39816 38784
rect 39880 38720 39896 38784
rect 39960 38720 39976 38784
rect 40040 38720 40056 38784
rect 40120 38720 40136 38784
rect 40200 38720 40216 38784
rect 40280 38720 40296 38784
rect 40360 38720 40368 38784
rect 36368 38704 40368 38720
rect 36368 38640 36376 38704
rect 36440 38640 36456 38704
rect 36520 38640 36536 38704
rect 36600 38640 36616 38704
rect 36680 38640 36696 38704
rect 36760 38640 36776 38704
rect 36840 38640 36856 38704
rect 36920 38640 36936 38704
rect 37000 38640 37016 38704
rect 37080 38640 37096 38704
rect 37160 38640 37176 38704
rect 37240 38640 37256 38704
rect 37320 38640 37336 38704
rect 37400 38640 37416 38704
rect 37480 38640 37496 38704
rect 37560 38640 37576 38704
rect 37640 38640 37656 38704
rect 37720 38640 37736 38704
rect 37800 38640 37816 38704
rect 37880 38640 37896 38704
rect 37960 38640 37976 38704
rect 38040 38640 38056 38704
rect 38120 38640 38136 38704
rect 38200 38640 38216 38704
rect 38280 38640 38296 38704
rect 38360 38640 38376 38704
rect 38440 38640 38456 38704
rect 38520 38640 38536 38704
rect 38600 38640 38616 38704
rect 38680 38640 38696 38704
rect 38760 38640 38776 38704
rect 38840 38640 38856 38704
rect 38920 38640 38936 38704
rect 39000 38640 39016 38704
rect 39080 38640 39096 38704
rect 39160 38640 39176 38704
rect 39240 38640 39256 38704
rect 39320 38640 39336 38704
rect 39400 38640 39416 38704
rect 39480 38640 39496 38704
rect 39560 38640 39576 38704
rect 39640 38640 39656 38704
rect 39720 38640 39736 38704
rect 39800 38640 39816 38704
rect 39880 38640 39896 38704
rect 39960 38640 39976 38704
rect 40040 38640 40056 38704
rect 40120 38640 40136 38704
rect 40200 38640 40216 38704
rect 40280 38640 40296 38704
rect 40360 38640 40368 38704
rect 36368 38624 40368 38640
rect 36368 38560 36376 38624
rect 36440 38560 36456 38624
rect 36520 38560 36536 38624
rect 36600 38560 36616 38624
rect 36680 38560 36696 38624
rect 36760 38560 36776 38624
rect 36840 38560 36856 38624
rect 36920 38560 36936 38624
rect 37000 38560 37016 38624
rect 37080 38560 37096 38624
rect 37160 38560 37176 38624
rect 37240 38560 37256 38624
rect 37320 38560 37336 38624
rect 37400 38560 37416 38624
rect 37480 38560 37496 38624
rect 37560 38560 37576 38624
rect 37640 38560 37656 38624
rect 37720 38560 37736 38624
rect 37800 38560 37816 38624
rect 37880 38560 37896 38624
rect 37960 38560 37976 38624
rect 38040 38560 38056 38624
rect 38120 38560 38136 38624
rect 38200 38560 38216 38624
rect 38280 38560 38296 38624
rect 38360 38560 38376 38624
rect 38440 38560 38456 38624
rect 38520 38560 38536 38624
rect 38600 38560 38616 38624
rect 38680 38560 38696 38624
rect 38760 38560 38776 38624
rect 38840 38560 38856 38624
rect 38920 38560 38936 38624
rect 39000 38560 39016 38624
rect 39080 38560 39096 38624
rect 39160 38560 39176 38624
rect 39240 38560 39256 38624
rect 39320 38560 39336 38624
rect 39400 38560 39416 38624
rect 39480 38560 39496 38624
rect 39560 38560 39576 38624
rect 39640 38560 39656 38624
rect 39720 38560 39736 38624
rect 39800 38560 39816 38624
rect 39880 38560 39896 38624
rect 39960 38560 39976 38624
rect 40040 38560 40056 38624
rect 40120 38560 40136 38624
rect 40200 38560 40216 38624
rect 40280 38560 40296 38624
rect 40360 38560 40368 38624
rect 36368 38544 40368 38560
rect 36368 38480 36376 38544
rect 36440 38480 36456 38544
rect 36520 38480 36536 38544
rect 36600 38480 36616 38544
rect 36680 38480 36696 38544
rect 36760 38480 36776 38544
rect 36840 38480 36856 38544
rect 36920 38480 36936 38544
rect 37000 38480 37016 38544
rect 37080 38480 37096 38544
rect 37160 38480 37176 38544
rect 37240 38480 37256 38544
rect 37320 38480 37336 38544
rect 37400 38480 37416 38544
rect 37480 38480 37496 38544
rect 37560 38480 37576 38544
rect 37640 38480 37656 38544
rect 37720 38480 37736 38544
rect 37800 38480 37816 38544
rect 37880 38480 37896 38544
rect 37960 38480 37976 38544
rect 38040 38480 38056 38544
rect 38120 38480 38136 38544
rect 38200 38480 38216 38544
rect 38280 38480 38296 38544
rect 38360 38480 38376 38544
rect 38440 38480 38456 38544
rect 38520 38480 38536 38544
rect 38600 38480 38616 38544
rect 38680 38480 38696 38544
rect 38760 38480 38776 38544
rect 38840 38480 38856 38544
rect 38920 38480 38936 38544
rect 39000 38480 39016 38544
rect 39080 38480 39096 38544
rect 39160 38480 39176 38544
rect 39240 38480 39256 38544
rect 39320 38480 39336 38544
rect 39400 38480 39416 38544
rect 39480 38480 39496 38544
rect 39560 38480 39576 38544
rect 39640 38480 39656 38544
rect 39720 38480 39736 38544
rect 39800 38480 39816 38544
rect 39880 38480 39896 38544
rect 39960 38480 39976 38544
rect 40040 38480 40056 38544
rect 40120 38480 40136 38544
rect 40200 38480 40216 38544
rect 40280 38480 40296 38544
rect 40360 38480 40368 38544
rect 36368 38464 40368 38480
rect 36368 38400 36376 38464
rect 36440 38400 36456 38464
rect 36520 38400 36536 38464
rect 36600 38400 36616 38464
rect 36680 38400 36696 38464
rect 36760 38400 36776 38464
rect 36840 38400 36856 38464
rect 36920 38400 36936 38464
rect 37000 38400 37016 38464
rect 37080 38400 37096 38464
rect 37160 38400 37176 38464
rect 37240 38400 37256 38464
rect 37320 38400 37336 38464
rect 37400 38400 37416 38464
rect 37480 38400 37496 38464
rect 37560 38400 37576 38464
rect 37640 38400 37656 38464
rect 37720 38400 37736 38464
rect 37800 38400 37816 38464
rect 37880 38400 37896 38464
rect 37960 38400 37976 38464
rect 38040 38400 38056 38464
rect 38120 38400 38136 38464
rect 38200 38400 38216 38464
rect 38280 38400 38296 38464
rect 38360 38400 38376 38464
rect 38440 38400 38456 38464
rect 38520 38400 38536 38464
rect 38600 38400 38616 38464
rect 38680 38400 38696 38464
rect 38760 38400 38776 38464
rect 38840 38400 38856 38464
rect 38920 38400 38936 38464
rect 39000 38400 39016 38464
rect 39080 38400 39096 38464
rect 39160 38400 39176 38464
rect 39240 38400 39256 38464
rect 39320 38400 39336 38464
rect 39400 38400 39416 38464
rect 39480 38400 39496 38464
rect 39560 38400 39576 38464
rect 39640 38400 39656 38464
rect 39720 38400 39736 38464
rect 39800 38400 39816 38464
rect 39880 38400 39896 38464
rect 39960 38400 39976 38464
rect 40040 38400 40056 38464
rect 40120 38400 40136 38464
rect 40200 38400 40216 38464
rect 40280 38400 40296 38464
rect 40360 38400 40368 38464
rect 36368 38384 40368 38400
rect 36368 38320 36376 38384
rect 36440 38320 36456 38384
rect 36520 38320 36536 38384
rect 36600 38320 36616 38384
rect 36680 38320 36696 38384
rect 36760 38320 36776 38384
rect 36840 38320 36856 38384
rect 36920 38320 36936 38384
rect 37000 38320 37016 38384
rect 37080 38320 37096 38384
rect 37160 38320 37176 38384
rect 37240 38320 37256 38384
rect 37320 38320 37336 38384
rect 37400 38320 37416 38384
rect 37480 38320 37496 38384
rect 37560 38320 37576 38384
rect 37640 38320 37656 38384
rect 37720 38320 37736 38384
rect 37800 38320 37816 38384
rect 37880 38320 37896 38384
rect 37960 38320 37976 38384
rect 38040 38320 38056 38384
rect 38120 38320 38136 38384
rect 38200 38320 38216 38384
rect 38280 38320 38296 38384
rect 38360 38320 38376 38384
rect 38440 38320 38456 38384
rect 38520 38320 38536 38384
rect 38600 38320 38616 38384
rect 38680 38320 38696 38384
rect 38760 38320 38776 38384
rect 38840 38320 38856 38384
rect 38920 38320 38936 38384
rect 39000 38320 39016 38384
rect 39080 38320 39096 38384
rect 39160 38320 39176 38384
rect 39240 38320 39256 38384
rect 39320 38320 39336 38384
rect 39400 38320 39416 38384
rect 39480 38320 39496 38384
rect 39560 38320 39576 38384
rect 39640 38320 39656 38384
rect 39720 38320 39736 38384
rect 39800 38320 39816 38384
rect 39880 38320 39896 38384
rect 39960 38320 39976 38384
rect 40040 38320 40056 38384
rect 40120 38320 40136 38384
rect 40200 38320 40216 38384
rect 40280 38320 40296 38384
rect 40360 38320 40368 38384
rect 36368 38304 40368 38320
rect 36368 38240 36376 38304
rect 36440 38240 36456 38304
rect 36520 38240 36536 38304
rect 36600 38240 36616 38304
rect 36680 38240 36696 38304
rect 36760 38240 36776 38304
rect 36840 38240 36856 38304
rect 36920 38240 36936 38304
rect 37000 38240 37016 38304
rect 37080 38240 37096 38304
rect 37160 38240 37176 38304
rect 37240 38240 37256 38304
rect 37320 38240 37336 38304
rect 37400 38240 37416 38304
rect 37480 38240 37496 38304
rect 37560 38240 37576 38304
rect 37640 38240 37656 38304
rect 37720 38240 37736 38304
rect 37800 38240 37816 38304
rect 37880 38240 37896 38304
rect 37960 38240 37976 38304
rect 38040 38240 38056 38304
rect 38120 38240 38136 38304
rect 38200 38240 38216 38304
rect 38280 38240 38296 38304
rect 38360 38240 38376 38304
rect 38440 38240 38456 38304
rect 38520 38240 38536 38304
rect 38600 38240 38616 38304
rect 38680 38240 38696 38304
rect 38760 38240 38776 38304
rect 38840 38240 38856 38304
rect 38920 38240 38936 38304
rect 39000 38240 39016 38304
rect 39080 38240 39096 38304
rect 39160 38240 39176 38304
rect 39240 38240 39256 38304
rect 39320 38240 39336 38304
rect 39400 38240 39416 38304
rect 39480 38240 39496 38304
rect 39560 38240 39576 38304
rect 39640 38240 39656 38304
rect 39720 38240 39736 38304
rect 39800 38240 39816 38304
rect 39880 38240 39896 38304
rect 39960 38240 39976 38304
rect 40040 38240 40056 38304
rect 40120 38240 40136 38304
rect 40200 38240 40216 38304
rect 40280 38240 40296 38304
rect 40360 38240 40368 38304
rect 36368 38224 40368 38240
rect 36368 38160 36376 38224
rect 36440 38160 36456 38224
rect 36520 38160 36536 38224
rect 36600 38160 36616 38224
rect 36680 38160 36696 38224
rect 36760 38160 36776 38224
rect 36840 38160 36856 38224
rect 36920 38160 36936 38224
rect 37000 38160 37016 38224
rect 37080 38160 37096 38224
rect 37160 38160 37176 38224
rect 37240 38160 37256 38224
rect 37320 38160 37336 38224
rect 37400 38160 37416 38224
rect 37480 38160 37496 38224
rect 37560 38160 37576 38224
rect 37640 38160 37656 38224
rect 37720 38160 37736 38224
rect 37800 38160 37816 38224
rect 37880 38160 37896 38224
rect 37960 38160 37976 38224
rect 38040 38160 38056 38224
rect 38120 38160 38136 38224
rect 38200 38160 38216 38224
rect 38280 38160 38296 38224
rect 38360 38160 38376 38224
rect 38440 38160 38456 38224
rect 38520 38160 38536 38224
rect 38600 38160 38616 38224
rect 38680 38160 38696 38224
rect 38760 38160 38776 38224
rect 38840 38160 38856 38224
rect 38920 38160 38936 38224
rect 39000 38160 39016 38224
rect 39080 38160 39096 38224
rect 39160 38160 39176 38224
rect 39240 38160 39256 38224
rect 39320 38160 39336 38224
rect 39400 38160 39416 38224
rect 39480 38160 39496 38224
rect 39560 38160 39576 38224
rect 39640 38160 39656 38224
rect 39720 38160 39736 38224
rect 39800 38160 39816 38224
rect 39880 38160 39896 38224
rect 39960 38160 39976 38224
rect 40040 38160 40056 38224
rect 40120 38160 40136 38224
rect 40200 38160 40216 38224
rect 40280 38160 40296 38224
rect 40360 38160 40368 38224
rect 36368 38144 40368 38160
rect 36368 38080 36376 38144
rect 36440 38080 36456 38144
rect 36520 38080 36536 38144
rect 36600 38080 36616 38144
rect 36680 38080 36696 38144
rect 36760 38080 36776 38144
rect 36840 38080 36856 38144
rect 36920 38080 36936 38144
rect 37000 38080 37016 38144
rect 37080 38080 37096 38144
rect 37160 38080 37176 38144
rect 37240 38080 37256 38144
rect 37320 38080 37336 38144
rect 37400 38080 37416 38144
rect 37480 38080 37496 38144
rect 37560 38080 37576 38144
rect 37640 38080 37656 38144
rect 37720 38080 37736 38144
rect 37800 38080 37816 38144
rect 37880 38080 37896 38144
rect 37960 38080 37976 38144
rect 38040 38080 38056 38144
rect 38120 38080 38136 38144
rect 38200 38080 38216 38144
rect 38280 38080 38296 38144
rect 38360 38080 38376 38144
rect 38440 38080 38456 38144
rect 38520 38080 38536 38144
rect 38600 38080 38616 38144
rect 38680 38080 38696 38144
rect 38760 38080 38776 38144
rect 38840 38080 38856 38144
rect 38920 38080 38936 38144
rect 39000 38080 39016 38144
rect 39080 38080 39096 38144
rect 39160 38080 39176 38144
rect 39240 38080 39256 38144
rect 39320 38080 39336 38144
rect 39400 38080 39416 38144
rect 39480 38080 39496 38144
rect 39560 38080 39576 38144
rect 39640 38080 39656 38144
rect 39720 38080 39736 38144
rect 39800 38080 39816 38144
rect 39880 38080 39896 38144
rect 39960 38080 39976 38144
rect 40040 38080 40056 38144
rect 40120 38080 40136 38144
rect 40200 38080 40216 38144
rect 40280 38080 40296 38144
rect 40360 38080 40368 38144
rect 36368 38064 40368 38080
rect 36368 38000 36376 38064
rect 36440 38000 36456 38064
rect 36520 38000 36536 38064
rect 36600 38000 36616 38064
rect 36680 38000 36696 38064
rect 36760 38000 36776 38064
rect 36840 38000 36856 38064
rect 36920 38000 36936 38064
rect 37000 38000 37016 38064
rect 37080 38000 37096 38064
rect 37160 38000 37176 38064
rect 37240 38000 37256 38064
rect 37320 38000 37336 38064
rect 37400 38000 37416 38064
rect 37480 38000 37496 38064
rect 37560 38000 37576 38064
rect 37640 38000 37656 38064
rect 37720 38000 37736 38064
rect 37800 38000 37816 38064
rect 37880 38000 37896 38064
rect 37960 38000 37976 38064
rect 38040 38000 38056 38064
rect 38120 38000 38136 38064
rect 38200 38000 38216 38064
rect 38280 38000 38296 38064
rect 38360 38000 38376 38064
rect 38440 38000 38456 38064
rect 38520 38000 38536 38064
rect 38600 38000 38616 38064
rect 38680 38000 38696 38064
rect 38760 38000 38776 38064
rect 38840 38000 38856 38064
rect 38920 38000 38936 38064
rect 39000 38000 39016 38064
rect 39080 38000 39096 38064
rect 39160 38000 39176 38064
rect 39240 38000 39256 38064
rect 39320 38000 39336 38064
rect 39400 38000 39416 38064
rect 39480 38000 39496 38064
rect 39560 38000 39576 38064
rect 39640 38000 39656 38064
rect 39720 38000 39736 38064
rect 39800 38000 39816 38064
rect 39880 38000 39896 38064
rect 39960 38000 39976 38064
rect 40040 38000 40056 38064
rect 40120 38000 40136 38064
rect 40200 38000 40216 38064
rect 40280 38000 40296 38064
rect 40360 38000 40368 38064
rect 36368 37984 40368 38000
rect 36368 37920 36376 37984
rect 36440 37920 36456 37984
rect 36520 37920 36536 37984
rect 36600 37920 36616 37984
rect 36680 37920 36696 37984
rect 36760 37920 36776 37984
rect 36840 37920 36856 37984
rect 36920 37920 36936 37984
rect 37000 37920 37016 37984
rect 37080 37920 37096 37984
rect 37160 37920 37176 37984
rect 37240 37920 37256 37984
rect 37320 37920 37336 37984
rect 37400 37920 37416 37984
rect 37480 37920 37496 37984
rect 37560 37920 37576 37984
rect 37640 37920 37656 37984
rect 37720 37920 37736 37984
rect 37800 37920 37816 37984
rect 37880 37920 37896 37984
rect 37960 37920 37976 37984
rect 38040 37920 38056 37984
rect 38120 37920 38136 37984
rect 38200 37920 38216 37984
rect 38280 37920 38296 37984
rect 38360 37920 38376 37984
rect 38440 37920 38456 37984
rect 38520 37920 38536 37984
rect 38600 37920 38616 37984
rect 38680 37920 38696 37984
rect 38760 37920 38776 37984
rect 38840 37920 38856 37984
rect 38920 37920 38936 37984
rect 39000 37920 39016 37984
rect 39080 37920 39096 37984
rect 39160 37920 39176 37984
rect 39240 37920 39256 37984
rect 39320 37920 39336 37984
rect 39400 37920 39416 37984
rect 39480 37920 39496 37984
rect 39560 37920 39576 37984
rect 39640 37920 39656 37984
rect 39720 37920 39736 37984
rect 39800 37920 39816 37984
rect 39880 37920 39896 37984
rect 39960 37920 39976 37984
rect 40040 37920 40056 37984
rect 40120 37920 40136 37984
rect 40200 37920 40216 37984
rect 40280 37920 40296 37984
rect 40360 37920 40368 37984
rect 36368 37904 40368 37920
rect 36368 37840 36376 37904
rect 36440 37840 36456 37904
rect 36520 37840 36536 37904
rect 36600 37840 36616 37904
rect 36680 37840 36696 37904
rect 36760 37840 36776 37904
rect 36840 37840 36856 37904
rect 36920 37840 36936 37904
rect 37000 37840 37016 37904
rect 37080 37840 37096 37904
rect 37160 37840 37176 37904
rect 37240 37840 37256 37904
rect 37320 37840 37336 37904
rect 37400 37840 37416 37904
rect 37480 37840 37496 37904
rect 37560 37840 37576 37904
rect 37640 37840 37656 37904
rect 37720 37840 37736 37904
rect 37800 37840 37816 37904
rect 37880 37840 37896 37904
rect 37960 37840 37976 37904
rect 38040 37840 38056 37904
rect 38120 37840 38136 37904
rect 38200 37840 38216 37904
rect 38280 37840 38296 37904
rect 38360 37840 38376 37904
rect 38440 37840 38456 37904
rect 38520 37840 38536 37904
rect 38600 37840 38616 37904
rect 38680 37840 38696 37904
rect 38760 37840 38776 37904
rect 38840 37840 38856 37904
rect 38920 37840 38936 37904
rect 39000 37840 39016 37904
rect 39080 37840 39096 37904
rect 39160 37840 39176 37904
rect 39240 37840 39256 37904
rect 39320 37840 39336 37904
rect 39400 37840 39416 37904
rect 39480 37840 39496 37904
rect 39560 37840 39576 37904
rect 39640 37840 39656 37904
rect 39720 37840 39736 37904
rect 39800 37840 39816 37904
rect 39880 37840 39896 37904
rect 39960 37840 39976 37904
rect 40040 37840 40056 37904
rect 40120 37840 40136 37904
rect 40200 37840 40216 37904
rect 40280 37840 40296 37904
rect 40360 37840 40368 37904
rect 36368 37824 40368 37840
rect 36368 37760 36376 37824
rect 36440 37760 36456 37824
rect 36520 37760 36536 37824
rect 36600 37760 36616 37824
rect 36680 37760 36696 37824
rect 36760 37760 36776 37824
rect 36840 37760 36856 37824
rect 36920 37760 36936 37824
rect 37000 37760 37016 37824
rect 37080 37760 37096 37824
rect 37160 37760 37176 37824
rect 37240 37760 37256 37824
rect 37320 37760 37336 37824
rect 37400 37760 37416 37824
rect 37480 37760 37496 37824
rect 37560 37760 37576 37824
rect 37640 37760 37656 37824
rect 37720 37760 37736 37824
rect 37800 37760 37816 37824
rect 37880 37760 37896 37824
rect 37960 37760 37976 37824
rect 38040 37760 38056 37824
rect 38120 37760 38136 37824
rect 38200 37760 38216 37824
rect 38280 37760 38296 37824
rect 38360 37760 38376 37824
rect 38440 37760 38456 37824
rect 38520 37760 38536 37824
rect 38600 37760 38616 37824
rect 38680 37760 38696 37824
rect 38760 37760 38776 37824
rect 38840 37760 38856 37824
rect 38920 37760 38936 37824
rect 39000 37760 39016 37824
rect 39080 37760 39096 37824
rect 39160 37760 39176 37824
rect 39240 37760 39256 37824
rect 39320 37760 39336 37824
rect 39400 37760 39416 37824
rect 39480 37760 39496 37824
rect 39560 37760 39576 37824
rect 39640 37760 39656 37824
rect 39720 37760 39736 37824
rect 39800 37760 39816 37824
rect 39880 37760 39896 37824
rect 39960 37760 39976 37824
rect 40040 37760 40056 37824
rect 40120 37760 40136 37824
rect 40200 37760 40216 37824
rect 40280 37760 40296 37824
rect 40360 37760 40368 37824
rect 36368 37744 40368 37760
rect 36368 37680 36376 37744
rect 36440 37680 36456 37744
rect 36520 37680 36536 37744
rect 36600 37680 36616 37744
rect 36680 37680 36696 37744
rect 36760 37680 36776 37744
rect 36840 37680 36856 37744
rect 36920 37680 36936 37744
rect 37000 37680 37016 37744
rect 37080 37680 37096 37744
rect 37160 37680 37176 37744
rect 37240 37680 37256 37744
rect 37320 37680 37336 37744
rect 37400 37680 37416 37744
rect 37480 37680 37496 37744
rect 37560 37680 37576 37744
rect 37640 37680 37656 37744
rect 37720 37680 37736 37744
rect 37800 37680 37816 37744
rect 37880 37680 37896 37744
rect 37960 37680 37976 37744
rect 38040 37680 38056 37744
rect 38120 37680 38136 37744
rect 38200 37680 38216 37744
rect 38280 37680 38296 37744
rect 38360 37680 38376 37744
rect 38440 37680 38456 37744
rect 38520 37680 38536 37744
rect 38600 37680 38616 37744
rect 38680 37680 38696 37744
rect 38760 37680 38776 37744
rect 38840 37680 38856 37744
rect 38920 37680 38936 37744
rect 39000 37680 39016 37744
rect 39080 37680 39096 37744
rect 39160 37680 39176 37744
rect 39240 37680 39256 37744
rect 39320 37680 39336 37744
rect 39400 37680 39416 37744
rect 39480 37680 39496 37744
rect 39560 37680 39576 37744
rect 39640 37680 39656 37744
rect 39720 37680 39736 37744
rect 39800 37680 39816 37744
rect 39880 37680 39896 37744
rect 39960 37680 39976 37744
rect 40040 37680 40056 37744
rect 40120 37680 40136 37744
rect 40200 37680 40216 37744
rect 40280 37680 40296 37744
rect 40360 37680 40368 37744
rect 36368 37664 40368 37680
rect 36368 37600 36376 37664
rect 36440 37600 36456 37664
rect 36520 37600 36536 37664
rect 36600 37600 36616 37664
rect 36680 37600 36696 37664
rect 36760 37600 36776 37664
rect 36840 37600 36856 37664
rect 36920 37600 36936 37664
rect 37000 37600 37016 37664
rect 37080 37600 37096 37664
rect 37160 37600 37176 37664
rect 37240 37600 37256 37664
rect 37320 37600 37336 37664
rect 37400 37600 37416 37664
rect 37480 37600 37496 37664
rect 37560 37600 37576 37664
rect 37640 37600 37656 37664
rect 37720 37600 37736 37664
rect 37800 37600 37816 37664
rect 37880 37600 37896 37664
rect 37960 37600 37976 37664
rect 38040 37600 38056 37664
rect 38120 37600 38136 37664
rect 38200 37600 38216 37664
rect 38280 37600 38296 37664
rect 38360 37600 38376 37664
rect 38440 37600 38456 37664
rect 38520 37600 38536 37664
rect 38600 37600 38616 37664
rect 38680 37600 38696 37664
rect 38760 37600 38776 37664
rect 38840 37600 38856 37664
rect 38920 37600 38936 37664
rect 39000 37600 39016 37664
rect 39080 37600 39096 37664
rect 39160 37600 39176 37664
rect 39240 37600 39256 37664
rect 39320 37600 39336 37664
rect 39400 37600 39416 37664
rect 39480 37600 39496 37664
rect 39560 37600 39576 37664
rect 39640 37600 39656 37664
rect 39720 37600 39736 37664
rect 39800 37600 39816 37664
rect 39880 37600 39896 37664
rect 39960 37600 39976 37664
rect 40040 37600 40056 37664
rect 40120 37600 40136 37664
rect 40200 37600 40216 37664
rect 40280 37600 40296 37664
rect 40360 37600 40368 37664
rect 36368 37584 40368 37600
rect 36368 37520 36376 37584
rect 36440 37520 36456 37584
rect 36520 37520 36536 37584
rect 36600 37520 36616 37584
rect 36680 37520 36696 37584
rect 36760 37520 36776 37584
rect 36840 37520 36856 37584
rect 36920 37520 36936 37584
rect 37000 37520 37016 37584
rect 37080 37520 37096 37584
rect 37160 37520 37176 37584
rect 37240 37520 37256 37584
rect 37320 37520 37336 37584
rect 37400 37520 37416 37584
rect 37480 37520 37496 37584
rect 37560 37520 37576 37584
rect 37640 37520 37656 37584
rect 37720 37520 37736 37584
rect 37800 37520 37816 37584
rect 37880 37520 37896 37584
rect 37960 37520 37976 37584
rect 38040 37520 38056 37584
rect 38120 37520 38136 37584
rect 38200 37520 38216 37584
rect 38280 37520 38296 37584
rect 38360 37520 38376 37584
rect 38440 37520 38456 37584
rect 38520 37520 38536 37584
rect 38600 37520 38616 37584
rect 38680 37520 38696 37584
rect 38760 37520 38776 37584
rect 38840 37520 38856 37584
rect 38920 37520 38936 37584
rect 39000 37520 39016 37584
rect 39080 37520 39096 37584
rect 39160 37520 39176 37584
rect 39240 37520 39256 37584
rect 39320 37520 39336 37584
rect 39400 37520 39416 37584
rect 39480 37520 39496 37584
rect 39560 37520 39576 37584
rect 39640 37520 39656 37584
rect 39720 37520 39736 37584
rect 39800 37520 39816 37584
rect 39880 37520 39896 37584
rect 39960 37520 39976 37584
rect 40040 37520 40056 37584
rect 40120 37520 40136 37584
rect 40200 37520 40216 37584
rect 40280 37520 40296 37584
rect 40360 37520 40368 37584
rect 36368 37504 40368 37520
rect 36368 37440 36376 37504
rect 36440 37440 36456 37504
rect 36520 37440 36536 37504
rect 36600 37440 36616 37504
rect 36680 37440 36696 37504
rect 36760 37440 36776 37504
rect 36840 37440 36856 37504
rect 36920 37440 36936 37504
rect 37000 37440 37016 37504
rect 37080 37440 37096 37504
rect 37160 37440 37176 37504
rect 37240 37440 37256 37504
rect 37320 37440 37336 37504
rect 37400 37440 37416 37504
rect 37480 37440 37496 37504
rect 37560 37440 37576 37504
rect 37640 37440 37656 37504
rect 37720 37440 37736 37504
rect 37800 37440 37816 37504
rect 37880 37440 37896 37504
rect 37960 37440 37976 37504
rect 38040 37440 38056 37504
rect 38120 37440 38136 37504
rect 38200 37440 38216 37504
rect 38280 37440 38296 37504
rect 38360 37440 38376 37504
rect 38440 37440 38456 37504
rect 38520 37440 38536 37504
rect 38600 37440 38616 37504
rect 38680 37440 38696 37504
rect 38760 37440 38776 37504
rect 38840 37440 38856 37504
rect 38920 37440 38936 37504
rect 39000 37440 39016 37504
rect 39080 37440 39096 37504
rect 39160 37440 39176 37504
rect 39240 37440 39256 37504
rect 39320 37440 39336 37504
rect 39400 37440 39416 37504
rect 39480 37440 39496 37504
rect 39560 37440 39576 37504
rect 39640 37440 39656 37504
rect 39720 37440 39736 37504
rect 39800 37440 39816 37504
rect 39880 37440 39896 37504
rect 39960 37440 39976 37504
rect 40040 37440 40056 37504
rect 40120 37440 40136 37504
rect 40200 37440 40216 37504
rect 40280 37440 40296 37504
rect 40360 37440 40368 37504
rect 36368 37424 40368 37440
rect 36368 37360 36376 37424
rect 36440 37360 36456 37424
rect 36520 37360 36536 37424
rect 36600 37360 36616 37424
rect 36680 37360 36696 37424
rect 36760 37360 36776 37424
rect 36840 37360 36856 37424
rect 36920 37360 36936 37424
rect 37000 37360 37016 37424
rect 37080 37360 37096 37424
rect 37160 37360 37176 37424
rect 37240 37360 37256 37424
rect 37320 37360 37336 37424
rect 37400 37360 37416 37424
rect 37480 37360 37496 37424
rect 37560 37360 37576 37424
rect 37640 37360 37656 37424
rect 37720 37360 37736 37424
rect 37800 37360 37816 37424
rect 37880 37360 37896 37424
rect 37960 37360 37976 37424
rect 38040 37360 38056 37424
rect 38120 37360 38136 37424
rect 38200 37360 38216 37424
rect 38280 37360 38296 37424
rect 38360 37360 38376 37424
rect 38440 37360 38456 37424
rect 38520 37360 38536 37424
rect 38600 37360 38616 37424
rect 38680 37360 38696 37424
rect 38760 37360 38776 37424
rect 38840 37360 38856 37424
rect 38920 37360 38936 37424
rect 39000 37360 39016 37424
rect 39080 37360 39096 37424
rect 39160 37360 39176 37424
rect 39240 37360 39256 37424
rect 39320 37360 39336 37424
rect 39400 37360 39416 37424
rect 39480 37360 39496 37424
rect 39560 37360 39576 37424
rect 39640 37360 39656 37424
rect 39720 37360 39736 37424
rect 39800 37360 39816 37424
rect 39880 37360 39896 37424
rect 39960 37360 39976 37424
rect 40040 37360 40056 37424
rect 40120 37360 40136 37424
rect 40200 37360 40216 37424
rect 40280 37360 40296 37424
rect 40360 37360 40368 37424
rect 36368 37344 40368 37360
rect 36368 37280 36376 37344
rect 36440 37280 36456 37344
rect 36520 37280 36536 37344
rect 36600 37280 36616 37344
rect 36680 37280 36696 37344
rect 36760 37280 36776 37344
rect 36840 37280 36856 37344
rect 36920 37280 36936 37344
rect 37000 37280 37016 37344
rect 37080 37280 37096 37344
rect 37160 37280 37176 37344
rect 37240 37280 37256 37344
rect 37320 37280 37336 37344
rect 37400 37280 37416 37344
rect 37480 37280 37496 37344
rect 37560 37280 37576 37344
rect 37640 37280 37656 37344
rect 37720 37280 37736 37344
rect 37800 37280 37816 37344
rect 37880 37280 37896 37344
rect 37960 37280 37976 37344
rect 38040 37280 38056 37344
rect 38120 37280 38136 37344
rect 38200 37280 38216 37344
rect 38280 37280 38296 37344
rect 38360 37280 38376 37344
rect 38440 37280 38456 37344
rect 38520 37280 38536 37344
rect 38600 37280 38616 37344
rect 38680 37280 38696 37344
rect 38760 37280 38776 37344
rect 38840 37280 38856 37344
rect 38920 37280 38936 37344
rect 39000 37280 39016 37344
rect 39080 37280 39096 37344
rect 39160 37280 39176 37344
rect 39240 37280 39256 37344
rect 39320 37280 39336 37344
rect 39400 37280 39416 37344
rect 39480 37280 39496 37344
rect 39560 37280 39576 37344
rect 39640 37280 39656 37344
rect 39720 37280 39736 37344
rect 39800 37280 39816 37344
rect 39880 37280 39896 37344
rect 39960 37280 39976 37344
rect 40040 37280 40056 37344
rect 40120 37280 40136 37344
rect 40200 37280 40216 37344
rect 40280 37280 40296 37344
rect 40360 37280 40368 37344
rect 36368 37264 40368 37280
rect 36368 37200 36376 37264
rect 36440 37200 36456 37264
rect 36520 37200 36536 37264
rect 36600 37200 36616 37264
rect 36680 37200 36696 37264
rect 36760 37200 36776 37264
rect 36840 37200 36856 37264
rect 36920 37200 36936 37264
rect 37000 37200 37016 37264
rect 37080 37200 37096 37264
rect 37160 37200 37176 37264
rect 37240 37200 37256 37264
rect 37320 37200 37336 37264
rect 37400 37200 37416 37264
rect 37480 37200 37496 37264
rect 37560 37200 37576 37264
rect 37640 37200 37656 37264
rect 37720 37200 37736 37264
rect 37800 37200 37816 37264
rect 37880 37200 37896 37264
rect 37960 37200 37976 37264
rect 38040 37200 38056 37264
rect 38120 37200 38136 37264
rect 38200 37200 38216 37264
rect 38280 37200 38296 37264
rect 38360 37200 38376 37264
rect 38440 37200 38456 37264
rect 38520 37200 38536 37264
rect 38600 37200 38616 37264
rect 38680 37200 38696 37264
rect 38760 37200 38776 37264
rect 38840 37200 38856 37264
rect 38920 37200 38936 37264
rect 39000 37200 39016 37264
rect 39080 37200 39096 37264
rect 39160 37200 39176 37264
rect 39240 37200 39256 37264
rect 39320 37200 39336 37264
rect 39400 37200 39416 37264
rect 39480 37200 39496 37264
rect 39560 37200 39576 37264
rect 39640 37200 39656 37264
rect 39720 37200 39736 37264
rect 39800 37200 39816 37264
rect 39880 37200 39896 37264
rect 39960 37200 39976 37264
rect 40040 37200 40056 37264
rect 40120 37200 40136 37264
rect 40200 37200 40216 37264
rect 40280 37200 40296 37264
rect 40360 37200 40368 37264
rect 36368 37184 40368 37200
rect 36368 37120 36376 37184
rect 36440 37120 36456 37184
rect 36520 37120 36536 37184
rect 36600 37120 36616 37184
rect 36680 37120 36696 37184
rect 36760 37120 36776 37184
rect 36840 37120 36856 37184
rect 36920 37120 36936 37184
rect 37000 37120 37016 37184
rect 37080 37120 37096 37184
rect 37160 37120 37176 37184
rect 37240 37120 37256 37184
rect 37320 37120 37336 37184
rect 37400 37120 37416 37184
rect 37480 37120 37496 37184
rect 37560 37120 37576 37184
rect 37640 37120 37656 37184
rect 37720 37120 37736 37184
rect 37800 37120 37816 37184
rect 37880 37120 37896 37184
rect 37960 37120 37976 37184
rect 38040 37120 38056 37184
rect 38120 37120 38136 37184
rect 38200 37120 38216 37184
rect 38280 37120 38296 37184
rect 38360 37120 38376 37184
rect 38440 37120 38456 37184
rect 38520 37120 38536 37184
rect 38600 37120 38616 37184
rect 38680 37120 38696 37184
rect 38760 37120 38776 37184
rect 38840 37120 38856 37184
rect 38920 37120 38936 37184
rect 39000 37120 39016 37184
rect 39080 37120 39096 37184
rect 39160 37120 39176 37184
rect 39240 37120 39256 37184
rect 39320 37120 39336 37184
rect 39400 37120 39416 37184
rect 39480 37120 39496 37184
rect 39560 37120 39576 37184
rect 39640 37120 39656 37184
rect 39720 37120 39736 37184
rect 39800 37120 39816 37184
rect 39880 37120 39896 37184
rect 39960 37120 39976 37184
rect 40040 37120 40056 37184
rect 40120 37120 40136 37184
rect 40200 37120 40216 37184
rect 40280 37120 40296 37184
rect 40360 37120 40368 37184
rect 36368 37104 40368 37120
rect 36368 37040 36376 37104
rect 36440 37040 36456 37104
rect 36520 37040 36536 37104
rect 36600 37040 36616 37104
rect 36680 37040 36696 37104
rect 36760 37040 36776 37104
rect 36840 37040 36856 37104
rect 36920 37040 36936 37104
rect 37000 37040 37016 37104
rect 37080 37040 37096 37104
rect 37160 37040 37176 37104
rect 37240 37040 37256 37104
rect 37320 37040 37336 37104
rect 37400 37040 37416 37104
rect 37480 37040 37496 37104
rect 37560 37040 37576 37104
rect 37640 37040 37656 37104
rect 37720 37040 37736 37104
rect 37800 37040 37816 37104
rect 37880 37040 37896 37104
rect 37960 37040 37976 37104
rect 38040 37040 38056 37104
rect 38120 37040 38136 37104
rect 38200 37040 38216 37104
rect 38280 37040 38296 37104
rect 38360 37040 38376 37104
rect 38440 37040 38456 37104
rect 38520 37040 38536 37104
rect 38600 37040 38616 37104
rect 38680 37040 38696 37104
rect 38760 37040 38776 37104
rect 38840 37040 38856 37104
rect 38920 37040 38936 37104
rect 39000 37040 39016 37104
rect 39080 37040 39096 37104
rect 39160 37040 39176 37104
rect 39240 37040 39256 37104
rect 39320 37040 39336 37104
rect 39400 37040 39416 37104
rect 39480 37040 39496 37104
rect 39560 37040 39576 37104
rect 39640 37040 39656 37104
rect 39720 37040 39736 37104
rect 39800 37040 39816 37104
rect 39880 37040 39896 37104
rect 39960 37040 39976 37104
rect 40040 37040 40056 37104
rect 40120 37040 40136 37104
rect 40200 37040 40216 37104
rect 40280 37040 40296 37104
rect 40360 37040 40368 37104
rect 36368 37024 40368 37040
rect 36368 36960 36376 37024
rect 36440 36960 36456 37024
rect 36520 36960 36536 37024
rect 36600 36960 36616 37024
rect 36680 36960 36696 37024
rect 36760 36960 36776 37024
rect 36840 36960 36856 37024
rect 36920 36960 36936 37024
rect 37000 36960 37016 37024
rect 37080 36960 37096 37024
rect 37160 36960 37176 37024
rect 37240 36960 37256 37024
rect 37320 36960 37336 37024
rect 37400 36960 37416 37024
rect 37480 36960 37496 37024
rect 37560 36960 37576 37024
rect 37640 36960 37656 37024
rect 37720 36960 37736 37024
rect 37800 36960 37816 37024
rect 37880 36960 37896 37024
rect 37960 36960 37976 37024
rect 38040 36960 38056 37024
rect 38120 36960 38136 37024
rect 38200 36960 38216 37024
rect 38280 36960 38296 37024
rect 38360 36960 38376 37024
rect 38440 36960 38456 37024
rect 38520 36960 38536 37024
rect 38600 36960 38616 37024
rect 38680 36960 38696 37024
rect 38760 36960 38776 37024
rect 38840 36960 38856 37024
rect 38920 36960 38936 37024
rect 39000 36960 39016 37024
rect 39080 36960 39096 37024
rect 39160 36960 39176 37024
rect 39240 36960 39256 37024
rect 39320 36960 39336 37024
rect 39400 36960 39416 37024
rect 39480 36960 39496 37024
rect 39560 36960 39576 37024
rect 39640 36960 39656 37024
rect 39720 36960 39736 37024
rect 39800 36960 39816 37024
rect 39880 36960 39896 37024
rect 39960 36960 39976 37024
rect 40040 36960 40056 37024
rect 40120 36960 40136 37024
rect 40200 36960 40216 37024
rect 40280 36960 40296 37024
rect 40360 36960 40368 37024
rect 36368 36944 40368 36960
rect 36368 36880 36376 36944
rect 36440 36880 36456 36944
rect 36520 36880 36536 36944
rect 36600 36880 36616 36944
rect 36680 36880 36696 36944
rect 36760 36880 36776 36944
rect 36840 36880 36856 36944
rect 36920 36880 36936 36944
rect 37000 36880 37016 36944
rect 37080 36880 37096 36944
rect 37160 36880 37176 36944
rect 37240 36880 37256 36944
rect 37320 36880 37336 36944
rect 37400 36880 37416 36944
rect 37480 36880 37496 36944
rect 37560 36880 37576 36944
rect 37640 36880 37656 36944
rect 37720 36880 37736 36944
rect 37800 36880 37816 36944
rect 37880 36880 37896 36944
rect 37960 36880 37976 36944
rect 38040 36880 38056 36944
rect 38120 36880 38136 36944
rect 38200 36880 38216 36944
rect 38280 36880 38296 36944
rect 38360 36880 38376 36944
rect 38440 36880 38456 36944
rect 38520 36880 38536 36944
rect 38600 36880 38616 36944
rect 38680 36880 38696 36944
rect 38760 36880 38776 36944
rect 38840 36880 38856 36944
rect 38920 36880 38936 36944
rect 39000 36880 39016 36944
rect 39080 36880 39096 36944
rect 39160 36880 39176 36944
rect 39240 36880 39256 36944
rect 39320 36880 39336 36944
rect 39400 36880 39416 36944
rect 39480 36880 39496 36944
rect 39560 36880 39576 36944
rect 39640 36880 39656 36944
rect 39720 36880 39736 36944
rect 39800 36880 39816 36944
rect 39880 36880 39896 36944
rect 39960 36880 39976 36944
rect 40040 36880 40056 36944
rect 40120 36880 40136 36944
rect 40200 36880 40216 36944
rect 40280 36880 40296 36944
rect 40360 36880 40368 36944
rect 36368 36864 40368 36880
rect 36368 36800 36376 36864
rect 36440 36800 36456 36864
rect 36520 36800 36536 36864
rect 36600 36800 36616 36864
rect 36680 36800 36696 36864
rect 36760 36800 36776 36864
rect 36840 36800 36856 36864
rect 36920 36800 36936 36864
rect 37000 36800 37016 36864
rect 37080 36800 37096 36864
rect 37160 36800 37176 36864
rect 37240 36800 37256 36864
rect 37320 36800 37336 36864
rect 37400 36800 37416 36864
rect 37480 36800 37496 36864
rect 37560 36800 37576 36864
rect 37640 36800 37656 36864
rect 37720 36800 37736 36864
rect 37800 36800 37816 36864
rect 37880 36800 37896 36864
rect 37960 36800 37976 36864
rect 38040 36800 38056 36864
rect 38120 36800 38136 36864
rect 38200 36800 38216 36864
rect 38280 36800 38296 36864
rect 38360 36800 38376 36864
rect 38440 36800 38456 36864
rect 38520 36800 38536 36864
rect 38600 36800 38616 36864
rect 38680 36800 38696 36864
rect 38760 36800 38776 36864
rect 38840 36800 38856 36864
rect 38920 36800 38936 36864
rect 39000 36800 39016 36864
rect 39080 36800 39096 36864
rect 39160 36800 39176 36864
rect 39240 36800 39256 36864
rect 39320 36800 39336 36864
rect 39400 36800 39416 36864
rect 39480 36800 39496 36864
rect 39560 36800 39576 36864
rect 39640 36800 39656 36864
rect 39720 36800 39736 36864
rect 39800 36800 39816 36864
rect 39880 36800 39896 36864
rect 39960 36800 39976 36864
rect 40040 36800 40056 36864
rect 40120 36800 40136 36864
rect 40200 36800 40216 36864
rect 40280 36800 40296 36864
rect 40360 36800 40368 36864
rect 36368 36784 40368 36800
rect 36368 36720 36376 36784
rect 36440 36720 36456 36784
rect 36520 36720 36536 36784
rect 36600 36720 36616 36784
rect 36680 36720 36696 36784
rect 36760 36720 36776 36784
rect 36840 36720 36856 36784
rect 36920 36720 36936 36784
rect 37000 36720 37016 36784
rect 37080 36720 37096 36784
rect 37160 36720 37176 36784
rect 37240 36720 37256 36784
rect 37320 36720 37336 36784
rect 37400 36720 37416 36784
rect 37480 36720 37496 36784
rect 37560 36720 37576 36784
rect 37640 36720 37656 36784
rect 37720 36720 37736 36784
rect 37800 36720 37816 36784
rect 37880 36720 37896 36784
rect 37960 36720 37976 36784
rect 38040 36720 38056 36784
rect 38120 36720 38136 36784
rect 38200 36720 38216 36784
rect 38280 36720 38296 36784
rect 38360 36720 38376 36784
rect 38440 36720 38456 36784
rect 38520 36720 38536 36784
rect 38600 36720 38616 36784
rect 38680 36720 38696 36784
rect 38760 36720 38776 36784
rect 38840 36720 38856 36784
rect 38920 36720 38936 36784
rect 39000 36720 39016 36784
rect 39080 36720 39096 36784
rect 39160 36720 39176 36784
rect 39240 36720 39256 36784
rect 39320 36720 39336 36784
rect 39400 36720 39416 36784
rect 39480 36720 39496 36784
rect 39560 36720 39576 36784
rect 39640 36720 39656 36784
rect 39720 36720 39736 36784
rect 39800 36720 39816 36784
rect 39880 36720 39896 36784
rect 39960 36720 39976 36784
rect 40040 36720 40056 36784
rect 40120 36720 40136 36784
rect 40200 36720 40216 36784
rect 40280 36720 40296 36784
rect 40360 36720 40368 36784
rect 36368 36704 40368 36720
rect 36368 36640 36376 36704
rect 36440 36640 36456 36704
rect 36520 36640 36536 36704
rect 36600 36640 36616 36704
rect 36680 36640 36696 36704
rect 36760 36640 36776 36704
rect 36840 36640 36856 36704
rect 36920 36640 36936 36704
rect 37000 36640 37016 36704
rect 37080 36640 37096 36704
rect 37160 36640 37176 36704
rect 37240 36640 37256 36704
rect 37320 36640 37336 36704
rect 37400 36640 37416 36704
rect 37480 36640 37496 36704
rect 37560 36640 37576 36704
rect 37640 36640 37656 36704
rect 37720 36640 37736 36704
rect 37800 36640 37816 36704
rect 37880 36640 37896 36704
rect 37960 36640 37976 36704
rect 38040 36640 38056 36704
rect 38120 36640 38136 36704
rect 38200 36640 38216 36704
rect 38280 36640 38296 36704
rect 38360 36640 38376 36704
rect 38440 36640 38456 36704
rect 38520 36640 38536 36704
rect 38600 36640 38616 36704
rect 38680 36640 38696 36704
rect 38760 36640 38776 36704
rect 38840 36640 38856 36704
rect 38920 36640 38936 36704
rect 39000 36640 39016 36704
rect 39080 36640 39096 36704
rect 39160 36640 39176 36704
rect 39240 36640 39256 36704
rect 39320 36640 39336 36704
rect 39400 36640 39416 36704
rect 39480 36640 39496 36704
rect 39560 36640 39576 36704
rect 39640 36640 39656 36704
rect 39720 36640 39736 36704
rect 39800 36640 39816 36704
rect 39880 36640 39896 36704
rect 39960 36640 39976 36704
rect 40040 36640 40056 36704
rect 40120 36640 40136 36704
rect 40200 36640 40216 36704
rect 40280 36640 40296 36704
rect 40360 36640 40368 36704
rect 36368 36624 40368 36640
rect 36368 36560 36376 36624
rect 36440 36560 36456 36624
rect 36520 36560 36536 36624
rect 36600 36560 36616 36624
rect 36680 36560 36696 36624
rect 36760 36560 36776 36624
rect 36840 36560 36856 36624
rect 36920 36560 36936 36624
rect 37000 36560 37016 36624
rect 37080 36560 37096 36624
rect 37160 36560 37176 36624
rect 37240 36560 37256 36624
rect 37320 36560 37336 36624
rect 37400 36560 37416 36624
rect 37480 36560 37496 36624
rect 37560 36560 37576 36624
rect 37640 36560 37656 36624
rect 37720 36560 37736 36624
rect 37800 36560 37816 36624
rect 37880 36560 37896 36624
rect 37960 36560 37976 36624
rect 38040 36560 38056 36624
rect 38120 36560 38136 36624
rect 38200 36560 38216 36624
rect 38280 36560 38296 36624
rect 38360 36560 38376 36624
rect 38440 36560 38456 36624
rect 38520 36560 38536 36624
rect 38600 36560 38616 36624
rect 38680 36560 38696 36624
rect 38760 36560 38776 36624
rect 38840 36560 38856 36624
rect 38920 36560 38936 36624
rect 39000 36560 39016 36624
rect 39080 36560 39096 36624
rect 39160 36560 39176 36624
rect 39240 36560 39256 36624
rect 39320 36560 39336 36624
rect 39400 36560 39416 36624
rect 39480 36560 39496 36624
rect 39560 36560 39576 36624
rect 39640 36560 39656 36624
rect 39720 36560 39736 36624
rect 39800 36560 39816 36624
rect 39880 36560 39896 36624
rect 39960 36560 39976 36624
rect 40040 36560 40056 36624
rect 40120 36560 40136 36624
rect 40200 36560 40216 36624
rect 40280 36560 40296 36624
rect 40360 36560 40368 36624
rect 36368 36544 40368 36560
rect 36368 36480 36376 36544
rect 36440 36480 36456 36544
rect 36520 36480 36536 36544
rect 36600 36480 36616 36544
rect 36680 36480 36696 36544
rect 36760 36480 36776 36544
rect 36840 36480 36856 36544
rect 36920 36480 36936 36544
rect 37000 36480 37016 36544
rect 37080 36480 37096 36544
rect 37160 36480 37176 36544
rect 37240 36480 37256 36544
rect 37320 36480 37336 36544
rect 37400 36480 37416 36544
rect 37480 36480 37496 36544
rect 37560 36480 37576 36544
rect 37640 36480 37656 36544
rect 37720 36480 37736 36544
rect 37800 36480 37816 36544
rect 37880 36480 37896 36544
rect 37960 36480 37976 36544
rect 38040 36480 38056 36544
rect 38120 36480 38136 36544
rect 38200 36480 38216 36544
rect 38280 36480 38296 36544
rect 38360 36480 38376 36544
rect 38440 36480 38456 36544
rect 38520 36480 38536 36544
rect 38600 36480 38616 36544
rect 38680 36480 38696 36544
rect 38760 36480 38776 36544
rect 38840 36480 38856 36544
rect 38920 36480 38936 36544
rect 39000 36480 39016 36544
rect 39080 36480 39096 36544
rect 39160 36480 39176 36544
rect 39240 36480 39256 36544
rect 39320 36480 39336 36544
rect 39400 36480 39416 36544
rect 39480 36480 39496 36544
rect 39560 36480 39576 36544
rect 39640 36480 39656 36544
rect 39720 36480 39736 36544
rect 39800 36480 39816 36544
rect 39880 36480 39896 36544
rect 39960 36480 39976 36544
rect 40040 36480 40056 36544
rect 40120 36480 40136 36544
rect 40200 36480 40216 36544
rect 40280 36480 40296 36544
rect 40360 36480 40368 36544
rect 36368 36464 40368 36480
rect 36368 36400 36376 36464
rect 36440 36400 36456 36464
rect 36520 36400 36536 36464
rect 36600 36400 36616 36464
rect 36680 36400 36696 36464
rect 36760 36400 36776 36464
rect 36840 36400 36856 36464
rect 36920 36400 36936 36464
rect 37000 36400 37016 36464
rect 37080 36400 37096 36464
rect 37160 36400 37176 36464
rect 37240 36400 37256 36464
rect 37320 36400 37336 36464
rect 37400 36400 37416 36464
rect 37480 36400 37496 36464
rect 37560 36400 37576 36464
rect 37640 36400 37656 36464
rect 37720 36400 37736 36464
rect 37800 36400 37816 36464
rect 37880 36400 37896 36464
rect 37960 36400 37976 36464
rect 38040 36400 38056 36464
rect 38120 36400 38136 36464
rect 38200 36400 38216 36464
rect 38280 36400 38296 36464
rect 38360 36400 38376 36464
rect 38440 36400 38456 36464
rect 38520 36400 38536 36464
rect 38600 36400 38616 36464
rect 38680 36400 38696 36464
rect 38760 36400 38776 36464
rect 38840 36400 38856 36464
rect 38920 36400 38936 36464
rect 39000 36400 39016 36464
rect 39080 36400 39096 36464
rect 39160 36400 39176 36464
rect 39240 36400 39256 36464
rect 39320 36400 39336 36464
rect 39400 36400 39416 36464
rect 39480 36400 39496 36464
rect 39560 36400 39576 36464
rect 39640 36400 39656 36464
rect 39720 36400 39736 36464
rect 39800 36400 39816 36464
rect 39880 36400 39896 36464
rect 39960 36400 39976 36464
rect 40040 36400 40056 36464
rect 40120 36400 40136 36464
rect 40200 36400 40216 36464
rect 40280 36400 40296 36464
rect 40360 36400 40368 36464
rect 36368 8992 40368 36400
rect 36368 8928 36376 8992
rect 36440 8928 36456 8992
rect 36520 8928 36536 8992
rect 36600 8928 36616 8992
rect 36680 8928 36696 8992
rect 36760 8928 36776 8992
rect 36840 8928 36856 8992
rect 36920 8928 36936 8992
rect 37000 8928 37016 8992
rect 37080 8928 37096 8992
rect 37160 8928 37176 8992
rect 37240 8928 37256 8992
rect 37320 8928 37336 8992
rect 37400 8928 37416 8992
rect 37480 8928 37496 8992
rect 37560 8928 37576 8992
rect 37640 8928 37656 8992
rect 37720 8928 37736 8992
rect 37800 8928 37816 8992
rect 37880 8928 37896 8992
rect 37960 8928 37976 8992
rect 38040 8928 38056 8992
rect 38120 8928 38136 8992
rect 38200 8928 38216 8992
rect 38280 8928 38296 8992
rect 38360 8928 38376 8992
rect 38440 8928 38456 8992
rect 38520 8928 38536 8992
rect 38600 8928 38616 8992
rect 38680 8928 38696 8992
rect 38760 8928 38776 8992
rect 38840 8928 38856 8992
rect 38920 8928 38936 8992
rect 39000 8928 39016 8992
rect 39080 8928 39096 8992
rect 39160 8928 39176 8992
rect 39240 8928 39256 8992
rect 39320 8928 39336 8992
rect 39400 8928 39416 8992
rect 39480 8928 39496 8992
rect 39560 8928 39576 8992
rect 39640 8928 39656 8992
rect 39720 8928 39736 8992
rect 39800 8928 39816 8992
rect 39880 8928 39896 8992
rect 39960 8928 39976 8992
rect 40040 8928 40056 8992
rect 40120 8928 40136 8992
rect 40200 8928 40216 8992
rect 40280 8928 40296 8992
rect 40360 8928 40368 8992
rect 36368 8912 40368 8928
rect 36368 8848 36376 8912
rect 36440 8848 36456 8912
rect 36520 8848 36536 8912
rect 36600 8848 36616 8912
rect 36680 8848 36696 8912
rect 36760 8848 36776 8912
rect 36840 8848 36856 8912
rect 36920 8848 36936 8912
rect 37000 8848 37016 8912
rect 37080 8848 37096 8912
rect 37160 8848 37176 8912
rect 37240 8848 37256 8912
rect 37320 8848 37336 8912
rect 37400 8848 37416 8912
rect 37480 8848 37496 8912
rect 37560 8848 37576 8912
rect 37640 8848 37656 8912
rect 37720 8848 37736 8912
rect 37800 8848 37816 8912
rect 37880 8848 37896 8912
rect 37960 8848 37976 8912
rect 38040 8848 38056 8912
rect 38120 8848 38136 8912
rect 38200 8848 38216 8912
rect 38280 8848 38296 8912
rect 38360 8848 38376 8912
rect 38440 8848 38456 8912
rect 38520 8848 38536 8912
rect 38600 8848 38616 8912
rect 38680 8848 38696 8912
rect 38760 8848 38776 8912
rect 38840 8848 38856 8912
rect 38920 8848 38936 8912
rect 39000 8848 39016 8912
rect 39080 8848 39096 8912
rect 39160 8848 39176 8912
rect 39240 8848 39256 8912
rect 39320 8848 39336 8912
rect 39400 8848 39416 8912
rect 39480 8848 39496 8912
rect 39560 8848 39576 8912
rect 39640 8848 39656 8912
rect 39720 8848 39736 8912
rect 39800 8848 39816 8912
rect 39880 8848 39896 8912
rect 39960 8848 39976 8912
rect 40040 8848 40056 8912
rect 40120 8848 40136 8912
rect 40200 8848 40216 8912
rect 40280 8848 40296 8912
rect 40360 8848 40368 8912
rect 36368 8832 40368 8848
rect 36368 8768 36376 8832
rect 36440 8768 36456 8832
rect 36520 8768 36536 8832
rect 36600 8768 36616 8832
rect 36680 8768 36696 8832
rect 36760 8768 36776 8832
rect 36840 8768 36856 8832
rect 36920 8768 36936 8832
rect 37000 8768 37016 8832
rect 37080 8768 37096 8832
rect 37160 8768 37176 8832
rect 37240 8768 37256 8832
rect 37320 8768 37336 8832
rect 37400 8768 37416 8832
rect 37480 8768 37496 8832
rect 37560 8768 37576 8832
rect 37640 8768 37656 8832
rect 37720 8768 37736 8832
rect 37800 8768 37816 8832
rect 37880 8768 37896 8832
rect 37960 8768 37976 8832
rect 38040 8768 38056 8832
rect 38120 8768 38136 8832
rect 38200 8768 38216 8832
rect 38280 8768 38296 8832
rect 38360 8768 38376 8832
rect 38440 8768 38456 8832
rect 38520 8768 38536 8832
rect 38600 8768 38616 8832
rect 38680 8768 38696 8832
rect 38760 8768 38776 8832
rect 38840 8768 38856 8832
rect 38920 8768 38936 8832
rect 39000 8768 39016 8832
rect 39080 8768 39096 8832
rect 39160 8768 39176 8832
rect 39240 8768 39256 8832
rect 39320 8768 39336 8832
rect 39400 8768 39416 8832
rect 39480 8768 39496 8832
rect 39560 8768 39576 8832
rect 39640 8768 39656 8832
rect 39720 8768 39736 8832
rect 39800 8768 39816 8832
rect 39880 8768 39896 8832
rect 39960 8768 39976 8832
rect 40040 8768 40056 8832
rect 40120 8768 40136 8832
rect 40200 8768 40216 8832
rect 40280 8768 40296 8832
rect 40360 8768 40368 8832
rect 36368 8752 40368 8768
rect 36368 8688 36376 8752
rect 36440 8688 36456 8752
rect 36520 8688 36536 8752
rect 36600 8688 36616 8752
rect 36680 8688 36696 8752
rect 36760 8688 36776 8752
rect 36840 8688 36856 8752
rect 36920 8688 36936 8752
rect 37000 8688 37016 8752
rect 37080 8688 37096 8752
rect 37160 8688 37176 8752
rect 37240 8688 37256 8752
rect 37320 8688 37336 8752
rect 37400 8688 37416 8752
rect 37480 8688 37496 8752
rect 37560 8688 37576 8752
rect 37640 8688 37656 8752
rect 37720 8688 37736 8752
rect 37800 8688 37816 8752
rect 37880 8688 37896 8752
rect 37960 8688 37976 8752
rect 38040 8688 38056 8752
rect 38120 8688 38136 8752
rect 38200 8688 38216 8752
rect 38280 8688 38296 8752
rect 38360 8688 38376 8752
rect 38440 8688 38456 8752
rect 38520 8688 38536 8752
rect 38600 8688 38616 8752
rect 38680 8688 38696 8752
rect 38760 8688 38776 8752
rect 38840 8688 38856 8752
rect 38920 8688 38936 8752
rect 39000 8688 39016 8752
rect 39080 8688 39096 8752
rect 39160 8688 39176 8752
rect 39240 8688 39256 8752
rect 39320 8688 39336 8752
rect 39400 8688 39416 8752
rect 39480 8688 39496 8752
rect 39560 8688 39576 8752
rect 39640 8688 39656 8752
rect 39720 8688 39736 8752
rect 39800 8688 39816 8752
rect 39880 8688 39896 8752
rect 39960 8688 39976 8752
rect 40040 8688 40056 8752
rect 40120 8688 40136 8752
rect 40200 8688 40216 8752
rect 40280 8688 40296 8752
rect 40360 8688 40368 8752
rect 36368 8672 40368 8688
rect 36368 8608 36376 8672
rect 36440 8608 36456 8672
rect 36520 8608 36536 8672
rect 36600 8608 36616 8672
rect 36680 8608 36696 8672
rect 36760 8608 36776 8672
rect 36840 8608 36856 8672
rect 36920 8608 36936 8672
rect 37000 8608 37016 8672
rect 37080 8608 37096 8672
rect 37160 8608 37176 8672
rect 37240 8608 37256 8672
rect 37320 8608 37336 8672
rect 37400 8608 37416 8672
rect 37480 8608 37496 8672
rect 37560 8608 37576 8672
rect 37640 8608 37656 8672
rect 37720 8608 37736 8672
rect 37800 8608 37816 8672
rect 37880 8608 37896 8672
rect 37960 8608 37976 8672
rect 38040 8608 38056 8672
rect 38120 8608 38136 8672
rect 38200 8608 38216 8672
rect 38280 8608 38296 8672
rect 38360 8608 38376 8672
rect 38440 8608 38456 8672
rect 38520 8608 38536 8672
rect 38600 8608 38616 8672
rect 38680 8608 38696 8672
rect 38760 8608 38776 8672
rect 38840 8608 38856 8672
rect 38920 8608 38936 8672
rect 39000 8608 39016 8672
rect 39080 8608 39096 8672
rect 39160 8608 39176 8672
rect 39240 8608 39256 8672
rect 39320 8608 39336 8672
rect 39400 8608 39416 8672
rect 39480 8608 39496 8672
rect 39560 8608 39576 8672
rect 39640 8608 39656 8672
rect 39720 8608 39736 8672
rect 39800 8608 39816 8672
rect 39880 8608 39896 8672
rect 39960 8608 39976 8672
rect 40040 8608 40056 8672
rect 40120 8608 40136 8672
rect 40200 8608 40216 8672
rect 40280 8608 40296 8672
rect 40360 8608 40368 8672
rect 36368 8592 40368 8608
rect 36368 8528 36376 8592
rect 36440 8528 36456 8592
rect 36520 8528 36536 8592
rect 36600 8528 36616 8592
rect 36680 8528 36696 8592
rect 36760 8528 36776 8592
rect 36840 8528 36856 8592
rect 36920 8528 36936 8592
rect 37000 8528 37016 8592
rect 37080 8528 37096 8592
rect 37160 8528 37176 8592
rect 37240 8528 37256 8592
rect 37320 8528 37336 8592
rect 37400 8528 37416 8592
rect 37480 8528 37496 8592
rect 37560 8528 37576 8592
rect 37640 8528 37656 8592
rect 37720 8528 37736 8592
rect 37800 8528 37816 8592
rect 37880 8528 37896 8592
rect 37960 8528 37976 8592
rect 38040 8528 38056 8592
rect 38120 8528 38136 8592
rect 38200 8528 38216 8592
rect 38280 8528 38296 8592
rect 38360 8528 38376 8592
rect 38440 8528 38456 8592
rect 38520 8528 38536 8592
rect 38600 8528 38616 8592
rect 38680 8528 38696 8592
rect 38760 8528 38776 8592
rect 38840 8528 38856 8592
rect 38920 8528 38936 8592
rect 39000 8528 39016 8592
rect 39080 8528 39096 8592
rect 39160 8528 39176 8592
rect 39240 8528 39256 8592
rect 39320 8528 39336 8592
rect 39400 8528 39416 8592
rect 39480 8528 39496 8592
rect 39560 8528 39576 8592
rect 39640 8528 39656 8592
rect 39720 8528 39736 8592
rect 39800 8528 39816 8592
rect 39880 8528 39896 8592
rect 39960 8528 39976 8592
rect 40040 8528 40056 8592
rect 40120 8528 40136 8592
rect 40200 8528 40216 8592
rect 40280 8528 40296 8592
rect 40360 8528 40368 8592
rect 36368 8512 40368 8528
rect 36368 8448 36376 8512
rect 36440 8448 36456 8512
rect 36520 8448 36536 8512
rect 36600 8448 36616 8512
rect 36680 8448 36696 8512
rect 36760 8448 36776 8512
rect 36840 8448 36856 8512
rect 36920 8448 36936 8512
rect 37000 8448 37016 8512
rect 37080 8448 37096 8512
rect 37160 8448 37176 8512
rect 37240 8448 37256 8512
rect 37320 8448 37336 8512
rect 37400 8448 37416 8512
rect 37480 8448 37496 8512
rect 37560 8448 37576 8512
rect 37640 8448 37656 8512
rect 37720 8448 37736 8512
rect 37800 8448 37816 8512
rect 37880 8448 37896 8512
rect 37960 8448 37976 8512
rect 38040 8448 38056 8512
rect 38120 8448 38136 8512
rect 38200 8448 38216 8512
rect 38280 8448 38296 8512
rect 38360 8448 38376 8512
rect 38440 8448 38456 8512
rect 38520 8448 38536 8512
rect 38600 8448 38616 8512
rect 38680 8448 38696 8512
rect 38760 8448 38776 8512
rect 38840 8448 38856 8512
rect 38920 8448 38936 8512
rect 39000 8448 39016 8512
rect 39080 8448 39096 8512
rect 39160 8448 39176 8512
rect 39240 8448 39256 8512
rect 39320 8448 39336 8512
rect 39400 8448 39416 8512
rect 39480 8448 39496 8512
rect 39560 8448 39576 8512
rect 39640 8448 39656 8512
rect 39720 8448 39736 8512
rect 39800 8448 39816 8512
rect 39880 8448 39896 8512
rect 39960 8448 39976 8512
rect 40040 8448 40056 8512
rect 40120 8448 40136 8512
rect 40200 8448 40216 8512
rect 40280 8448 40296 8512
rect 40360 8448 40368 8512
rect 36368 8432 40368 8448
rect 36368 8368 36376 8432
rect 36440 8368 36456 8432
rect 36520 8368 36536 8432
rect 36600 8368 36616 8432
rect 36680 8368 36696 8432
rect 36760 8368 36776 8432
rect 36840 8368 36856 8432
rect 36920 8368 36936 8432
rect 37000 8368 37016 8432
rect 37080 8368 37096 8432
rect 37160 8368 37176 8432
rect 37240 8368 37256 8432
rect 37320 8368 37336 8432
rect 37400 8368 37416 8432
rect 37480 8368 37496 8432
rect 37560 8368 37576 8432
rect 37640 8368 37656 8432
rect 37720 8368 37736 8432
rect 37800 8368 37816 8432
rect 37880 8368 37896 8432
rect 37960 8368 37976 8432
rect 38040 8368 38056 8432
rect 38120 8368 38136 8432
rect 38200 8368 38216 8432
rect 38280 8368 38296 8432
rect 38360 8368 38376 8432
rect 38440 8368 38456 8432
rect 38520 8368 38536 8432
rect 38600 8368 38616 8432
rect 38680 8368 38696 8432
rect 38760 8368 38776 8432
rect 38840 8368 38856 8432
rect 38920 8368 38936 8432
rect 39000 8368 39016 8432
rect 39080 8368 39096 8432
rect 39160 8368 39176 8432
rect 39240 8368 39256 8432
rect 39320 8368 39336 8432
rect 39400 8368 39416 8432
rect 39480 8368 39496 8432
rect 39560 8368 39576 8432
rect 39640 8368 39656 8432
rect 39720 8368 39736 8432
rect 39800 8368 39816 8432
rect 39880 8368 39896 8432
rect 39960 8368 39976 8432
rect 40040 8368 40056 8432
rect 40120 8368 40136 8432
rect 40200 8368 40216 8432
rect 40280 8368 40296 8432
rect 40360 8368 40368 8432
rect 36368 8352 40368 8368
rect 36368 8288 36376 8352
rect 36440 8288 36456 8352
rect 36520 8288 36536 8352
rect 36600 8288 36616 8352
rect 36680 8288 36696 8352
rect 36760 8288 36776 8352
rect 36840 8288 36856 8352
rect 36920 8288 36936 8352
rect 37000 8288 37016 8352
rect 37080 8288 37096 8352
rect 37160 8288 37176 8352
rect 37240 8288 37256 8352
rect 37320 8288 37336 8352
rect 37400 8288 37416 8352
rect 37480 8288 37496 8352
rect 37560 8288 37576 8352
rect 37640 8288 37656 8352
rect 37720 8288 37736 8352
rect 37800 8288 37816 8352
rect 37880 8288 37896 8352
rect 37960 8288 37976 8352
rect 38040 8288 38056 8352
rect 38120 8288 38136 8352
rect 38200 8288 38216 8352
rect 38280 8288 38296 8352
rect 38360 8288 38376 8352
rect 38440 8288 38456 8352
rect 38520 8288 38536 8352
rect 38600 8288 38616 8352
rect 38680 8288 38696 8352
rect 38760 8288 38776 8352
rect 38840 8288 38856 8352
rect 38920 8288 38936 8352
rect 39000 8288 39016 8352
rect 39080 8288 39096 8352
rect 39160 8288 39176 8352
rect 39240 8288 39256 8352
rect 39320 8288 39336 8352
rect 39400 8288 39416 8352
rect 39480 8288 39496 8352
rect 39560 8288 39576 8352
rect 39640 8288 39656 8352
rect 39720 8288 39736 8352
rect 39800 8288 39816 8352
rect 39880 8288 39896 8352
rect 39960 8288 39976 8352
rect 40040 8288 40056 8352
rect 40120 8288 40136 8352
rect 40200 8288 40216 8352
rect 40280 8288 40296 8352
rect 40360 8288 40368 8352
rect 36368 8272 40368 8288
rect 36368 8208 36376 8272
rect 36440 8208 36456 8272
rect 36520 8208 36536 8272
rect 36600 8208 36616 8272
rect 36680 8208 36696 8272
rect 36760 8208 36776 8272
rect 36840 8208 36856 8272
rect 36920 8208 36936 8272
rect 37000 8208 37016 8272
rect 37080 8208 37096 8272
rect 37160 8208 37176 8272
rect 37240 8208 37256 8272
rect 37320 8208 37336 8272
rect 37400 8208 37416 8272
rect 37480 8208 37496 8272
rect 37560 8208 37576 8272
rect 37640 8208 37656 8272
rect 37720 8208 37736 8272
rect 37800 8208 37816 8272
rect 37880 8208 37896 8272
rect 37960 8208 37976 8272
rect 38040 8208 38056 8272
rect 38120 8208 38136 8272
rect 38200 8208 38216 8272
rect 38280 8208 38296 8272
rect 38360 8208 38376 8272
rect 38440 8208 38456 8272
rect 38520 8208 38536 8272
rect 38600 8208 38616 8272
rect 38680 8208 38696 8272
rect 38760 8208 38776 8272
rect 38840 8208 38856 8272
rect 38920 8208 38936 8272
rect 39000 8208 39016 8272
rect 39080 8208 39096 8272
rect 39160 8208 39176 8272
rect 39240 8208 39256 8272
rect 39320 8208 39336 8272
rect 39400 8208 39416 8272
rect 39480 8208 39496 8272
rect 39560 8208 39576 8272
rect 39640 8208 39656 8272
rect 39720 8208 39736 8272
rect 39800 8208 39816 8272
rect 39880 8208 39896 8272
rect 39960 8208 39976 8272
rect 40040 8208 40056 8272
rect 40120 8208 40136 8272
rect 40200 8208 40216 8272
rect 40280 8208 40296 8272
rect 40360 8208 40368 8272
rect 36368 8192 40368 8208
rect 36368 8128 36376 8192
rect 36440 8128 36456 8192
rect 36520 8128 36536 8192
rect 36600 8128 36616 8192
rect 36680 8128 36696 8192
rect 36760 8128 36776 8192
rect 36840 8128 36856 8192
rect 36920 8128 36936 8192
rect 37000 8128 37016 8192
rect 37080 8128 37096 8192
rect 37160 8128 37176 8192
rect 37240 8128 37256 8192
rect 37320 8128 37336 8192
rect 37400 8128 37416 8192
rect 37480 8128 37496 8192
rect 37560 8128 37576 8192
rect 37640 8128 37656 8192
rect 37720 8128 37736 8192
rect 37800 8128 37816 8192
rect 37880 8128 37896 8192
rect 37960 8128 37976 8192
rect 38040 8128 38056 8192
rect 38120 8128 38136 8192
rect 38200 8128 38216 8192
rect 38280 8128 38296 8192
rect 38360 8128 38376 8192
rect 38440 8128 38456 8192
rect 38520 8128 38536 8192
rect 38600 8128 38616 8192
rect 38680 8128 38696 8192
rect 38760 8128 38776 8192
rect 38840 8128 38856 8192
rect 38920 8128 38936 8192
rect 39000 8128 39016 8192
rect 39080 8128 39096 8192
rect 39160 8128 39176 8192
rect 39240 8128 39256 8192
rect 39320 8128 39336 8192
rect 39400 8128 39416 8192
rect 39480 8128 39496 8192
rect 39560 8128 39576 8192
rect 39640 8128 39656 8192
rect 39720 8128 39736 8192
rect 39800 8128 39816 8192
rect 39880 8128 39896 8192
rect 39960 8128 39976 8192
rect 40040 8128 40056 8192
rect 40120 8128 40136 8192
rect 40200 8128 40216 8192
rect 40280 8128 40296 8192
rect 40360 8128 40368 8192
rect 36368 8112 40368 8128
rect 36368 8048 36376 8112
rect 36440 8048 36456 8112
rect 36520 8048 36536 8112
rect 36600 8048 36616 8112
rect 36680 8048 36696 8112
rect 36760 8048 36776 8112
rect 36840 8048 36856 8112
rect 36920 8048 36936 8112
rect 37000 8048 37016 8112
rect 37080 8048 37096 8112
rect 37160 8048 37176 8112
rect 37240 8048 37256 8112
rect 37320 8048 37336 8112
rect 37400 8048 37416 8112
rect 37480 8048 37496 8112
rect 37560 8048 37576 8112
rect 37640 8048 37656 8112
rect 37720 8048 37736 8112
rect 37800 8048 37816 8112
rect 37880 8048 37896 8112
rect 37960 8048 37976 8112
rect 38040 8048 38056 8112
rect 38120 8048 38136 8112
rect 38200 8048 38216 8112
rect 38280 8048 38296 8112
rect 38360 8048 38376 8112
rect 38440 8048 38456 8112
rect 38520 8048 38536 8112
rect 38600 8048 38616 8112
rect 38680 8048 38696 8112
rect 38760 8048 38776 8112
rect 38840 8048 38856 8112
rect 38920 8048 38936 8112
rect 39000 8048 39016 8112
rect 39080 8048 39096 8112
rect 39160 8048 39176 8112
rect 39240 8048 39256 8112
rect 39320 8048 39336 8112
rect 39400 8048 39416 8112
rect 39480 8048 39496 8112
rect 39560 8048 39576 8112
rect 39640 8048 39656 8112
rect 39720 8048 39736 8112
rect 39800 8048 39816 8112
rect 39880 8048 39896 8112
rect 39960 8048 39976 8112
rect 40040 8048 40056 8112
rect 40120 8048 40136 8112
rect 40200 8048 40216 8112
rect 40280 8048 40296 8112
rect 40360 8048 40368 8112
rect 36368 8032 40368 8048
rect 36368 7968 36376 8032
rect 36440 7968 36456 8032
rect 36520 7968 36536 8032
rect 36600 7968 36616 8032
rect 36680 7968 36696 8032
rect 36760 7968 36776 8032
rect 36840 7968 36856 8032
rect 36920 7968 36936 8032
rect 37000 7968 37016 8032
rect 37080 7968 37096 8032
rect 37160 7968 37176 8032
rect 37240 7968 37256 8032
rect 37320 7968 37336 8032
rect 37400 7968 37416 8032
rect 37480 7968 37496 8032
rect 37560 7968 37576 8032
rect 37640 7968 37656 8032
rect 37720 7968 37736 8032
rect 37800 7968 37816 8032
rect 37880 7968 37896 8032
rect 37960 7968 37976 8032
rect 38040 7968 38056 8032
rect 38120 7968 38136 8032
rect 38200 7968 38216 8032
rect 38280 7968 38296 8032
rect 38360 7968 38376 8032
rect 38440 7968 38456 8032
rect 38520 7968 38536 8032
rect 38600 7968 38616 8032
rect 38680 7968 38696 8032
rect 38760 7968 38776 8032
rect 38840 7968 38856 8032
rect 38920 7968 38936 8032
rect 39000 7968 39016 8032
rect 39080 7968 39096 8032
rect 39160 7968 39176 8032
rect 39240 7968 39256 8032
rect 39320 7968 39336 8032
rect 39400 7968 39416 8032
rect 39480 7968 39496 8032
rect 39560 7968 39576 8032
rect 39640 7968 39656 8032
rect 39720 7968 39736 8032
rect 39800 7968 39816 8032
rect 39880 7968 39896 8032
rect 39960 7968 39976 8032
rect 40040 7968 40056 8032
rect 40120 7968 40136 8032
rect 40200 7968 40216 8032
rect 40280 7968 40296 8032
rect 40360 7968 40368 8032
rect 36368 7952 40368 7968
rect 36368 7888 36376 7952
rect 36440 7888 36456 7952
rect 36520 7888 36536 7952
rect 36600 7888 36616 7952
rect 36680 7888 36696 7952
rect 36760 7888 36776 7952
rect 36840 7888 36856 7952
rect 36920 7888 36936 7952
rect 37000 7888 37016 7952
rect 37080 7888 37096 7952
rect 37160 7888 37176 7952
rect 37240 7888 37256 7952
rect 37320 7888 37336 7952
rect 37400 7888 37416 7952
rect 37480 7888 37496 7952
rect 37560 7888 37576 7952
rect 37640 7888 37656 7952
rect 37720 7888 37736 7952
rect 37800 7888 37816 7952
rect 37880 7888 37896 7952
rect 37960 7888 37976 7952
rect 38040 7888 38056 7952
rect 38120 7888 38136 7952
rect 38200 7888 38216 7952
rect 38280 7888 38296 7952
rect 38360 7888 38376 7952
rect 38440 7888 38456 7952
rect 38520 7888 38536 7952
rect 38600 7888 38616 7952
rect 38680 7888 38696 7952
rect 38760 7888 38776 7952
rect 38840 7888 38856 7952
rect 38920 7888 38936 7952
rect 39000 7888 39016 7952
rect 39080 7888 39096 7952
rect 39160 7888 39176 7952
rect 39240 7888 39256 7952
rect 39320 7888 39336 7952
rect 39400 7888 39416 7952
rect 39480 7888 39496 7952
rect 39560 7888 39576 7952
rect 39640 7888 39656 7952
rect 39720 7888 39736 7952
rect 39800 7888 39816 7952
rect 39880 7888 39896 7952
rect 39960 7888 39976 7952
rect 40040 7888 40056 7952
rect 40120 7888 40136 7952
rect 40200 7888 40216 7952
rect 40280 7888 40296 7952
rect 40360 7888 40368 7952
rect 36368 7872 40368 7888
rect 36368 7808 36376 7872
rect 36440 7808 36456 7872
rect 36520 7808 36536 7872
rect 36600 7808 36616 7872
rect 36680 7808 36696 7872
rect 36760 7808 36776 7872
rect 36840 7808 36856 7872
rect 36920 7808 36936 7872
rect 37000 7808 37016 7872
rect 37080 7808 37096 7872
rect 37160 7808 37176 7872
rect 37240 7808 37256 7872
rect 37320 7808 37336 7872
rect 37400 7808 37416 7872
rect 37480 7808 37496 7872
rect 37560 7808 37576 7872
rect 37640 7808 37656 7872
rect 37720 7808 37736 7872
rect 37800 7808 37816 7872
rect 37880 7808 37896 7872
rect 37960 7808 37976 7872
rect 38040 7808 38056 7872
rect 38120 7808 38136 7872
rect 38200 7808 38216 7872
rect 38280 7808 38296 7872
rect 38360 7808 38376 7872
rect 38440 7808 38456 7872
rect 38520 7808 38536 7872
rect 38600 7808 38616 7872
rect 38680 7808 38696 7872
rect 38760 7808 38776 7872
rect 38840 7808 38856 7872
rect 38920 7808 38936 7872
rect 39000 7808 39016 7872
rect 39080 7808 39096 7872
rect 39160 7808 39176 7872
rect 39240 7808 39256 7872
rect 39320 7808 39336 7872
rect 39400 7808 39416 7872
rect 39480 7808 39496 7872
rect 39560 7808 39576 7872
rect 39640 7808 39656 7872
rect 39720 7808 39736 7872
rect 39800 7808 39816 7872
rect 39880 7808 39896 7872
rect 39960 7808 39976 7872
rect 40040 7808 40056 7872
rect 40120 7808 40136 7872
rect 40200 7808 40216 7872
rect 40280 7808 40296 7872
rect 40360 7808 40368 7872
rect 36368 7792 40368 7808
rect 36368 7728 36376 7792
rect 36440 7728 36456 7792
rect 36520 7728 36536 7792
rect 36600 7728 36616 7792
rect 36680 7728 36696 7792
rect 36760 7728 36776 7792
rect 36840 7728 36856 7792
rect 36920 7728 36936 7792
rect 37000 7728 37016 7792
rect 37080 7728 37096 7792
rect 37160 7728 37176 7792
rect 37240 7728 37256 7792
rect 37320 7728 37336 7792
rect 37400 7728 37416 7792
rect 37480 7728 37496 7792
rect 37560 7728 37576 7792
rect 37640 7728 37656 7792
rect 37720 7728 37736 7792
rect 37800 7728 37816 7792
rect 37880 7728 37896 7792
rect 37960 7728 37976 7792
rect 38040 7728 38056 7792
rect 38120 7728 38136 7792
rect 38200 7728 38216 7792
rect 38280 7728 38296 7792
rect 38360 7728 38376 7792
rect 38440 7728 38456 7792
rect 38520 7728 38536 7792
rect 38600 7728 38616 7792
rect 38680 7728 38696 7792
rect 38760 7728 38776 7792
rect 38840 7728 38856 7792
rect 38920 7728 38936 7792
rect 39000 7728 39016 7792
rect 39080 7728 39096 7792
rect 39160 7728 39176 7792
rect 39240 7728 39256 7792
rect 39320 7728 39336 7792
rect 39400 7728 39416 7792
rect 39480 7728 39496 7792
rect 39560 7728 39576 7792
rect 39640 7728 39656 7792
rect 39720 7728 39736 7792
rect 39800 7728 39816 7792
rect 39880 7728 39896 7792
rect 39960 7728 39976 7792
rect 40040 7728 40056 7792
rect 40120 7728 40136 7792
rect 40200 7728 40216 7792
rect 40280 7728 40296 7792
rect 40360 7728 40368 7792
rect 36368 7712 40368 7728
rect 36368 7648 36376 7712
rect 36440 7648 36456 7712
rect 36520 7648 36536 7712
rect 36600 7648 36616 7712
rect 36680 7648 36696 7712
rect 36760 7648 36776 7712
rect 36840 7648 36856 7712
rect 36920 7648 36936 7712
rect 37000 7648 37016 7712
rect 37080 7648 37096 7712
rect 37160 7648 37176 7712
rect 37240 7648 37256 7712
rect 37320 7648 37336 7712
rect 37400 7648 37416 7712
rect 37480 7648 37496 7712
rect 37560 7648 37576 7712
rect 37640 7648 37656 7712
rect 37720 7648 37736 7712
rect 37800 7648 37816 7712
rect 37880 7648 37896 7712
rect 37960 7648 37976 7712
rect 38040 7648 38056 7712
rect 38120 7648 38136 7712
rect 38200 7648 38216 7712
rect 38280 7648 38296 7712
rect 38360 7648 38376 7712
rect 38440 7648 38456 7712
rect 38520 7648 38536 7712
rect 38600 7648 38616 7712
rect 38680 7648 38696 7712
rect 38760 7648 38776 7712
rect 38840 7648 38856 7712
rect 38920 7648 38936 7712
rect 39000 7648 39016 7712
rect 39080 7648 39096 7712
rect 39160 7648 39176 7712
rect 39240 7648 39256 7712
rect 39320 7648 39336 7712
rect 39400 7648 39416 7712
rect 39480 7648 39496 7712
rect 39560 7648 39576 7712
rect 39640 7648 39656 7712
rect 39720 7648 39736 7712
rect 39800 7648 39816 7712
rect 39880 7648 39896 7712
rect 39960 7648 39976 7712
rect 40040 7648 40056 7712
rect 40120 7648 40136 7712
rect 40200 7648 40216 7712
rect 40280 7648 40296 7712
rect 40360 7648 40368 7712
rect 36368 7632 40368 7648
rect 36368 7568 36376 7632
rect 36440 7568 36456 7632
rect 36520 7568 36536 7632
rect 36600 7568 36616 7632
rect 36680 7568 36696 7632
rect 36760 7568 36776 7632
rect 36840 7568 36856 7632
rect 36920 7568 36936 7632
rect 37000 7568 37016 7632
rect 37080 7568 37096 7632
rect 37160 7568 37176 7632
rect 37240 7568 37256 7632
rect 37320 7568 37336 7632
rect 37400 7568 37416 7632
rect 37480 7568 37496 7632
rect 37560 7568 37576 7632
rect 37640 7568 37656 7632
rect 37720 7568 37736 7632
rect 37800 7568 37816 7632
rect 37880 7568 37896 7632
rect 37960 7568 37976 7632
rect 38040 7568 38056 7632
rect 38120 7568 38136 7632
rect 38200 7568 38216 7632
rect 38280 7568 38296 7632
rect 38360 7568 38376 7632
rect 38440 7568 38456 7632
rect 38520 7568 38536 7632
rect 38600 7568 38616 7632
rect 38680 7568 38696 7632
rect 38760 7568 38776 7632
rect 38840 7568 38856 7632
rect 38920 7568 38936 7632
rect 39000 7568 39016 7632
rect 39080 7568 39096 7632
rect 39160 7568 39176 7632
rect 39240 7568 39256 7632
rect 39320 7568 39336 7632
rect 39400 7568 39416 7632
rect 39480 7568 39496 7632
rect 39560 7568 39576 7632
rect 39640 7568 39656 7632
rect 39720 7568 39736 7632
rect 39800 7568 39816 7632
rect 39880 7568 39896 7632
rect 39960 7568 39976 7632
rect 40040 7568 40056 7632
rect 40120 7568 40136 7632
rect 40200 7568 40216 7632
rect 40280 7568 40296 7632
rect 40360 7568 40368 7632
rect 36368 7552 40368 7568
rect 36368 7488 36376 7552
rect 36440 7488 36456 7552
rect 36520 7488 36536 7552
rect 36600 7488 36616 7552
rect 36680 7488 36696 7552
rect 36760 7488 36776 7552
rect 36840 7488 36856 7552
rect 36920 7488 36936 7552
rect 37000 7488 37016 7552
rect 37080 7488 37096 7552
rect 37160 7488 37176 7552
rect 37240 7488 37256 7552
rect 37320 7488 37336 7552
rect 37400 7488 37416 7552
rect 37480 7488 37496 7552
rect 37560 7488 37576 7552
rect 37640 7488 37656 7552
rect 37720 7488 37736 7552
rect 37800 7488 37816 7552
rect 37880 7488 37896 7552
rect 37960 7488 37976 7552
rect 38040 7488 38056 7552
rect 38120 7488 38136 7552
rect 38200 7488 38216 7552
rect 38280 7488 38296 7552
rect 38360 7488 38376 7552
rect 38440 7488 38456 7552
rect 38520 7488 38536 7552
rect 38600 7488 38616 7552
rect 38680 7488 38696 7552
rect 38760 7488 38776 7552
rect 38840 7488 38856 7552
rect 38920 7488 38936 7552
rect 39000 7488 39016 7552
rect 39080 7488 39096 7552
rect 39160 7488 39176 7552
rect 39240 7488 39256 7552
rect 39320 7488 39336 7552
rect 39400 7488 39416 7552
rect 39480 7488 39496 7552
rect 39560 7488 39576 7552
rect 39640 7488 39656 7552
rect 39720 7488 39736 7552
rect 39800 7488 39816 7552
rect 39880 7488 39896 7552
rect 39960 7488 39976 7552
rect 40040 7488 40056 7552
rect 40120 7488 40136 7552
rect 40200 7488 40216 7552
rect 40280 7488 40296 7552
rect 40360 7488 40368 7552
rect 36368 7472 40368 7488
rect 36368 7408 36376 7472
rect 36440 7408 36456 7472
rect 36520 7408 36536 7472
rect 36600 7408 36616 7472
rect 36680 7408 36696 7472
rect 36760 7408 36776 7472
rect 36840 7408 36856 7472
rect 36920 7408 36936 7472
rect 37000 7408 37016 7472
rect 37080 7408 37096 7472
rect 37160 7408 37176 7472
rect 37240 7408 37256 7472
rect 37320 7408 37336 7472
rect 37400 7408 37416 7472
rect 37480 7408 37496 7472
rect 37560 7408 37576 7472
rect 37640 7408 37656 7472
rect 37720 7408 37736 7472
rect 37800 7408 37816 7472
rect 37880 7408 37896 7472
rect 37960 7408 37976 7472
rect 38040 7408 38056 7472
rect 38120 7408 38136 7472
rect 38200 7408 38216 7472
rect 38280 7408 38296 7472
rect 38360 7408 38376 7472
rect 38440 7408 38456 7472
rect 38520 7408 38536 7472
rect 38600 7408 38616 7472
rect 38680 7408 38696 7472
rect 38760 7408 38776 7472
rect 38840 7408 38856 7472
rect 38920 7408 38936 7472
rect 39000 7408 39016 7472
rect 39080 7408 39096 7472
rect 39160 7408 39176 7472
rect 39240 7408 39256 7472
rect 39320 7408 39336 7472
rect 39400 7408 39416 7472
rect 39480 7408 39496 7472
rect 39560 7408 39576 7472
rect 39640 7408 39656 7472
rect 39720 7408 39736 7472
rect 39800 7408 39816 7472
rect 39880 7408 39896 7472
rect 39960 7408 39976 7472
rect 40040 7408 40056 7472
rect 40120 7408 40136 7472
rect 40200 7408 40216 7472
rect 40280 7408 40296 7472
rect 40360 7408 40368 7472
rect 36368 7392 40368 7408
rect 36368 7328 36376 7392
rect 36440 7328 36456 7392
rect 36520 7328 36536 7392
rect 36600 7328 36616 7392
rect 36680 7328 36696 7392
rect 36760 7328 36776 7392
rect 36840 7328 36856 7392
rect 36920 7328 36936 7392
rect 37000 7328 37016 7392
rect 37080 7328 37096 7392
rect 37160 7328 37176 7392
rect 37240 7328 37256 7392
rect 37320 7328 37336 7392
rect 37400 7328 37416 7392
rect 37480 7328 37496 7392
rect 37560 7328 37576 7392
rect 37640 7328 37656 7392
rect 37720 7328 37736 7392
rect 37800 7328 37816 7392
rect 37880 7328 37896 7392
rect 37960 7328 37976 7392
rect 38040 7328 38056 7392
rect 38120 7328 38136 7392
rect 38200 7328 38216 7392
rect 38280 7328 38296 7392
rect 38360 7328 38376 7392
rect 38440 7328 38456 7392
rect 38520 7328 38536 7392
rect 38600 7328 38616 7392
rect 38680 7328 38696 7392
rect 38760 7328 38776 7392
rect 38840 7328 38856 7392
rect 38920 7328 38936 7392
rect 39000 7328 39016 7392
rect 39080 7328 39096 7392
rect 39160 7328 39176 7392
rect 39240 7328 39256 7392
rect 39320 7328 39336 7392
rect 39400 7328 39416 7392
rect 39480 7328 39496 7392
rect 39560 7328 39576 7392
rect 39640 7328 39656 7392
rect 39720 7328 39736 7392
rect 39800 7328 39816 7392
rect 39880 7328 39896 7392
rect 39960 7328 39976 7392
rect 40040 7328 40056 7392
rect 40120 7328 40136 7392
rect 40200 7328 40216 7392
rect 40280 7328 40296 7392
rect 40360 7328 40368 7392
rect 36368 7312 40368 7328
rect 36368 7248 36376 7312
rect 36440 7248 36456 7312
rect 36520 7248 36536 7312
rect 36600 7248 36616 7312
rect 36680 7248 36696 7312
rect 36760 7248 36776 7312
rect 36840 7248 36856 7312
rect 36920 7248 36936 7312
rect 37000 7248 37016 7312
rect 37080 7248 37096 7312
rect 37160 7248 37176 7312
rect 37240 7248 37256 7312
rect 37320 7248 37336 7312
rect 37400 7248 37416 7312
rect 37480 7248 37496 7312
rect 37560 7248 37576 7312
rect 37640 7248 37656 7312
rect 37720 7248 37736 7312
rect 37800 7248 37816 7312
rect 37880 7248 37896 7312
rect 37960 7248 37976 7312
rect 38040 7248 38056 7312
rect 38120 7248 38136 7312
rect 38200 7248 38216 7312
rect 38280 7248 38296 7312
rect 38360 7248 38376 7312
rect 38440 7248 38456 7312
rect 38520 7248 38536 7312
rect 38600 7248 38616 7312
rect 38680 7248 38696 7312
rect 38760 7248 38776 7312
rect 38840 7248 38856 7312
rect 38920 7248 38936 7312
rect 39000 7248 39016 7312
rect 39080 7248 39096 7312
rect 39160 7248 39176 7312
rect 39240 7248 39256 7312
rect 39320 7248 39336 7312
rect 39400 7248 39416 7312
rect 39480 7248 39496 7312
rect 39560 7248 39576 7312
rect 39640 7248 39656 7312
rect 39720 7248 39736 7312
rect 39800 7248 39816 7312
rect 39880 7248 39896 7312
rect 39960 7248 39976 7312
rect 40040 7248 40056 7312
rect 40120 7248 40136 7312
rect 40200 7248 40216 7312
rect 40280 7248 40296 7312
rect 40360 7248 40368 7312
rect 36368 7232 40368 7248
rect 36368 7168 36376 7232
rect 36440 7168 36456 7232
rect 36520 7168 36536 7232
rect 36600 7168 36616 7232
rect 36680 7168 36696 7232
rect 36760 7168 36776 7232
rect 36840 7168 36856 7232
rect 36920 7168 36936 7232
rect 37000 7168 37016 7232
rect 37080 7168 37096 7232
rect 37160 7168 37176 7232
rect 37240 7168 37256 7232
rect 37320 7168 37336 7232
rect 37400 7168 37416 7232
rect 37480 7168 37496 7232
rect 37560 7168 37576 7232
rect 37640 7168 37656 7232
rect 37720 7168 37736 7232
rect 37800 7168 37816 7232
rect 37880 7168 37896 7232
rect 37960 7168 37976 7232
rect 38040 7168 38056 7232
rect 38120 7168 38136 7232
rect 38200 7168 38216 7232
rect 38280 7168 38296 7232
rect 38360 7168 38376 7232
rect 38440 7168 38456 7232
rect 38520 7168 38536 7232
rect 38600 7168 38616 7232
rect 38680 7168 38696 7232
rect 38760 7168 38776 7232
rect 38840 7168 38856 7232
rect 38920 7168 38936 7232
rect 39000 7168 39016 7232
rect 39080 7168 39096 7232
rect 39160 7168 39176 7232
rect 39240 7168 39256 7232
rect 39320 7168 39336 7232
rect 39400 7168 39416 7232
rect 39480 7168 39496 7232
rect 39560 7168 39576 7232
rect 39640 7168 39656 7232
rect 39720 7168 39736 7232
rect 39800 7168 39816 7232
rect 39880 7168 39896 7232
rect 39960 7168 39976 7232
rect 40040 7168 40056 7232
rect 40120 7168 40136 7232
rect 40200 7168 40216 7232
rect 40280 7168 40296 7232
rect 40360 7168 40368 7232
rect 36368 7152 40368 7168
rect 36368 7088 36376 7152
rect 36440 7088 36456 7152
rect 36520 7088 36536 7152
rect 36600 7088 36616 7152
rect 36680 7088 36696 7152
rect 36760 7088 36776 7152
rect 36840 7088 36856 7152
rect 36920 7088 36936 7152
rect 37000 7088 37016 7152
rect 37080 7088 37096 7152
rect 37160 7088 37176 7152
rect 37240 7088 37256 7152
rect 37320 7088 37336 7152
rect 37400 7088 37416 7152
rect 37480 7088 37496 7152
rect 37560 7088 37576 7152
rect 37640 7088 37656 7152
rect 37720 7088 37736 7152
rect 37800 7088 37816 7152
rect 37880 7088 37896 7152
rect 37960 7088 37976 7152
rect 38040 7088 38056 7152
rect 38120 7088 38136 7152
rect 38200 7088 38216 7152
rect 38280 7088 38296 7152
rect 38360 7088 38376 7152
rect 38440 7088 38456 7152
rect 38520 7088 38536 7152
rect 38600 7088 38616 7152
rect 38680 7088 38696 7152
rect 38760 7088 38776 7152
rect 38840 7088 38856 7152
rect 38920 7088 38936 7152
rect 39000 7088 39016 7152
rect 39080 7088 39096 7152
rect 39160 7088 39176 7152
rect 39240 7088 39256 7152
rect 39320 7088 39336 7152
rect 39400 7088 39416 7152
rect 39480 7088 39496 7152
rect 39560 7088 39576 7152
rect 39640 7088 39656 7152
rect 39720 7088 39736 7152
rect 39800 7088 39816 7152
rect 39880 7088 39896 7152
rect 39960 7088 39976 7152
rect 40040 7088 40056 7152
rect 40120 7088 40136 7152
rect 40200 7088 40216 7152
rect 40280 7088 40296 7152
rect 40360 7088 40368 7152
rect 36368 7072 40368 7088
rect 36368 7008 36376 7072
rect 36440 7008 36456 7072
rect 36520 7008 36536 7072
rect 36600 7008 36616 7072
rect 36680 7008 36696 7072
rect 36760 7008 36776 7072
rect 36840 7008 36856 7072
rect 36920 7008 36936 7072
rect 37000 7008 37016 7072
rect 37080 7008 37096 7072
rect 37160 7008 37176 7072
rect 37240 7008 37256 7072
rect 37320 7008 37336 7072
rect 37400 7008 37416 7072
rect 37480 7008 37496 7072
rect 37560 7008 37576 7072
rect 37640 7008 37656 7072
rect 37720 7008 37736 7072
rect 37800 7008 37816 7072
rect 37880 7008 37896 7072
rect 37960 7008 37976 7072
rect 38040 7008 38056 7072
rect 38120 7008 38136 7072
rect 38200 7008 38216 7072
rect 38280 7008 38296 7072
rect 38360 7008 38376 7072
rect 38440 7008 38456 7072
rect 38520 7008 38536 7072
rect 38600 7008 38616 7072
rect 38680 7008 38696 7072
rect 38760 7008 38776 7072
rect 38840 7008 38856 7072
rect 38920 7008 38936 7072
rect 39000 7008 39016 7072
rect 39080 7008 39096 7072
rect 39160 7008 39176 7072
rect 39240 7008 39256 7072
rect 39320 7008 39336 7072
rect 39400 7008 39416 7072
rect 39480 7008 39496 7072
rect 39560 7008 39576 7072
rect 39640 7008 39656 7072
rect 39720 7008 39736 7072
rect 39800 7008 39816 7072
rect 39880 7008 39896 7072
rect 39960 7008 39976 7072
rect 40040 7008 40056 7072
rect 40120 7008 40136 7072
rect 40200 7008 40216 7072
rect 40280 7008 40296 7072
rect 40360 7008 40368 7072
rect 36368 6992 40368 7008
rect 36368 6928 36376 6992
rect 36440 6928 36456 6992
rect 36520 6928 36536 6992
rect 36600 6928 36616 6992
rect 36680 6928 36696 6992
rect 36760 6928 36776 6992
rect 36840 6928 36856 6992
rect 36920 6928 36936 6992
rect 37000 6928 37016 6992
rect 37080 6928 37096 6992
rect 37160 6928 37176 6992
rect 37240 6928 37256 6992
rect 37320 6928 37336 6992
rect 37400 6928 37416 6992
rect 37480 6928 37496 6992
rect 37560 6928 37576 6992
rect 37640 6928 37656 6992
rect 37720 6928 37736 6992
rect 37800 6928 37816 6992
rect 37880 6928 37896 6992
rect 37960 6928 37976 6992
rect 38040 6928 38056 6992
rect 38120 6928 38136 6992
rect 38200 6928 38216 6992
rect 38280 6928 38296 6992
rect 38360 6928 38376 6992
rect 38440 6928 38456 6992
rect 38520 6928 38536 6992
rect 38600 6928 38616 6992
rect 38680 6928 38696 6992
rect 38760 6928 38776 6992
rect 38840 6928 38856 6992
rect 38920 6928 38936 6992
rect 39000 6928 39016 6992
rect 39080 6928 39096 6992
rect 39160 6928 39176 6992
rect 39240 6928 39256 6992
rect 39320 6928 39336 6992
rect 39400 6928 39416 6992
rect 39480 6928 39496 6992
rect 39560 6928 39576 6992
rect 39640 6928 39656 6992
rect 39720 6928 39736 6992
rect 39800 6928 39816 6992
rect 39880 6928 39896 6992
rect 39960 6928 39976 6992
rect 40040 6928 40056 6992
rect 40120 6928 40136 6992
rect 40200 6928 40216 6992
rect 40280 6928 40296 6992
rect 40360 6928 40368 6992
rect 36368 6912 40368 6928
rect 36368 6848 36376 6912
rect 36440 6848 36456 6912
rect 36520 6848 36536 6912
rect 36600 6848 36616 6912
rect 36680 6848 36696 6912
rect 36760 6848 36776 6912
rect 36840 6848 36856 6912
rect 36920 6848 36936 6912
rect 37000 6848 37016 6912
rect 37080 6848 37096 6912
rect 37160 6848 37176 6912
rect 37240 6848 37256 6912
rect 37320 6848 37336 6912
rect 37400 6848 37416 6912
rect 37480 6848 37496 6912
rect 37560 6848 37576 6912
rect 37640 6848 37656 6912
rect 37720 6848 37736 6912
rect 37800 6848 37816 6912
rect 37880 6848 37896 6912
rect 37960 6848 37976 6912
rect 38040 6848 38056 6912
rect 38120 6848 38136 6912
rect 38200 6848 38216 6912
rect 38280 6848 38296 6912
rect 38360 6848 38376 6912
rect 38440 6848 38456 6912
rect 38520 6848 38536 6912
rect 38600 6848 38616 6912
rect 38680 6848 38696 6912
rect 38760 6848 38776 6912
rect 38840 6848 38856 6912
rect 38920 6848 38936 6912
rect 39000 6848 39016 6912
rect 39080 6848 39096 6912
rect 39160 6848 39176 6912
rect 39240 6848 39256 6912
rect 39320 6848 39336 6912
rect 39400 6848 39416 6912
rect 39480 6848 39496 6912
rect 39560 6848 39576 6912
rect 39640 6848 39656 6912
rect 39720 6848 39736 6912
rect 39800 6848 39816 6912
rect 39880 6848 39896 6912
rect 39960 6848 39976 6912
rect 40040 6848 40056 6912
rect 40120 6848 40136 6912
rect 40200 6848 40216 6912
rect 40280 6848 40296 6912
rect 40360 6848 40368 6912
rect 36368 6832 40368 6848
rect 36368 6768 36376 6832
rect 36440 6768 36456 6832
rect 36520 6768 36536 6832
rect 36600 6768 36616 6832
rect 36680 6768 36696 6832
rect 36760 6768 36776 6832
rect 36840 6768 36856 6832
rect 36920 6768 36936 6832
rect 37000 6768 37016 6832
rect 37080 6768 37096 6832
rect 37160 6768 37176 6832
rect 37240 6768 37256 6832
rect 37320 6768 37336 6832
rect 37400 6768 37416 6832
rect 37480 6768 37496 6832
rect 37560 6768 37576 6832
rect 37640 6768 37656 6832
rect 37720 6768 37736 6832
rect 37800 6768 37816 6832
rect 37880 6768 37896 6832
rect 37960 6768 37976 6832
rect 38040 6768 38056 6832
rect 38120 6768 38136 6832
rect 38200 6768 38216 6832
rect 38280 6768 38296 6832
rect 38360 6768 38376 6832
rect 38440 6768 38456 6832
rect 38520 6768 38536 6832
rect 38600 6768 38616 6832
rect 38680 6768 38696 6832
rect 38760 6768 38776 6832
rect 38840 6768 38856 6832
rect 38920 6768 38936 6832
rect 39000 6768 39016 6832
rect 39080 6768 39096 6832
rect 39160 6768 39176 6832
rect 39240 6768 39256 6832
rect 39320 6768 39336 6832
rect 39400 6768 39416 6832
rect 39480 6768 39496 6832
rect 39560 6768 39576 6832
rect 39640 6768 39656 6832
rect 39720 6768 39736 6832
rect 39800 6768 39816 6832
rect 39880 6768 39896 6832
rect 39960 6768 39976 6832
rect 40040 6768 40056 6832
rect 40120 6768 40136 6832
rect 40200 6768 40216 6832
rect 40280 6768 40296 6832
rect 40360 6768 40368 6832
rect 36368 6752 40368 6768
rect 36368 6688 36376 6752
rect 36440 6688 36456 6752
rect 36520 6688 36536 6752
rect 36600 6688 36616 6752
rect 36680 6688 36696 6752
rect 36760 6688 36776 6752
rect 36840 6688 36856 6752
rect 36920 6688 36936 6752
rect 37000 6688 37016 6752
rect 37080 6688 37096 6752
rect 37160 6688 37176 6752
rect 37240 6688 37256 6752
rect 37320 6688 37336 6752
rect 37400 6688 37416 6752
rect 37480 6688 37496 6752
rect 37560 6688 37576 6752
rect 37640 6688 37656 6752
rect 37720 6688 37736 6752
rect 37800 6688 37816 6752
rect 37880 6688 37896 6752
rect 37960 6688 37976 6752
rect 38040 6688 38056 6752
rect 38120 6688 38136 6752
rect 38200 6688 38216 6752
rect 38280 6688 38296 6752
rect 38360 6688 38376 6752
rect 38440 6688 38456 6752
rect 38520 6688 38536 6752
rect 38600 6688 38616 6752
rect 38680 6688 38696 6752
rect 38760 6688 38776 6752
rect 38840 6688 38856 6752
rect 38920 6688 38936 6752
rect 39000 6688 39016 6752
rect 39080 6688 39096 6752
rect 39160 6688 39176 6752
rect 39240 6688 39256 6752
rect 39320 6688 39336 6752
rect 39400 6688 39416 6752
rect 39480 6688 39496 6752
rect 39560 6688 39576 6752
rect 39640 6688 39656 6752
rect 39720 6688 39736 6752
rect 39800 6688 39816 6752
rect 39880 6688 39896 6752
rect 39960 6688 39976 6752
rect 40040 6688 40056 6752
rect 40120 6688 40136 6752
rect 40200 6688 40216 6752
rect 40280 6688 40296 6752
rect 40360 6688 40368 6752
rect 36368 6672 40368 6688
rect 36368 6608 36376 6672
rect 36440 6608 36456 6672
rect 36520 6608 36536 6672
rect 36600 6608 36616 6672
rect 36680 6608 36696 6672
rect 36760 6608 36776 6672
rect 36840 6608 36856 6672
rect 36920 6608 36936 6672
rect 37000 6608 37016 6672
rect 37080 6608 37096 6672
rect 37160 6608 37176 6672
rect 37240 6608 37256 6672
rect 37320 6608 37336 6672
rect 37400 6608 37416 6672
rect 37480 6608 37496 6672
rect 37560 6608 37576 6672
rect 37640 6608 37656 6672
rect 37720 6608 37736 6672
rect 37800 6608 37816 6672
rect 37880 6608 37896 6672
rect 37960 6608 37976 6672
rect 38040 6608 38056 6672
rect 38120 6608 38136 6672
rect 38200 6608 38216 6672
rect 38280 6608 38296 6672
rect 38360 6608 38376 6672
rect 38440 6608 38456 6672
rect 38520 6608 38536 6672
rect 38600 6608 38616 6672
rect 38680 6608 38696 6672
rect 38760 6608 38776 6672
rect 38840 6608 38856 6672
rect 38920 6608 38936 6672
rect 39000 6608 39016 6672
rect 39080 6608 39096 6672
rect 39160 6608 39176 6672
rect 39240 6608 39256 6672
rect 39320 6608 39336 6672
rect 39400 6608 39416 6672
rect 39480 6608 39496 6672
rect 39560 6608 39576 6672
rect 39640 6608 39656 6672
rect 39720 6608 39736 6672
rect 39800 6608 39816 6672
rect 39880 6608 39896 6672
rect 39960 6608 39976 6672
rect 40040 6608 40056 6672
rect 40120 6608 40136 6672
rect 40200 6608 40216 6672
rect 40280 6608 40296 6672
rect 40360 6608 40368 6672
rect 36368 6592 40368 6608
rect 36368 6528 36376 6592
rect 36440 6528 36456 6592
rect 36520 6528 36536 6592
rect 36600 6528 36616 6592
rect 36680 6528 36696 6592
rect 36760 6528 36776 6592
rect 36840 6528 36856 6592
rect 36920 6528 36936 6592
rect 37000 6528 37016 6592
rect 37080 6528 37096 6592
rect 37160 6528 37176 6592
rect 37240 6528 37256 6592
rect 37320 6528 37336 6592
rect 37400 6528 37416 6592
rect 37480 6528 37496 6592
rect 37560 6528 37576 6592
rect 37640 6528 37656 6592
rect 37720 6528 37736 6592
rect 37800 6528 37816 6592
rect 37880 6528 37896 6592
rect 37960 6528 37976 6592
rect 38040 6528 38056 6592
rect 38120 6528 38136 6592
rect 38200 6528 38216 6592
rect 38280 6528 38296 6592
rect 38360 6528 38376 6592
rect 38440 6528 38456 6592
rect 38520 6528 38536 6592
rect 38600 6528 38616 6592
rect 38680 6528 38696 6592
rect 38760 6528 38776 6592
rect 38840 6528 38856 6592
rect 38920 6528 38936 6592
rect 39000 6528 39016 6592
rect 39080 6528 39096 6592
rect 39160 6528 39176 6592
rect 39240 6528 39256 6592
rect 39320 6528 39336 6592
rect 39400 6528 39416 6592
rect 39480 6528 39496 6592
rect 39560 6528 39576 6592
rect 39640 6528 39656 6592
rect 39720 6528 39736 6592
rect 39800 6528 39816 6592
rect 39880 6528 39896 6592
rect 39960 6528 39976 6592
rect 40040 6528 40056 6592
rect 40120 6528 40136 6592
rect 40200 6528 40216 6592
rect 40280 6528 40296 6592
rect 40360 6528 40368 6592
rect 36368 6512 40368 6528
rect 36368 6448 36376 6512
rect 36440 6448 36456 6512
rect 36520 6448 36536 6512
rect 36600 6448 36616 6512
rect 36680 6448 36696 6512
rect 36760 6448 36776 6512
rect 36840 6448 36856 6512
rect 36920 6448 36936 6512
rect 37000 6448 37016 6512
rect 37080 6448 37096 6512
rect 37160 6448 37176 6512
rect 37240 6448 37256 6512
rect 37320 6448 37336 6512
rect 37400 6448 37416 6512
rect 37480 6448 37496 6512
rect 37560 6448 37576 6512
rect 37640 6448 37656 6512
rect 37720 6448 37736 6512
rect 37800 6448 37816 6512
rect 37880 6448 37896 6512
rect 37960 6448 37976 6512
rect 38040 6448 38056 6512
rect 38120 6448 38136 6512
rect 38200 6448 38216 6512
rect 38280 6448 38296 6512
rect 38360 6448 38376 6512
rect 38440 6448 38456 6512
rect 38520 6448 38536 6512
rect 38600 6448 38616 6512
rect 38680 6448 38696 6512
rect 38760 6448 38776 6512
rect 38840 6448 38856 6512
rect 38920 6448 38936 6512
rect 39000 6448 39016 6512
rect 39080 6448 39096 6512
rect 39160 6448 39176 6512
rect 39240 6448 39256 6512
rect 39320 6448 39336 6512
rect 39400 6448 39416 6512
rect 39480 6448 39496 6512
rect 39560 6448 39576 6512
rect 39640 6448 39656 6512
rect 39720 6448 39736 6512
rect 39800 6448 39816 6512
rect 39880 6448 39896 6512
rect 39960 6448 39976 6512
rect 40040 6448 40056 6512
rect 40120 6448 40136 6512
rect 40200 6448 40216 6512
rect 40280 6448 40296 6512
rect 40360 6448 40368 6512
rect 36368 6432 40368 6448
rect 36368 6368 36376 6432
rect 36440 6368 36456 6432
rect 36520 6368 36536 6432
rect 36600 6368 36616 6432
rect 36680 6368 36696 6432
rect 36760 6368 36776 6432
rect 36840 6368 36856 6432
rect 36920 6368 36936 6432
rect 37000 6368 37016 6432
rect 37080 6368 37096 6432
rect 37160 6368 37176 6432
rect 37240 6368 37256 6432
rect 37320 6368 37336 6432
rect 37400 6368 37416 6432
rect 37480 6368 37496 6432
rect 37560 6368 37576 6432
rect 37640 6368 37656 6432
rect 37720 6368 37736 6432
rect 37800 6368 37816 6432
rect 37880 6368 37896 6432
rect 37960 6368 37976 6432
rect 38040 6368 38056 6432
rect 38120 6368 38136 6432
rect 38200 6368 38216 6432
rect 38280 6368 38296 6432
rect 38360 6368 38376 6432
rect 38440 6368 38456 6432
rect 38520 6368 38536 6432
rect 38600 6368 38616 6432
rect 38680 6368 38696 6432
rect 38760 6368 38776 6432
rect 38840 6368 38856 6432
rect 38920 6368 38936 6432
rect 39000 6368 39016 6432
rect 39080 6368 39096 6432
rect 39160 6368 39176 6432
rect 39240 6368 39256 6432
rect 39320 6368 39336 6432
rect 39400 6368 39416 6432
rect 39480 6368 39496 6432
rect 39560 6368 39576 6432
rect 39640 6368 39656 6432
rect 39720 6368 39736 6432
rect 39800 6368 39816 6432
rect 39880 6368 39896 6432
rect 39960 6368 39976 6432
rect 40040 6368 40056 6432
rect 40120 6368 40136 6432
rect 40200 6368 40216 6432
rect 40280 6368 40296 6432
rect 40360 6368 40368 6432
rect 36368 6352 40368 6368
rect 36368 6288 36376 6352
rect 36440 6288 36456 6352
rect 36520 6288 36536 6352
rect 36600 6288 36616 6352
rect 36680 6288 36696 6352
rect 36760 6288 36776 6352
rect 36840 6288 36856 6352
rect 36920 6288 36936 6352
rect 37000 6288 37016 6352
rect 37080 6288 37096 6352
rect 37160 6288 37176 6352
rect 37240 6288 37256 6352
rect 37320 6288 37336 6352
rect 37400 6288 37416 6352
rect 37480 6288 37496 6352
rect 37560 6288 37576 6352
rect 37640 6288 37656 6352
rect 37720 6288 37736 6352
rect 37800 6288 37816 6352
rect 37880 6288 37896 6352
rect 37960 6288 37976 6352
rect 38040 6288 38056 6352
rect 38120 6288 38136 6352
rect 38200 6288 38216 6352
rect 38280 6288 38296 6352
rect 38360 6288 38376 6352
rect 38440 6288 38456 6352
rect 38520 6288 38536 6352
rect 38600 6288 38616 6352
rect 38680 6288 38696 6352
rect 38760 6288 38776 6352
rect 38840 6288 38856 6352
rect 38920 6288 38936 6352
rect 39000 6288 39016 6352
rect 39080 6288 39096 6352
rect 39160 6288 39176 6352
rect 39240 6288 39256 6352
rect 39320 6288 39336 6352
rect 39400 6288 39416 6352
rect 39480 6288 39496 6352
rect 39560 6288 39576 6352
rect 39640 6288 39656 6352
rect 39720 6288 39736 6352
rect 39800 6288 39816 6352
rect 39880 6288 39896 6352
rect 39960 6288 39976 6352
rect 40040 6288 40056 6352
rect 40120 6288 40136 6352
rect 40200 6288 40216 6352
rect 40280 6288 40296 6352
rect 40360 6288 40368 6352
rect 36368 6272 40368 6288
rect 36368 6208 36376 6272
rect 36440 6208 36456 6272
rect 36520 6208 36536 6272
rect 36600 6208 36616 6272
rect 36680 6208 36696 6272
rect 36760 6208 36776 6272
rect 36840 6208 36856 6272
rect 36920 6208 36936 6272
rect 37000 6208 37016 6272
rect 37080 6208 37096 6272
rect 37160 6208 37176 6272
rect 37240 6208 37256 6272
rect 37320 6208 37336 6272
rect 37400 6208 37416 6272
rect 37480 6208 37496 6272
rect 37560 6208 37576 6272
rect 37640 6208 37656 6272
rect 37720 6208 37736 6272
rect 37800 6208 37816 6272
rect 37880 6208 37896 6272
rect 37960 6208 37976 6272
rect 38040 6208 38056 6272
rect 38120 6208 38136 6272
rect 38200 6208 38216 6272
rect 38280 6208 38296 6272
rect 38360 6208 38376 6272
rect 38440 6208 38456 6272
rect 38520 6208 38536 6272
rect 38600 6208 38616 6272
rect 38680 6208 38696 6272
rect 38760 6208 38776 6272
rect 38840 6208 38856 6272
rect 38920 6208 38936 6272
rect 39000 6208 39016 6272
rect 39080 6208 39096 6272
rect 39160 6208 39176 6272
rect 39240 6208 39256 6272
rect 39320 6208 39336 6272
rect 39400 6208 39416 6272
rect 39480 6208 39496 6272
rect 39560 6208 39576 6272
rect 39640 6208 39656 6272
rect 39720 6208 39736 6272
rect 39800 6208 39816 6272
rect 39880 6208 39896 6272
rect 39960 6208 39976 6272
rect 40040 6208 40056 6272
rect 40120 6208 40136 6272
rect 40200 6208 40216 6272
rect 40280 6208 40296 6272
rect 40360 6208 40368 6272
rect 36368 6192 40368 6208
rect 36368 6128 36376 6192
rect 36440 6128 36456 6192
rect 36520 6128 36536 6192
rect 36600 6128 36616 6192
rect 36680 6128 36696 6192
rect 36760 6128 36776 6192
rect 36840 6128 36856 6192
rect 36920 6128 36936 6192
rect 37000 6128 37016 6192
rect 37080 6128 37096 6192
rect 37160 6128 37176 6192
rect 37240 6128 37256 6192
rect 37320 6128 37336 6192
rect 37400 6128 37416 6192
rect 37480 6128 37496 6192
rect 37560 6128 37576 6192
rect 37640 6128 37656 6192
rect 37720 6128 37736 6192
rect 37800 6128 37816 6192
rect 37880 6128 37896 6192
rect 37960 6128 37976 6192
rect 38040 6128 38056 6192
rect 38120 6128 38136 6192
rect 38200 6128 38216 6192
rect 38280 6128 38296 6192
rect 38360 6128 38376 6192
rect 38440 6128 38456 6192
rect 38520 6128 38536 6192
rect 38600 6128 38616 6192
rect 38680 6128 38696 6192
rect 38760 6128 38776 6192
rect 38840 6128 38856 6192
rect 38920 6128 38936 6192
rect 39000 6128 39016 6192
rect 39080 6128 39096 6192
rect 39160 6128 39176 6192
rect 39240 6128 39256 6192
rect 39320 6128 39336 6192
rect 39400 6128 39416 6192
rect 39480 6128 39496 6192
rect 39560 6128 39576 6192
rect 39640 6128 39656 6192
rect 39720 6128 39736 6192
rect 39800 6128 39816 6192
rect 39880 6128 39896 6192
rect 39960 6128 39976 6192
rect 40040 6128 40056 6192
rect 40120 6128 40136 6192
rect 40200 6128 40216 6192
rect 40280 6128 40296 6192
rect 40360 6128 40368 6192
rect 36368 6112 40368 6128
rect 36368 6048 36376 6112
rect 36440 6048 36456 6112
rect 36520 6048 36536 6112
rect 36600 6048 36616 6112
rect 36680 6048 36696 6112
rect 36760 6048 36776 6112
rect 36840 6048 36856 6112
rect 36920 6048 36936 6112
rect 37000 6048 37016 6112
rect 37080 6048 37096 6112
rect 37160 6048 37176 6112
rect 37240 6048 37256 6112
rect 37320 6048 37336 6112
rect 37400 6048 37416 6112
rect 37480 6048 37496 6112
rect 37560 6048 37576 6112
rect 37640 6048 37656 6112
rect 37720 6048 37736 6112
rect 37800 6048 37816 6112
rect 37880 6048 37896 6112
rect 37960 6048 37976 6112
rect 38040 6048 38056 6112
rect 38120 6048 38136 6112
rect 38200 6048 38216 6112
rect 38280 6048 38296 6112
rect 38360 6048 38376 6112
rect 38440 6048 38456 6112
rect 38520 6048 38536 6112
rect 38600 6048 38616 6112
rect 38680 6048 38696 6112
rect 38760 6048 38776 6112
rect 38840 6048 38856 6112
rect 38920 6048 38936 6112
rect 39000 6048 39016 6112
rect 39080 6048 39096 6112
rect 39160 6048 39176 6112
rect 39240 6048 39256 6112
rect 39320 6048 39336 6112
rect 39400 6048 39416 6112
rect 39480 6048 39496 6112
rect 39560 6048 39576 6112
rect 39640 6048 39656 6112
rect 39720 6048 39736 6112
rect 39800 6048 39816 6112
rect 39880 6048 39896 6112
rect 39960 6048 39976 6112
rect 40040 6048 40056 6112
rect 40120 6048 40136 6112
rect 40200 6048 40216 6112
rect 40280 6048 40296 6112
rect 40360 6048 40368 6112
rect 36368 6032 40368 6048
rect 36368 5968 36376 6032
rect 36440 5968 36456 6032
rect 36520 5968 36536 6032
rect 36600 5968 36616 6032
rect 36680 5968 36696 6032
rect 36760 5968 36776 6032
rect 36840 5968 36856 6032
rect 36920 5968 36936 6032
rect 37000 5968 37016 6032
rect 37080 5968 37096 6032
rect 37160 5968 37176 6032
rect 37240 5968 37256 6032
rect 37320 5968 37336 6032
rect 37400 5968 37416 6032
rect 37480 5968 37496 6032
rect 37560 5968 37576 6032
rect 37640 5968 37656 6032
rect 37720 5968 37736 6032
rect 37800 5968 37816 6032
rect 37880 5968 37896 6032
rect 37960 5968 37976 6032
rect 38040 5968 38056 6032
rect 38120 5968 38136 6032
rect 38200 5968 38216 6032
rect 38280 5968 38296 6032
rect 38360 5968 38376 6032
rect 38440 5968 38456 6032
rect 38520 5968 38536 6032
rect 38600 5968 38616 6032
rect 38680 5968 38696 6032
rect 38760 5968 38776 6032
rect 38840 5968 38856 6032
rect 38920 5968 38936 6032
rect 39000 5968 39016 6032
rect 39080 5968 39096 6032
rect 39160 5968 39176 6032
rect 39240 5968 39256 6032
rect 39320 5968 39336 6032
rect 39400 5968 39416 6032
rect 39480 5968 39496 6032
rect 39560 5968 39576 6032
rect 39640 5968 39656 6032
rect 39720 5968 39736 6032
rect 39800 5968 39816 6032
rect 39880 5968 39896 6032
rect 39960 5968 39976 6032
rect 40040 5968 40056 6032
rect 40120 5968 40136 6032
rect 40200 5968 40216 6032
rect 40280 5968 40296 6032
rect 40360 5968 40368 6032
rect 36368 5952 40368 5968
rect 36368 5888 36376 5952
rect 36440 5888 36456 5952
rect 36520 5888 36536 5952
rect 36600 5888 36616 5952
rect 36680 5888 36696 5952
rect 36760 5888 36776 5952
rect 36840 5888 36856 5952
rect 36920 5888 36936 5952
rect 37000 5888 37016 5952
rect 37080 5888 37096 5952
rect 37160 5888 37176 5952
rect 37240 5888 37256 5952
rect 37320 5888 37336 5952
rect 37400 5888 37416 5952
rect 37480 5888 37496 5952
rect 37560 5888 37576 5952
rect 37640 5888 37656 5952
rect 37720 5888 37736 5952
rect 37800 5888 37816 5952
rect 37880 5888 37896 5952
rect 37960 5888 37976 5952
rect 38040 5888 38056 5952
rect 38120 5888 38136 5952
rect 38200 5888 38216 5952
rect 38280 5888 38296 5952
rect 38360 5888 38376 5952
rect 38440 5888 38456 5952
rect 38520 5888 38536 5952
rect 38600 5888 38616 5952
rect 38680 5888 38696 5952
rect 38760 5888 38776 5952
rect 38840 5888 38856 5952
rect 38920 5888 38936 5952
rect 39000 5888 39016 5952
rect 39080 5888 39096 5952
rect 39160 5888 39176 5952
rect 39240 5888 39256 5952
rect 39320 5888 39336 5952
rect 39400 5888 39416 5952
rect 39480 5888 39496 5952
rect 39560 5888 39576 5952
rect 39640 5888 39656 5952
rect 39720 5888 39736 5952
rect 39800 5888 39816 5952
rect 39880 5888 39896 5952
rect 39960 5888 39976 5952
rect 40040 5888 40056 5952
rect 40120 5888 40136 5952
rect 40200 5888 40216 5952
rect 40280 5888 40296 5952
rect 40360 5888 40368 5952
rect 36368 5872 40368 5888
rect 36368 5808 36376 5872
rect 36440 5808 36456 5872
rect 36520 5808 36536 5872
rect 36600 5808 36616 5872
rect 36680 5808 36696 5872
rect 36760 5808 36776 5872
rect 36840 5808 36856 5872
rect 36920 5808 36936 5872
rect 37000 5808 37016 5872
rect 37080 5808 37096 5872
rect 37160 5808 37176 5872
rect 37240 5808 37256 5872
rect 37320 5808 37336 5872
rect 37400 5808 37416 5872
rect 37480 5808 37496 5872
rect 37560 5808 37576 5872
rect 37640 5808 37656 5872
rect 37720 5808 37736 5872
rect 37800 5808 37816 5872
rect 37880 5808 37896 5872
rect 37960 5808 37976 5872
rect 38040 5808 38056 5872
rect 38120 5808 38136 5872
rect 38200 5808 38216 5872
rect 38280 5808 38296 5872
rect 38360 5808 38376 5872
rect 38440 5808 38456 5872
rect 38520 5808 38536 5872
rect 38600 5808 38616 5872
rect 38680 5808 38696 5872
rect 38760 5808 38776 5872
rect 38840 5808 38856 5872
rect 38920 5808 38936 5872
rect 39000 5808 39016 5872
rect 39080 5808 39096 5872
rect 39160 5808 39176 5872
rect 39240 5808 39256 5872
rect 39320 5808 39336 5872
rect 39400 5808 39416 5872
rect 39480 5808 39496 5872
rect 39560 5808 39576 5872
rect 39640 5808 39656 5872
rect 39720 5808 39736 5872
rect 39800 5808 39816 5872
rect 39880 5808 39896 5872
rect 39960 5808 39976 5872
rect 40040 5808 40056 5872
rect 40120 5808 40136 5872
rect 40200 5808 40216 5872
rect 40280 5808 40296 5872
rect 40360 5808 40368 5872
rect 36368 5792 40368 5808
rect 36368 5728 36376 5792
rect 36440 5728 36456 5792
rect 36520 5728 36536 5792
rect 36600 5728 36616 5792
rect 36680 5728 36696 5792
rect 36760 5728 36776 5792
rect 36840 5728 36856 5792
rect 36920 5728 36936 5792
rect 37000 5728 37016 5792
rect 37080 5728 37096 5792
rect 37160 5728 37176 5792
rect 37240 5728 37256 5792
rect 37320 5728 37336 5792
rect 37400 5728 37416 5792
rect 37480 5728 37496 5792
rect 37560 5728 37576 5792
rect 37640 5728 37656 5792
rect 37720 5728 37736 5792
rect 37800 5728 37816 5792
rect 37880 5728 37896 5792
rect 37960 5728 37976 5792
rect 38040 5728 38056 5792
rect 38120 5728 38136 5792
rect 38200 5728 38216 5792
rect 38280 5728 38296 5792
rect 38360 5728 38376 5792
rect 38440 5728 38456 5792
rect 38520 5728 38536 5792
rect 38600 5728 38616 5792
rect 38680 5728 38696 5792
rect 38760 5728 38776 5792
rect 38840 5728 38856 5792
rect 38920 5728 38936 5792
rect 39000 5728 39016 5792
rect 39080 5728 39096 5792
rect 39160 5728 39176 5792
rect 39240 5728 39256 5792
rect 39320 5728 39336 5792
rect 39400 5728 39416 5792
rect 39480 5728 39496 5792
rect 39560 5728 39576 5792
rect 39640 5728 39656 5792
rect 39720 5728 39736 5792
rect 39800 5728 39816 5792
rect 39880 5728 39896 5792
rect 39960 5728 39976 5792
rect 40040 5728 40056 5792
rect 40120 5728 40136 5792
rect 40200 5728 40216 5792
rect 40280 5728 40296 5792
rect 40360 5728 40368 5792
rect 36368 5712 40368 5728
rect 36368 5648 36376 5712
rect 36440 5648 36456 5712
rect 36520 5648 36536 5712
rect 36600 5648 36616 5712
rect 36680 5648 36696 5712
rect 36760 5648 36776 5712
rect 36840 5648 36856 5712
rect 36920 5648 36936 5712
rect 37000 5648 37016 5712
rect 37080 5648 37096 5712
rect 37160 5648 37176 5712
rect 37240 5648 37256 5712
rect 37320 5648 37336 5712
rect 37400 5648 37416 5712
rect 37480 5648 37496 5712
rect 37560 5648 37576 5712
rect 37640 5648 37656 5712
rect 37720 5648 37736 5712
rect 37800 5648 37816 5712
rect 37880 5648 37896 5712
rect 37960 5648 37976 5712
rect 38040 5648 38056 5712
rect 38120 5648 38136 5712
rect 38200 5648 38216 5712
rect 38280 5648 38296 5712
rect 38360 5648 38376 5712
rect 38440 5648 38456 5712
rect 38520 5648 38536 5712
rect 38600 5648 38616 5712
rect 38680 5648 38696 5712
rect 38760 5648 38776 5712
rect 38840 5648 38856 5712
rect 38920 5648 38936 5712
rect 39000 5648 39016 5712
rect 39080 5648 39096 5712
rect 39160 5648 39176 5712
rect 39240 5648 39256 5712
rect 39320 5648 39336 5712
rect 39400 5648 39416 5712
rect 39480 5648 39496 5712
rect 39560 5648 39576 5712
rect 39640 5648 39656 5712
rect 39720 5648 39736 5712
rect 39800 5648 39816 5712
rect 39880 5648 39896 5712
rect 39960 5648 39976 5712
rect 40040 5648 40056 5712
rect 40120 5648 40136 5712
rect 40200 5648 40216 5712
rect 40280 5648 40296 5712
rect 40360 5648 40368 5712
rect 36368 5632 40368 5648
rect 36368 5568 36376 5632
rect 36440 5568 36456 5632
rect 36520 5568 36536 5632
rect 36600 5568 36616 5632
rect 36680 5568 36696 5632
rect 36760 5568 36776 5632
rect 36840 5568 36856 5632
rect 36920 5568 36936 5632
rect 37000 5568 37016 5632
rect 37080 5568 37096 5632
rect 37160 5568 37176 5632
rect 37240 5568 37256 5632
rect 37320 5568 37336 5632
rect 37400 5568 37416 5632
rect 37480 5568 37496 5632
rect 37560 5568 37576 5632
rect 37640 5568 37656 5632
rect 37720 5568 37736 5632
rect 37800 5568 37816 5632
rect 37880 5568 37896 5632
rect 37960 5568 37976 5632
rect 38040 5568 38056 5632
rect 38120 5568 38136 5632
rect 38200 5568 38216 5632
rect 38280 5568 38296 5632
rect 38360 5568 38376 5632
rect 38440 5568 38456 5632
rect 38520 5568 38536 5632
rect 38600 5568 38616 5632
rect 38680 5568 38696 5632
rect 38760 5568 38776 5632
rect 38840 5568 38856 5632
rect 38920 5568 38936 5632
rect 39000 5568 39016 5632
rect 39080 5568 39096 5632
rect 39160 5568 39176 5632
rect 39240 5568 39256 5632
rect 39320 5568 39336 5632
rect 39400 5568 39416 5632
rect 39480 5568 39496 5632
rect 39560 5568 39576 5632
rect 39640 5568 39656 5632
rect 39720 5568 39736 5632
rect 39800 5568 39816 5632
rect 39880 5568 39896 5632
rect 39960 5568 39976 5632
rect 40040 5568 40056 5632
rect 40120 5568 40136 5632
rect 40200 5568 40216 5632
rect 40280 5568 40296 5632
rect 40360 5568 40368 5632
rect 36368 5552 40368 5568
rect 36368 5488 36376 5552
rect 36440 5488 36456 5552
rect 36520 5488 36536 5552
rect 36600 5488 36616 5552
rect 36680 5488 36696 5552
rect 36760 5488 36776 5552
rect 36840 5488 36856 5552
rect 36920 5488 36936 5552
rect 37000 5488 37016 5552
rect 37080 5488 37096 5552
rect 37160 5488 37176 5552
rect 37240 5488 37256 5552
rect 37320 5488 37336 5552
rect 37400 5488 37416 5552
rect 37480 5488 37496 5552
rect 37560 5488 37576 5552
rect 37640 5488 37656 5552
rect 37720 5488 37736 5552
rect 37800 5488 37816 5552
rect 37880 5488 37896 5552
rect 37960 5488 37976 5552
rect 38040 5488 38056 5552
rect 38120 5488 38136 5552
rect 38200 5488 38216 5552
rect 38280 5488 38296 5552
rect 38360 5488 38376 5552
rect 38440 5488 38456 5552
rect 38520 5488 38536 5552
rect 38600 5488 38616 5552
rect 38680 5488 38696 5552
rect 38760 5488 38776 5552
rect 38840 5488 38856 5552
rect 38920 5488 38936 5552
rect 39000 5488 39016 5552
rect 39080 5488 39096 5552
rect 39160 5488 39176 5552
rect 39240 5488 39256 5552
rect 39320 5488 39336 5552
rect 39400 5488 39416 5552
rect 39480 5488 39496 5552
rect 39560 5488 39576 5552
rect 39640 5488 39656 5552
rect 39720 5488 39736 5552
rect 39800 5488 39816 5552
rect 39880 5488 39896 5552
rect 39960 5488 39976 5552
rect 40040 5488 40056 5552
rect 40120 5488 40136 5552
rect 40200 5488 40216 5552
rect 40280 5488 40296 5552
rect 40360 5488 40368 5552
rect 36368 5472 40368 5488
rect 36368 5408 36376 5472
rect 36440 5408 36456 5472
rect 36520 5408 36536 5472
rect 36600 5408 36616 5472
rect 36680 5408 36696 5472
rect 36760 5408 36776 5472
rect 36840 5408 36856 5472
rect 36920 5408 36936 5472
rect 37000 5408 37016 5472
rect 37080 5408 37096 5472
rect 37160 5408 37176 5472
rect 37240 5408 37256 5472
rect 37320 5408 37336 5472
rect 37400 5408 37416 5472
rect 37480 5408 37496 5472
rect 37560 5408 37576 5472
rect 37640 5408 37656 5472
rect 37720 5408 37736 5472
rect 37800 5408 37816 5472
rect 37880 5408 37896 5472
rect 37960 5408 37976 5472
rect 38040 5408 38056 5472
rect 38120 5408 38136 5472
rect 38200 5408 38216 5472
rect 38280 5408 38296 5472
rect 38360 5408 38376 5472
rect 38440 5408 38456 5472
rect 38520 5408 38536 5472
rect 38600 5408 38616 5472
rect 38680 5408 38696 5472
rect 38760 5408 38776 5472
rect 38840 5408 38856 5472
rect 38920 5408 38936 5472
rect 39000 5408 39016 5472
rect 39080 5408 39096 5472
rect 39160 5408 39176 5472
rect 39240 5408 39256 5472
rect 39320 5408 39336 5472
rect 39400 5408 39416 5472
rect 39480 5408 39496 5472
rect 39560 5408 39576 5472
rect 39640 5408 39656 5472
rect 39720 5408 39736 5472
rect 39800 5408 39816 5472
rect 39880 5408 39896 5472
rect 39960 5408 39976 5472
rect 40040 5408 40056 5472
rect 40120 5408 40136 5472
rect 40200 5408 40216 5472
rect 40280 5408 40296 5472
rect 40360 5408 40368 5472
rect 36368 5392 40368 5408
rect 36368 5328 36376 5392
rect 36440 5328 36456 5392
rect 36520 5328 36536 5392
rect 36600 5328 36616 5392
rect 36680 5328 36696 5392
rect 36760 5328 36776 5392
rect 36840 5328 36856 5392
rect 36920 5328 36936 5392
rect 37000 5328 37016 5392
rect 37080 5328 37096 5392
rect 37160 5328 37176 5392
rect 37240 5328 37256 5392
rect 37320 5328 37336 5392
rect 37400 5328 37416 5392
rect 37480 5328 37496 5392
rect 37560 5328 37576 5392
rect 37640 5328 37656 5392
rect 37720 5328 37736 5392
rect 37800 5328 37816 5392
rect 37880 5328 37896 5392
rect 37960 5328 37976 5392
rect 38040 5328 38056 5392
rect 38120 5328 38136 5392
rect 38200 5328 38216 5392
rect 38280 5328 38296 5392
rect 38360 5328 38376 5392
rect 38440 5328 38456 5392
rect 38520 5328 38536 5392
rect 38600 5328 38616 5392
rect 38680 5328 38696 5392
rect 38760 5328 38776 5392
rect 38840 5328 38856 5392
rect 38920 5328 38936 5392
rect 39000 5328 39016 5392
rect 39080 5328 39096 5392
rect 39160 5328 39176 5392
rect 39240 5328 39256 5392
rect 39320 5328 39336 5392
rect 39400 5328 39416 5392
rect 39480 5328 39496 5392
rect 39560 5328 39576 5392
rect 39640 5328 39656 5392
rect 39720 5328 39736 5392
rect 39800 5328 39816 5392
rect 39880 5328 39896 5392
rect 39960 5328 39976 5392
rect 40040 5328 40056 5392
rect 40120 5328 40136 5392
rect 40200 5328 40216 5392
rect 40280 5328 40296 5392
rect 40360 5328 40368 5392
rect 36368 5312 40368 5328
rect 36368 5248 36376 5312
rect 36440 5248 36456 5312
rect 36520 5248 36536 5312
rect 36600 5248 36616 5312
rect 36680 5248 36696 5312
rect 36760 5248 36776 5312
rect 36840 5248 36856 5312
rect 36920 5248 36936 5312
rect 37000 5248 37016 5312
rect 37080 5248 37096 5312
rect 37160 5248 37176 5312
rect 37240 5248 37256 5312
rect 37320 5248 37336 5312
rect 37400 5248 37416 5312
rect 37480 5248 37496 5312
rect 37560 5248 37576 5312
rect 37640 5248 37656 5312
rect 37720 5248 37736 5312
rect 37800 5248 37816 5312
rect 37880 5248 37896 5312
rect 37960 5248 37976 5312
rect 38040 5248 38056 5312
rect 38120 5248 38136 5312
rect 38200 5248 38216 5312
rect 38280 5248 38296 5312
rect 38360 5248 38376 5312
rect 38440 5248 38456 5312
rect 38520 5248 38536 5312
rect 38600 5248 38616 5312
rect 38680 5248 38696 5312
rect 38760 5248 38776 5312
rect 38840 5248 38856 5312
rect 38920 5248 38936 5312
rect 39000 5248 39016 5312
rect 39080 5248 39096 5312
rect 39160 5248 39176 5312
rect 39240 5248 39256 5312
rect 39320 5248 39336 5312
rect 39400 5248 39416 5312
rect 39480 5248 39496 5312
rect 39560 5248 39576 5312
rect 39640 5248 39656 5312
rect 39720 5248 39736 5312
rect 39800 5248 39816 5312
rect 39880 5248 39896 5312
rect 39960 5248 39976 5312
rect 40040 5248 40056 5312
rect 40120 5248 40136 5312
rect 40200 5248 40216 5312
rect 40280 5248 40296 5312
rect 40360 5248 40368 5312
rect 36368 5232 40368 5248
rect 36368 5168 36376 5232
rect 36440 5168 36456 5232
rect 36520 5168 36536 5232
rect 36600 5168 36616 5232
rect 36680 5168 36696 5232
rect 36760 5168 36776 5232
rect 36840 5168 36856 5232
rect 36920 5168 36936 5232
rect 37000 5168 37016 5232
rect 37080 5168 37096 5232
rect 37160 5168 37176 5232
rect 37240 5168 37256 5232
rect 37320 5168 37336 5232
rect 37400 5168 37416 5232
rect 37480 5168 37496 5232
rect 37560 5168 37576 5232
rect 37640 5168 37656 5232
rect 37720 5168 37736 5232
rect 37800 5168 37816 5232
rect 37880 5168 37896 5232
rect 37960 5168 37976 5232
rect 38040 5168 38056 5232
rect 38120 5168 38136 5232
rect 38200 5168 38216 5232
rect 38280 5168 38296 5232
rect 38360 5168 38376 5232
rect 38440 5168 38456 5232
rect 38520 5168 38536 5232
rect 38600 5168 38616 5232
rect 38680 5168 38696 5232
rect 38760 5168 38776 5232
rect 38840 5168 38856 5232
rect 38920 5168 38936 5232
rect 39000 5168 39016 5232
rect 39080 5168 39096 5232
rect 39160 5168 39176 5232
rect 39240 5168 39256 5232
rect 39320 5168 39336 5232
rect 39400 5168 39416 5232
rect 39480 5168 39496 5232
rect 39560 5168 39576 5232
rect 39640 5168 39656 5232
rect 39720 5168 39736 5232
rect 39800 5168 39816 5232
rect 39880 5168 39896 5232
rect 39960 5168 39976 5232
rect 40040 5168 40056 5232
rect 40120 5168 40136 5232
rect 40200 5168 40216 5232
rect 40280 5168 40296 5232
rect 40360 5168 40368 5232
rect 36368 5152 40368 5168
rect 36368 5088 36376 5152
rect 36440 5088 36456 5152
rect 36520 5088 36536 5152
rect 36600 5088 36616 5152
rect 36680 5088 36696 5152
rect 36760 5088 36776 5152
rect 36840 5088 36856 5152
rect 36920 5088 36936 5152
rect 37000 5088 37016 5152
rect 37080 5088 37096 5152
rect 37160 5088 37176 5152
rect 37240 5088 37256 5152
rect 37320 5088 37336 5152
rect 37400 5088 37416 5152
rect 37480 5088 37496 5152
rect 37560 5088 37576 5152
rect 37640 5088 37656 5152
rect 37720 5088 37736 5152
rect 37800 5088 37816 5152
rect 37880 5088 37896 5152
rect 37960 5088 37976 5152
rect 38040 5088 38056 5152
rect 38120 5088 38136 5152
rect 38200 5088 38216 5152
rect 38280 5088 38296 5152
rect 38360 5088 38376 5152
rect 38440 5088 38456 5152
rect 38520 5088 38536 5152
rect 38600 5088 38616 5152
rect 38680 5088 38696 5152
rect 38760 5088 38776 5152
rect 38840 5088 38856 5152
rect 38920 5088 38936 5152
rect 39000 5088 39016 5152
rect 39080 5088 39096 5152
rect 39160 5088 39176 5152
rect 39240 5088 39256 5152
rect 39320 5088 39336 5152
rect 39400 5088 39416 5152
rect 39480 5088 39496 5152
rect 39560 5088 39576 5152
rect 39640 5088 39656 5152
rect 39720 5088 39736 5152
rect 39800 5088 39816 5152
rect 39880 5088 39896 5152
rect 39960 5088 39976 5152
rect 40040 5088 40056 5152
rect 40120 5088 40136 5152
rect 40200 5088 40216 5152
rect 40280 5088 40296 5152
rect 40360 5088 40368 5152
rect 36368 5072 40368 5088
rect 36368 5008 36376 5072
rect 36440 5008 36456 5072
rect 36520 5008 36536 5072
rect 36600 5008 36616 5072
rect 36680 5008 36696 5072
rect 36760 5008 36776 5072
rect 36840 5008 36856 5072
rect 36920 5008 36936 5072
rect 37000 5008 37016 5072
rect 37080 5008 37096 5072
rect 37160 5008 37176 5072
rect 37240 5008 37256 5072
rect 37320 5008 37336 5072
rect 37400 5008 37416 5072
rect 37480 5008 37496 5072
rect 37560 5008 37576 5072
rect 37640 5008 37656 5072
rect 37720 5008 37736 5072
rect 37800 5008 37816 5072
rect 37880 5008 37896 5072
rect 37960 5008 37976 5072
rect 38040 5008 38056 5072
rect 38120 5008 38136 5072
rect 38200 5008 38216 5072
rect 38280 5008 38296 5072
rect 38360 5008 38376 5072
rect 38440 5008 38456 5072
rect 38520 5008 38536 5072
rect 38600 5008 38616 5072
rect 38680 5008 38696 5072
rect 38760 5008 38776 5072
rect 38840 5008 38856 5072
rect 38920 5008 38936 5072
rect 39000 5008 39016 5072
rect 39080 5008 39096 5072
rect 39160 5008 39176 5072
rect 39240 5008 39256 5072
rect 39320 5008 39336 5072
rect 39400 5008 39416 5072
rect 39480 5008 39496 5072
rect 39560 5008 39576 5072
rect 39640 5008 39656 5072
rect 39720 5008 39736 5072
rect 39800 5008 39816 5072
rect 39880 5008 39896 5072
rect 39960 5008 39976 5072
rect 40040 5008 40056 5072
rect 40120 5008 40136 5072
rect 40200 5008 40216 5072
rect 40280 5008 40296 5072
rect 40360 5008 40368 5072
rect 36368 5000 40368 5008
rect 29104 3928 29112 3992
rect 29176 3928 29192 3992
rect 29256 3928 29272 3992
rect 29336 3928 29352 3992
rect 29416 3928 29424 3992
rect 29104 3912 29424 3928
rect 29104 3848 29112 3912
rect 29176 3848 29192 3912
rect 29256 3848 29272 3912
rect 29336 3848 29352 3912
rect 29416 3848 29424 3912
rect 29104 3832 29424 3848
rect 29104 3768 29112 3832
rect 29176 3768 29192 3832
rect 29256 3768 29272 3832
rect 29336 3768 29352 3832
rect 29416 3768 29424 3832
rect 29104 3752 29424 3768
rect 29104 3688 29112 3752
rect 29176 3688 29192 3752
rect 29256 3688 29272 3752
rect 29336 3688 29352 3752
rect 29416 3688 29424 3752
rect 29104 3672 29424 3688
rect 29104 3608 29112 3672
rect 29176 3608 29192 3672
rect 29256 3608 29272 3672
rect 29336 3608 29352 3672
rect 29416 3608 29424 3672
rect 29104 3592 29424 3608
rect 29104 3528 29112 3592
rect 29176 3528 29192 3592
rect 29256 3528 29272 3592
rect 29336 3528 29352 3592
rect 29416 3528 29424 3592
rect 29104 3512 29424 3528
rect 29104 3448 29112 3512
rect 29176 3448 29192 3512
rect 29256 3448 29272 3512
rect 29336 3448 29352 3512
rect 29416 3448 29424 3512
rect 29104 3432 29424 3448
rect 29104 3368 29112 3432
rect 29176 3368 29192 3432
rect 29256 3368 29272 3432
rect 29336 3368 29352 3432
rect 29416 3368 29424 3432
rect 29104 3352 29424 3368
rect 29104 3288 29112 3352
rect 29176 3288 29192 3352
rect 29256 3288 29272 3352
rect 29336 3288 29352 3352
rect 29416 3288 29424 3352
rect 29104 3272 29424 3288
rect 29104 3208 29112 3272
rect 29176 3208 29192 3272
rect 29256 3208 29272 3272
rect 29336 3208 29352 3272
rect 29416 3208 29424 3272
rect 29104 3192 29424 3208
rect 29104 3128 29112 3192
rect 29176 3128 29192 3192
rect 29256 3128 29272 3192
rect 29336 3128 29352 3192
rect 29416 3128 29424 3192
rect 29104 3112 29424 3128
rect 29104 3048 29112 3112
rect 29176 3048 29192 3112
rect 29256 3048 29272 3112
rect 29336 3048 29352 3112
rect 29416 3048 29424 3112
rect 29104 3032 29424 3048
rect 29104 2968 29112 3032
rect 29176 2968 29192 3032
rect 29256 2968 29272 3032
rect 29336 2968 29352 3032
rect 29416 2968 29424 3032
rect 29104 2952 29424 2968
rect 29104 2888 29112 2952
rect 29176 2888 29192 2952
rect 29256 2888 29272 2952
rect 29336 2888 29352 2952
rect 29416 2888 29424 2952
rect 29104 2872 29424 2888
rect 29104 2808 29112 2872
rect 29176 2808 29192 2872
rect 29256 2808 29272 2872
rect 29336 2808 29352 2872
rect 29416 2808 29424 2872
rect 29104 2792 29424 2808
rect 29104 2728 29112 2792
rect 29176 2728 29192 2792
rect 29256 2728 29272 2792
rect 29336 2728 29352 2792
rect 29416 2728 29424 2792
rect 29104 2712 29424 2728
rect 29104 2648 29112 2712
rect 29176 2648 29192 2712
rect 29256 2648 29272 2712
rect 29336 2648 29352 2712
rect 29416 2648 29424 2712
rect 29104 2632 29424 2648
rect 29104 2568 29112 2632
rect 29176 2568 29192 2632
rect 29256 2568 29272 2632
rect 29336 2568 29352 2632
rect 29416 2568 29424 2632
rect 29104 2552 29424 2568
rect 29104 2488 29112 2552
rect 29176 2488 29192 2552
rect 29256 2488 29272 2552
rect 29336 2488 29352 2552
rect 29416 2488 29424 2552
rect 29104 2472 29424 2488
rect 29104 2408 29112 2472
rect 29176 2408 29192 2472
rect 29256 2408 29272 2472
rect 29336 2408 29352 2472
rect 29416 2408 29424 2472
rect 29104 2392 29424 2408
rect 29104 2328 29112 2392
rect 29176 2328 29192 2392
rect 29256 2328 29272 2392
rect 29336 2328 29352 2392
rect 29416 2328 29424 2392
rect 29104 2312 29424 2328
rect 29104 2248 29112 2312
rect 29176 2248 29192 2312
rect 29256 2248 29272 2312
rect 29336 2248 29352 2312
rect 29416 2248 29424 2312
rect 29104 2232 29424 2248
rect 29104 2168 29112 2232
rect 29176 2168 29192 2232
rect 29256 2168 29272 2232
rect 29336 2168 29352 2232
rect 29416 2168 29424 2232
rect 29104 2152 29424 2168
rect 29104 2088 29112 2152
rect 29176 2088 29192 2152
rect 29256 2088 29272 2152
rect 29336 2088 29352 2152
rect 29416 2088 29424 2152
rect 29104 2072 29424 2088
rect 29104 2008 29112 2072
rect 29176 2008 29192 2072
rect 29256 2008 29272 2072
rect 29336 2008 29352 2072
rect 29416 2008 29424 2072
rect 29104 1992 29424 2008
rect 29104 1928 29112 1992
rect 29176 1928 29192 1992
rect 29256 1928 29272 1992
rect 29336 1928 29352 1992
rect 29416 1928 29424 1992
rect 29104 1912 29424 1928
rect 29104 1848 29112 1912
rect 29176 1848 29192 1912
rect 29256 1848 29272 1912
rect 29336 1848 29352 1912
rect 29416 1848 29424 1912
rect 29104 1832 29424 1848
rect 29104 1768 29112 1832
rect 29176 1768 29192 1832
rect 29256 1768 29272 1832
rect 29336 1768 29352 1832
rect 29416 1768 29424 1832
rect 29104 1752 29424 1768
rect 29104 1688 29112 1752
rect 29176 1688 29192 1752
rect 29256 1688 29272 1752
rect 29336 1688 29352 1752
rect 29416 1688 29424 1752
rect 29104 1672 29424 1688
rect 29104 1608 29112 1672
rect 29176 1608 29192 1672
rect 29256 1608 29272 1672
rect 29336 1608 29352 1672
rect 29416 1608 29424 1672
rect 29104 1592 29424 1608
rect 29104 1528 29112 1592
rect 29176 1528 29192 1592
rect 29256 1528 29272 1592
rect 29336 1528 29352 1592
rect 29416 1528 29424 1592
rect 29104 1512 29424 1528
rect 29104 1448 29112 1512
rect 29176 1448 29192 1512
rect 29256 1448 29272 1512
rect 29336 1448 29352 1512
rect 29416 1448 29424 1512
rect 29104 1432 29424 1448
rect 29104 1368 29112 1432
rect 29176 1368 29192 1432
rect 29256 1368 29272 1432
rect 29336 1368 29352 1432
rect 29416 1368 29424 1432
rect 29104 1352 29424 1368
rect 29104 1288 29112 1352
rect 29176 1288 29192 1352
rect 29256 1288 29272 1352
rect 29336 1288 29352 1352
rect 29416 1288 29424 1352
rect 29104 1272 29424 1288
rect 29104 1208 29112 1272
rect 29176 1208 29192 1272
rect 29256 1208 29272 1272
rect 29336 1208 29352 1272
rect 29416 1208 29424 1272
rect 29104 1192 29424 1208
rect 29104 1128 29112 1192
rect 29176 1128 29192 1192
rect 29256 1128 29272 1192
rect 29336 1128 29352 1192
rect 29416 1128 29424 1192
rect 29104 1112 29424 1128
rect 29104 1048 29112 1112
rect 29176 1048 29192 1112
rect 29256 1048 29272 1112
rect 29336 1048 29352 1112
rect 29416 1048 29424 1112
rect 29104 1032 29424 1048
rect 29104 968 29112 1032
rect 29176 968 29192 1032
rect 29256 968 29272 1032
rect 29336 968 29352 1032
rect 29416 968 29424 1032
rect 29104 952 29424 968
rect 29104 888 29112 952
rect 29176 888 29192 952
rect 29256 888 29272 952
rect 29336 888 29352 952
rect 29416 888 29424 952
rect 29104 872 29424 888
rect 29104 808 29112 872
rect 29176 808 29192 872
rect 29256 808 29272 872
rect 29336 808 29352 872
rect 29416 808 29424 872
rect 29104 792 29424 808
rect 29104 728 29112 792
rect 29176 728 29192 792
rect 29256 728 29272 792
rect 29336 728 29352 792
rect 29416 728 29424 792
rect 29104 712 29424 728
rect 29104 648 29112 712
rect 29176 648 29192 712
rect 29256 648 29272 712
rect 29336 648 29352 712
rect 29416 648 29424 712
rect 29104 632 29424 648
rect 29104 568 29112 632
rect 29176 568 29192 632
rect 29256 568 29272 632
rect 29336 568 29352 632
rect 29416 568 29424 632
rect 29104 552 29424 568
rect 29104 488 29112 552
rect 29176 488 29192 552
rect 29256 488 29272 552
rect 29336 488 29352 552
rect 29416 488 29424 552
rect 29104 472 29424 488
rect 29104 408 29112 472
rect 29176 408 29192 472
rect 29256 408 29272 472
rect 29336 408 29352 472
rect 29416 408 29424 472
rect 29104 392 29424 408
rect 29104 328 29112 392
rect 29176 328 29192 392
rect 29256 328 29272 392
rect 29336 328 29352 392
rect 29416 328 29424 392
rect 29104 312 29424 328
rect 29104 248 29112 312
rect 29176 248 29192 312
rect 29256 248 29272 312
rect 29336 248 29352 312
rect 29416 248 29424 312
rect 29104 232 29424 248
rect 29104 168 29112 232
rect 29176 168 29192 232
rect 29256 168 29272 232
rect 29336 168 29352 232
rect 29416 168 29424 232
rect 29104 152 29424 168
rect 29104 88 29112 152
rect 29176 88 29192 152
rect 29256 88 29272 152
rect 29336 88 29352 152
rect 29416 88 29424 152
rect 29104 72 29424 88
rect 29104 8 29112 72
rect 29176 8 29192 72
rect 29256 8 29272 72
rect 29336 8 29352 72
rect 29416 8 29424 72
rect 29104 0 29424 8
rect 41368 3992 45368 41400
rect 41368 3928 41376 3992
rect 41440 3928 41456 3992
rect 41520 3928 41536 3992
rect 41600 3928 41616 3992
rect 41680 3928 41696 3992
rect 41760 3928 41776 3992
rect 41840 3928 41856 3992
rect 41920 3928 41936 3992
rect 42000 3928 42016 3992
rect 42080 3928 42096 3992
rect 42160 3928 42176 3992
rect 42240 3928 42256 3992
rect 42320 3928 42336 3992
rect 42400 3928 42416 3992
rect 42480 3928 42496 3992
rect 42560 3928 42576 3992
rect 42640 3928 42656 3992
rect 42720 3928 42736 3992
rect 42800 3928 42816 3992
rect 42880 3928 42896 3992
rect 42960 3928 42976 3992
rect 43040 3928 43056 3992
rect 43120 3928 43136 3992
rect 43200 3928 43216 3992
rect 43280 3928 43296 3992
rect 43360 3928 43376 3992
rect 43440 3928 43456 3992
rect 43520 3928 43536 3992
rect 43600 3928 43616 3992
rect 43680 3928 43696 3992
rect 43760 3928 43776 3992
rect 43840 3928 43856 3992
rect 43920 3928 43936 3992
rect 44000 3928 44016 3992
rect 44080 3928 44096 3992
rect 44160 3928 44176 3992
rect 44240 3928 44256 3992
rect 44320 3928 44336 3992
rect 44400 3928 44416 3992
rect 44480 3928 44496 3992
rect 44560 3928 44576 3992
rect 44640 3928 44656 3992
rect 44720 3928 44736 3992
rect 44800 3928 44816 3992
rect 44880 3928 44896 3992
rect 44960 3928 44976 3992
rect 45040 3928 45056 3992
rect 45120 3928 45136 3992
rect 45200 3928 45216 3992
rect 45280 3928 45296 3992
rect 45360 3928 45368 3992
rect 41368 3912 45368 3928
rect 41368 3848 41376 3912
rect 41440 3848 41456 3912
rect 41520 3848 41536 3912
rect 41600 3848 41616 3912
rect 41680 3848 41696 3912
rect 41760 3848 41776 3912
rect 41840 3848 41856 3912
rect 41920 3848 41936 3912
rect 42000 3848 42016 3912
rect 42080 3848 42096 3912
rect 42160 3848 42176 3912
rect 42240 3848 42256 3912
rect 42320 3848 42336 3912
rect 42400 3848 42416 3912
rect 42480 3848 42496 3912
rect 42560 3848 42576 3912
rect 42640 3848 42656 3912
rect 42720 3848 42736 3912
rect 42800 3848 42816 3912
rect 42880 3848 42896 3912
rect 42960 3848 42976 3912
rect 43040 3848 43056 3912
rect 43120 3848 43136 3912
rect 43200 3848 43216 3912
rect 43280 3848 43296 3912
rect 43360 3848 43376 3912
rect 43440 3848 43456 3912
rect 43520 3848 43536 3912
rect 43600 3848 43616 3912
rect 43680 3848 43696 3912
rect 43760 3848 43776 3912
rect 43840 3848 43856 3912
rect 43920 3848 43936 3912
rect 44000 3848 44016 3912
rect 44080 3848 44096 3912
rect 44160 3848 44176 3912
rect 44240 3848 44256 3912
rect 44320 3848 44336 3912
rect 44400 3848 44416 3912
rect 44480 3848 44496 3912
rect 44560 3848 44576 3912
rect 44640 3848 44656 3912
rect 44720 3848 44736 3912
rect 44800 3848 44816 3912
rect 44880 3848 44896 3912
rect 44960 3848 44976 3912
rect 45040 3848 45056 3912
rect 45120 3848 45136 3912
rect 45200 3848 45216 3912
rect 45280 3848 45296 3912
rect 45360 3848 45368 3912
rect 41368 3832 45368 3848
rect 41368 3768 41376 3832
rect 41440 3768 41456 3832
rect 41520 3768 41536 3832
rect 41600 3768 41616 3832
rect 41680 3768 41696 3832
rect 41760 3768 41776 3832
rect 41840 3768 41856 3832
rect 41920 3768 41936 3832
rect 42000 3768 42016 3832
rect 42080 3768 42096 3832
rect 42160 3768 42176 3832
rect 42240 3768 42256 3832
rect 42320 3768 42336 3832
rect 42400 3768 42416 3832
rect 42480 3768 42496 3832
rect 42560 3768 42576 3832
rect 42640 3768 42656 3832
rect 42720 3768 42736 3832
rect 42800 3768 42816 3832
rect 42880 3768 42896 3832
rect 42960 3768 42976 3832
rect 43040 3768 43056 3832
rect 43120 3768 43136 3832
rect 43200 3768 43216 3832
rect 43280 3768 43296 3832
rect 43360 3768 43376 3832
rect 43440 3768 43456 3832
rect 43520 3768 43536 3832
rect 43600 3768 43616 3832
rect 43680 3768 43696 3832
rect 43760 3768 43776 3832
rect 43840 3768 43856 3832
rect 43920 3768 43936 3832
rect 44000 3768 44016 3832
rect 44080 3768 44096 3832
rect 44160 3768 44176 3832
rect 44240 3768 44256 3832
rect 44320 3768 44336 3832
rect 44400 3768 44416 3832
rect 44480 3768 44496 3832
rect 44560 3768 44576 3832
rect 44640 3768 44656 3832
rect 44720 3768 44736 3832
rect 44800 3768 44816 3832
rect 44880 3768 44896 3832
rect 44960 3768 44976 3832
rect 45040 3768 45056 3832
rect 45120 3768 45136 3832
rect 45200 3768 45216 3832
rect 45280 3768 45296 3832
rect 45360 3768 45368 3832
rect 41368 3752 45368 3768
rect 41368 3688 41376 3752
rect 41440 3688 41456 3752
rect 41520 3688 41536 3752
rect 41600 3688 41616 3752
rect 41680 3688 41696 3752
rect 41760 3688 41776 3752
rect 41840 3688 41856 3752
rect 41920 3688 41936 3752
rect 42000 3688 42016 3752
rect 42080 3688 42096 3752
rect 42160 3688 42176 3752
rect 42240 3688 42256 3752
rect 42320 3688 42336 3752
rect 42400 3688 42416 3752
rect 42480 3688 42496 3752
rect 42560 3688 42576 3752
rect 42640 3688 42656 3752
rect 42720 3688 42736 3752
rect 42800 3688 42816 3752
rect 42880 3688 42896 3752
rect 42960 3688 42976 3752
rect 43040 3688 43056 3752
rect 43120 3688 43136 3752
rect 43200 3688 43216 3752
rect 43280 3688 43296 3752
rect 43360 3688 43376 3752
rect 43440 3688 43456 3752
rect 43520 3688 43536 3752
rect 43600 3688 43616 3752
rect 43680 3688 43696 3752
rect 43760 3688 43776 3752
rect 43840 3688 43856 3752
rect 43920 3688 43936 3752
rect 44000 3688 44016 3752
rect 44080 3688 44096 3752
rect 44160 3688 44176 3752
rect 44240 3688 44256 3752
rect 44320 3688 44336 3752
rect 44400 3688 44416 3752
rect 44480 3688 44496 3752
rect 44560 3688 44576 3752
rect 44640 3688 44656 3752
rect 44720 3688 44736 3752
rect 44800 3688 44816 3752
rect 44880 3688 44896 3752
rect 44960 3688 44976 3752
rect 45040 3688 45056 3752
rect 45120 3688 45136 3752
rect 45200 3688 45216 3752
rect 45280 3688 45296 3752
rect 45360 3688 45368 3752
rect 41368 3672 45368 3688
rect 41368 3608 41376 3672
rect 41440 3608 41456 3672
rect 41520 3608 41536 3672
rect 41600 3608 41616 3672
rect 41680 3608 41696 3672
rect 41760 3608 41776 3672
rect 41840 3608 41856 3672
rect 41920 3608 41936 3672
rect 42000 3608 42016 3672
rect 42080 3608 42096 3672
rect 42160 3608 42176 3672
rect 42240 3608 42256 3672
rect 42320 3608 42336 3672
rect 42400 3608 42416 3672
rect 42480 3608 42496 3672
rect 42560 3608 42576 3672
rect 42640 3608 42656 3672
rect 42720 3608 42736 3672
rect 42800 3608 42816 3672
rect 42880 3608 42896 3672
rect 42960 3608 42976 3672
rect 43040 3608 43056 3672
rect 43120 3608 43136 3672
rect 43200 3608 43216 3672
rect 43280 3608 43296 3672
rect 43360 3608 43376 3672
rect 43440 3608 43456 3672
rect 43520 3608 43536 3672
rect 43600 3608 43616 3672
rect 43680 3608 43696 3672
rect 43760 3608 43776 3672
rect 43840 3608 43856 3672
rect 43920 3608 43936 3672
rect 44000 3608 44016 3672
rect 44080 3608 44096 3672
rect 44160 3608 44176 3672
rect 44240 3608 44256 3672
rect 44320 3608 44336 3672
rect 44400 3608 44416 3672
rect 44480 3608 44496 3672
rect 44560 3608 44576 3672
rect 44640 3608 44656 3672
rect 44720 3608 44736 3672
rect 44800 3608 44816 3672
rect 44880 3608 44896 3672
rect 44960 3608 44976 3672
rect 45040 3608 45056 3672
rect 45120 3608 45136 3672
rect 45200 3608 45216 3672
rect 45280 3608 45296 3672
rect 45360 3608 45368 3672
rect 41368 3592 45368 3608
rect 41368 3528 41376 3592
rect 41440 3528 41456 3592
rect 41520 3528 41536 3592
rect 41600 3528 41616 3592
rect 41680 3528 41696 3592
rect 41760 3528 41776 3592
rect 41840 3528 41856 3592
rect 41920 3528 41936 3592
rect 42000 3528 42016 3592
rect 42080 3528 42096 3592
rect 42160 3528 42176 3592
rect 42240 3528 42256 3592
rect 42320 3528 42336 3592
rect 42400 3528 42416 3592
rect 42480 3528 42496 3592
rect 42560 3528 42576 3592
rect 42640 3528 42656 3592
rect 42720 3528 42736 3592
rect 42800 3528 42816 3592
rect 42880 3528 42896 3592
rect 42960 3528 42976 3592
rect 43040 3528 43056 3592
rect 43120 3528 43136 3592
rect 43200 3528 43216 3592
rect 43280 3528 43296 3592
rect 43360 3528 43376 3592
rect 43440 3528 43456 3592
rect 43520 3528 43536 3592
rect 43600 3528 43616 3592
rect 43680 3528 43696 3592
rect 43760 3528 43776 3592
rect 43840 3528 43856 3592
rect 43920 3528 43936 3592
rect 44000 3528 44016 3592
rect 44080 3528 44096 3592
rect 44160 3528 44176 3592
rect 44240 3528 44256 3592
rect 44320 3528 44336 3592
rect 44400 3528 44416 3592
rect 44480 3528 44496 3592
rect 44560 3528 44576 3592
rect 44640 3528 44656 3592
rect 44720 3528 44736 3592
rect 44800 3528 44816 3592
rect 44880 3528 44896 3592
rect 44960 3528 44976 3592
rect 45040 3528 45056 3592
rect 45120 3528 45136 3592
rect 45200 3528 45216 3592
rect 45280 3528 45296 3592
rect 45360 3528 45368 3592
rect 41368 3512 45368 3528
rect 41368 3448 41376 3512
rect 41440 3448 41456 3512
rect 41520 3448 41536 3512
rect 41600 3448 41616 3512
rect 41680 3448 41696 3512
rect 41760 3448 41776 3512
rect 41840 3448 41856 3512
rect 41920 3448 41936 3512
rect 42000 3448 42016 3512
rect 42080 3448 42096 3512
rect 42160 3448 42176 3512
rect 42240 3448 42256 3512
rect 42320 3448 42336 3512
rect 42400 3448 42416 3512
rect 42480 3448 42496 3512
rect 42560 3448 42576 3512
rect 42640 3448 42656 3512
rect 42720 3448 42736 3512
rect 42800 3448 42816 3512
rect 42880 3448 42896 3512
rect 42960 3448 42976 3512
rect 43040 3448 43056 3512
rect 43120 3448 43136 3512
rect 43200 3448 43216 3512
rect 43280 3448 43296 3512
rect 43360 3448 43376 3512
rect 43440 3448 43456 3512
rect 43520 3448 43536 3512
rect 43600 3448 43616 3512
rect 43680 3448 43696 3512
rect 43760 3448 43776 3512
rect 43840 3448 43856 3512
rect 43920 3448 43936 3512
rect 44000 3448 44016 3512
rect 44080 3448 44096 3512
rect 44160 3448 44176 3512
rect 44240 3448 44256 3512
rect 44320 3448 44336 3512
rect 44400 3448 44416 3512
rect 44480 3448 44496 3512
rect 44560 3448 44576 3512
rect 44640 3448 44656 3512
rect 44720 3448 44736 3512
rect 44800 3448 44816 3512
rect 44880 3448 44896 3512
rect 44960 3448 44976 3512
rect 45040 3448 45056 3512
rect 45120 3448 45136 3512
rect 45200 3448 45216 3512
rect 45280 3448 45296 3512
rect 45360 3448 45368 3512
rect 41368 3432 45368 3448
rect 41368 3368 41376 3432
rect 41440 3368 41456 3432
rect 41520 3368 41536 3432
rect 41600 3368 41616 3432
rect 41680 3368 41696 3432
rect 41760 3368 41776 3432
rect 41840 3368 41856 3432
rect 41920 3368 41936 3432
rect 42000 3368 42016 3432
rect 42080 3368 42096 3432
rect 42160 3368 42176 3432
rect 42240 3368 42256 3432
rect 42320 3368 42336 3432
rect 42400 3368 42416 3432
rect 42480 3368 42496 3432
rect 42560 3368 42576 3432
rect 42640 3368 42656 3432
rect 42720 3368 42736 3432
rect 42800 3368 42816 3432
rect 42880 3368 42896 3432
rect 42960 3368 42976 3432
rect 43040 3368 43056 3432
rect 43120 3368 43136 3432
rect 43200 3368 43216 3432
rect 43280 3368 43296 3432
rect 43360 3368 43376 3432
rect 43440 3368 43456 3432
rect 43520 3368 43536 3432
rect 43600 3368 43616 3432
rect 43680 3368 43696 3432
rect 43760 3368 43776 3432
rect 43840 3368 43856 3432
rect 43920 3368 43936 3432
rect 44000 3368 44016 3432
rect 44080 3368 44096 3432
rect 44160 3368 44176 3432
rect 44240 3368 44256 3432
rect 44320 3368 44336 3432
rect 44400 3368 44416 3432
rect 44480 3368 44496 3432
rect 44560 3368 44576 3432
rect 44640 3368 44656 3432
rect 44720 3368 44736 3432
rect 44800 3368 44816 3432
rect 44880 3368 44896 3432
rect 44960 3368 44976 3432
rect 45040 3368 45056 3432
rect 45120 3368 45136 3432
rect 45200 3368 45216 3432
rect 45280 3368 45296 3432
rect 45360 3368 45368 3432
rect 41368 3352 45368 3368
rect 41368 3288 41376 3352
rect 41440 3288 41456 3352
rect 41520 3288 41536 3352
rect 41600 3288 41616 3352
rect 41680 3288 41696 3352
rect 41760 3288 41776 3352
rect 41840 3288 41856 3352
rect 41920 3288 41936 3352
rect 42000 3288 42016 3352
rect 42080 3288 42096 3352
rect 42160 3288 42176 3352
rect 42240 3288 42256 3352
rect 42320 3288 42336 3352
rect 42400 3288 42416 3352
rect 42480 3288 42496 3352
rect 42560 3288 42576 3352
rect 42640 3288 42656 3352
rect 42720 3288 42736 3352
rect 42800 3288 42816 3352
rect 42880 3288 42896 3352
rect 42960 3288 42976 3352
rect 43040 3288 43056 3352
rect 43120 3288 43136 3352
rect 43200 3288 43216 3352
rect 43280 3288 43296 3352
rect 43360 3288 43376 3352
rect 43440 3288 43456 3352
rect 43520 3288 43536 3352
rect 43600 3288 43616 3352
rect 43680 3288 43696 3352
rect 43760 3288 43776 3352
rect 43840 3288 43856 3352
rect 43920 3288 43936 3352
rect 44000 3288 44016 3352
rect 44080 3288 44096 3352
rect 44160 3288 44176 3352
rect 44240 3288 44256 3352
rect 44320 3288 44336 3352
rect 44400 3288 44416 3352
rect 44480 3288 44496 3352
rect 44560 3288 44576 3352
rect 44640 3288 44656 3352
rect 44720 3288 44736 3352
rect 44800 3288 44816 3352
rect 44880 3288 44896 3352
rect 44960 3288 44976 3352
rect 45040 3288 45056 3352
rect 45120 3288 45136 3352
rect 45200 3288 45216 3352
rect 45280 3288 45296 3352
rect 45360 3288 45368 3352
rect 41368 3272 45368 3288
rect 41368 3208 41376 3272
rect 41440 3208 41456 3272
rect 41520 3208 41536 3272
rect 41600 3208 41616 3272
rect 41680 3208 41696 3272
rect 41760 3208 41776 3272
rect 41840 3208 41856 3272
rect 41920 3208 41936 3272
rect 42000 3208 42016 3272
rect 42080 3208 42096 3272
rect 42160 3208 42176 3272
rect 42240 3208 42256 3272
rect 42320 3208 42336 3272
rect 42400 3208 42416 3272
rect 42480 3208 42496 3272
rect 42560 3208 42576 3272
rect 42640 3208 42656 3272
rect 42720 3208 42736 3272
rect 42800 3208 42816 3272
rect 42880 3208 42896 3272
rect 42960 3208 42976 3272
rect 43040 3208 43056 3272
rect 43120 3208 43136 3272
rect 43200 3208 43216 3272
rect 43280 3208 43296 3272
rect 43360 3208 43376 3272
rect 43440 3208 43456 3272
rect 43520 3208 43536 3272
rect 43600 3208 43616 3272
rect 43680 3208 43696 3272
rect 43760 3208 43776 3272
rect 43840 3208 43856 3272
rect 43920 3208 43936 3272
rect 44000 3208 44016 3272
rect 44080 3208 44096 3272
rect 44160 3208 44176 3272
rect 44240 3208 44256 3272
rect 44320 3208 44336 3272
rect 44400 3208 44416 3272
rect 44480 3208 44496 3272
rect 44560 3208 44576 3272
rect 44640 3208 44656 3272
rect 44720 3208 44736 3272
rect 44800 3208 44816 3272
rect 44880 3208 44896 3272
rect 44960 3208 44976 3272
rect 45040 3208 45056 3272
rect 45120 3208 45136 3272
rect 45200 3208 45216 3272
rect 45280 3208 45296 3272
rect 45360 3208 45368 3272
rect 41368 3192 45368 3208
rect 41368 3128 41376 3192
rect 41440 3128 41456 3192
rect 41520 3128 41536 3192
rect 41600 3128 41616 3192
rect 41680 3128 41696 3192
rect 41760 3128 41776 3192
rect 41840 3128 41856 3192
rect 41920 3128 41936 3192
rect 42000 3128 42016 3192
rect 42080 3128 42096 3192
rect 42160 3128 42176 3192
rect 42240 3128 42256 3192
rect 42320 3128 42336 3192
rect 42400 3128 42416 3192
rect 42480 3128 42496 3192
rect 42560 3128 42576 3192
rect 42640 3128 42656 3192
rect 42720 3128 42736 3192
rect 42800 3128 42816 3192
rect 42880 3128 42896 3192
rect 42960 3128 42976 3192
rect 43040 3128 43056 3192
rect 43120 3128 43136 3192
rect 43200 3128 43216 3192
rect 43280 3128 43296 3192
rect 43360 3128 43376 3192
rect 43440 3128 43456 3192
rect 43520 3128 43536 3192
rect 43600 3128 43616 3192
rect 43680 3128 43696 3192
rect 43760 3128 43776 3192
rect 43840 3128 43856 3192
rect 43920 3128 43936 3192
rect 44000 3128 44016 3192
rect 44080 3128 44096 3192
rect 44160 3128 44176 3192
rect 44240 3128 44256 3192
rect 44320 3128 44336 3192
rect 44400 3128 44416 3192
rect 44480 3128 44496 3192
rect 44560 3128 44576 3192
rect 44640 3128 44656 3192
rect 44720 3128 44736 3192
rect 44800 3128 44816 3192
rect 44880 3128 44896 3192
rect 44960 3128 44976 3192
rect 45040 3128 45056 3192
rect 45120 3128 45136 3192
rect 45200 3128 45216 3192
rect 45280 3128 45296 3192
rect 45360 3128 45368 3192
rect 41368 3112 45368 3128
rect 41368 3048 41376 3112
rect 41440 3048 41456 3112
rect 41520 3048 41536 3112
rect 41600 3048 41616 3112
rect 41680 3048 41696 3112
rect 41760 3048 41776 3112
rect 41840 3048 41856 3112
rect 41920 3048 41936 3112
rect 42000 3048 42016 3112
rect 42080 3048 42096 3112
rect 42160 3048 42176 3112
rect 42240 3048 42256 3112
rect 42320 3048 42336 3112
rect 42400 3048 42416 3112
rect 42480 3048 42496 3112
rect 42560 3048 42576 3112
rect 42640 3048 42656 3112
rect 42720 3048 42736 3112
rect 42800 3048 42816 3112
rect 42880 3048 42896 3112
rect 42960 3048 42976 3112
rect 43040 3048 43056 3112
rect 43120 3048 43136 3112
rect 43200 3048 43216 3112
rect 43280 3048 43296 3112
rect 43360 3048 43376 3112
rect 43440 3048 43456 3112
rect 43520 3048 43536 3112
rect 43600 3048 43616 3112
rect 43680 3048 43696 3112
rect 43760 3048 43776 3112
rect 43840 3048 43856 3112
rect 43920 3048 43936 3112
rect 44000 3048 44016 3112
rect 44080 3048 44096 3112
rect 44160 3048 44176 3112
rect 44240 3048 44256 3112
rect 44320 3048 44336 3112
rect 44400 3048 44416 3112
rect 44480 3048 44496 3112
rect 44560 3048 44576 3112
rect 44640 3048 44656 3112
rect 44720 3048 44736 3112
rect 44800 3048 44816 3112
rect 44880 3048 44896 3112
rect 44960 3048 44976 3112
rect 45040 3048 45056 3112
rect 45120 3048 45136 3112
rect 45200 3048 45216 3112
rect 45280 3048 45296 3112
rect 45360 3048 45368 3112
rect 41368 3032 45368 3048
rect 41368 2968 41376 3032
rect 41440 2968 41456 3032
rect 41520 2968 41536 3032
rect 41600 2968 41616 3032
rect 41680 2968 41696 3032
rect 41760 2968 41776 3032
rect 41840 2968 41856 3032
rect 41920 2968 41936 3032
rect 42000 2968 42016 3032
rect 42080 2968 42096 3032
rect 42160 2968 42176 3032
rect 42240 2968 42256 3032
rect 42320 2968 42336 3032
rect 42400 2968 42416 3032
rect 42480 2968 42496 3032
rect 42560 2968 42576 3032
rect 42640 2968 42656 3032
rect 42720 2968 42736 3032
rect 42800 2968 42816 3032
rect 42880 2968 42896 3032
rect 42960 2968 42976 3032
rect 43040 2968 43056 3032
rect 43120 2968 43136 3032
rect 43200 2968 43216 3032
rect 43280 2968 43296 3032
rect 43360 2968 43376 3032
rect 43440 2968 43456 3032
rect 43520 2968 43536 3032
rect 43600 2968 43616 3032
rect 43680 2968 43696 3032
rect 43760 2968 43776 3032
rect 43840 2968 43856 3032
rect 43920 2968 43936 3032
rect 44000 2968 44016 3032
rect 44080 2968 44096 3032
rect 44160 2968 44176 3032
rect 44240 2968 44256 3032
rect 44320 2968 44336 3032
rect 44400 2968 44416 3032
rect 44480 2968 44496 3032
rect 44560 2968 44576 3032
rect 44640 2968 44656 3032
rect 44720 2968 44736 3032
rect 44800 2968 44816 3032
rect 44880 2968 44896 3032
rect 44960 2968 44976 3032
rect 45040 2968 45056 3032
rect 45120 2968 45136 3032
rect 45200 2968 45216 3032
rect 45280 2968 45296 3032
rect 45360 2968 45368 3032
rect 41368 2952 45368 2968
rect 41368 2888 41376 2952
rect 41440 2888 41456 2952
rect 41520 2888 41536 2952
rect 41600 2888 41616 2952
rect 41680 2888 41696 2952
rect 41760 2888 41776 2952
rect 41840 2888 41856 2952
rect 41920 2888 41936 2952
rect 42000 2888 42016 2952
rect 42080 2888 42096 2952
rect 42160 2888 42176 2952
rect 42240 2888 42256 2952
rect 42320 2888 42336 2952
rect 42400 2888 42416 2952
rect 42480 2888 42496 2952
rect 42560 2888 42576 2952
rect 42640 2888 42656 2952
rect 42720 2888 42736 2952
rect 42800 2888 42816 2952
rect 42880 2888 42896 2952
rect 42960 2888 42976 2952
rect 43040 2888 43056 2952
rect 43120 2888 43136 2952
rect 43200 2888 43216 2952
rect 43280 2888 43296 2952
rect 43360 2888 43376 2952
rect 43440 2888 43456 2952
rect 43520 2888 43536 2952
rect 43600 2888 43616 2952
rect 43680 2888 43696 2952
rect 43760 2888 43776 2952
rect 43840 2888 43856 2952
rect 43920 2888 43936 2952
rect 44000 2888 44016 2952
rect 44080 2888 44096 2952
rect 44160 2888 44176 2952
rect 44240 2888 44256 2952
rect 44320 2888 44336 2952
rect 44400 2888 44416 2952
rect 44480 2888 44496 2952
rect 44560 2888 44576 2952
rect 44640 2888 44656 2952
rect 44720 2888 44736 2952
rect 44800 2888 44816 2952
rect 44880 2888 44896 2952
rect 44960 2888 44976 2952
rect 45040 2888 45056 2952
rect 45120 2888 45136 2952
rect 45200 2888 45216 2952
rect 45280 2888 45296 2952
rect 45360 2888 45368 2952
rect 41368 2872 45368 2888
rect 41368 2808 41376 2872
rect 41440 2808 41456 2872
rect 41520 2808 41536 2872
rect 41600 2808 41616 2872
rect 41680 2808 41696 2872
rect 41760 2808 41776 2872
rect 41840 2808 41856 2872
rect 41920 2808 41936 2872
rect 42000 2808 42016 2872
rect 42080 2808 42096 2872
rect 42160 2808 42176 2872
rect 42240 2808 42256 2872
rect 42320 2808 42336 2872
rect 42400 2808 42416 2872
rect 42480 2808 42496 2872
rect 42560 2808 42576 2872
rect 42640 2808 42656 2872
rect 42720 2808 42736 2872
rect 42800 2808 42816 2872
rect 42880 2808 42896 2872
rect 42960 2808 42976 2872
rect 43040 2808 43056 2872
rect 43120 2808 43136 2872
rect 43200 2808 43216 2872
rect 43280 2808 43296 2872
rect 43360 2808 43376 2872
rect 43440 2808 43456 2872
rect 43520 2808 43536 2872
rect 43600 2808 43616 2872
rect 43680 2808 43696 2872
rect 43760 2808 43776 2872
rect 43840 2808 43856 2872
rect 43920 2808 43936 2872
rect 44000 2808 44016 2872
rect 44080 2808 44096 2872
rect 44160 2808 44176 2872
rect 44240 2808 44256 2872
rect 44320 2808 44336 2872
rect 44400 2808 44416 2872
rect 44480 2808 44496 2872
rect 44560 2808 44576 2872
rect 44640 2808 44656 2872
rect 44720 2808 44736 2872
rect 44800 2808 44816 2872
rect 44880 2808 44896 2872
rect 44960 2808 44976 2872
rect 45040 2808 45056 2872
rect 45120 2808 45136 2872
rect 45200 2808 45216 2872
rect 45280 2808 45296 2872
rect 45360 2808 45368 2872
rect 41368 2792 45368 2808
rect 41368 2728 41376 2792
rect 41440 2728 41456 2792
rect 41520 2728 41536 2792
rect 41600 2728 41616 2792
rect 41680 2728 41696 2792
rect 41760 2728 41776 2792
rect 41840 2728 41856 2792
rect 41920 2728 41936 2792
rect 42000 2728 42016 2792
rect 42080 2728 42096 2792
rect 42160 2728 42176 2792
rect 42240 2728 42256 2792
rect 42320 2728 42336 2792
rect 42400 2728 42416 2792
rect 42480 2728 42496 2792
rect 42560 2728 42576 2792
rect 42640 2728 42656 2792
rect 42720 2728 42736 2792
rect 42800 2728 42816 2792
rect 42880 2728 42896 2792
rect 42960 2728 42976 2792
rect 43040 2728 43056 2792
rect 43120 2728 43136 2792
rect 43200 2728 43216 2792
rect 43280 2728 43296 2792
rect 43360 2728 43376 2792
rect 43440 2728 43456 2792
rect 43520 2728 43536 2792
rect 43600 2728 43616 2792
rect 43680 2728 43696 2792
rect 43760 2728 43776 2792
rect 43840 2728 43856 2792
rect 43920 2728 43936 2792
rect 44000 2728 44016 2792
rect 44080 2728 44096 2792
rect 44160 2728 44176 2792
rect 44240 2728 44256 2792
rect 44320 2728 44336 2792
rect 44400 2728 44416 2792
rect 44480 2728 44496 2792
rect 44560 2728 44576 2792
rect 44640 2728 44656 2792
rect 44720 2728 44736 2792
rect 44800 2728 44816 2792
rect 44880 2728 44896 2792
rect 44960 2728 44976 2792
rect 45040 2728 45056 2792
rect 45120 2728 45136 2792
rect 45200 2728 45216 2792
rect 45280 2728 45296 2792
rect 45360 2728 45368 2792
rect 41368 2712 45368 2728
rect 41368 2648 41376 2712
rect 41440 2648 41456 2712
rect 41520 2648 41536 2712
rect 41600 2648 41616 2712
rect 41680 2648 41696 2712
rect 41760 2648 41776 2712
rect 41840 2648 41856 2712
rect 41920 2648 41936 2712
rect 42000 2648 42016 2712
rect 42080 2648 42096 2712
rect 42160 2648 42176 2712
rect 42240 2648 42256 2712
rect 42320 2648 42336 2712
rect 42400 2648 42416 2712
rect 42480 2648 42496 2712
rect 42560 2648 42576 2712
rect 42640 2648 42656 2712
rect 42720 2648 42736 2712
rect 42800 2648 42816 2712
rect 42880 2648 42896 2712
rect 42960 2648 42976 2712
rect 43040 2648 43056 2712
rect 43120 2648 43136 2712
rect 43200 2648 43216 2712
rect 43280 2648 43296 2712
rect 43360 2648 43376 2712
rect 43440 2648 43456 2712
rect 43520 2648 43536 2712
rect 43600 2648 43616 2712
rect 43680 2648 43696 2712
rect 43760 2648 43776 2712
rect 43840 2648 43856 2712
rect 43920 2648 43936 2712
rect 44000 2648 44016 2712
rect 44080 2648 44096 2712
rect 44160 2648 44176 2712
rect 44240 2648 44256 2712
rect 44320 2648 44336 2712
rect 44400 2648 44416 2712
rect 44480 2648 44496 2712
rect 44560 2648 44576 2712
rect 44640 2648 44656 2712
rect 44720 2648 44736 2712
rect 44800 2648 44816 2712
rect 44880 2648 44896 2712
rect 44960 2648 44976 2712
rect 45040 2648 45056 2712
rect 45120 2648 45136 2712
rect 45200 2648 45216 2712
rect 45280 2648 45296 2712
rect 45360 2648 45368 2712
rect 41368 2632 45368 2648
rect 41368 2568 41376 2632
rect 41440 2568 41456 2632
rect 41520 2568 41536 2632
rect 41600 2568 41616 2632
rect 41680 2568 41696 2632
rect 41760 2568 41776 2632
rect 41840 2568 41856 2632
rect 41920 2568 41936 2632
rect 42000 2568 42016 2632
rect 42080 2568 42096 2632
rect 42160 2568 42176 2632
rect 42240 2568 42256 2632
rect 42320 2568 42336 2632
rect 42400 2568 42416 2632
rect 42480 2568 42496 2632
rect 42560 2568 42576 2632
rect 42640 2568 42656 2632
rect 42720 2568 42736 2632
rect 42800 2568 42816 2632
rect 42880 2568 42896 2632
rect 42960 2568 42976 2632
rect 43040 2568 43056 2632
rect 43120 2568 43136 2632
rect 43200 2568 43216 2632
rect 43280 2568 43296 2632
rect 43360 2568 43376 2632
rect 43440 2568 43456 2632
rect 43520 2568 43536 2632
rect 43600 2568 43616 2632
rect 43680 2568 43696 2632
rect 43760 2568 43776 2632
rect 43840 2568 43856 2632
rect 43920 2568 43936 2632
rect 44000 2568 44016 2632
rect 44080 2568 44096 2632
rect 44160 2568 44176 2632
rect 44240 2568 44256 2632
rect 44320 2568 44336 2632
rect 44400 2568 44416 2632
rect 44480 2568 44496 2632
rect 44560 2568 44576 2632
rect 44640 2568 44656 2632
rect 44720 2568 44736 2632
rect 44800 2568 44816 2632
rect 44880 2568 44896 2632
rect 44960 2568 44976 2632
rect 45040 2568 45056 2632
rect 45120 2568 45136 2632
rect 45200 2568 45216 2632
rect 45280 2568 45296 2632
rect 45360 2568 45368 2632
rect 41368 2552 45368 2568
rect 41368 2488 41376 2552
rect 41440 2488 41456 2552
rect 41520 2488 41536 2552
rect 41600 2488 41616 2552
rect 41680 2488 41696 2552
rect 41760 2488 41776 2552
rect 41840 2488 41856 2552
rect 41920 2488 41936 2552
rect 42000 2488 42016 2552
rect 42080 2488 42096 2552
rect 42160 2488 42176 2552
rect 42240 2488 42256 2552
rect 42320 2488 42336 2552
rect 42400 2488 42416 2552
rect 42480 2488 42496 2552
rect 42560 2488 42576 2552
rect 42640 2488 42656 2552
rect 42720 2488 42736 2552
rect 42800 2488 42816 2552
rect 42880 2488 42896 2552
rect 42960 2488 42976 2552
rect 43040 2488 43056 2552
rect 43120 2488 43136 2552
rect 43200 2488 43216 2552
rect 43280 2488 43296 2552
rect 43360 2488 43376 2552
rect 43440 2488 43456 2552
rect 43520 2488 43536 2552
rect 43600 2488 43616 2552
rect 43680 2488 43696 2552
rect 43760 2488 43776 2552
rect 43840 2488 43856 2552
rect 43920 2488 43936 2552
rect 44000 2488 44016 2552
rect 44080 2488 44096 2552
rect 44160 2488 44176 2552
rect 44240 2488 44256 2552
rect 44320 2488 44336 2552
rect 44400 2488 44416 2552
rect 44480 2488 44496 2552
rect 44560 2488 44576 2552
rect 44640 2488 44656 2552
rect 44720 2488 44736 2552
rect 44800 2488 44816 2552
rect 44880 2488 44896 2552
rect 44960 2488 44976 2552
rect 45040 2488 45056 2552
rect 45120 2488 45136 2552
rect 45200 2488 45216 2552
rect 45280 2488 45296 2552
rect 45360 2488 45368 2552
rect 41368 2472 45368 2488
rect 41368 2408 41376 2472
rect 41440 2408 41456 2472
rect 41520 2408 41536 2472
rect 41600 2408 41616 2472
rect 41680 2408 41696 2472
rect 41760 2408 41776 2472
rect 41840 2408 41856 2472
rect 41920 2408 41936 2472
rect 42000 2408 42016 2472
rect 42080 2408 42096 2472
rect 42160 2408 42176 2472
rect 42240 2408 42256 2472
rect 42320 2408 42336 2472
rect 42400 2408 42416 2472
rect 42480 2408 42496 2472
rect 42560 2408 42576 2472
rect 42640 2408 42656 2472
rect 42720 2408 42736 2472
rect 42800 2408 42816 2472
rect 42880 2408 42896 2472
rect 42960 2408 42976 2472
rect 43040 2408 43056 2472
rect 43120 2408 43136 2472
rect 43200 2408 43216 2472
rect 43280 2408 43296 2472
rect 43360 2408 43376 2472
rect 43440 2408 43456 2472
rect 43520 2408 43536 2472
rect 43600 2408 43616 2472
rect 43680 2408 43696 2472
rect 43760 2408 43776 2472
rect 43840 2408 43856 2472
rect 43920 2408 43936 2472
rect 44000 2408 44016 2472
rect 44080 2408 44096 2472
rect 44160 2408 44176 2472
rect 44240 2408 44256 2472
rect 44320 2408 44336 2472
rect 44400 2408 44416 2472
rect 44480 2408 44496 2472
rect 44560 2408 44576 2472
rect 44640 2408 44656 2472
rect 44720 2408 44736 2472
rect 44800 2408 44816 2472
rect 44880 2408 44896 2472
rect 44960 2408 44976 2472
rect 45040 2408 45056 2472
rect 45120 2408 45136 2472
rect 45200 2408 45216 2472
rect 45280 2408 45296 2472
rect 45360 2408 45368 2472
rect 41368 2392 45368 2408
rect 41368 2328 41376 2392
rect 41440 2328 41456 2392
rect 41520 2328 41536 2392
rect 41600 2328 41616 2392
rect 41680 2328 41696 2392
rect 41760 2328 41776 2392
rect 41840 2328 41856 2392
rect 41920 2328 41936 2392
rect 42000 2328 42016 2392
rect 42080 2328 42096 2392
rect 42160 2328 42176 2392
rect 42240 2328 42256 2392
rect 42320 2328 42336 2392
rect 42400 2328 42416 2392
rect 42480 2328 42496 2392
rect 42560 2328 42576 2392
rect 42640 2328 42656 2392
rect 42720 2328 42736 2392
rect 42800 2328 42816 2392
rect 42880 2328 42896 2392
rect 42960 2328 42976 2392
rect 43040 2328 43056 2392
rect 43120 2328 43136 2392
rect 43200 2328 43216 2392
rect 43280 2328 43296 2392
rect 43360 2328 43376 2392
rect 43440 2328 43456 2392
rect 43520 2328 43536 2392
rect 43600 2328 43616 2392
rect 43680 2328 43696 2392
rect 43760 2328 43776 2392
rect 43840 2328 43856 2392
rect 43920 2328 43936 2392
rect 44000 2328 44016 2392
rect 44080 2328 44096 2392
rect 44160 2328 44176 2392
rect 44240 2328 44256 2392
rect 44320 2328 44336 2392
rect 44400 2328 44416 2392
rect 44480 2328 44496 2392
rect 44560 2328 44576 2392
rect 44640 2328 44656 2392
rect 44720 2328 44736 2392
rect 44800 2328 44816 2392
rect 44880 2328 44896 2392
rect 44960 2328 44976 2392
rect 45040 2328 45056 2392
rect 45120 2328 45136 2392
rect 45200 2328 45216 2392
rect 45280 2328 45296 2392
rect 45360 2328 45368 2392
rect 41368 2312 45368 2328
rect 41368 2248 41376 2312
rect 41440 2248 41456 2312
rect 41520 2248 41536 2312
rect 41600 2248 41616 2312
rect 41680 2248 41696 2312
rect 41760 2248 41776 2312
rect 41840 2248 41856 2312
rect 41920 2248 41936 2312
rect 42000 2248 42016 2312
rect 42080 2248 42096 2312
rect 42160 2248 42176 2312
rect 42240 2248 42256 2312
rect 42320 2248 42336 2312
rect 42400 2248 42416 2312
rect 42480 2248 42496 2312
rect 42560 2248 42576 2312
rect 42640 2248 42656 2312
rect 42720 2248 42736 2312
rect 42800 2248 42816 2312
rect 42880 2248 42896 2312
rect 42960 2248 42976 2312
rect 43040 2248 43056 2312
rect 43120 2248 43136 2312
rect 43200 2248 43216 2312
rect 43280 2248 43296 2312
rect 43360 2248 43376 2312
rect 43440 2248 43456 2312
rect 43520 2248 43536 2312
rect 43600 2248 43616 2312
rect 43680 2248 43696 2312
rect 43760 2248 43776 2312
rect 43840 2248 43856 2312
rect 43920 2248 43936 2312
rect 44000 2248 44016 2312
rect 44080 2248 44096 2312
rect 44160 2248 44176 2312
rect 44240 2248 44256 2312
rect 44320 2248 44336 2312
rect 44400 2248 44416 2312
rect 44480 2248 44496 2312
rect 44560 2248 44576 2312
rect 44640 2248 44656 2312
rect 44720 2248 44736 2312
rect 44800 2248 44816 2312
rect 44880 2248 44896 2312
rect 44960 2248 44976 2312
rect 45040 2248 45056 2312
rect 45120 2248 45136 2312
rect 45200 2248 45216 2312
rect 45280 2248 45296 2312
rect 45360 2248 45368 2312
rect 41368 2232 45368 2248
rect 41368 2168 41376 2232
rect 41440 2168 41456 2232
rect 41520 2168 41536 2232
rect 41600 2168 41616 2232
rect 41680 2168 41696 2232
rect 41760 2168 41776 2232
rect 41840 2168 41856 2232
rect 41920 2168 41936 2232
rect 42000 2168 42016 2232
rect 42080 2168 42096 2232
rect 42160 2168 42176 2232
rect 42240 2168 42256 2232
rect 42320 2168 42336 2232
rect 42400 2168 42416 2232
rect 42480 2168 42496 2232
rect 42560 2168 42576 2232
rect 42640 2168 42656 2232
rect 42720 2168 42736 2232
rect 42800 2168 42816 2232
rect 42880 2168 42896 2232
rect 42960 2168 42976 2232
rect 43040 2168 43056 2232
rect 43120 2168 43136 2232
rect 43200 2168 43216 2232
rect 43280 2168 43296 2232
rect 43360 2168 43376 2232
rect 43440 2168 43456 2232
rect 43520 2168 43536 2232
rect 43600 2168 43616 2232
rect 43680 2168 43696 2232
rect 43760 2168 43776 2232
rect 43840 2168 43856 2232
rect 43920 2168 43936 2232
rect 44000 2168 44016 2232
rect 44080 2168 44096 2232
rect 44160 2168 44176 2232
rect 44240 2168 44256 2232
rect 44320 2168 44336 2232
rect 44400 2168 44416 2232
rect 44480 2168 44496 2232
rect 44560 2168 44576 2232
rect 44640 2168 44656 2232
rect 44720 2168 44736 2232
rect 44800 2168 44816 2232
rect 44880 2168 44896 2232
rect 44960 2168 44976 2232
rect 45040 2168 45056 2232
rect 45120 2168 45136 2232
rect 45200 2168 45216 2232
rect 45280 2168 45296 2232
rect 45360 2168 45368 2232
rect 41368 2152 45368 2168
rect 41368 2088 41376 2152
rect 41440 2088 41456 2152
rect 41520 2088 41536 2152
rect 41600 2088 41616 2152
rect 41680 2088 41696 2152
rect 41760 2088 41776 2152
rect 41840 2088 41856 2152
rect 41920 2088 41936 2152
rect 42000 2088 42016 2152
rect 42080 2088 42096 2152
rect 42160 2088 42176 2152
rect 42240 2088 42256 2152
rect 42320 2088 42336 2152
rect 42400 2088 42416 2152
rect 42480 2088 42496 2152
rect 42560 2088 42576 2152
rect 42640 2088 42656 2152
rect 42720 2088 42736 2152
rect 42800 2088 42816 2152
rect 42880 2088 42896 2152
rect 42960 2088 42976 2152
rect 43040 2088 43056 2152
rect 43120 2088 43136 2152
rect 43200 2088 43216 2152
rect 43280 2088 43296 2152
rect 43360 2088 43376 2152
rect 43440 2088 43456 2152
rect 43520 2088 43536 2152
rect 43600 2088 43616 2152
rect 43680 2088 43696 2152
rect 43760 2088 43776 2152
rect 43840 2088 43856 2152
rect 43920 2088 43936 2152
rect 44000 2088 44016 2152
rect 44080 2088 44096 2152
rect 44160 2088 44176 2152
rect 44240 2088 44256 2152
rect 44320 2088 44336 2152
rect 44400 2088 44416 2152
rect 44480 2088 44496 2152
rect 44560 2088 44576 2152
rect 44640 2088 44656 2152
rect 44720 2088 44736 2152
rect 44800 2088 44816 2152
rect 44880 2088 44896 2152
rect 44960 2088 44976 2152
rect 45040 2088 45056 2152
rect 45120 2088 45136 2152
rect 45200 2088 45216 2152
rect 45280 2088 45296 2152
rect 45360 2088 45368 2152
rect 41368 2072 45368 2088
rect 41368 2008 41376 2072
rect 41440 2008 41456 2072
rect 41520 2008 41536 2072
rect 41600 2008 41616 2072
rect 41680 2008 41696 2072
rect 41760 2008 41776 2072
rect 41840 2008 41856 2072
rect 41920 2008 41936 2072
rect 42000 2008 42016 2072
rect 42080 2008 42096 2072
rect 42160 2008 42176 2072
rect 42240 2008 42256 2072
rect 42320 2008 42336 2072
rect 42400 2008 42416 2072
rect 42480 2008 42496 2072
rect 42560 2008 42576 2072
rect 42640 2008 42656 2072
rect 42720 2008 42736 2072
rect 42800 2008 42816 2072
rect 42880 2008 42896 2072
rect 42960 2008 42976 2072
rect 43040 2008 43056 2072
rect 43120 2008 43136 2072
rect 43200 2008 43216 2072
rect 43280 2008 43296 2072
rect 43360 2008 43376 2072
rect 43440 2008 43456 2072
rect 43520 2008 43536 2072
rect 43600 2008 43616 2072
rect 43680 2008 43696 2072
rect 43760 2008 43776 2072
rect 43840 2008 43856 2072
rect 43920 2008 43936 2072
rect 44000 2008 44016 2072
rect 44080 2008 44096 2072
rect 44160 2008 44176 2072
rect 44240 2008 44256 2072
rect 44320 2008 44336 2072
rect 44400 2008 44416 2072
rect 44480 2008 44496 2072
rect 44560 2008 44576 2072
rect 44640 2008 44656 2072
rect 44720 2008 44736 2072
rect 44800 2008 44816 2072
rect 44880 2008 44896 2072
rect 44960 2008 44976 2072
rect 45040 2008 45056 2072
rect 45120 2008 45136 2072
rect 45200 2008 45216 2072
rect 45280 2008 45296 2072
rect 45360 2008 45368 2072
rect 41368 1992 45368 2008
rect 41368 1928 41376 1992
rect 41440 1928 41456 1992
rect 41520 1928 41536 1992
rect 41600 1928 41616 1992
rect 41680 1928 41696 1992
rect 41760 1928 41776 1992
rect 41840 1928 41856 1992
rect 41920 1928 41936 1992
rect 42000 1928 42016 1992
rect 42080 1928 42096 1992
rect 42160 1928 42176 1992
rect 42240 1928 42256 1992
rect 42320 1928 42336 1992
rect 42400 1928 42416 1992
rect 42480 1928 42496 1992
rect 42560 1928 42576 1992
rect 42640 1928 42656 1992
rect 42720 1928 42736 1992
rect 42800 1928 42816 1992
rect 42880 1928 42896 1992
rect 42960 1928 42976 1992
rect 43040 1928 43056 1992
rect 43120 1928 43136 1992
rect 43200 1928 43216 1992
rect 43280 1928 43296 1992
rect 43360 1928 43376 1992
rect 43440 1928 43456 1992
rect 43520 1928 43536 1992
rect 43600 1928 43616 1992
rect 43680 1928 43696 1992
rect 43760 1928 43776 1992
rect 43840 1928 43856 1992
rect 43920 1928 43936 1992
rect 44000 1928 44016 1992
rect 44080 1928 44096 1992
rect 44160 1928 44176 1992
rect 44240 1928 44256 1992
rect 44320 1928 44336 1992
rect 44400 1928 44416 1992
rect 44480 1928 44496 1992
rect 44560 1928 44576 1992
rect 44640 1928 44656 1992
rect 44720 1928 44736 1992
rect 44800 1928 44816 1992
rect 44880 1928 44896 1992
rect 44960 1928 44976 1992
rect 45040 1928 45056 1992
rect 45120 1928 45136 1992
rect 45200 1928 45216 1992
rect 45280 1928 45296 1992
rect 45360 1928 45368 1992
rect 41368 1912 45368 1928
rect 41368 1848 41376 1912
rect 41440 1848 41456 1912
rect 41520 1848 41536 1912
rect 41600 1848 41616 1912
rect 41680 1848 41696 1912
rect 41760 1848 41776 1912
rect 41840 1848 41856 1912
rect 41920 1848 41936 1912
rect 42000 1848 42016 1912
rect 42080 1848 42096 1912
rect 42160 1848 42176 1912
rect 42240 1848 42256 1912
rect 42320 1848 42336 1912
rect 42400 1848 42416 1912
rect 42480 1848 42496 1912
rect 42560 1848 42576 1912
rect 42640 1848 42656 1912
rect 42720 1848 42736 1912
rect 42800 1848 42816 1912
rect 42880 1848 42896 1912
rect 42960 1848 42976 1912
rect 43040 1848 43056 1912
rect 43120 1848 43136 1912
rect 43200 1848 43216 1912
rect 43280 1848 43296 1912
rect 43360 1848 43376 1912
rect 43440 1848 43456 1912
rect 43520 1848 43536 1912
rect 43600 1848 43616 1912
rect 43680 1848 43696 1912
rect 43760 1848 43776 1912
rect 43840 1848 43856 1912
rect 43920 1848 43936 1912
rect 44000 1848 44016 1912
rect 44080 1848 44096 1912
rect 44160 1848 44176 1912
rect 44240 1848 44256 1912
rect 44320 1848 44336 1912
rect 44400 1848 44416 1912
rect 44480 1848 44496 1912
rect 44560 1848 44576 1912
rect 44640 1848 44656 1912
rect 44720 1848 44736 1912
rect 44800 1848 44816 1912
rect 44880 1848 44896 1912
rect 44960 1848 44976 1912
rect 45040 1848 45056 1912
rect 45120 1848 45136 1912
rect 45200 1848 45216 1912
rect 45280 1848 45296 1912
rect 45360 1848 45368 1912
rect 41368 1832 45368 1848
rect 41368 1768 41376 1832
rect 41440 1768 41456 1832
rect 41520 1768 41536 1832
rect 41600 1768 41616 1832
rect 41680 1768 41696 1832
rect 41760 1768 41776 1832
rect 41840 1768 41856 1832
rect 41920 1768 41936 1832
rect 42000 1768 42016 1832
rect 42080 1768 42096 1832
rect 42160 1768 42176 1832
rect 42240 1768 42256 1832
rect 42320 1768 42336 1832
rect 42400 1768 42416 1832
rect 42480 1768 42496 1832
rect 42560 1768 42576 1832
rect 42640 1768 42656 1832
rect 42720 1768 42736 1832
rect 42800 1768 42816 1832
rect 42880 1768 42896 1832
rect 42960 1768 42976 1832
rect 43040 1768 43056 1832
rect 43120 1768 43136 1832
rect 43200 1768 43216 1832
rect 43280 1768 43296 1832
rect 43360 1768 43376 1832
rect 43440 1768 43456 1832
rect 43520 1768 43536 1832
rect 43600 1768 43616 1832
rect 43680 1768 43696 1832
rect 43760 1768 43776 1832
rect 43840 1768 43856 1832
rect 43920 1768 43936 1832
rect 44000 1768 44016 1832
rect 44080 1768 44096 1832
rect 44160 1768 44176 1832
rect 44240 1768 44256 1832
rect 44320 1768 44336 1832
rect 44400 1768 44416 1832
rect 44480 1768 44496 1832
rect 44560 1768 44576 1832
rect 44640 1768 44656 1832
rect 44720 1768 44736 1832
rect 44800 1768 44816 1832
rect 44880 1768 44896 1832
rect 44960 1768 44976 1832
rect 45040 1768 45056 1832
rect 45120 1768 45136 1832
rect 45200 1768 45216 1832
rect 45280 1768 45296 1832
rect 45360 1768 45368 1832
rect 41368 1752 45368 1768
rect 41368 1688 41376 1752
rect 41440 1688 41456 1752
rect 41520 1688 41536 1752
rect 41600 1688 41616 1752
rect 41680 1688 41696 1752
rect 41760 1688 41776 1752
rect 41840 1688 41856 1752
rect 41920 1688 41936 1752
rect 42000 1688 42016 1752
rect 42080 1688 42096 1752
rect 42160 1688 42176 1752
rect 42240 1688 42256 1752
rect 42320 1688 42336 1752
rect 42400 1688 42416 1752
rect 42480 1688 42496 1752
rect 42560 1688 42576 1752
rect 42640 1688 42656 1752
rect 42720 1688 42736 1752
rect 42800 1688 42816 1752
rect 42880 1688 42896 1752
rect 42960 1688 42976 1752
rect 43040 1688 43056 1752
rect 43120 1688 43136 1752
rect 43200 1688 43216 1752
rect 43280 1688 43296 1752
rect 43360 1688 43376 1752
rect 43440 1688 43456 1752
rect 43520 1688 43536 1752
rect 43600 1688 43616 1752
rect 43680 1688 43696 1752
rect 43760 1688 43776 1752
rect 43840 1688 43856 1752
rect 43920 1688 43936 1752
rect 44000 1688 44016 1752
rect 44080 1688 44096 1752
rect 44160 1688 44176 1752
rect 44240 1688 44256 1752
rect 44320 1688 44336 1752
rect 44400 1688 44416 1752
rect 44480 1688 44496 1752
rect 44560 1688 44576 1752
rect 44640 1688 44656 1752
rect 44720 1688 44736 1752
rect 44800 1688 44816 1752
rect 44880 1688 44896 1752
rect 44960 1688 44976 1752
rect 45040 1688 45056 1752
rect 45120 1688 45136 1752
rect 45200 1688 45216 1752
rect 45280 1688 45296 1752
rect 45360 1688 45368 1752
rect 41368 1672 45368 1688
rect 41368 1608 41376 1672
rect 41440 1608 41456 1672
rect 41520 1608 41536 1672
rect 41600 1608 41616 1672
rect 41680 1608 41696 1672
rect 41760 1608 41776 1672
rect 41840 1608 41856 1672
rect 41920 1608 41936 1672
rect 42000 1608 42016 1672
rect 42080 1608 42096 1672
rect 42160 1608 42176 1672
rect 42240 1608 42256 1672
rect 42320 1608 42336 1672
rect 42400 1608 42416 1672
rect 42480 1608 42496 1672
rect 42560 1608 42576 1672
rect 42640 1608 42656 1672
rect 42720 1608 42736 1672
rect 42800 1608 42816 1672
rect 42880 1608 42896 1672
rect 42960 1608 42976 1672
rect 43040 1608 43056 1672
rect 43120 1608 43136 1672
rect 43200 1608 43216 1672
rect 43280 1608 43296 1672
rect 43360 1608 43376 1672
rect 43440 1608 43456 1672
rect 43520 1608 43536 1672
rect 43600 1608 43616 1672
rect 43680 1608 43696 1672
rect 43760 1608 43776 1672
rect 43840 1608 43856 1672
rect 43920 1608 43936 1672
rect 44000 1608 44016 1672
rect 44080 1608 44096 1672
rect 44160 1608 44176 1672
rect 44240 1608 44256 1672
rect 44320 1608 44336 1672
rect 44400 1608 44416 1672
rect 44480 1608 44496 1672
rect 44560 1608 44576 1672
rect 44640 1608 44656 1672
rect 44720 1608 44736 1672
rect 44800 1608 44816 1672
rect 44880 1608 44896 1672
rect 44960 1608 44976 1672
rect 45040 1608 45056 1672
rect 45120 1608 45136 1672
rect 45200 1608 45216 1672
rect 45280 1608 45296 1672
rect 45360 1608 45368 1672
rect 41368 1592 45368 1608
rect 41368 1528 41376 1592
rect 41440 1528 41456 1592
rect 41520 1528 41536 1592
rect 41600 1528 41616 1592
rect 41680 1528 41696 1592
rect 41760 1528 41776 1592
rect 41840 1528 41856 1592
rect 41920 1528 41936 1592
rect 42000 1528 42016 1592
rect 42080 1528 42096 1592
rect 42160 1528 42176 1592
rect 42240 1528 42256 1592
rect 42320 1528 42336 1592
rect 42400 1528 42416 1592
rect 42480 1528 42496 1592
rect 42560 1528 42576 1592
rect 42640 1528 42656 1592
rect 42720 1528 42736 1592
rect 42800 1528 42816 1592
rect 42880 1528 42896 1592
rect 42960 1528 42976 1592
rect 43040 1528 43056 1592
rect 43120 1528 43136 1592
rect 43200 1528 43216 1592
rect 43280 1528 43296 1592
rect 43360 1528 43376 1592
rect 43440 1528 43456 1592
rect 43520 1528 43536 1592
rect 43600 1528 43616 1592
rect 43680 1528 43696 1592
rect 43760 1528 43776 1592
rect 43840 1528 43856 1592
rect 43920 1528 43936 1592
rect 44000 1528 44016 1592
rect 44080 1528 44096 1592
rect 44160 1528 44176 1592
rect 44240 1528 44256 1592
rect 44320 1528 44336 1592
rect 44400 1528 44416 1592
rect 44480 1528 44496 1592
rect 44560 1528 44576 1592
rect 44640 1528 44656 1592
rect 44720 1528 44736 1592
rect 44800 1528 44816 1592
rect 44880 1528 44896 1592
rect 44960 1528 44976 1592
rect 45040 1528 45056 1592
rect 45120 1528 45136 1592
rect 45200 1528 45216 1592
rect 45280 1528 45296 1592
rect 45360 1528 45368 1592
rect 41368 1512 45368 1528
rect 41368 1448 41376 1512
rect 41440 1448 41456 1512
rect 41520 1448 41536 1512
rect 41600 1448 41616 1512
rect 41680 1448 41696 1512
rect 41760 1448 41776 1512
rect 41840 1448 41856 1512
rect 41920 1448 41936 1512
rect 42000 1448 42016 1512
rect 42080 1448 42096 1512
rect 42160 1448 42176 1512
rect 42240 1448 42256 1512
rect 42320 1448 42336 1512
rect 42400 1448 42416 1512
rect 42480 1448 42496 1512
rect 42560 1448 42576 1512
rect 42640 1448 42656 1512
rect 42720 1448 42736 1512
rect 42800 1448 42816 1512
rect 42880 1448 42896 1512
rect 42960 1448 42976 1512
rect 43040 1448 43056 1512
rect 43120 1448 43136 1512
rect 43200 1448 43216 1512
rect 43280 1448 43296 1512
rect 43360 1448 43376 1512
rect 43440 1448 43456 1512
rect 43520 1448 43536 1512
rect 43600 1448 43616 1512
rect 43680 1448 43696 1512
rect 43760 1448 43776 1512
rect 43840 1448 43856 1512
rect 43920 1448 43936 1512
rect 44000 1448 44016 1512
rect 44080 1448 44096 1512
rect 44160 1448 44176 1512
rect 44240 1448 44256 1512
rect 44320 1448 44336 1512
rect 44400 1448 44416 1512
rect 44480 1448 44496 1512
rect 44560 1448 44576 1512
rect 44640 1448 44656 1512
rect 44720 1448 44736 1512
rect 44800 1448 44816 1512
rect 44880 1448 44896 1512
rect 44960 1448 44976 1512
rect 45040 1448 45056 1512
rect 45120 1448 45136 1512
rect 45200 1448 45216 1512
rect 45280 1448 45296 1512
rect 45360 1448 45368 1512
rect 41368 1432 45368 1448
rect 41368 1368 41376 1432
rect 41440 1368 41456 1432
rect 41520 1368 41536 1432
rect 41600 1368 41616 1432
rect 41680 1368 41696 1432
rect 41760 1368 41776 1432
rect 41840 1368 41856 1432
rect 41920 1368 41936 1432
rect 42000 1368 42016 1432
rect 42080 1368 42096 1432
rect 42160 1368 42176 1432
rect 42240 1368 42256 1432
rect 42320 1368 42336 1432
rect 42400 1368 42416 1432
rect 42480 1368 42496 1432
rect 42560 1368 42576 1432
rect 42640 1368 42656 1432
rect 42720 1368 42736 1432
rect 42800 1368 42816 1432
rect 42880 1368 42896 1432
rect 42960 1368 42976 1432
rect 43040 1368 43056 1432
rect 43120 1368 43136 1432
rect 43200 1368 43216 1432
rect 43280 1368 43296 1432
rect 43360 1368 43376 1432
rect 43440 1368 43456 1432
rect 43520 1368 43536 1432
rect 43600 1368 43616 1432
rect 43680 1368 43696 1432
rect 43760 1368 43776 1432
rect 43840 1368 43856 1432
rect 43920 1368 43936 1432
rect 44000 1368 44016 1432
rect 44080 1368 44096 1432
rect 44160 1368 44176 1432
rect 44240 1368 44256 1432
rect 44320 1368 44336 1432
rect 44400 1368 44416 1432
rect 44480 1368 44496 1432
rect 44560 1368 44576 1432
rect 44640 1368 44656 1432
rect 44720 1368 44736 1432
rect 44800 1368 44816 1432
rect 44880 1368 44896 1432
rect 44960 1368 44976 1432
rect 45040 1368 45056 1432
rect 45120 1368 45136 1432
rect 45200 1368 45216 1432
rect 45280 1368 45296 1432
rect 45360 1368 45368 1432
rect 41368 1352 45368 1368
rect 41368 1288 41376 1352
rect 41440 1288 41456 1352
rect 41520 1288 41536 1352
rect 41600 1288 41616 1352
rect 41680 1288 41696 1352
rect 41760 1288 41776 1352
rect 41840 1288 41856 1352
rect 41920 1288 41936 1352
rect 42000 1288 42016 1352
rect 42080 1288 42096 1352
rect 42160 1288 42176 1352
rect 42240 1288 42256 1352
rect 42320 1288 42336 1352
rect 42400 1288 42416 1352
rect 42480 1288 42496 1352
rect 42560 1288 42576 1352
rect 42640 1288 42656 1352
rect 42720 1288 42736 1352
rect 42800 1288 42816 1352
rect 42880 1288 42896 1352
rect 42960 1288 42976 1352
rect 43040 1288 43056 1352
rect 43120 1288 43136 1352
rect 43200 1288 43216 1352
rect 43280 1288 43296 1352
rect 43360 1288 43376 1352
rect 43440 1288 43456 1352
rect 43520 1288 43536 1352
rect 43600 1288 43616 1352
rect 43680 1288 43696 1352
rect 43760 1288 43776 1352
rect 43840 1288 43856 1352
rect 43920 1288 43936 1352
rect 44000 1288 44016 1352
rect 44080 1288 44096 1352
rect 44160 1288 44176 1352
rect 44240 1288 44256 1352
rect 44320 1288 44336 1352
rect 44400 1288 44416 1352
rect 44480 1288 44496 1352
rect 44560 1288 44576 1352
rect 44640 1288 44656 1352
rect 44720 1288 44736 1352
rect 44800 1288 44816 1352
rect 44880 1288 44896 1352
rect 44960 1288 44976 1352
rect 45040 1288 45056 1352
rect 45120 1288 45136 1352
rect 45200 1288 45216 1352
rect 45280 1288 45296 1352
rect 45360 1288 45368 1352
rect 41368 1272 45368 1288
rect 41368 1208 41376 1272
rect 41440 1208 41456 1272
rect 41520 1208 41536 1272
rect 41600 1208 41616 1272
rect 41680 1208 41696 1272
rect 41760 1208 41776 1272
rect 41840 1208 41856 1272
rect 41920 1208 41936 1272
rect 42000 1208 42016 1272
rect 42080 1208 42096 1272
rect 42160 1208 42176 1272
rect 42240 1208 42256 1272
rect 42320 1208 42336 1272
rect 42400 1208 42416 1272
rect 42480 1208 42496 1272
rect 42560 1208 42576 1272
rect 42640 1208 42656 1272
rect 42720 1208 42736 1272
rect 42800 1208 42816 1272
rect 42880 1208 42896 1272
rect 42960 1208 42976 1272
rect 43040 1208 43056 1272
rect 43120 1208 43136 1272
rect 43200 1208 43216 1272
rect 43280 1208 43296 1272
rect 43360 1208 43376 1272
rect 43440 1208 43456 1272
rect 43520 1208 43536 1272
rect 43600 1208 43616 1272
rect 43680 1208 43696 1272
rect 43760 1208 43776 1272
rect 43840 1208 43856 1272
rect 43920 1208 43936 1272
rect 44000 1208 44016 1272
rect 44080 1208 44096 1272
rect 44160 1208 44176 1272
rect 44240 1208 44256 1272
rect 44320 1208 44336 1272
rect 44400 1208 44416 1272
rect 44480 1208 44496 1272
rect 44560 1208 44576 1272
rect 44640 1208 44656 1272
rect 44720 1208 44736 1272
rect 44800 1208 44816 1272
rect 44880 1208 44896 1272
rect 44960 1208 44976 1272
rect 45040 1208 45056 1272
rect 45120 1208 45136 1272
rect 45200 1208 45216 1272
rect 45280 1208 45296 1272
rect 45360 1208 45368 1272
rect 41368 1192 45368 1208
rect 41368 1128 41376 1192
rect 41440 1128 41456 1192
rect 41520 1128 41536 1192
rect 41600 1128 41616 1192
rect 41680 1128 41696 1192
rect 41760 1128 41776 1192
rect 41840 1128 41856 1192
rect 41920 1128 41936 1192
rect 42000 1128 42016 1192
rect 42080 1128 42096 1192
rect 42160 1128 42176 1192
rect 42240 1128 42256 1192
rect 42320 1128 42336 1192
rect 42400 1128 42416 1192
rect 42480 1128 42496 1192
rect 42560 1128 42576 1192
rect 42640 1128 42656 1192
rect 42720 1128 42736 1192
rect 42800 1128 42816 1192
rect 42880 1128 42896 1192
rect 42960 1128 42976 1192
rect 43040 1128 43056 1192
rect 43120 1128 43136 1192
rect 43200 1128 43216 1192
rect 43280 1128 43296 1192
rect 43360 1128 43376 1192
rect 43440 1128 43456 1192
rect 43520 1128 43536 1192
rect 43600 1128 43616 1192
rect 43680 1128 43696 1192
rect 43760 1128 43776 1192
rect 43840 1128 43856 1192
rect 43920 1128 43936 1192
rect 44000 1128 44016 1192
rect 44080 1128 44096 1192
rect 44160 1128 44176 1192
rect 44240 1128 44256 1192
rect 44320 1128 44336 1192
rect 44400 1128 44416 1192
rect 44480 1128 44496 1192
rect 44560 1128 44576 1192
rect 44640 1128 44656 1192
rect 44720 1128 44736 1192
rect 44800 1128 44816 1192
rect 44880 1128 44896 1192
rect 44960 1128 44976 1192
rect 45040 1128 45056 1192
rect 45120 1128 45136 1192
rect 45200 1128 45216 1192
rect 45280 1128 45296 1192
rect 45360 1128 45368 1192
rect 41368 1112 45368 1128
rect 41368 1048 41376 1112
rect 41440 1048 41456 1112
rect 41520 1048 41536 1112
rect 41600 1048 41616 1112
rect 41680 1048 41696 1112
rect 41760 1048 41776 1112
rect 41840 1048 41856 1112
rect 41920 1048 41936 1112
rect 42000 1048 42016 1112
rect 42080 1048 42096 1112
rect 42160 1048 42176 1112
rect 42240 1048 42256 1112
rect 42320 1048 42336 1112
rect 42400 1048 42416 1112
rect 42480 1048 42496 1112
rect 42560 1048 42576 1112
rect 42640 1048 42656 1112
rect 42720 1048 42736 1112
rect 42800 1048 42816 1112
rect 42880 1048 42896 1112
rect 42960 1048 42976 1112
rect 43040 1048 43056 1112
rect 43120 1048 43136 1112
rect 43200 1048 43216 1112
rect 43280 1048 43296 1112
rect 43360 1048 43376 1112
rect 43440 1048 43456 1112
rect 43520 1048 43536 1112
rect 43600 1048 43616 1112
rect 43680 1048 43696 1112
rect 43760 1048 43776 1112
rect 43840 1048 43856 1112
rect 43920 1048 43936 1112
rect 44000 1048 44016 1112
rect 44080 1048 44096 1112
rect 44160 1048 44176 1112
rect 44240 1048 44256 1112
rect 44320 1048 44336 1112
rect 44400 1048 44416 1112
rect 44480 1048 44496 1112
rect 44560 1048 44576 1112
rect 44640 1048 44656 1112
rect 44720 1048 44736 1112
rect 44800 1048 44816 1112
rect 44880 1048 44896 1112
rect 44960 1048 44976 1112
rect 45040 1048 45056 1112
rect 45120 1048 45136 1112
rect 45200 1048 45216 1112
rect 45280 1048 45296 1112
rect 45360 1048 45368 1112
rect 41368 1032 45368 1048
rect 41368 968 41376 1032
rect 41440 968 41456 1032
rect 41520 968 41536 1032
rect 41600 968 41616 1032
rect 41680 968 41696 1032
rect 41760 968 41776 1032
rect 41840 968 41856 1032
rect 41920 968 41936 1032
rect 42000 968 42016 1032
rect 42080 968 42096 1032
rect 42160 968 42176 1032
rect 42240 968 42256 1032
rect 42320 968 42336 1032
rect 42400 968 42416 1032
rect 42480 968 42496 1032
rect 42560 968 42576 1032
rect 42640 968 42656 1032
rect 42720 968 42736 1032
rect 42800 968 42816 1032
rect 42880 968 42896 1032
rect 42960 968 42976 1032
rect 43040 968 43056 1032
rect 43120 968 43136 1032
rect 43200 968 43216 1032
rect 43280 968 43296 1032
rect 43360 968 43376 1032
rect 43440 968 43456 1032
rect 43520 968 43536 1032
rect 43600 968 43616 1032
rect 43680 968 43696 1032
rect 43760 968 43776 1032
rect 43840 968 43856 1032
rect 43920 968 43936 1032
rect 44000 968 44016 1032
rect 44080 968 44096 1032
rect 44160 968 44176 1032
rect 44240 968 44256 1032
rect 44320 968 44336 1032
rect 44400 968 44416 1032
rect 44480 968 44496 1032
rect 44560 968 44576 1032
rect 44640 968 44656 1032
rect 44720 968 44736 1032
rect 44800 968 44816 1032
rect 44880 968 44896 1032
rect 44960 968 44976 1032
rect 45040 968 45056 1032
rect 45120 968 45136 1032
rect 45200 968 45216 1032
rect 45280 968 45296 1032
rect 45360 968 45368 1032
rect 41368 952 45368 968
rect 41368 888 41376 952
rect 41440 888 41456 952
rect 41520 888 41536 952
rect 41600 888 41616 952
rect 41680 888 41696 952
rect 41760 888 41776 952
rect 41840 888 41856 952
rect 41920 888 41936 952
rect 42000 888 42016 952
rect 42080 888 42096 952
rect 42160 888 42176 952
rect 42240 888 42256 952
rect 42320 888 42336 952
rect 42400 888 42416 952
rect 42480 888 42496 952
rect 42560 888 42576 952
rect 42640 888 42656 952
rect 42720 888 42736 952
rect 42800 888 42816 952
rect 42880 888 42896 952
rect 42960 888 42976 952
rect 43040 888 43056 952
rect 43120 888 43136 952
rect 43200 888 43216 952
rect 43280 888 43296 952
rect 43360 888 43376 952
rect 43440 888 43456 952
rect 43520 888 43536 952
rect 43600 888 43616 952
rect 43680 888 43696 952
rect 43760 888 43776 952
rect 43840 888 43856 952
rect 43920 888 43936 952
rect 44000 888 44016 952
rect 44080 888 44096 952
rect 44160 888 44176 952
rect 44240 888 44256 952
rect 44320 888 44336 952
rect 44400 888 44416 952
rect 44480 888 44496 952
rect 44560 888 44576 952
rect 44640 888 44656 952
rect 44720 888 44736 952
rect 44800 888 44816 952
rect 44880 888 44896 952
rect 44960 888 44976 952
rect 45040 888 45056 952
rect 45120 888 45136 952
rect 45200 888 45216 952
rect 45280 888 45296 952
rect 45360 888 45368 952
rect 41368 872 45368 888
rect 41368 808 41376 872
rect 41440 808 41456 872
rect 41520 808 41536 872
rect 41600 808 41616 872
rect 41680 808 41696 872
rect 41760 808 41776 872
rect 41840 808 41856 872
rect 41920 808 41936 872
rect 42000 808 42016 872
rect 42080 808 42096 872
rect 42160 808 42176 872
rect 42240 808 42256 872
rect 42320 808 42336 872
rect 42400 808 42416 872
rect 42480 808 42496 872
rect 42560 808 42576 872
rect 42640 808 42656 872
rect 42720 808 42736 872
rect 42800 808 42816 872
rect 42880 808 42896 872
rect 42960 808 42976 872
rect 43040 808 43056 872
rect 43120 808 43136 872
rect 43200 808 43216 872
rect 43280 808 43296 872
rect 43360 808 43376 872
rect 43440 808 43456 872
rect 43520 808 43536 872
rect 43600 808 43616 872
rect 43680 808 43696 872
rect 43760 808 43776 872
rect 43840 808 43856 872
rect 43920 808 43936 872
rect 44000 808 44016 872
rect 44080 808 44096 872
rect 44160 808 44176 872
rect 44240 808 44256 872
rect 44320 808 44336 872
rect 44400 808 44416 872
rect 44480 808 44496 872
rect 44560 808 44576 872
rect 44640 808 44656 872
rect 44720 808 44736 872
rect 44800 808 44816 872
rect 44880 808 44896 872
rect 44960 808 44976 872
rect 45040 808 45056 872
rect 45120 808 45136 872
rect 45200 808 45216 872
rect 45280 808 45296 872
rect 45360 808 45368 872
rect 41368 792 45368 808
rect 41368 728 41376 792
rect 41440 728 41456 792
rect 41520 728 41536 792
rect 41600 728 41616 792
rect 41680 728 41696 792
rect 41760 728 41776 792
rect 41840 728 41856 792
rect 41920 728 41936 792
rect 42000 728 42016 792
rect 42080 728 42096 792
rect 42160 728 42176 792
rect 42240 728 42256 792
rect 42320 728 42336 792
rect 42400 728 42416 792
rect 42480 728 42496 792
rect 42560 728 42576 792
rect 42640 728 42656 792
rect 42720 728 42736 792
rect 42800 728 42816 792
rect 42880 728 42896 792
rect 42960 728 42976 792
rect 43040 728 43056 792
rect 43120 728 43136 792
rect 43200 728 43216 792
rect 43280 728 43296 792
rect 43360 728 43376 792
rect 43440 728 43456 792
rect 43520 728 43536 792
rect 43600 728 43616 792
rect 43680 728 43696 792
rect 43760 728 43776 792
rect 43840 728 43856 792
rect 43920 728 43936 792
rect 44000 728 44016 792
rect 44080 728 44096 792
rect 44160 728 44176 792
rect 44240 728 44256 792
rect 44320 728 44336 792
rect 44400 728 44416 792
rect 44480 728 44496 792
rect 44560 728 44576 792
rect 44640 728 44656 792
rect 44720 728 44736 792
rect 44800 728 44816 792
rect 44880 728 44896 792
rect 44960 728 44976 792
rect 45040 728 45056 792
rect 45120 728 45136 792
rect 45200 728 45216 792
rect 45280 728 45296 792
rect 45360 728 45368 792
rect 41368 712 45368 728
rect 41368 648 41376 712
rect 41440 648 41456 712
rect 41520 648 41536 712
rect 41600 648 41616 712
rect 41680 648 41696 712
rect 41760 648 41776 712
rect 41840 648 41856 712
rect 41920 648 41936 712
rect 42000 648 42016 712
rect 42080 648 42096 712
rect 42160 648 42176 712
rect 42240 648 42256 712
rect 42320 648 42336 712
rect 42400 648 42416 712
rect 42480 648 42496 712
rect 42560 648 42576 712
rect 42640 648 42656 712
rect 42720 648 42736 712
rect 42800 648 42816 712
rect 42880 648 42896 712
rect 42960 648 42976 712
rect 43040 648 43056 712
rect 43120 648 43136 712
rect 43200 648 43216 712
rect 43280 648 43296 712
rect 43360 648 43376 712
rect 43440 648 43456 712
rect 43520 648 43536 712
rect 43600 648 43616 712
rect 43680 648 43696 712
rect 43760 648 43776 712
rect 43840 648 43856 712
rect 43920 648 43936 712
rect 44000 648 44016 712
rect 44080 648 44096 712
rect 44160 648 44176 712
rect 44240 648 44256 712
rect 44320 648 44336 712
rect 44400 648 44416 712
rect 44480 648 44496 712
rect 44560 648 44576 712
rect 44640 648 44656 712
rect 44720 648 44736 712
rect 44800 648 44816 712
rect 44880 648 44896 712
rect 44960 648 44976 712
rect 45040 648 45056 712
rect 45120 648 45136 712
rect 45200 648 45216 712
rect 45280 648 45296 712
rect 45360 648 45368 712
rect 41368 632 45368 648
rect 41368 568 41376 632
rect 41440 568 41456 632
rect 41520 568 41536 632
rect 41600 568 41616 632
rect 41680 568 41696 632
rect 41760 568 41776 632
rect 41840 568 41856 632
rect 41920 568 41936 632
rect 42000 568 42016 632
rect 42080 568 42096 632
rect 42160 568 42176 632
rect 42240 568 42256 632
rect 42320 568 42336 632
rect 42400 568 42416 632
rect 42480 568 42496 632
rect 42560 568 42576 632
rect 42640 568 42656 632
rect 42720 568 42736 632
rect 42800 568 42816 632
rect 42880 568 42896 632
rect 42960 568 42976 632
rect 43040 568 43056 632
rect 43120 568 43136 632
rect 43200 568 43216 632
rect 43280 568 43296 632
rect 43360 568 43376 632
rect 43440 568 43456 632
rect 43520 568 43536 632
rect 43600 568 43616 632
rect 43680 568 43696 632
rect 43760 568 43776 632
rect 43840 568 43856 632
rect 43920 568 43936 632
rect 44000 568 44016 632
rect 44080 568 44096 632
rect 44160 568 44176 632
rect 44240 568 44256 632
rect 44320 568 44336 632
rect 44400 568 44416 632
rect 44480 568 44496 632
rect 44560 568 44576 632
rect 44640 568 44656 632
rect 44720 568 44736 632
rect 44800 568 44816 632
rect 44880 568 44896 632
rect 44960 568 44976 632
rect 45040 568 45056 632
rect 45120 568 45136 632
rect 45200 568 45216 632
rect 45280 568 45296 632
rect 45360 568 45368 632
rect 41368 552 45368 568
rect 41368 488 41376 552
rect 41440 488 41456 552
rect 41520 488 41536 552
rect 41600 488 41616 552
rect 41680 488 41696 552
rect 41760 488 41776 552
rect 41840 488 41856 552
rect 41920 488 41936 552
rect 42000 488 42016 552
rect 42080 488 42096 552
rect 42160 488 42176 552
rect 42240 488 42256 552
rect 42320 488 42336 552
rect 42400 488 42416 552
rect 42480 488 42496 552
rect 42560 488 42576 552
rect 42640 488 42656 552
rect 42720 488 42736 552
rect 42800 488 42816 552
rect 42880 488 42896 552
rect 42960 488 42976 552
rect 43040 488 43056 552
rect 43120 488 43136 552
rect 43200 488 43216 552
rect 43280 488 43296 552
rect 43360 488 43376 552
rect 43440 488 43456 552
rect 43520 488 43536 552
rect 43600 488 43616 552
rect 43680 488 43696 552
rect 43760 488 43776 552
rect 43840 488 43856 552
rect 43920 488 43936 552
rect 44000 488 44016 552
rect 44080 488 44096 552
rect 44160 488 44176 552
rect 44240 488 44256 552
rect 44320 488 44336 552
rect 44400 488 44416 552
rect 44480 488 44496 552
rect 44560 488 44576 552
rect 44640 488 44656 552
rect 44720 488 44736 552
rect 44800 488 44816 552
rect 44880 488 44896 552
rect 44960 488 44976 552
rect 45040 488 45056 552
rect 45120 488 45136 552
rect 45200 488 45216 552
rect 45280 488 45296 552
rect 45360 488 45368 552
rect 41368 472 45368 488
rect 41368 408 41376 472
rect 41440 408 41456 472
rect 41520 408 41536 472
rect 41600 408 41616 472
rect 41680 408 41696 472
rect 41760 408 41776 472
rect 41840 408 41856 472
rect 41920 408 41936 472
rect 42000 408 42016 472
rect 42080 408 42096 472
rect 42160 408 42176 472
rect 42240 408 42256 472
rect 42320 408 42336 472
rect 42400 408 42416 472
rect 42480 408 42496 472
rect 42560 408 42576 472
rect 42640 408 42656 472
rect 42720 408 42736 472
rect 42800 408 42816 472
rect 42880 408 42896 472
rect 42960 408 42976 472
rect 43040 408 43056 472
rect 43120 408 43136 472
rect 43200 408 43216 472
rect 43280 408 43296 472
rect 43360 408 43376 472
rect 43440 408 43456 472
rect 43520 408 43536 472
rect 43600 408 43616 472
rect 43680 408 43696 472
rect 43760 408 43776 472
rect 43840 408 43856 472
rect 43920 408 43936 472
rect 44000 408 44016 472
rect 44080 408 44096 472
rect 44160 408 44176 472
rect 44240 408 44256 472
rect 44320 408 44336 472
rect 44400 408 44416 472
rect 44480 408 44496 472
rect 44560 408 44576 472
rect 44640 408 44656 472
rect 44720 408 44736 472
rect 44800 408 44816 472
rect 44880 408 44896 472
rect 44960 408 44976 472
rect 45040 408 45056 472
rect 45120 408 45136 472
rect 45200 408 45216 472
rect 45280 408 45296 472
rect 45360 408 45368 472
rect 41368 392 45368 408
rect 41368 328 41376 392
rect 41440 328 41456 392
rect 41520 328 41536 392
rect 41600 328 41616 392
rect 41680 328 41696 392
rect 41760 328 41776 392
rect 41840 328 41856 392
rect 41920 328 41936 392
rect 42000 328 42016 392
rect 42080 328 42096 392
rect 42160 328 42176 392
rect 42240 328 42256 392
rect 42320 328 42336 392
rect 42400 328 42416 392
rect 42480 328 42496 392
rect 42560 328 42576 392
rect 42640 328 42656 392
rect 42720 328 42736 392
rect 42800 328 42816 392
rect 42880 328 42896 392
rect 42960 328 42976 392
rect 43040 328 43056 392
rect 43120 328 43136 392
rect 43200 328 43216 392
rect 43280 328 43296 392
rect 43360 328 43376 392
rect 43440 328 43456 392
rect 43520 328 43536 392
rect 43600 328 43616 392
rect 43680 328 43696 392
rect 43760 328 43776 392
rect 43840 328 43856 392
rect 43920 328 43936 392
rect 44000 328 44016 392
rect 44080 328 44096 392
rect 44160 328 44176 392
rect 44240 328 44256 392
rect 44320 328 44336 392
rect 44400 328 44416 392
rect 44480 328 44496 392
rect 44560 328 44576 392
rect 44640 328 44656 392
rect 44720 328 44736 392
rect 44800 328 44816 392
rect 44880 328 44896 392
rect 44960 328 44976 392
rect 45040 328 45056 392
rect 45120 328 45136 392
rect 45200 328 45216 392
rect 45280 328 45296 392
rect 45360 328 45368 392
rect 41368 312 45368 328
rect 41368 248 41376 312
rect 41440 248 41456 312
rect 41520 248 41536 312
rect 41600 248 41616 312
rect 41680 248 41696 312
rect 41760 248 41776 312
rect 41840 248 41856 312
rect 41920 248 41936 312
rect 42000 248 42016 312
rect 42080 248 42096 312
rect 42160 248 42176 312
rect 42240 248 42256 312
rect 42320 248 42336 312
rect 42400 248 42416 312
rect 42480 248 42496 312
rect 42560 248 42576 312
rect 42640 248 42656 312
rect 42720 248 42736 312
rect 42800 248 42816 312
rect 42880 248 42896 312
rect 42960 248 42976 312
rect 43040 248 43056 312
rect 43120 248 43136 312
rect 43200 248 43216 312
rect 43280 248 43296 312
rect 43360 248 43376 312
rect 43440 248 43456 312
rect 43520 248 43536 312
rect 43600 248 43616 312
rect 43680 248 43696 312
rect 43760 248 43776 312
rect 43840 248 43856 312
rect 43920 248 43936 312
rect 44000 248 44016 312
rect 44080 248 44096 312
rect 44160 248 44176 312
rect 44240 248 44256 312
rect 44320 248 44336 312
rect 44400 248 44416 312
rect 44480 248 44496 312
rect 44560 248 44576 312
rect 44640 248 44656 312
rect 44720 248 44736 312
rect 44800 248 44816 312
rect 44880 248 44896 312
rect 44960 248 44976 312
rect 45040 248 45056 312
rect 45120 248 45136 312
rect 45200 248 45216 312
rect 45280 248 45296 312
rect 45360 248 45368 312
rect 41368 232 45368 248
rect 41368 168 41376 232
rect 41440 168 41456 232
rect 41520 168 41536 232
rect 41600 168 41616 232
rect 41680 168 41696 232
rect 41760 168 41776 232
rect 41840 168 41856 232
rect 41920 168 41936 232
rect 42000 168 42016 232
rect 42080 168 42096 232
rect 42160 168 42176 232
rect 42240 168 42256 232
rect 42320 168 42336 232
rect 42400 168 42416 232
rect 42480 168 42496 232
rect 42560 168 42576 232
rect 42640 168 42656 232
rect 42720 168 42736 232
rect 42800 168 42816 232
rect 42880 168 42896 232
rect 42960 168 42976 232
rect 43040 168 43056 232
rect 43120 168 43136 232
rect 43200 168 43216 232
rect 43280 168 43296 232
rect 43360 168 43376 232
rect 43440 168 43456 232
rect 43520 168 43536 232
rect 43600 168 43616 232
rect 43680 168 43696 232
rect 43760 168 43776 232
rect 43840 168 43856 232
rect 43920 168 43936 232
rect 44000 168 44016 232
rect 44080 168 44096 232
rect 44160 168 44176 232
rect 44240 168 44256 232
rect 44320 168 44336 232
rect 44400 168 44416 232
rect 44480 168 44496 232
rect 44560 168 44576 232
rect 44640 168 44656 232
rect 44720 168 44736 232
rect 44800 168 44816 232
rect 44880 168 44896 232
rect 44960 168 44976 232
rect 45040 168 45056 232
rect 45120 168 45136 232
rect 45200 168 45216 232
rect 45280 168 45296 232
rect 45360 168 45368 232
rect 41368 152 45368 168
rect 41368 88 41376 152
rect 41440 88 41456 152
rect 41520 88 41536 152
rect 41600 88 41616 152
rect 41680 88 41696 152
rect 41760 88 41776 152
rect 41840 88 41856 152
rect 41920 88 41936 152
rect 42000 88 42016 152
rect 42080 88 42096 152
rect 42160 88 42176 152
rect 42240 88 42256 152
rect 42320 88 42336 152
rect 42400 88 42416 152
rect 42480 88 42496 152
rect 42560 88 42576 152
rect 42640 88 42656 152
rect 42720 88 42736 152
rect 42800 88 42816 152
rect 42880 88 42896 152
rect 42960 88 42976 152
rect 43040 88 43056 152
rect 43120 88 43136 152
rect 43200 88 43216 152
rect 43280 88 43296 152
rect 43360 88 43376 152
rect 43440 88 43456 152
rect 43520 88 43536 152
rect 43600 88 43616 152
rect 43680 88 43696 152
rect 43760 88 43776 152
rect 43840 88 43856 152
rect 43920 88 43936 152
rect 44000 88 44016 152
rect 44080 88 44096 152
rect 44160 88 44176 152
rect 44240 88 44256 152
rect 44320 88 44336 152
rect 44400 88 44416 152
rect 44480 88 44496 152
rect 44560 88 44576 152
rect 44640 88 44656 152
rect 44720 88 44736 152
rect 44800 88 44816 152
rect 44880 88 44896 152
rect 44960 88 44976 152
rect 45040 88 45056 152
rect 45120 88 45136 152
rect 45200 88 45216 152
rect 45280 88 45296 152
rect 45360 88 45368 152
rect 41368 72 45368 88
rect 41368 8 41376 72
rect 41440 8 41456 72
rect 41520 8 41536 72
rect 41600 8 41616 72
rect 41680 8 41696 72
rect 41760 8 41776 72
rect 41840 8 41856 72
rect 41920 8 41936 72
rect 42000 8 42016 72
rect 42080 8 42096 72
rect 42160 8 42176 72
rect 42240 8 42256 72
rect 42320 8 42336 72
rect 42400 8 42416 72
rect 42480 8 42496 72
rect 42560 8 42576 72
rect 42640 8 42656 72
rect 42720 8 42736 72
rect 42800 8 42816 72
rect 42880 8 42896 72
rect 42960 8 42976 72
rect 43040 8 43056 72
rect 43120 8 43136 72
rect 43200 8 43216 72
rect 43280 8 43296 72
rect 43360 8 43376 72
rect 43440 8 43456 72
rect 43520 8 43536 72
rect 43600 8 43616 72
rect 43680 8 43696 72
rect 43760 8 43776 72
rect 43840 8 43856 72
rect 43920 8 43936 72
rect 44000 8 44016 72
rect 44080 8 44096 72
rect 44160 8 44176 72
rect 44240 8 44256 72
rect 44320 8 44336 72
rect 44400 8 44416 72
rect 44480 8 44496 72
rect 44560 8 44576 72
rect 44640 8 44656 72
rect 44720 8 44736 72
rect 44800 8 44816 72
rect 44880 8 44896 72
rect 44960 8 44976 72
rect 45040 8 45056 72
rect 45120 8 45136 72
rect 45200 8 45216 72
rect 45280 8 45296 72
rect 45360 8 45368 72
rect 41368 0 45368 8
use sky130_fd_sc_hd__decap_3  PHY_0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 11000 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1600868798
transform 1 0 11000 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 11276 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1600868798
transform 1 0 12380 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1600868798
transform 1 0 11276 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1600868798
transform 1 0 12380 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _244_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 14680 0 -1 11544
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _536_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 14128 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13852 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13484 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13944 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_27 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13484 0 1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_33 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 14036 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1600868798
transform 1 0 16244 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1600868798
transform 1 0 16152 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49
timestamp 1600868798
transform 1 0 15508 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _512_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 15876 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1600868798
transform 1 0 17072 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1600868798
transform 1 0 16704 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1600868798
transform 1 0 17164 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1600868798
transform 1 0 16796 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1600868798
transform 1 0 16612 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1600868798
transform 1 0 16704 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _504_
timestamp 1600868798
transform 1 0 17256 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _243_
timestamp 1600868798
transform 1 0 17164 0 1 11544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1600868798
transform 1 0 17532 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _505_
timestamp 1600868798
transform 1 0 19648 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _520_
timestamp 1600868798
transform 1 0 18360 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1600868798
transform 1 0 19556 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83
timestamp 1600868798
transform 1 0 18636 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 19372 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1600868798
transform 1 0 17992 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _245_
timestamp 1600868798
transform 1 0 20844 0 1 11544
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _246_
timestamp 1600868798
transform 1 0 20844 0 -1 11544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1600868798
transform 1 0 19924 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1600868798
transform 1 0 20660 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1600868798
transform 1 0 21672 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1600868798
transform 1 0 20476 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1600868798
transform 1 0 21672 0 1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _511_
timestamp 1600868798
transform 1 0 22960 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _514_
timestamp 1600868798
transform 1 0 22316 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1600868798
transform 1 0 22408 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1600868798
transform 1 0 22224 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1600868798
transform 1 0 22500 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1600868798
transform 1 0 22868 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_133
timestamp 1600868798
transform 1 0 23236 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _260_
timestamp 1600868798
transform 1 0 25352 0 -1 11544
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _510_
timestamp 1600868798
transform 1 0 24524 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1600868798
transform 1 0 24800 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1600868798
transform 1 0 25260 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1600868798
transform 1 0 24340 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1600868798
transform 1 0 24800 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1600868798
transform 1 0 25168 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_165
timestamp 1600868798
transform 1 0 26180 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1600868798
transform 1 0 24432 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1600868798
transform 1 0 28112 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1600868798
transform 1 0 27836 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1600868798
transform 1 0 27284 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1600868798
transform 1 0 28020 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1600868798
transform 1 0 28204 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_173
timestamp 1600868798
transform 1 0 26916 0 1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1600868798
transform 1 0 27652 0 1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1600868798
transform 1 0 27928 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1600868798
transform 1 0 29308 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1600868798
transform 1 0 30412 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1600868798
transform 1 0 29032 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1600868798
transform 1 0 30136 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1600868798
transform 1 0 30964 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1600868798
transform 1 0 31056 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1600868798
transform 1 0 32160 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1600868798
transform 1 0 31240 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1600868798
transform 1 0 32344 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1600868798
transform -1 0 34368 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1600868798
transform -1 0 34368 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1600868798
transform 1 0 33816 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1600868798
transform 1 0 33448 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1600868798
transform 1 0 33264 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_249
timestamp 1600868798
transform 1 0 33908 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_245
timestamp 1600868798
transform 1 0 33540 0 1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _303_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 12196 0 -1 12632
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1600868798
transform 1 0 11000 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1600868798
transform 1 0 11276 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1600868798
transform 1 0 12012 0 -1 12632
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _265_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 14496 0 -1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1600868798
transform 1 0 13852 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1600868798
transform 1 0 13484 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1600868798
transform 1 0 13944 0 -1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1600868798
transform 1 0 16336 0 -1 12632
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1600868798
transform 1 0 15968 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _364_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 19556 0 -1 12632
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1600868798
transform 1 0 19464 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1600868798
transform 1 0 18452 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1600868798
transform 1 0 19188 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _535_
timestamp 1600868798
transform 1 0 21396 0 -1 12632
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_2_106
timestamp 1600868798
transform 1 0 20752 0 -1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1600868798
transform 1 0 21304 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_136
timestamp 1600868798
transform 1 0 23512 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 25168 0 -1 12632
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1600868798
transform 1 0 25076 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1600868798
transform 1 0 24616 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1600868798
transform 1 0 24984 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_167
timestamp 1600868798
transform 1 0 26364 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_179
timestamp 1600868798
transform 1 0 27468 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1600868798
transform 1 0 30688 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_191
timestamp 1600868798
transform 1 0 28572 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1600868798
transform 1 0 29676 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1600868798
transform 1 0 30412 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1600868798
transform 1 0 30780 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1600868798
transform 1 0 31884 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1600868798
transform -1 0 34368 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1600868798
transform 1 0 32988 0 -1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _304_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 12564 0 1 12632
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1600868798
transform 1 0 11000 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1600868798
transform 1 0 11276 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1600868798
transform 1 0 12380 0 1 12632
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _297_
timestamp 1600868798
transform 1 0 14128 0 1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1600868798
transform 1 0 13760 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1600868798
transform 1 0 16612 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_50
timestamp 1600868798
transform 1 0 15600 0 1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1600868798
transform 1 0 16336 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1600868798
transform 1 0 16704 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _363_
timestamp 1600868798
transform 1 0 17900 0 1 12632
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_3_74
timestamp 1600868798
transform 1 0 17808 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_88
timestamp 1600868798
transform 1 0 19096 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _268_
timestamp 1600868798
transform 1 0 20384 0 1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1600868798
transform 1 0 20200 0 1 12632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1600868798
transform 1 0 21856 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _284_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 22316 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1600868798
transform 1 0 22224 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1600868798
transform 1 0 23420 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _509_
timestamp 1600868798
transform 1 0 24984 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 25628 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1600868798
transform 1 0 24524 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1600868798
transform 1 0 24892 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1600868798
transform 1 0 25260 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_163
timestamp 1600868798
transform 1 0 25996 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1600868798
transform 1 0 27836 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1600868798
transform 1 0 27100 0 1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1600868798
transform 1 0 27928 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1600868798
transform 1 0 29032 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1600868798
transform 1 0 30136 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1600868798
transform 1 0 31240 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1600868798
transform 1 0 32344 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1600868798
transform -1 0 34368 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1600868798
transform 1 0 33448 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_245
timestamp 1600868798
transform 1 0 33540 0 1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _300_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 12840 0 -1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1600868798
transform 1 0 11000 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1600868798
transform 1 0 11276 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1600868798
transform 1 0 12380 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1600868798
transform 1 0 12748 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _299_
timestamp 1600868798
transform 1 0 13944 0 -1 13720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1600868798
transform 1 0 13852 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1600868798
transform 1 0 13484 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _362_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 16980 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_48
timestamp 1600868798
transform 1 0 15416 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1600868798
transform 1 0 16520 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1600868798
transform 1 0 16888 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _283_
timestamp 1600868798
transform 1 0 19648 0 -1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _361_
timestamp 1600868798
transform 1 0 18452 0 -1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1600868798
transform 1 0 19464 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_77
timestamp 1600868798
transform 1 0 18084 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1600868798
transform 1 0 19096 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1600868798
transform 1 0 19556 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _288_
timestamp 1600868798
transform 1 0 20660 0 -1 13720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 1600868798
transform 1 0 20292 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _301_
timestamp 1600868798
transform 1 0 23236 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1600868798
transform 1 0 22132 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _516_
timestamp 1600868798
transform 1 0 25168 0 -1 13720
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1600868798
transform 1 0 25076 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1600868798
transform 1 0 24340 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1600868798
transform 1 0 27284 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_189
timestamp 1600868798
transform 1 0 28388 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1600868798
transform 1 0 30688 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1600868798
transform 1 0 29492 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1600868798
transform 1 0 30596 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1600868798
transform 1 0 30780 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1600868798
transform 1 0 31884 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1600868798
transform -1 0 34368 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1600868798
transform 1 0 32988 0 -1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _261_
timestamp 1600868798
transform 1 0 11552 0 1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _281_
timestamp 1600868798
transform 1 0 12748 0 1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1600868798
transform 1 0 11000 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1600868798
transform 1 0 11276 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1600868798
transform 1 0 12380 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _305_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13944 0 1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_26
timestamp 1600868798
transform 1 0 13392 0 1 13720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1600868798
transform 1 0 14588 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _372_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 17072 0 1 13720
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1600868798
transform 1 0 16612 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1600868798
transform 1 0 15692 0 1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1600868798
transform 1 0 16428 0 1 13720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1600868798
transform 1 0 16704 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _365_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 18728 0 1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1600868798
transform 1 0 18360 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1600868798
transform 1 0 19556 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _298_
timestamp 1600868798
transform 1 0 20016 0 1 13720
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1600868798
transform 1 0 19924 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_112
timestamp 1600868798
transform 1 0 21304 0 1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _292_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 23512 0 1 13720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1600868798
transform 1 0 22224 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1600868798
transform 1 0 22040 0 1 13720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1600868798
transform 1 0 22316 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_135
timestamp 1600868798
transform 1 0 23420 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_4  _263_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 25076 0 1 13720
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1600868798
transform 1 0 24708 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1600868798
transform 1 0 27836 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1600868798
transform 1 0 27100 0 1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1600868798
transform 1 0 27928 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1600868798
transform 1 0 29032 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1600868798
transform 1 0 30136 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1600868798
transform 1 0 31240 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1600868798
transform 1 0 32344 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1600868798
transform -1 0 34368 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1600868798
transform 1 0 33448 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_245
timestamp 1600868798
transform 1 0 33540 0 1 13720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  _295_
timestamp 1600868798
transform 1 0 11276 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _312_
timestamp 1600868798
transform 1 0 11920 0 -1 14808
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _313_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 12472 0 1 14808
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1600868798
transform 1 0 11000 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1600868798
transform 1 0 11000 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1600868798
transform 1 0 11276 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1600868798
transform 1 0 11828 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1600868798
transform 1 0 13116 0 -1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1600868798
transform 1 0 12104 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _271_
timestamp 1600868798
transform 1 0 14772 0 1 14808
box -38 -48 1510 592
use sky130_fd_sc_hd__nor3_4  _302_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 13944 0 -1 14808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1600868798
transform 1 0 13852 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1600868798
transform 1 0 15140 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_33
timestamp 1600868798
transform 1 0 14036 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _251_
timestamp 1600868798
transform 1 0 16704 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _493_
timestamp 1600868798
transform 1 0 15508 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _517_
timestamp 1600868798
transform 1 0 16704 0 -1 14808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1600868798
transform 1 0 16612 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_52
timestamp 1600868798
transform 1 0 15784 0 -1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1600868798
transform 1 0 16520 0 -1 14808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1600868798
transform 1 0 16244 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1600868798
transform 1 0 17532 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _368_
timestamp 1600868798
transform 1 0 18820 0 1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _508_
timestamp 1600868798
transform 1 0 17900 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1600868798
transform 1 0 19464 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1600868798
transform 1 0 18820 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1600868798
transform 1 0 19372 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1600868798
transform 1 0 19556 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_78
timestamp 1600868798
transform 1 0 18176 0 1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1600868798
transform 1 0 18728 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_92
timestamp 1600868798
transform 1 0 19464 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _247_
timestamp 1600868798
transform 1 0 20200 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _289_
timestamp 1600868798
transform 1 0 21304 0 -1 14808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_6_105
timestamp 1600868798
transform 1 0 20660 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 1600868798
transform 1 0 21212 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_109
timestamp 1600868798
transform 1 0 21028 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _248_
timestamp 1600868798
transform 1 0 22316 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _293_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 23788 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _294_
timestamp 1600868798
transform 1 0 23144 0 -1 14808
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1600868798
transform 1 0 22224 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_125
timestamp 1600868798
transform 1 0 22500 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1600868798
transform 1 0 23052 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1600868798
transform 1 0 22132 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_132
timestamp 1600868798
transform 1 0 23144 0 1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1600868798
transform 1 0 23696 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _291_
timestamp 1600868798
transform 1 0 25168 0 -1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1600868798
transform 1 0 25076 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1600868798
transform 1 0 24432 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1600868798
transform 1 0 24984 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_161
timestamp 1600868798
transform 1 0 25812 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_148
timestamp 1600868798
transform 1 0 24616 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_160
timestamp 1600868798
transform 1 0 25720 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1600868798
transform 1 0 27836 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_173
timestamp 1600868798
transform 1 0 26916 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_185
timestamp 1600868798
transform 1 0 28020 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_172
timestamp 1600868798
transform 1 0 26824 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1600868798
transform 1 0 27560 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1600868798
transform 1 0 27928 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1600868798
transform 1 0 30688 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1600868798
transform 1 0 29124 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1600868798
transform 1 0 30228 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1600868798
transform 1 0 30596 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1600868798
transform 1 0 29032 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1600868798
transform 1 0 30136 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1600868798
transform 1 0 30780 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1600868798
transform 1 0 31884 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1600868798
transform 1 0 31240 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1600868798
transform 1 0 32344 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1600868798
transform -1 0 34368 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1600868798
transform -1 0 34368 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1600868798
transform 1 0 33448 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1600868798
transform 1 0 32988 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_245
timestamp 1600868798
transform 1 0 33540 0 1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _282_
timestamp 1600868798
transform 1 0 11920 0 -1 15896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1600868798
transform 1 0 11000 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1600868798
transform 1 0 11276 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1600868798
transform 1 0 11828 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1600868798
transform 1 0 13116 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _532_
timestamp 1600868798
transform 1 0 14312 0 -1 15896
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1600868798
transform 1 0 13852 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1600868798
transform 1 0 13944 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _276_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 16796 0 -1 15896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1600868798
transform 1 0 16428 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _360_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 18268 0 -1 15896
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _519_
timestamp 1600868798
transform 1 0 19556 0 -1 15896
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1600868798
transform 1 0 19464 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_72
timestamp 1600868798
transform 1 0 17624 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1600868798
transform 1 0 18176 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1600868798
transform 1 0 19096 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp 1600868798
transform 1 0 21672 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _290_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 22040 0 -1 15896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_8_142
timestamp 1600868798
transform 1 0 24064 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1600868798
transform 1 0 25076 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1600868798
transform 1 0 24800 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1600868798
transform 1 0 25168 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1600868798
transform 1 0 26272 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1600868798
transform 1 0 27376 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1600868798
transform 1 0 28480 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1600868798
transform 1 0 30688 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1600868798
transform 1 0 29584 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1600868798
transform 1 0 30780 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1600868798
transform 1 0 31884 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1600868798
transform -1 0 34368 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1600868798
transform 1 0 32988 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _296_
timestamp 1600868798
transform 1 0 11828 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1600868798
transform 1 0 11000 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1600868798
transform 1 0 11276 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_21
timestamp 1600868798
transform 1 0 12932 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _280_
timestamp 1600868798
transform 1 0 14772 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_33
timestamp 1600868798
transform 1 0 14036 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _359_
timestamp 1600868798
transform 1 0 17164 0 1 15896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1600868798
transform 1 0 16612 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1600868798
transform 1 0 15876 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1600868798
transform 1 0 16704 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1600868798
transform 1 0 17072 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _367_
timestamp 1600868798
transform 1 0 18176 0 1 15896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1600868798
transform 1 0 17808 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_91
timestamp 1600868798
transform 1 0 19372 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _287_
timestamp 1600868798
transform 1 0 20568 0 1 15896
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _506_
timestamp 1600868798
transform 1 0 19924 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_100
timestamp 1600868798
transform 1 0 20200 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1600868798
transform 1 0 21856 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _534_
timestamp 1600868798
transform 1 0 23236 0 1 15896
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1600868798
transform 1 0 22224 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1600868798
transform 1 0 22316 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1600868798
transform 1 0 23052 0 1 15896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1600868798
transform 1 0 25352 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1600868798
transform 1 0 27836 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_168
timestamp 1600868798
transform 1 0 26456 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1600868798
transform 1 0 27560 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1600868798
transform 1 0 27928 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1600868798
transform 1 0 29032 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1600868798
transform 1 0 30136 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1600868798
transform 1 0 31240 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1600868798
transform 1 0 32344 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1600868798
transform -1 0 34368 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1600868798
transform 1 0 33448 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1600868798
transform 1 0 33540 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _279_
timestamp 1600868798
transform 1 0 11828 0 -1 16984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1600868798
transform 1 0 11000 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1600868798
transform 1 0 11276 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_18
timestamp 1600868798
transform 1 0 12656 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1600868798
transform 1 0 13852 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1600868798
transform 1 0 13760 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1600868798
transform 1 0 13944 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_44
timestamp 1600868798
transform 1 0 15048 0 -1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _275_
timestamp 1600868798
transform 1 0 15416 0 -1 16984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_64
timestamp 1600868798
transform 1 0 16888 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _369_
timestamp 1600868798
transform 1 0 19556 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _370_
timestamp 1600868798
transform 1 0 18084 0 -1 16984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1600868798
transform 1 0 19464 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1600868798
transform 1 0 17992 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_86
timestamp 1600868798
transform 1 0 18912 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _285_
timestamp 1600868798
transform 1 0 21028 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_10_100
timestamp 1600868798
transform 1 0 20200 0 -1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_108
timestamp 1600868798
transform 1 0 20936 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1600868798
transform 1 0 21672 0 -1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _269_
timestamp 1600868798
transform 1 0 22040 0 -1 16984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_136
timestamp 1600868798
transform 1 0 23512 0 -1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _491_
timestamp 1600868798
transform 1 0 24248 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1600868798
transform 1 0 25076 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1600868798
transform 1 0 24524 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1600868798
transform 1 0 25168 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1600868798
transform 1 0 26272 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1600868798
transform 1 0 27376 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1600868798
transform 1 0 28480 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1600868798
transform 1 0 30688 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1600868798
transform 1 0 29584 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1600868798
transform 1 0 30780 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1600868798
transform 1 0 31884 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1600868798
transform -1 0 34368 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1600868798
transform 1 0 32988 0 -1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _278_
timestamp 1600868798
transform 1 0 11920 0 1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1600868798
transform 1 0 11000 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1600868798
transform 1 0 11276 0 1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1600868798
transform 1 0 11828 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_17
timestamp 1600868798
transform 1 0 12564 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _277_
timestamp 1600868798
transform 1 0 14772 0 1 16984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1600868798
transform 1 0 13668 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _286_
timestamp 1600868798
transform 1 0 16704 0 1 16984
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1600868798
transform 1 0 16612 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1600868798
transform 1 0 16244 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _366_
timestamp 1600868798
transform 1 0 18636 0 1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _371_
timestamp 1600868798
transform 1 0 19648 0 1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_11_76
timestamp 1600868798
transform 1 0 17992 0 1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_82
timestamp 1600868798
transform 1 0 18544 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1600868798
transform 1 0 19280 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_101
timestamp 1600868798
transform 1 0 20292 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1600868798
transform 1 0 21396 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _531_
timestamp 1600868798
transform 1 0 23512 0 1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1600868798
transform 1 0 22224 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1600868798
transform 1 0 22132 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1600868798
transform 1 0 22316 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1600868798
transform 1 0 23420 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1600868798
transform 1 0 25628 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1600868798
transform 1 0 27836 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1600868798
transform 1 0 26732 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1600868798
transform 1 0 27928 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1600868798
transform 1 0 29032 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1600868798
transform 1 0 30136 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1600868798
transform 1 0 31240 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1600868798
transform 1 0 32344 0 1 16984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1600868798
transform -1 0 34368 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1600868798
transform 1 0 33448 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_245
timestamp 1600868798
transform 1 0 33540 0 1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1600868798
transform 1 0 11000 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1600868798
transform 1 0 11276 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1600868798
transform 1 0 12380 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _533_
timestamp 1600868798
transform 1 0 13944 0 -1 18072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1600868798
transform 1 0 13852 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1600868798
transform 1 0 13484 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _270_
timestamp 1600868798
transform 1 0 16428 0 -1 18072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1600868798
transform 1 0 16060 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _249_
timestamp 1600868798
transform 1 0 18268 0 -1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _264_
timestamp 1600868798
transform 1 0 19740 0 -1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1600868798
transform 1 0 19464 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1600868798
transform 1 0 17900 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1600868798
transform 1 0 19096 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1600868798
transform 1 0 19556 0 -1 18072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _507_
timestamp 1600868798
transform 1 0 20936 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_104
timestamp 1600868798
transform 1 0 20568 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1600868798
transform 1 0 21212 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _272_
timestamp 1600868798
transform 1 0 22316 0 -1 18072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_139
timestamp 1600868798
transform 1 0 23788 0 -1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _494_
timestamp 1600868798
transform 1 0 24432 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1600868798
transform 1 0 25076 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1600868798
transform 1 0 24340 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1600868798
transform 1 0 24708 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1600868798
transform 1 0 25168 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_166
timestamp 1600868798
transform 1 0 26272 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _490_
timestamp 1600868798
transform 1 0 26548 0 -1 18072
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 28112 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1600868798
transform 1 0 27744 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_189
timestamp 1600868798
transform 1 0 28388 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1600868798
transform 1 0 30688 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1600868798
transform 1 0 29492 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1600868798
transform 1 0 30596 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1600868798
transform 1 0 30780 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1600868798
transform 1 0 31884 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1600868798
transform -1 0 34368 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1600868798
transform 1 0 32988 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1600868798
transform 1 0 11000 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1600868798
transform 1 0 11000 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1600868798
transform 1 0 11276 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1600868798
transform 1 0 12380 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1600868798
transform 1 0 11276 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1600868798
transform 1 0 12380 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1600868798
transform 1 0 13484 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1600868798
transform 1 0 14220 0 1 18072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1600868798
transform 1 0 13484 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1600868798
transform 1 0 13852 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 1600868798
transform 1 0 15048 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1600868798
transform 1 0 14680 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _492_
timestamp 1600868798
transform 1 0 14404 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _250_
timestamp 1600868798
transform 1 0 15140 0 1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1600868798
transform 1 0 15048 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1600868798
transform 1 0 13944 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1600868798
transform 1 0 16612 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_54
timestamp 1600868798
transform 1 0 15968 0 1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1600868798
transform 1 0 16520 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1600868798
transform 1 0 16704 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_70
timestamp 1600868798
transform 1 0 17440 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1600868798
transform 1 0 16152 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_68
timestamp 1600868798
transform 1 0 17256 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _315_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 18268 0 -1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _518_
timestamp 1600868798
transform 1 0 17716 0 1 18072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1600868798
transform 1 0 19464 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_76
timestamp 1600868798
transform 1 0 17992 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1600868798
transform 1 0 19096 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1600868798
transform 1 0 19556 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _274_
timestamp 1600868798
transform 1 0 20568 0 1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _496_
timestamp 1600868798
transform 1 0 21580 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _529_
timestamp 1600868798
transform 1 0 19924 0 -1 19160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_13_96
timestamp 1600868798
transform 1 0 19832 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_111
timestamp 1600868798
transform 1 0 21212 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1600868798
transform 1 0 21856 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _314_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 22408 0 -1 19160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_4  _530_
timestamp 1600868798
transform 1 0 23052 0 1 18072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1600868798
transform 1 0 22224 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1600868798
transform 1 0 22316 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_120
timestamp 1600868798
transform 1 0 22040 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1600868798
transform 1 0 23972 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _495_
timestamp 1600868798
transform 1 0 24340 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 26180 0 -1 19160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1600868798
transform 1 0 25076 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1600868798
transform 1 0 25168 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1600868798
transform 1 0 26272 0 1 18072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1600868798
transform 1 0 24616 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1600868798
transform 1 0 24984 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1600868798
transform 1 0 25168 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_162
timestamp 1600868798
transform 1 0 25904 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _425_
timestamp 1600868798
transform 1 0 27192 0 -1 19160
box -38 -48 1234 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1600868798
transform 1 0 27928 0 1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 26456 0 1 18072
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1600868798
transform 1 0 27836 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1600868798
transform 1 0 27468 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1600868798
transform 1 0 26824 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_189
timestamp 1600868798
transform 1 0 28388 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 28756 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 29400 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1600868798
transform 1 0 30688 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_191
timestamp 1600868798
transform 1 0 28572 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_203
timestamp 1600868798
transform 1 0 29676 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_196
timestamp 1600868798
transform 1 0 29032 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_203
timestamp 1600868798
transform 1 0 29676 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1600868798
transform 1 0 30412 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1600868798
transform 1 0 30780 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1600868798
transform 1 0 31884 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1600868798
transform 1 0 30780 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1600868798
transform 1 0 31884 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1600868798
transform -1 0 34368 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1600868798
transform -1 0 34368 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1600868798
transform 1 0 33448 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1600868798
transform 1 0 32988 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1600868798
transform 1 0 33356 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_245
timestamp 1600868798
transform 1 0 33540 0 1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1600868798
transform 1 0 32988 0 -1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1600868798
transform 1 0 11000 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1600868798
transform 1 0 11276 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1600868798
transform 1 0 12380 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _322_
timestamp 1600868798
transform 1 0 15140 0 1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _502_
timestamp 1600868798
transform 1 0 14312 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_27
timestamp 1600868798
transform 1 0 13484 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_35
timestamp 1600868798
transform 1 0 14220 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1600868798
transform 1 0 14588 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1600868798
transform 1 0 16612 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1600868798
transform 1 0 15968 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1600868798
transform 1 0 16520 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1600868798
transform 1 0 16704 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1600868798
transform 1 0 17440 0 1 19160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _259_
timestamp 1600868798
transform 1 0 17624 0 1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _357_
timestamp 1600868798
transform 1 0 18820 0 1 19160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1600868798
transform 1 0 18452 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1600868798
transform 1 0 19464 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _503_
timestamp 1600868798
transform 1 0 19832 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_99
timestamp 1600868798
transform 1 0 20108 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_111
timestamp 1600868798
transform 1 0 21212 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1600868798
transform 1 0 21948 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _273_
timestamp 1600868798
transform 1 0 22316 0 1 19160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1600868798
transform 1 0 22224 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1600868798
transform 1 0 23788 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1600868798
transform 1 0 25536 0 1 19160
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1600868798
transform 1 0 24892 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1600868798
transform 1 0 25168 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_165
timestamp 1600868798
transform 1 0 26180 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 27928 0 1 19160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1600868798
transform 1 0 27836 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1600868798
transform 1 0 27284 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1600868798
transform 1 0 29952 0 1 19160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1600868798
transform 1 0 29584 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_219
timestamp 1600868798
transform 1 0 31148 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_231
timestamp 1600868798
transform 1 0 32252 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1600868798
transform -1 0 34368 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1600868798
transform 1 0 33448 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1600868798
transform 1 0 33356 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_245
timestamp 1600868798
transform 1 0 33540 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1600868798
transform 1 0 11000 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1600868798
transform 1 0 11276 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1600868798
transform 1 0 12380 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1600868798
transform 1 0 13944 0 -1 20248
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1600868798
transform 1 0 13852 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1600868798
transform 1 0 13484 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _355_
timestamp 1600868798
transform 1 0 16428 0 -1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1600868798
transform 1 0 16060 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_66
timestamp 1600868798
transform 1 0 17072 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _358_
timestamp 1600868798
transform 1 0 17624 0 -1 20248
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1600868798
transform 1 0 19464 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1600868798
transform 1 0 18820 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1600868798
transform 1 0 19372 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1600868798
transform 1 0 19556 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _266_
timestamp 1600868798
transform 1 0 21396 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 1600868798
transform 1 0 20660 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _252_
timestamp 1600868798
transform 1 0 22960 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_122
timestamp 1600868798
transform 1 0 22224 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_139
timestamp 1600868798
transform 1 0 23788 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1600868798
transform 1 0 24432 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1600868798
transform 1 0 25260 0 -1 20248
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1600868798
transform 1 0 25076 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1600868798
transform 1 0 24340 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1600868798
transform 1 0 24708 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1600868798
transform 1 0 25168 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 27284 0 -1 20248
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 28112 0 -1 20248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1600868798
transform 1 0 26916 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1600868798
transform 1 0 27744 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1600868798
transform 1 0 29492 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1600868798
transform 1 0 30688 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_191
timestamp 1600868798
transform 1 0 28572 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1600868798
transform 1 0 29308 0 -1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1600868798
transform 1 0 29860 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1600868798
transform 1 0 30596 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1600868798
transform 1 0 30780 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1600868798
transform 1 0 31884 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1600868798
transform -1 0 34368 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1600868798
transform 1 0 32988 0 -1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1600868798
transform 1 0 11000 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1600868798
transform 1 0 11276 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1600868798
transform 1 0 12380 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _356_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 14404 0 1 20248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1600868798
transform 1 0 13484 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1600868798
transform 1 0 14220 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _258_
timestamp 1600868798
transform 1 0 16704 0 1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1600868798
transform 1 0 16612 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_54
timestamp 1600868798
transform 1 0 15968 0 1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1600868798
transform 1 0 16520 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1600868798
transform 1 0 17532 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _522_
timestamp 1600868798
transform 1 0 17992 0 1 20248
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1600868798
transform 1 0 17900 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _262_
timestamp 1600868798
transform 1 0 21028 0 1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_99
timestamp 1600868798
transform 1 0 20108 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1600868798
transform 1 0 20844 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1600868798
transform 1 0 21856 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _267_
timestamp 1600868798
transform 1 0 22316 0 1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _487_
timestamp 1600868798
transform 1 0 23512 0 1 20248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1600868798
transform 1 0 22224 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1600868798
transform 1 0 23144 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1600868798
transform 1 0 25444 0 1 20248
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1600868798
transform 1 0 25076 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1600868798
transform 1 0 26824 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1600868798
transform 1 0 27836 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_168
timestamp 1600868798
transform 1 0 26456 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1600868798
transform 1 0 27468 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1600868798
transform 1 0 27928 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 29584 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_196
timestamp 1600868798
transform 1 0 29032 0 1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_206
timestamp 1600868798
transform 1 0 29952 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_218
timestamp 1600868798
transform 1 0 31056 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_230
timestamp 1600868798
transform 1 0 32160 0 1 20248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1600868798
transform -1 0 34368 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1600868798
transform 1 0 33448 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1600868798
transform 1 0 33264 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_245
timestamp 1600868798
transform 1 0 33540 0 1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1600868798
transform 1 0 11000 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1600868798
transform 1 0 11276 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1600868798
transform 1 0 12380 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _321_
timestamp 1600868798
transform 1 0 15140 0 -1 21336
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1600868798
transform 1 0 13852 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1600868798
transform 1 0 13484 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1600868798
transform 1 0 13944 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_44
timestamp 1600868798
transform 1 0 15048 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _306_
timestamp 1600868798
transform 1 0 16796 0 -1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1600868798
transform 1 0 16428 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _311_
timestamp 1600868798
transform 1 0 17992 0 -1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _319_
timestamp 1600868798
transform 1 0 19556 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1600868798
transform 1 0 19464 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_72
timestamp 1600868798
transform 1 0 17624 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1600868798
transform 1 0 18820 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1600868798
transform 1 0 19372 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _484_
timestamp 1600868798
transform 1 0 20844 0 -1 21336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_18_100
timestamp 1600868798
transform 1 0 20200 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_106
timestamp 1600868798
transform 1 0 20752 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _436_
timestamp 1600868798
transform 1 0 22500 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _473_
timestamp 1600868798
transform 1 0 23696 0 -1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1600868798
transform 1 0 22132 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_132
timestamp 1600868798
transform 1 0 23144 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1600868798
transform 1 0 25168 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1600868798
transform 1 0 25076 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1600868798
transform 1 0 24524 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_161
timestamp 1600868798
transform 1 0 25812 0 -1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1600868798
transform 1 0 26548 0 -1 21336
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1600868798
transform 1 0 27928 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1600868798
transform 1 0 27560 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_188
timestamp 1600868798
transform 1 0 28296 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1600868798
transform 1 0 29584 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1600868798
transform 1 0 28664 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1600868798
transform 1 0 30688 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_195
timestamp 1600868798
transform 1 0 28940 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1600868798
transform 1 0 29492 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1600868798
transform 1 0 30228 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1600868798
transform 1 0 30596 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1600868798
transform 1 0 30780 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1600868798
transform 1 0 31884 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1600868798
transform -1 0 34368 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1600868798
transform 1 0 32988 0 -1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1600868798
transform 1 0 11000 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1600868798
transform 1 0 11000 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1600868798
transform 1 0 11276 0 1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1600868798
transform 1 0 12380 0 1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1600868798
transform 1 0 11276 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1600868798
transform 1 0 12380 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1600868798
transform 1 0 13484 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_33
timestamp 1600868798
transform 1 0 14036 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1600868798
transform 1 0 13484 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1600868798
transform 1 0 13852 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _501_
timestamp 1600868798
transform 1 0 14128 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _348_
timestamp 1600868798
transform 1 0 13944 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1600868798
transform 1 0 14772 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1600868798
transform 1 0 14956 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_37
timestamp 1600868798
transform 1 0 14404 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _347_
timestamp 1600868798
transform 1 0 15140 0 -1 22424
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _323_
timestamp 1600868798
transform 1 0 15048 0 1 21336
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  _320_
timestamp 1600868798
transform 1 0 16796 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1600868798
transform 1 0 16612 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1600868798
transform 1 0 16244 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1600868798
transform 1 0 16704 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_59
timestamp 1600868798
transform 1 0 16428 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_71
timestamp 1600868798
transform 1 0 17532 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _310_
timestamp 1600868798
transform 1 0 19740 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _316_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 17808 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _318_
timestamp 1600868798
transform 1 0 17992 0 1 21336
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1600868798
transform 1 0 19464 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_72
timestamp 1600868798
transform 1 0 17624 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_89
timestamp 1600868798
transform 1 0 19188 0 1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1600868798
transform 1 0 18636 0 -1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1600868798
transform 1 0 19372 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1600868798
transform 1 0 19556 0 -1 22424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _256_
timestamp 1600868798
transform 1 0 20016 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _373_
timestamp 1600868798
transform 1 0 21212 0 1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _435_
timestamp 1600868798
transform 1 0 21212 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1600868798
transform 1 0 19924 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1600868798
transform 1 0 20844 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1600868798
transform 1 0 21856 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_104
timestamp 1600868798
transform 1 0 20568 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1600868798
transform 1 0 21120 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _375_
timestamp 1600868798
transform 1 0 22868 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _426_
timestamp 1600868798
transform 1 0 22408 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _441_
timestamp 1600868798
transform 1 0 23604 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_4  _476_
timestamp 1600868798
transform 1 0 24064 0 1 21336
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1600868798
transform 1 0 22224 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1600868798
transform 1 0 22316 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1600868798
transform 1 0 23696 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 1600868798
transform 1 0 22040 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_133
timestamp 1600868798
transform 1 0 23236 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _469_
timestamp 1600868798
transform 1 0 25168 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1600868798
transform 1 0 26272 0 -1 22424
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1600868798
transform 1 0 25076 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_155
timestamp 1600868798
transform 1 0 25260 0 1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_146
timestamp 1600868798
transform 1 0 24432 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1600868798
transform 1 0 24984 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1600868798
transform 1 0 25812 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_165
timestamp 1600868798
transform 1 0 26180 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1600868798
transform 1 0 27928 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1600868798
transform 1 0 26640 0 1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1600868798
transform 1 0 27836 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_167
timestamp 1600868798
transform 1 0 26364 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1600868798
transform 1 0 27284 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1600868798
transform 1 0 28204 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_184
timestamp 1600868798
transform 1 0 27928 0 -1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _427_
timestamp 1600868798
transform 1 0 29216 0 1 21336
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1600868798
transform 1 0 28572 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1600868798
transform 1 0 29308 0 -1 22424
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1600868798
transform 1 0 28664 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1600868798
transform 1 0 30688 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1600868798
transform 1 0 28848 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_195
timestamp 1600868798
transform 1 0 28940 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1600868798
transform 1 0 30320 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _402_
timestamp 1600868798
transform 1 0 31148 0 1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1600868798
transform 1 0 30780 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1600868798
transform 1 0 30780 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_231
timestamp 1600868798
transform 1 0 32252 0 1 21336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_222
timestamp 1600868798
transform 1 0 31424 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_234
timestamp 1600868798
transform 1 0 32528 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1600868798
transform -1 0 34368 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1600868798
transform -1 0 34368 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1600868798
transform 1 0 33448 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 1600868798
transform 1 0 33356 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_245
timestamp 1600868798
transform 1 0 33540 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_246
timestamp 1600868798
transform 1 0 33632 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_250
timestamp 1600868798
transform 1 0 34000 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _524_
timestamp 1600868798
transform 1 0 13116 0 1 22424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1600868798
transform 1 0 11000 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1600868798
transform 1 0 11276 0 1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1600868798
transform 1 0 12380 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1600868798
transform 1 0 15232 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _257_
timestamp 1600868798
transform 1 0 16796 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _353_
timestamp 1600868798
transform 1 0 15600 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1600868798
transform 1 0 16612 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1600868798
transform 1 0 16244 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1600868798
transform 1 0 16704 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _317_
timestamp 1600868798
transform 1 0 18360 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _326_
timestamp 1600868798
transform 1 0 19556 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_72
timestamp 1600868798
transform 1 0 17624 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1600868798
transform 1 0 19188 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _474_
timestamp 1600868798
transform 1 0 21028 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_100
timestamp 1600868798
transform 1 0 20200 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_108
timestamp 1600868798
transform 1 0 20936 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1600868798
transform 1 0 21856 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _434_
timestamp 1600868798
transform 1 0 22316 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _475_
timestamp 1600868798
transform 1 0 23604 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1600868798
transform 1 0 22224 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1600868798
transform 1 0 23144 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1600868798
transform 1 0 23512 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _424_
timestamp 1600868798
transform 1 0 24892 0 1 22424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1600868798
transform 1 0 24432 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1600868798
transform 1 0 24800 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1600868798
transform 1 0 26088 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _472_
timestamp 1600868798
transform 1 0 26456 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1600868798
transform 1 0 27836 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1600868798
transform 1 0 27100 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_184
timestamp 1600868798
transform 1 0 27928 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1600868798
transform 1 0 28848 0 1 22424
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1600868798
transform 1 0 28664 0 1 22424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_212
timestamp 1600868798
transform 1 0 30504 0 1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_224
timestamp 1600868798
transform 1 0 31608 0 1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1600868798
transform 1 0 32712 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1600868798
transform -1 0 34368 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1600868798
transform 1 0 33448 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_245
timestamp 1600868798
transform 1 0 33540 0 1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1600868798
transform 1 0 11000 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1600868798
transform 1 0 11276 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1600868798
transform 1 0 12380 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _354_
timestamp 1600868798
transform 1 0 14128 0 -1 23512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1600868798
transform 1 0 13852 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1600868798
transform 1 0 13484 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1600868798
transform 1 0 13944 0 -1 23512
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _324_
timestamp 1600868798
transform 1 0 16796 0 -1 23512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_22_51
timestamp 1600868798
transform 1 0 15692 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _308_
timestamp 1600868798
transform 1 0 18452 0 -1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _309_
timestamp 1600868798
transform 1 0 19556 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1600868798
transform 1 0 19464 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_77
timestamp 1600868798
transform 1 0 18084 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1600868798
transform 1 0 19096 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _377_
timestamp 1600868798
transform 1 0 20752 0 -1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _437_
timestamp 1600868798
transform 1 0 21856 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1600868798
transform 1 0 20384 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1600868798
transform 1 0 21396 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1600868798
transform 1 0 21764 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _442_
timestamp 1600868798
transform 1 0 23052 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1600868798
transform 1 0 22684 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_140
timestamp 1600868798
transform 1 0 23880 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _423_
timestamp 1600868798
transform 1 0 25168 0 -1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1600868798
transform 1 0 25076 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1600868798
transform 1 0 24984 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_161
timestamp 1600868798
transform 1 0 25812 0 -1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_4  _374_
timestamp 1600868798
transform 1 0 26364 0 -1 23512
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  _376_
timestamp 1600868798
transform 1 0 27928 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1600868798
transform 1 0 27560 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _401_
timestamp 1600868798
transform 1 0 29124 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1600868798
transform 1 0 30688 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_193
timestamp 1600868798
transform 1 0 28756 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1600868798
transform 1 0 29952 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1600868798
transform 1 0 30780 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_219
timestamp 1600868798
transform 1 0 31148 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_231
timestamp 1600868798
transform 1 0 32252 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1600868798
transform -1 0 34368 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1600868798
transform 1 0 33356 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1600868798
transform 1 0 11000 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1600868798
transform 1 0 11276 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1600868798
transform 1 0 12380 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _349_
timestamp 1600868798
transform 1 0 14680 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1600868798
transform 1 0 13484 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp 1600868798
transform 1 0 14588 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1600868798
transform 1 0 16612 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_52
timestamp 1600868798
transform 1 0 15784 0 1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1600868798
transform 1 0 16520 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1600868798
transform 1 0 16704 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _328_
timestamp 1600868798
transform 1 0 17992 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_4  _439_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 19004 0 1 23512
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1600868798
transform 1 0 17808 0 1 23512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1600868798
transform 1 0 18636 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _440_
timestamp 1600868798
transform 1 0 21028 0 1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_105
timestamp 1600868798
transform 1 0 20660 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1600868798
transform 1 0 21856 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _327_
timestamp 1600868798
transform 1 0 22316 0 1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _486_
timestamp 1600868798
transform 1 0 23604 0 1 23512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1600868798
transform 1 0 22224 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1600868798
transform 1 0 23144 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_136
timestamp 1600868798
transform 1 0 23512 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _400_
timestamp 1600868798
transform 1 0 26272 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1600868798
transform 1 0 25168 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1600868798
transform 1 0 28204 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1600868798
transform 1 0 27836 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1600868798
transform 1 0 26916 0 1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1600868798
transform 1 0 27652 0 1 23512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1600868798
transform 1 0 27928 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1600868798
transform 1 0 28480 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1600868798
transform 1 0 30228 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1600868798
transform 1 0 28848 0 1 23512
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1600868798
transform 1 0 29860 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1600868798
transform 1 0 31240 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1600868798
transform 1 0 30872 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_227
timestamp 1600868798
transform 1 0 31884 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1600868798
transform -1 0 34368 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1600868798
transform 1 0 33448 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_239
timestamp 1600868798
transform 1 0 32988 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1600868798
transform 1 0 33356 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_245
timestamp 1600868798
transform 1 0 33540 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _351_
timestamp 1600868798
transform 1 0 12840 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1600868798
transform 1 0 11000 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1600868798
transform 1 0 11276 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1600868798
transform 1 0 12380 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_19
timestamp 1600868798
transform 1 0 12748 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _350_
timestamp 1600868798
transform 1 0 14404 0 -1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1600868798
transform 1 0 13852 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1600868798
transform 1 0 13484 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1600868798
transform 1 0 13944 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1600868798
transform 1 0 14312 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_46
timestamp 1600868798
transform 1 0 15232 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _331_
timestamp 1600868798
transform 1 0 16520 0 -1 24600
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1600868798
transform 1 0 16336 0 -1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _307_
timestamp 1600868798
transform 1 0 18452 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _330_
timestamp 1600868798
transform 1 0 19556 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1600868798
transform 1 0 19464 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1600868798
transform 1 0 18084 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1600868798
transform 1 0 19096 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _438_
timestamp 1600868798
transform 1 0 21856 0 -1 24600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_24_100
timestamp 1600868798
transform 1 0 20200 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_112
timestamp 1600868798
transform 1 0 21304 0 -1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _406_
timestamp 1600868798
transform 1 0 23512 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_132
timestamp 1600868798
transform 1 0 23144 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _481_
timestamp 1600868798
transform 1 0 25168 0 -1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1600868798
transform 1 0 25076 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1600868798
transform 1 0 24616 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1600868798
transform 1 0 24984 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_163
timestamp 1600868798
transform 1 0 25996 0 -1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _444_
timestamp 1600868798
transform 1 0 26916 0 -1 24600
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_4  _449_
timestamp 1600868798
transform 1 0 28480 0 -1 24600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_24_171
timestamp 1600868798
transform 1 0 26732 0 -1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1600868798
transform 1 0 28112 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1600868798
transform 1 0 30044 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1600868798
transform 1 0 30688 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1600868798
transform 1 0 29676 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1600868798
transform 1 0 30320 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1600868798
transform 1 0 31976 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1600868798
transform 1 0 30964 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1600868798
transform 1 0 30780 0 -1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_224
timestamp 1600868798
transform 1 0 31608 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_232
timestamp 1600868798
transform 1 0 32344 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1600868798
transform -1 0 34368 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_244
timestamp 1600868798
transform 1 0 33448 0 -1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_250
timestamp 1600868798
transform 1 0 34000 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1600868798
transform 1 0 11000 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1600868798
transform 1 0 11276 0 1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1600868798
transform 1 0 12380 0 1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _352_
timestamp 1600868798
transform 1 0 14128 0 1 24600
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1600868798
transform 1 0 13484 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1600868798
transform 1 0 14036 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _325_
timestamp 1600868798
transform 1 0 16704 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1600868798
transform 1 0 16612 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1600868798
transform 1 0 15692 0 1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1600868798
transform 1 0 16428 0 1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_71
timestamp 1600868798
transform 1 0 17532 0 1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_4  _383_
timestamp 1600868798
transform 1 0 19096 0 1 24600
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1600868798
transform 1 0 18636 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1600868798
transform 1 0 19004 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _471_
timestamp 1600868798
transform 1 0 21212 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_106
timestamp 1600868798
transform 1 0 20752 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_110
timestamp 1600868798
transform 1 0 21120 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1600868798
transform 1 0 21856 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _410_
timestamp 1600868798
transform 1 0 23420 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _452_
timestamp 1600868798
transform 1 0 22316 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1600868798
transform 1 0 22224 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1600868798
transform 1 0 22960 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_134
timestamp 1600868798
transform 1 0 23328 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_142
timestamp 1600868798
transform 1 0 24064 0 1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _443_
timestamp 1600868798
transform 1 0 26180 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _461_
timestamp 1600868798
transform 1 0 25168 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_161
timestamp 1600868798
transform 1 0 25812 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _477_
timestamp 1600868798
transform 1 0 27928 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1600868798
transform 1 0 27836 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_172
timestamp 1600868798
transform 1 0 26824 0 1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1600868798
transform 1 0 27560 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1600868798
transform 1 0 29400 0 1 24600
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1600868798
transform 1 0 28572 0 1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_199
timestamp 1600868798
transform 1 0 29308 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1600868798
transform 1 0 31424 0 1 24600
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1600868798
transform 1 0 31056 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1600868798
transform -1 0 34368 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1600868798
transform 1 0 33448 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1600868798
transform 1 0 33080 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_245
timestamp 1600868798
transform 1 0 33540 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1600868798
transform 1 0 11000 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1600868798
transform 1 0 11000 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1600868798
transform 1 0 11276 0 -1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1600868798
transform 1 0 12380 0 -1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1600868798
transform 1 0 11276 0 1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1600868798
transform 1 0 12380 0 1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _337_
timestamp 1600868798
transform 1 0 14404 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _500_
timestamp 1600868798
transform 1 0 13760 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _525_
timestamp 1600868798
transform 1 0 13944 0 -1 25688
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1600868798
transform 1 0 13852 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1600868798
transform 1 0 13484 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1600868798
transform 1 0 13484 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1600868798
transform 1 0 14036 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_44
timestamp 1600868798
transform 1 0 15048 0 1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _333_
timestamp 1600868798
transform 1 0 17072 0 -1 25688
box -38 -48 1326 592
use sky130_fd_sc_hd__a32o_4  _335_
timestamp 1600868798
transform 1 0 16704 0 1 25688
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_4  _345_
timestamp 1600868798
transform 1 0 15600 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1600868798
transform 1 0 16612 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_55
timestamp 1600868798
transform 1 0 16060 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_63
timestamp 1600868798
transform 1 0 16796 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1600868798
transform 1 0 16244 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _385_
timestamp 1600868798
transform 1 0 19372 0 1 25688
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _446_
timestamp 1600868798
transform 1 0 19556 0 -1 25688
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1600868798
transform 1 0 19464 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1600868798
transform 1 0 18360 0 -1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_79
timestamp 1600868798
transform 1 0 18268 0 1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _384_
timestamp 1600868798
transform 1 0 20936 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _445_
timestamp 1600868798
transform 1 0 21120 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1600868798
transform 1 0 20752 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1600868798
transform 1 0 21948 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_104
timestamp 1600868798
transform 1 0 20568 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1600868798
transform 1 0 21764 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1600868798
transform 1 0 22132 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1600868798
transform 1 0 22224 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _488_
timestamp 1600868798
transform 1 0 22316 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _447_
timestamp 1600868798
transform 1 0 22316 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1600868798
transform 1 0 23144 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1600868798
transform 1 0 23144 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _468_
timestamp 1600868798
transform 1 0 23512 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_140
timestamp 1600868798
transform 1 0 23880 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_143
timestamp 1600868798
transform 1 0 24156 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _386_
timestamp 1600868798
transform 1 0 23972 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _433_
timestamp 1600868798
transform 1 0 25536 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _482_
timestamp 1600868798
transform 1 0 25536 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1600868798
transform 1 0 25076 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1600868798
transform 1 0 24892 0 -1 25688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1600868798
transform 1 0 25168 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1600868798
transform 1 0 24616 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1600868798
transform 1 0 25352 0 1 25688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1600868798
transform 1 0 27376 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_167
timestamp 1600868798
transform 1 0 26364 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_178
timestamp 1600868798
transform 1 0 27376 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1600868798
transform 1 0 26364 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _451_
timestamp 1600868798
transform 1 0 26732 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _448_
timestamp 1600868798
transform 1 0 26732 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1600868798
transform 1 0 27928 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1600868798
transform 1 0 27744 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1600868798
transform 1 0 27836 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1600868798
transform 1 0 28296 0 1 25688
box -38 -48 1050 592
use sky130_fd_sc_hd__a21bo_4  _483_
timestamp 1600868798
transform 1 0 28112 0 -1 25688
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1600868798
transform 1 0 29676 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1600868798
transform 1 0 29676 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1600868798
transform 1 0 30688 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_199
timestamp 1600868798
transform 1 0 29308 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1600868798
transform 1 0 30044 0 -1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1600868798
transform 1 0 30596 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1600868798
transform 1 0 29308 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1600868798
transform 1 0 30320 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_214
timestamp 1600868798
transform 1 0 30688 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1600868798
transform 1 0 32160 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1600868798
transform 1 0 30780 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1600868798
transform 1 0 30780 0 -1 25688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1600868798
transform 1 0 31792 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1600868798
transform 1 0 31792 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1600868798
transform 1 0 32436 0 -1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_222
timestamp 1600868798
transform 1 0 31424 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1600868798
transform 1 0 32068 0 1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1600868798
transform -1 0 34368 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1600868798
transform -1 0 34368 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1600868798
transform 1 0 33448 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1600868798
transform 1 0 33540 0 -1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_241
timestamp 1600868798
transform 1 0 33172 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_245
timestamp 1600868798
transform 1 0 33540 0 1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1600868798
transform 1 0 11000 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1600868798
transform 1 0 11276 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1600868798
transform 1 0 12380 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _336_
timestamp 1600868798
transform 1 0 14588 0 -1 26776
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1600868798
transform 1 0 13852 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1600868798
transform 1 0 13484 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_32
timestamp 1600868798
transform 1 0 13944 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_38
timestamp 1600868798
transform 1 0 14496 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _332_
timestamp 1600868798
transform 1 0 17072 0 -1 26776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1600868798
transform 1 0 15876 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1600868798
transform 1 0 16980 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _458_
timestamp 1600868798
transform 1 0 19556 0 -1 26776
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1600868798
transform 1 0 19464 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1600868798
transform 1 0 18360 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1600868798
transform 1 0 21120 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _457_
timestamp 1600868798
transform 1 0 22316 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _460_
timestamp 1600868798
transform 1 0 23512 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_122
timestamp 1600868798
transform 1 0 22224 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_132
timestamp 1600868798
transform 1 0 23144 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _462_
timestamp 1600868798
transform 1 0 26088 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1600868798
transform 1 0 25076 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1600868798
transform 1 0 24340 0 -1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1600868798
transform 1 0 25168 0 -1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_162
timestamp 1600868798
transform 1 0 25904 0 -1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _453_
timestamp 1600868798
transform 1 0 28480 0 -1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _489_
timestamp 1600868798
transform 1 0 27284 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1600868798
transform 1 0 26916 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_186
timestamp 1600868798
transform 1 0 28112 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1600868798
transform 1 0 29492 0 -1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1600868798
transform 1 0 30688 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1600868798
transform 1 0 29124 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1600868798
transform 1 0 30136 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1600868798
transform 1 0 30780 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1600868798
transform 1 0 31424 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1600868798
transform 1 0 31056 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1600868798
transform 1 0 31700 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1600868798
transform 1 0 32804 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1600868798
transform -1 0 34368 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1600868798
transform 1 0 33908 0 -1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1600868798
transform 1 0 11000 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1600868798
transform 1 0 11276 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1600868798
transform 1 0 12380 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _338_
timestamp 1600868798
transform 1 0 14220 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1600868798
transform 1 0 13484 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_44
timestamp 1600868798
transform 1 0 15048 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _334_
timestamp 1600868798
transform 1 0 15416 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _341_
timestamp 1600868798
transform 1 0 16796 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1600868798
transform 1 0 16612 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1600868798
transform 1 0 16244 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1600868798
transform 1 0 16704 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _340_
timestamp 1600868798
transform 1 0 18268 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1600868798
transform 1 0 17900 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_88
timestamp 1600868798
transform 1 0 19096 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _432_
timestamp 1600868798
transform 1 0 20752 0 1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_29_100
timestamp 1600868798
transform 1 0 20200 0 1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1600868798
transform 1 0 21396 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _459_
timestamp 1600868798
transform 1 0 22408 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _464_
timestamp 1600868798
transform 1 0 23972 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1600868798
transform 1 0 22224 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1600868798
transform 1 0 22132 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1600868798
transform 1 0 22316 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_133
timestamp 1600868798
transform 1 0 23236 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _465_
timestamp 1600868798
transform 1 0 25720 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_150
timestamp 1600868798
transform 1 0 24800 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1600868798
transform 1 0 25536 0 1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1600868798
transform 1 0 28204 0 1 26776
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1600868798
transform 1 0 27836 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1600868798
transform 1 0 26548 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1600868798
transform 1 0 27652 0 1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1600868798
transform 1 0 27928 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _392_
timestamp 1600868798
transform 1 0 30228 0 1 26776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1600868798
transform 1 0 29860 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_222
timestamp 1600868798
transform 1 0 31424 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 1600868798
transform 1 0 32528 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1600868798
transform -1 0 34368 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1600868798
transform 1 0 33448 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 1600868798
transform 1 0 33264 0 1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_245
timestamp 1600868798
transform 1 0 33540 0 1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1600868798
transform 1 0 11000 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1600868798
transform 1 0 11276 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1600868798
transform 1 0 12380 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _339_
timestamp 1600868798
transform 1 0 14036 0 -1 27864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1600868798
transform 1 0 13852 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1600868798
transform 1 0 13484 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1600868798
transform 1 0 13944 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _346_
timestamp 1600868798
transform 1 0 16796 0 -1 27864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_30_50
timestamp 1600868798
transform 1 0 15600 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_62
timestamp 1600868798
transform 1 0 16704 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1600868798
transform 1 0 19464 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1600868798
transform 1 0 18360 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1600868798
transform 1 0 19556 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _412_
timestamp 1600868798
transform 1 0 21488 0 -1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _430_
timestamp 1600868798
transform 1 0 20016 0 -1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1600868798
transform 1 0 19924 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_107
timestamp 1600868798
transform 1 0 20844 0 -1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_113
timestamp 1600868798
transform 1 0 21396 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _394_
timestamp 1600868798
transform 1 0 24064 0 -1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _428_
timestamp 1600868798
transform 1 0 22684 0 -1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1600868798
transform 1 0 22316 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_136
timestamp 1600868798
transform 1 0 23512 0 -1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _399_
timestamp 1600868798
transform 1 0 25352 0 -1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1600868798
transform 1 0 25076 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1600868798
transform 1 0 24708 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1600868798
transform 1 0 25168 0 -1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1600868798
transform 1 0 25996 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _420_
timestamp 1600868798
transform 1 0 27744 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _454_
timestamp 1600868798
transform 1 0 26364 0 -1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_176
timestamp 1600868798
transform 1 0 27192 0 -1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _391_
timestamp 1600868798
transform 1 0 29216 0 -1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1600868798
transform 1 0 30688 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_194
timestamp 1600868798
transform 1 0 28848 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_205
timestamp 1600868798
transform 1 0 29860 0 -1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1600868798
transform 1 0 30596 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1600868798
transform 1 0 30780 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1600868798
transform 1 0 31884 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1600868798
transform -1 0 34368 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1600868798
transform 1 0 32988 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1600868798
transform 1 0 11000 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1600868798
transform 1 0 11276 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1600868798
transform 1 0 12380 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _528_
timestamp 1600868798
transform 1 0 13484 0 1 27864
box -38 -48 2154 592
use sky130_fd_sc_hd__a32o_4  _344_
timestamp 1600868798
transform 1 0 16704 0 1 27864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1600868798
transform 1 0 16612 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_50
timestamp 1600868798
transform 1 0 15600 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1600868798
transform 1 0 16336 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _253_
timestamp 1600868798
transform 1 0 18728 0 1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1600868798
transform 1 0 18268 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_83
timestamp 1600868798
transform 1 0 18636 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1600868798
transform 1 0 19556 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _329_
timestamp 1600868798
transform 1 0 19924 0 1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _414_
timestamp 1600868798
transform 1 0 21212 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_106
timestamp 1600868798
transform 1 0 20752 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_110
timestamp 1600868798
transform 1 0 21120 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1600868798
transform 1 0 21856 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _413_
timestamp 1600868798
transform 1 0 22316 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _456_
timestamp 1600868798
transform 1 0 23328 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1600868798
transform 1 0 22224 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1600868798
transform 1 0 22960 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_141
timestamp 1600868798
transform 1 0 23972 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _429_
timestamp 1600868798
transform 1 0 26272 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _485_
timestamp 1600868798
transform 1 0 24616 0 1 27864
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_31_147
timestamp 1600868798
transform 1 0 24524 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_162
timestamp 1600868798
transform 1 0 25904 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _421_
timestamp 1600868798
transform 1 0 28480 0 1 27864
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1600868798
transform 1 0 27836 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_173
timestamp 1600868798
transform 1 0 26916 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1600868798
transform 1 0 27652 0 1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp 1600868798
transform 1 0 27928 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_203
timestamp 1600868798
transform 1 0 29676 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_215
timestamp 1600868798
transform 1 0 30780 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_227
timestamp 1600868798
transform 1 0 31884 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1600868798
transform -1 0 34368 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1600868798
transform 1 0 33448 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_239
timestamp 1600868798
transform 1 0 32988 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1600868798
transform 1 0 33356 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_245
timestamp 1600868798
transform 1 0 33540 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1600868798
transform 1 0 11000 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1600868798
transform 1 0 11276 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1600868798
transform 1 0 12380 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _497_
timestamp 1600868798
transform 1 0 14404 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _527_
timestamp 1600868798
transform 1 0 15324 0 -1 28952
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1600868798
transform 1 0 13852 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1600868798
transform 1 0 13484 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1600868798
transform 1 0 13944 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1600868798
transform 1 0 14312 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_40
timestamp 1600868798
transform 1 0 14680 0 -1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_46
timestamp 1600868798
transform 1 0 15232 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1600868798
transform 1 0 17440 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _343_
timestamp 1600868798
transform 1 0 17808 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1600868798
transform 1 0 19464 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_81
timestamp 1600868798
transform 1 0 18452 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1600868798
transform 1 0 19188 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1600868798
transform 1 0 19556 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _378_
timestamp 1600868798
transform 1 0 19832 0 -1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _431_
timestamp 1600868798
transform 1 0 21028 0 -1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1600868798
transform 1 0 20660 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp 1600868798
transform 1 0 21856 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _381_
timestamp 1600868798
transform 1 0 22868 0 -1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _393_
timestamp 1600868798
transform 1 0 24064 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_32_126
timestamp 1600868798
transform 1 0 22592 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_138
timestamp 1600868798
transform 1 0 23696 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _382_
timestamp 1600868798
transform 1 0 25168 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1600868798
transform 1 0 25076 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1600868798
transform 1 0 24708 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_161
timestamp 1600868798
transform 1 0 25812 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _463_
timestamp 1600868798
transform 1 0 26916 0 -1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1600868798
transform 1 0 28112 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1600868798
transform 1 0 29124 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1600868798
transform 1 0 30688 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_194
timestamp 1600868798
transform 1 0 28848 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1600868798
transform 1 0 29400 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1600868798
transform 1 0 30504 0 -1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1600868798
transform 1 0 31424 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1600868798
transform 1 0 30780 0 -1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1600868798
transform 1 0 31332 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_226
timestamp 1600868798
transform 1 0 31792 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_238
timestamp 1600868798
transform 1 0 32896 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1600868798
transform -1 0 34368 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_250
timestamp 1600868798
transform 1 0 34000 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1600868798
transform 1 0 11000 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1600868798
transform 1 0 11000 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1600868798
transform 1 0 11276 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1600868798
transform 1 0 12380 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1600868798
transform 1 0 11276 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1600868798
transform 1 0 12380 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1600868798
transform 1 0 13852 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1600868798
transform 1 0 13484 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1600868798
transform 1 0 14588 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1600868798
transform 1 0 13484 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1600868798
transform 1 0 13944 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1600868798
transform 1 0 15048 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _342_
timestamp 1600868798
transform 1 0 16704 0 1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _498_
timestamp 1600868798
transform 1 0 16152 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _526_
timestamp 1600868798
transform 1 0 16796 0 -1 30040
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1600868798
transform 1 0 16612 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1600868798
transform 1 0 15692 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1600868798
transform 1 0 16428 0 1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_71
timestamp 1600868798
transform 1 0 17532 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1600868798
transform 1 0 16428 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _254_
timestamp 1600868798
transform 1 0 18452 0 1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1600868798
transform 1 0 19464 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1600868798
transform 1 0 18268 0 1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_90
timestamp 1600868798
transform 1 0 19280 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1600868798
transform 1 0 18912 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_93
timestamp 1600868798
transform 1 0 19556 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _379_
timestamp 1600868798
transform 1 0 20568 0 1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _397_
timestamp 1600868798
transform 1 0 21396 0 -1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _403_
timestamp 1600868798
transform 1 0 20200 0 -1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_102
timestamp 1600868798
transform 1 0 20384 0 1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1600868798
transform 1 0 21396 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_99
timestamp 1600868798
transform 1 0 20108 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1600868798
transform 1 0 21028 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_120
timestamp 1600868798
transform 1 0 22040 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1600868798
transform 1 0 22868 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1600868798
transform 1 0 22316 0 1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1600868798
transform 1 0 22132 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1600868798
transform 1 0 22224 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _395_
timestamp 1600868798
transform 1 0 22408 0 -1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1600868798
transform 1 0 23236 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _380_
timestamp 1600868798
transform 1 0 22960 0 1 28952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1600868798
transform 1 0 23788 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1600868798
transform 1 0 24156 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1600868798
transform 1 0 23788 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _479_
timestamp 1600868798
transform 1 0 23880 0 -1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1600868798
transform 1 0 24708 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _411_
timestamp 1600868798
transform 1 0 24248 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1600868798
transform 1 0 24892 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1600868798
transform 1 0 25076 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _389_
timestamp 1600868798
transform 1 0 25260 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _387_
timestamp 1600868798
transform 1 0 25168 0 -1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1600868798
transform 1 0 25812 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_162
timestamp 1600868798
transform 1 0 25904 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _450_
timestamp 1600868798
transform 1 0 26272 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _390_
timestamp 1600868798
transform 1 0 26180 0 -1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _407_
timestamp 1600868798
transform 1 0 27192 0 -1 30040
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _466_
timestamp 1600868798
transform 1 0 27928 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1600868798
transform 1 0 27836 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_173
timestamp 1600868798
transform 1 0 26916 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1600868798
transform 1 0 27652 0 1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1600868798
transform 1 0 26824 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1600868798
transform 1 0 28664 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_202
timestamp 1600868798
transform 1 0 29584 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1600868798
transform 1 0 28572 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1600868798
transform 1 0 29032 0 -1 30040
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1600868798
transform 1 0 28940 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1600868798
transform 1 0 30596 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_207
timestamp 1600868798
transform 1 0 30044 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_210
timestamp 1600868798
transform 1 0 30320 0 1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1600868798
transform 1 0 30688 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1600868798
transform 1 0 30504 0 1 28952
box -38 -48 1050 592
use sky130_fd_sc_hd__a21bo_4  _455_
timestamp 1600868798
transform 1 0 30780 0 -1 30040
box -38 -48 1234 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1600868798
transform 1 0 32344 0 -1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_33_223
timestamp 1600868798
transform 1 0 31516 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_235
timestamp 1600868798
transform 1 0 32620 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1600868798
transform 1 0 31976 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1600868798
transform -1 0 34368 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1600868798
transform -1 0 34368 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1600868798
transform 1 0 33448 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1600868798
transform 1 0 33356 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_245
timestamp 1600868798
transform 1 0 33540 0 1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1600868798
transform 1 0 32988 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1600868798
transform 1 0 11000 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1600868798
transform 1 0 11276 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1600868798
transform 1 0 12380 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1600868798
transform 1 0 13484 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1600868798
transform 1 0 14588 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1600868798
transform 1 0 16612 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1600868798
transform 1 0 15692 0 1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1600868798
transform 1 0 16428 0 1 30040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_62
timestamp 1600868798
transform 1 0 16704 0 1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_70
timestamp 1600868798
transform 1 0 17440 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _255_
timestamp 1600868798
transform 1 0 18452 0 1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _499_
timestamp 1600868798
transform 1 0 17716 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1600868798
transform 1 0 17992 0 1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_80
timestamp 1600868798
transform 1 0 18360 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_90
timestamp 1600868798
transform 1 0 19280 0 1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _415_
timestamp 1600868798
transform 1 0 20108 0 1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_98
timestamp 1600868798
transform 1 0 20016 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_108
timestamp 1600868798
transform 1 0 20936 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _396_
timestamp 1600868798
transform 1 0 22316 0 1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1600868798
transform 1 0 22224 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1600868798
transform 1 0 22040 0 1 30040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_132
timestamp 1600868798
transform 1 0 23144 0 1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _388_
timestamp 1600868798
transform 1 0 24432 0 1 30040
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_4  _408_
timestamp 1600868798
transform 1 0 25812 0 1 30040
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_35_144
timestamp 1600868798
transform 1 0 24248 0 1 30040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_155
timestamp 1600868798
transform 1 0 25260 0 1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1600868798
transform 1 0 28480 0 1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1600868798
transform 1 0 27836 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1600868798
transform 1 0 27008 0 1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1600868798
transform 1 0 27744 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_184
timestamp 1600868798
transform 1 0 27928 0 1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1600868798
transform 1 0 29860 0 1 30040
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_35_197
timestamp 1600868798
transform 1 0 29124 0 1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1600868798
transform 1 0 31884 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1600868798
transform 1 0 32528 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_223
timestamp 1600868798
transform 1 0 31516 0 1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1600868798
transform 1 0 32160 0 1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_237
timestamp 1600868798
transform 1 0 32804 0 1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1600868798
transform -1 0 34368 0 1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1600868798
transform 1 0 33448 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1600868798
transform 1 0 33356 0 1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_245
timestamp 1600868798
transform 1 0 33540 0 1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1600868798
transform 1 0 11000 0 -1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1600868798
transform 1 0 11276 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1600868798
transform 1 0 12380 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1600868798
transform 1 0 13852 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1600868798
transform 1 0 13484 0 -1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1600868798
transform 1 0 13944 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1600868798
transform 1 0 15048 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1600868798
transform 1 0 16152 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1600868798
transform 1 0 17256 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1600868798
transform 1 0 19464 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1600868798
transform 1 0 18360 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1600868798
transform 1 0 19556 0 -1 31128
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_4  _405_
timestamp 1600868798
transform 1 0 21120 0 -1 31128
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _416_
timestamp 1600868798
transform 1 0 20108 0 -1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_36_106
timestamp 1600868798
transform 1 0 20752 0 -1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _398_
timestamp 1600868798
transform 1 0 23880 0 -1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _417_
timestamp 1600868798
transform 1 0 22684 0 -1 31128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1600868798
transform 1 0 22316 0 -1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1600868798
transform 1 0 23512 0 -1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _422_
timestamp 1600868798
transform 1 0 25996 0 -1 31128
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1600868798
transform 1 0 25076 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_147
timestamp 1600868798
transform 1 0 24524 0 -1 31128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_154
timestamp 1600868798
transform 1 0 25168 0 -1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1600868798
transform 1 0 25904 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1600868798
transform 1 0 28204 0 -1 31128
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_36_176
timestamp 1600868798
transform 1 0 27192 0 -1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_184
timestamp 1600868798
transform 1 0 27928 0 -1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1600868798
transform 1 0 30688 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1600868798
transform 1 0 29860 0 -1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1600868798
transform 1 0 30596 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1600868798
transform 1 0 30780 0 -1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_36_222
timestamp 1600868798
transform 1 0 31424 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_234
timestamp 1600868798
transform 1 0 32528 0 -1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1600868798
transform -1 0 34368 0 -1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_246
timestamp 1600868798
transform 1 0 33632 0 -1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_250
timestamp 1600868798
transform 1 0 34000 0 -1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1600868798
transform 1 0 11000 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1600868798
transform 1 0 11276 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1600868798
transform 1 0 12380 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1600868798
transform 1 0 13484 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1600868798
transform 1 0 14588 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1600868798
transform 1 0 16612 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1600868798
transform 1 0 15692 0 1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1600868798
transform 1 0 16428 0 1 31128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1600868798
transform 1 0 16704 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1600868798
transform 1 0 17808 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1600868798
transform 1 0 18912 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _404_
timestamp 1600868798
transform 1 0 21028 0 1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1600868798
transform 1 0 20016 0 1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_37_105
timestamp 1600868798
transform 1 0 20660 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_116
timestamp 1600868798
transform 1 0 21672 0 1 31128
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _478_
timestamp 1600868798
transform 1 0 23972 0 1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1600868798
transform 1 0 22960 0 1 31128
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1600868798
transform 1 0 22316 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1600868798
transform 1 0 22224 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp 1600868798
transform 1 0 22592 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1600868798
transform 1 0 23604 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_148
timestamp 1600868798
transform 1 0 24616 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_160
timestamp 1600868798
transform 1 0 25720 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1600868798
transform 1 0 28204 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1600868798
transform 1 0 27836 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_172
timestamp 1600868798
transform 1 0 26824 0 1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_180
timestamp 1600868798
transform 1 0 27560 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_184
timestamp 1600868798
transform 1 0 27928 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1600868798
transform 1 0 30044 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1600868798
transform 1 0 28940 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1600868798
transform 1 0 28572 0 1 31128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_198
timestamp 1600868798
transform 1 0 29216 0 1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_206
timestamp 1600868798
transform 1 0 29952 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_211
timestamp 1600868798
transform 1 0 30412 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_223
timestamp 1600868798
transform 1 0 31516 0 1 31128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_235
timestamp 1600868798
transform 1 0 32620 0 1 31128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1600868798
transform -1 0 34368 0 1 31128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1600868798
transform 1 0 33448 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1600868798
transform 1 0 33356 0 1 31128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_245
timestamp 1600868798
transform 1 0 33540 0 1 31128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1600868798
transform 1 0 11000 0 -1 32216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1600868798
transform 1 0 11276 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1600868798
transform 1 0 12380 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1600868798
transform 1 0 13852 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1600868798
transform 1 0 13484 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1600868798
transform 1 0 13944 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1600868798
transform 1 0 15048 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1600868798
transform 1 0 16152 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1600868798
transform 1 0 17256 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _419_
timestamp 1600868798
transform 1 0 19740 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1600868798
transform 1 0 19464 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1600868798
transform 1 0 18360 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1600868798
transform 1 0 19556 0 -1 32216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1600868798
transform 1 0 21764 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_107
timestamp 1600868798
transform 1 0 20844 0 -1 32216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_115
timestamp 1600868798
transform 1 0 21580 0 -1 32216
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1600868798
transform 1 0 22776 0 -1 32216
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_38_121
timestamp 1600868798
transform 1 0 22132 0 -1 32216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_127
timestamp 1600868798
transform 1 0 22684 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_139
timestamp 1600868798
transform 1 0 23788 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_143
timestamp 1600868798
transform 1 0 24156 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1600868798
transform 1 0 26180 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1600868798
transform 1 0 25168 0 -1 32216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1600868798
transform 1 0 24248 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1600868798
transform 1 0 25076 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1600868798
transform 1 0 24616 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1600868798
transform 1 0 24984 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1600868798
transform 1 0 25812 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1600868798
transform 1 0 28480 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1600868798
transform 1 0 27376 0 -1 32216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_38_169
timestamp 1600868798
transform 1 0 26548 0 -1 32216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_177
timestamp 1600868798
transform 1 0 27284 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_185
timestamp 1600868798
transform 1 0 28020 0 -1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1600868798
transform 1 0 28388 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1600868798
transform 1 0 30688 0 -1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_194
timestamp 1600868798
transform 1 0 28848 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1600868798
transform 1 0 29952 0 -1 32216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1600868798
transform 1 0 30780 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1600868798
transform 1 0 31884 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1600868798
transform -1 0 34368 0 -1 32216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1600868798
transform 1 0 32988 0 -1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1600868798
transform 1 0 11000 0 1 32216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1600868798
transform 1 0 11000 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1600868798
transform 1 0 11276 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1600868798
transform 1 0 12380 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1600868798
transform 1 0 11276 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1600868798
transform 1 0 12380 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1600868798
transform 1 0 13852 0 -1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1600868798
transform 1 0 13484 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1600868798
transform 1 0 14588 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1600868798
transform 1 0 13484 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1600868798
transform 1 0 13944 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1600868798
transform 1 0 15048 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1600868798
transform 1 0 16612 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1600868798
transform 1 0 15692 0 1 32216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1600868798
transform 1 0 16428 0 1 32216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1600868798
transform 1 0 16704 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1600868798
transform 1 0 16152 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1600868798
transform 1 0 17256 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _480_
timestamp 1600868798
transform 1 0 19556 0 -1 33304
box -38 -48 1234 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1600868798
transform 1 0 19004 0 1 32216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1600868798
transform 1 0 19464 0 -1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1600868798
transform 1 0 17808 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_86
timestamp 1600868798
transform 1 0 18912 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_94
timestamp 1600868798
transform 1 0 19648 0 1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1600868798
transform 1 0 18360 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1600868798
transform 1 0 21764 0 -1 33304
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1600868798
transform 1 0 21120 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1600868798
transform 1 0 20016 0 1 32216
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_39_116
timestamp 1600868798
transform 1 0 21672 0 1 32216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1600868798
transform 1 0 20752 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_113
timestamp 1600868798
transform 1 0 21396 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _409_
timestamp 1600868798
transform 1 0 22776 0 1 32216
box -38 -48 1234 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1600868798
transform 1 0 23788 0 -1 33304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1600868798
transform 1 0 22224 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1600868798
transform 1 0 22316 0 1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1600868798
transform 1 0 22684 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1600868798
transform 1 0 23972 0 1 32216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1600868798
transform 1 0 23420 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1600868798
transform 1 0 25168 0 -1 33304
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1600868798
transform 1 0 24340 0 1 32216
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1600868798
transform 1 0 25076 0 -1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_163
timestamp 1600868798
transform 1 0 25996 0 1 32216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_146
timestamp 1600868798
transform 1 0 24432 0 -1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1600868798
transform 1 0 24984 0 -1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_161
timestamp 1600868798
transform 1 0 25812 0 -1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1600868798
transform 1 0 28388 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1600868798
transform 1 0 26640 0 1 32216
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1600868798
transform 1 0 26364 0 -1 33304
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1600868798
transform 1 0 27928 0 1 32216
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1600868798
transform 1 0 27836 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1600868798
transform 1 0 26548 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_177
timestamp 1600868798
transform 1 0 27284 0 1 32216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1600868798
transform 1 0 28020 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1600868798
transform 1 0 29032 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1600868798
transform 1 0 30688 0 -1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_195
timestamp 1600868798
transform 1 0 28940 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_207
timestamp 1600868798
transform 1 0 30044 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1600868798
transform 1 0 28664 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_199
timestamp 1600868798
transform 1 0 29308 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1600868798
transform 1 0 30412 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _513_ /home/ag/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1600868798
transform 1 0 30780 0 -1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_219
timestamp 1600868798
transform 1 0 31148 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_231
timestamp 1600868798
transform 1 0 32252 0 1 32216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1600868798
transform 1 0 31148 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1600868798
transform 1 0 32252 0 -1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1600868798
transform -1 0 34368 0 1 32216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1600868798
transform -1 0 34368 0 -1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1600868798
transform 1 0 33448 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1600868798
transform 1 0 33356 0 1 32216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_245
timestamp 1600868798
transform 1 0 33540 0 1 32216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1600868798
transform 1 0 33356 0 -1 33304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1600868798
transform 1 0 11000 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1600868798
transform 1 0 11276 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1600868798
transform 1 0 12380 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1600868798
transform 1 0 13484 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1600868798
transform 1 0 14588 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1600868798
transform 1 0 16612 0 1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1600868798
transform 1 0 15692 0 1 33304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1600868798
transform 1 0 16428 0 1 33304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1600868798
transform 1 0 16704 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1600868798
transform 1 0 17808 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_86
timestamp 1600868798
transform 1 0 18912 0 1 33304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_94
timestamp 1600868798
transform 1 0 19648 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1600868798
transform 1 0 19924 0 1 33304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1600868798
transform 1 0 21304 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1600868798
transform 1 0 20936 0 1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_115
timestamp 1600868798
transform 1 0 21580 0 1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_4  _418_
timestamp 1600868798
transform 1 0 22316 0 1 33304
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_4  _470_
timestamp 1600868798
transform 1 0 24064 0 1 33304
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1600868798
transform 1 0 22224 0 1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1600868798
transform 1 0 22132 0 1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_136
timestamp 1600868798
transform 1 0 23512 0 1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1600868798
transform 1 0 25628 0 1 33304
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1600868798
transform 1 0 25260 0 1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _467_
timestamp 1600868798
transform 1 0 27928 0 1 33304
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1600868798
transform 1 0 27008 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1600868798
transform 1 0 27836 0 1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_170
timestamp 1600868798
transform 1 0 26640 0 1 33304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_177
timestamp 1600868798
transform 1 0 27284 0 1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_197
timestamp 1600868798
transform 1 0 29124 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_209
timestamp 1600868798
transform 1 0 30228 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_221
timestamp 1600868798
transform 1 0 31332 0 1 33304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_233
timestamp 1600868798
transform 1 0 32436 0 1 33304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1600868798
transform -1 0 34368 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1600868798
transform 1 0 33448 0 1 33304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_241
timestamp 1600868798
transform 1 0 33172 0 1 33304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_245
timestamp 1600868798
transform 1 0 33540 0 1 33304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1600868798
transform 1 0 11000 0 -1 34392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1600868798
transform 1 0 11276 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1600868798
transform 1 0 12380 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1600868798
transform 1 0 13852 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1600868798
transform 1 0 13484 0 -1 34392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1600868798
transform 1 0 13944 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1600868798
transform 1 0 15048 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1600868798
transform 1 0 16704 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1600868798
transform 1 0 16152 0 -1 34392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1600868798
transform 1 0 16796 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1600868798
transform 1 0 19556 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1600868798
transform 1 0 17900 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1600868798
transform 1 0 19004 0 -1 34392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1600868798
transform 1 0 19648 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1600868798
transform 1 0 20752 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1600868798
transform 1 0 21856 0 -1 34392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1600868798
transform 1 0 23420 0 -1 34392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1600868798
transform 1 0 22408 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_125
timestamp 1600868798
transform 1 0 22500 0 -1 34392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_133
timestamp 1600868798
transform 1 0 23236 0 -1 34392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_138
timestamp 1600868798
transform 1 0 23696 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1600868798
transform 1 0 25536 0 -1 34392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1600868798
transform 1 0 25260 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_150
timestamp 1600868798
transform 1 0 24800 0 -1 34392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_154
timestamp 1600868798
transform 1 0 25168 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_156
timestamp 1600868798
transform 1 0 25352 0 -1 34392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_161
timestamp 1600868798
transform 1 0 25812 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1600868798
transform 1 0 28112 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_173
timestamp 1600868798
transform 1 0 26916 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_185
timestamp 1600868798
transform 1 0 28020 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1600868798
transform 1 0 28204 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1600868798
transform 1 0 29308 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1600868798
transform 1 0 30412 0 -1 34392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1600868798
transform 1 0 30964 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1600868798
transform 1 0 31056 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1600868798
transform 1 0 32160 0 -1 34392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1600868798
transform -1 0 34368 0 -1 34392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1600868798
transform 1 0 33816 0 -1 34392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1600868798
transform 1 0 33264 0 -1 34392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_249
timestamp 1600868798
transform 1 0 33908 0 -1 34392
box -38 -48 222 592
<< labels >>
rlabel metal2 s 31442 35809 31498 36609 6 clockp[0]
port 0 nsew default tristate
rlabel metal2 s 24082 8824 24138 9624 6 clockp[1]
port 1 nsew default tristate
rlabel metal2 s 12674 8824 12730 9624 6 dco
port 2 nsew default input
rlabel metal2 s 10466 8824 10522 9624 6 div[0]
port 3 nsew default input
rlabel metal3 s 9896 19712 10696 19832 6 div[1]
port 4 nsew default input
rlabel metal2 s 30890 8824 30946 9624 6 div[2]
port 5 nsew default input
rlabel metal3 s 34737 10464 35537 10584 6 div[3]
port 6 nsew default input
rlabel metal3 s 9896 12912 10696 13032 6 div[4]
port 7 nsew default input
rlabel metal2 s 22242 35809 22298 36609 6 enable
port 8 nsew default input
rlabel metal2 s 15434 35809 15490 36609 6 ext_trim[0]
port 9 nsew default input
rlabel metal2 s 26842 35809 26898 36609 6 ext_trim[10]
port 10 nsew default input
rlabel metal3 s 9896 26240 10696 26360 6 ext_trim[11]
port 11 nsew default input
rlabel metal3 s 34737 13728 35537 13848 6 ext_trim[12]
port 12 nsew default input
rlabel metal2 s 33098 8824 33154 9624 6 ext_trim[13]
port 13 nsew default input
rlabel metal3 s 9896 22976 10696 23096 6 ext_trim[14]
port 14 nsew default input
rlabel metal2 s 14882 8824 14938 9624 6 ext_trim[15]
port 15 nsew default input
rlabel metal3 s 34737 30592 35537 30712 6 ext_trim[16]
port 16 nsew default input
rlabel metal3 s 9896 29776 10696 29896 6 ext_trim[17]
port 17 nsew default input
rlabel metal2 s 33650 35809 33706 36609 6 ext_trim[18]
port 18 nsew default input
rlabel metal2 s 20034 35809 20090 36609 6 ext_trim[19]
port 19 nsew default input
rlabel metal3 s 34737 27328 35537 27448 6 ext_trim[1]
port 20 nsew default input
rlabel metal2 s 28682 8824 28738 9624 6 ext_trim[20]
port 21 nsew default input
rlabel metal3 s 9896 33040 10696 33160 6 ext_trim[21]
port 22 nsew default input
rlabel metal3 s 34737 23792 35537 23912 6 ext_trim[22]
port 23 nsew default input
rlabel metal3 s 9896 16176 10696 16296 6 ext_trim[23]
port 24 nsew default input
rlabel metal2 s 21690 8824 21746 9624 6 ext_trim[24]
port 25 nsew default input
rlabel metal3 s 34737 16992 35537 17112 6 ext_trim[25]
port 26 nsew default input
rlabel metal3 s 34737 20528 35537 20648 6 ext_trim[2]
port 27 nsew default input
rlabel metal2 s 13226 35809 13282 36609 6 ext_trim[3]
port 28 nsew default input
rlabel metal2 s 29234 35809 29290 36609 6 ext_trim[4]
port 29 nsew default input
rlabel metal2 s 26290 8824 26346 9624 6 ext_trim[5]
port 30 nsew default input
rlabel metal2 s 24634 35809 24690 36609 6 ext_trim[6]
port 31 nsew default input
rlabel metal2 s 11018 35809 11074 36609 6 ext_trim[7]
port 32 nsew default input
rlabel metal2 s 17826 35809 17882 36609 6 ext_trim[8]
port 33 nsew default input
rlabel metal3 s 34737 33856 35537 33976 6 ext_trim[9]
port 34 nsew default input
rlabel metal2 s 19482 8824 19538 9624 6 osc
port 35 nsew default input
rlabel metal2 s 17274 8824 17330 9624 6 resetb
port 36 nsew default input
rlabel metal4 s 5000 5000 9000 40392 4 VPWR
port 37 nsew default input
rlabel metal4 s 0 0 4000 45392 4 VGND
port 38 nsew default input
<< properties >>
string FIXED_BBOX 0 0 45368 45392
<< end >>
