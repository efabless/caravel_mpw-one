VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.190 BY 50.240 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 3.000 2000.190 3.600 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 9.120 2000.190 9.720 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 15.240 2000.190 15.840 ;
    END
  END caravel_rstn
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.080 47.840 313.360 50.240 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.920 47.840 752.200 50.240 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 756.520 47.840 756.800 50.240 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.660 47.840 760.940 50.240 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.260 47.840 765.540 50.240 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.400 47.840 769.680 50.240 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 774.000 47.840 774.280 50.240 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.140 47.840 778.420 50.240 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 782.740 47.840 783.020 50.240 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.880 47.840 787.160 50.240 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 791.480 47.840 791.760 50.240 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.240 47.840 357.520 50.240 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.620 47.840 795.900 50.240 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.220 47.840 800.500 50.240 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.360 47.840 804.640 50.240 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.960 47.840 809.240 50.240 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.100 47.840 813.380 50.240 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.700 47.840 817.980 50.240 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 822.300 47.840 822.580 50.240 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 826.440 47.840 826.720 50.240 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 831.040 47.840 831.320 50.240 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.180 47.840 835.460 50.240 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.380 47.840 361.660 50.240 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.780 47.840 840.060 50.240 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 843.920 47.840 844.200 50.240 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 848.520 47.840 848.800 50.240 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.660 47.840 852.940 50.240 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 857.260 47.840 857.540 50.240 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 861.400 47.840 861.680 50.240 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.000 47.840 866.280 50.240 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.140 47.840 870.420 50.240 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.980 47.840 366.260 50.240 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.120 47.840 370.400 50.240 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.720 47.840 375.000 50.240 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.320 47.840 379.600 50.240 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.460 47.840 383.740 50.240 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.060 47.840 388.340 50.240 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.200 47.840 392.480 50.240 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.800 47.840 397.080 50.240 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.680 47.840 317.960 50.240 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 400.940 47.840 401.220 50.240 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 405.540 47.840 405.820 50.240 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.680 47.840 409.960 50.240 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.280 47.840 414.560 50.240 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 418.420 47.840 418.700 50.240 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.020 47.840 423.300 50.240 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.160 47.840 427.440 50.240 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.760 47.840 432.040 50.240 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.900 47.840 436.180 50.240 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 440.500 47.840 440.780 50.240 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.280 47.840 322.560 50.240 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.100 47.840 445.380 50.240 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.240 47.840 449.520 50.240 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.840 47.840 454.120 50.240 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.980 47.840 458.260 50.240 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.580 47.840 462.860 50.240 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.720 47.840 467.000 50.240 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.320 47.840 471.600 50.240 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.460 47.840 475.740 50.240 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 480.060 47.840 480.340 50.240 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.200 47.840 484.480 50.240 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.420 47.840 326.700 50.240 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.800 47.840 489.080 50.240 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.940 47.840 493.220 50.240 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 497.540 47.840 497.820 50.240 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.140 47.840 502.420 50.240 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.280 47.840 506.560 50.240 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 510.880 47.840 511.160 50.240 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 515.020 47.840 515.300 50.240 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.620 47.840 519.900 50.240 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.760 47.840 524.040 50.240 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 528.360 47.840 528.640 50.240 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.020 47.840 331.300 50.240 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 532.500 47.840 532.780 50.240 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.100 47.840 537.380 50.240 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 541.240 47.840 541.520 50.240 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.840 47.840 546.120 50.240 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.980 47.840 550.260 50.240 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 554.580 47.840 554.860 50.240 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.720 47.840 559.000 50.240 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.320 47.840 563.600 50.240 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.920 47.840 568.200 50.240 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 572.060 47.840 572.340 50.240 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.160 47.840 335.440 50.240 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.660 47.840 576.940 50.240 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.800 47.840 581.080 50.240 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.400 47.840 585.680 50.240 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.540 47.840 589.820 50.240 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 594.140 47.840 594.420 50.240 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.280 47.840 598.560 50.240 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 602.880 47.840 603.160 50.240 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.020 47.840 607.300 50.240 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 611.620 47.840 611.900 50.240 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 615.760 47.840 616.040 50.240 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.760 47.840 340.040 50.240 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.360 47.840 620.640 50.240 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 624.500 47.840 624.780 50.240 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 629.100 47.840 629.380 50.240 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 633.700 47.840 633.980 50.240 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.840 47.840 638.120 50.240 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 642.440 47.840 642.720 50.240 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.580 47.840 646.860 50.240 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.180 47.840 651.460 50.240 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.320 47.840 655.600 50.240 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.920 47.840 660.200 50.240 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.900 47.840 344.180 50.240 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.060 47.840 664.340 50.240 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.660 47.840 668.940 50.240 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 672.800 47.840 673.080 50.240 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.400 47.840 677.680 50.240 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.540 47.840 681.820 50.240 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.140 47.840 686.420 50.240 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.740 47.840 691.020 50.240 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.880 47.840 695.160 50.240 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.480 47.840 699.760 50.240 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 703.620 47.840 703.900 50.240 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.500 47.840 348.780 50.240 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 708.220 47.840 708.500 50.240 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.360 47.840 712.640 50.240 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.960 47.840 717.240 50.240 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 721.100 47.840 721.380 50.240 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.700 47.840 725.980 50.240 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.840 47.840 730.120 50.240 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 734.440 47.840 734.720 50.240 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 738.580 47.840 738.860 50.240 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 743.180 47.840 743.460 50.240 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 747.320 47.840 747.600 50.240 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 352.640 47.840 352.920 50.240 ;
    END
  END la_data_in_mprj[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.740 47.840 875.020 50.240 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1313.120 47.840 1313.400 50.240 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.720 47.840 1318.000 50.240 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.320 47.840 1322.600 50.240 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1326.460 47.840 1326.740 50.240 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.060 47.840 1331.340 50.240 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.200 47.840 1335.480 50.240 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1339.800 47.840 1340.080 50.240 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1343.940 47.840 1344.220 50.240 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.540 47.840 1348.820 50.240 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1352.680 47.840 1352.960 50.240 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.440 47.840 918.720 50.240 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1357.280 47.840 1357.560 50.240 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1361.420 47.840 1361.700 50.240 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1366.020 47.840 1366.300 50.240 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1370.160 47.840 1370.440 50.240 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1374.760 47.840 1375.040 50.240 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1379.360 47.840 1379.640 50.240 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1383.500 47.840 1383.780 50.240 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1388.100 47.840 1388.380 50.240 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1392.240 47.840 1392.520 50.240 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1396.840 47.840 1397.120 50.240 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 923.040 47.840 923.320 50.240 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.980 47.840 1401.260 50.240 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1405.580 47.840 1405.860 50.240 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.720 47.840 1410.000 50.240 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.320 47.840 1414.600 50.240 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.460 47.840 1418.740 50.240 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1423.060 47.840 1423.340 50.240 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1427.200 47.840 1427.480 50.240 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1431.800 47.840 1432.080 50.240 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.180 47.840 927.460 50.240 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.780 47.840 932.060 50.240 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.920 47.840 936.200 50.240 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.520 47.840 940.800 50.240 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.120 47.840 945.400 50.240 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.260 47.840 949.540 50.240 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.860 47.840 954.140 50.240 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.000 47.840 958.280 50.240 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 879.340 47.840 879.620 50.240 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.600 47.840 962.880 50.240 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 966.740 47.840 967.020 50.240 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.340 47.840 971.620 50.240 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 975.480 47.840 975.760 50.240 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 980.080 47.840 980.360 50.240 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.220 47.840 984.500 50.240 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 988.820 47.840 989.100 50.240 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 992.960 47.840 993.240 50.240 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.560 47.840 997.840 50.240 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1002.160 47.840 1002.440 50.240 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 883.480 47.840 883.760 50.240 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.300 47.840 1006.580 50.240 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.900 47.840 1011.180 50.240 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.040 47.840 1015.320 50.240 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.640 47.840 1019.920 50.240 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.780 47.840 1024.060 50.240 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.380 47.840 1028.660 50.240 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.520 47.840 1032.800 50.240 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.120 47.840 1037.400 50.240 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.260 47.840 1041.540 50.240 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.860 47.840 1046.140 50.240 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.080 47.840 888.360 50.240 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.000 47.840 1050.280 50.240 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.600 47.840 1054.880 50.240 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.740 47.840 1059.020 50.240 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.340 47.840 1063.620 50.240 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.940 47.840 1068.220 50.240 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.080 47.840 1072.360 50.240 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.680 47.840 1076.960 50.240 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.820 47.840 1081.100 50.240 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1085.420 47.840 1085.700 50.240 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1089.560 47.840 1089.840 50.240 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.220 47.840 892.500 50.240 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.160 47.840 1094.440 50.240 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.300 47.840 1098.580 50.240 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1102.900 47.840 1103.180 50.240 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1107.040 47.840 1107.320 50.240 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1111.640 47.840 1111.920 50.240 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.780 47.840 1116.060 50.240 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1120.380 47.840 1120.660 50.240 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1124.520 47.840 1124.800 50.240 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1129.120 47.840 1129.400 50.240 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.720 47.840 1134.000 50.240 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.820 47.840 897.100 50.240 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.860 47.840 1138.140 50.240 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1142.460 47.840 1142.740 50.240 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1146.600 47.840 1146.880 50.240 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.200 47.840 1151.480 50.240 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1155.340 47.840 1155.620 50.240 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1159.940 47.840 1160.220 50.240 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1164.080 47.840 1164.360 50.240 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.680 47.840 1168.960 50.240 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.820 47.840 1173.100 50.240 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1177.420 47.840 1177.700 50.240 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.960 47.840 901.240 50.240 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1181.560 47.840 1181.840 50.240 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1186.160 47.840 1186.440 50.240 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.760 47.840 1191.040 50.240 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.900 47.840 1195.180 50.240 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.500 47.840 1199.780 50.240 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.640 47.840 1203.920 50.240 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.240 47.840 1208.520 50.240 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1212.380 47.840 1212.660 50.240 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1216.980 47.840 1217.260 50.240 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.120 47.840 1221.400 50.240 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 905.560 47.840 905.840 50.240 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.720 47.840 1226.000 50.240 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.860 47.840 1230.140 50.240 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.460 47.840 1234.740 50.240 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.600 47.840 1238.880 50.240 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.200 47.840 1243.480 50.240 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.340 47.840 1247.620 50.240 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.940 47.840 1252.220 50.240 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1256.540 47.840 1256.820 50.240 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.680 47.840 1260.960 50.240 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1265.280 47.840 1265.560 50.240 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.700 47.840 909.980 50.240 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.420 47.840 1269.700 50.240 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1274.020 47.840 1274.300 50.240 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1278.160 47.840 1278.440 50.240 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1282.760 47.840 1283.040 50.240 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1286.900 47.840 1287.180 50.240 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1291.500 47.840 1291.780 50.240 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1295.640 47.840 1295.920 50.240 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.240 47.840 1300.520 50.240 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.380 47.840 1304.660 50.240 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.980 47.840 1309.260 50.240 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 914.300 47.840 914.580 50.240 ;
    END
  END la_oen[9]
  PIN la_output_core[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.940 47.840 1436.220 50.240 ;
    END
  END la_output_core[0]
  PIN la_output_core[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1874.780 47.840 1875.060 50.240 ;
    END
  END la_output_core[100]
  PIN la_output_core[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1879.380 47.840 1879.660 50.240 ;
    END
  END la_output_core[101]
  PIN la_output_core[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1883.520 47.840 1883.800 50.240 ;
    END
  END la_output_core[102]
  PIN la_output_core[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1888.120 47.840 1888.400 50.240 ;
    END
  END la_output_core[103]
  PIN la_output_core[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1892.260 47.840 1892.540 50.240 ;
    END
  END la_output_core[104]
  PIN la_output_core[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1896.860 47.840 1897.140 50.240 ;
    END
  END la_output_core[105]
  PIN la_output_core[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1901.000 47.840 1901.280 50.240 ;
    END
  END la_output_core[106]
  PIN la_output_core[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1905.600 47.840 1905.880 50.240 ;
    END
  END la_output_core[107]
  PIN la_output_core[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1909.740 47.840 1910.020 50.240 ;
    END
  END la_output_core[108]
  PIN la_output_core[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1914.340 47.840 1914.620 50.240 ;
    END
  END la_output_core[109]
  PIN la_output_core[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1480.100 47.840 1480.380 50.240 ;
    END
  END la_output_core[10]
  PIN la_output_core[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.480 47.840 1918.760 50.240 ;
    END
  END la_output_core[110]
  PIN la_output_core[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1923.080 47.840 1923.360 50.240 ;
    END
  END la_output_core[111]
  PIN la_output_core[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1927.220 47.840 1927.500 50.240 ;
    END
  END la_output_core[112]
  PIN la_output_core[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1931.820 47.840 1932.100 50.240 ;
    END
  END la_output_core[113]
  PIN la_output_core[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.960 47.840 1936.240 50.240 ;
    END
  END la_output_core[114]
  PIN la_output_core[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1940.560 47.840 1940.840 50.240 ;
    END
  END la_output_core[115]
  PIN la_output_core[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1945.160 47.840 1945.440 50.240 ;
    END
  END la_output_core[116]
  PIN la_output_core[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1949.300 47.840 1949.580 50.240 ;
    END
  END la_output_core[117]
  PIN la_output_core[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.900 47.840 1954.180 50.240 ;
    END
  END la_output_core[118]
  PIN la_output_core[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1958.040 47.840 1958.320 50.240 ;
    END
  END la_output_core[119]
  PIN la_output_core[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1484.240 47.840 1484.520 50.240 ;
    END
  END la_output_core[11]
  PIN la_output_core[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1962.640 47.840 1962.920 50.240 ;
    END
  END la_output_core[120]
  PIN la_output_core[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1966.780 47.840 1967.060 50.240 ;
    END
  END la_output_core[121]
  PIN la_output_core[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.380 47.840 1971.660 50.240 ;
    END
  END la_output_core[122]
  PIN la_output_core[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1975.520 47.840 1975.800 50.240 ;
    END
  END la_output_core[123]
  PIN la_output_core[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1980.120 47.840 1980.400 50.240 ;
    END
  END la_output_core[124]
  PIN la_output_core[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1984.260 47.840 1984.540 50.240 ;
    END
  END la_output_core[125]
  PIN la_output_core[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.860 47.840 1989.140 50.240 ;
    END
  END la_output_core[126]
  PIN la_output_core[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1993.000 47.840 1993.280 50.240 ;
    END
  END la_output_core[127]
  PIN la_output_core[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1488.840 47.840 1489.120 50.240 ;
    END
  END la_output_core[12]
  PIN la_output_core[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.980 47.840 1493.260 50.240 ;
    END
  END la_output_core[13]
  PIN la_output_core[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1497.580 47.840 1497.860 50.240 ;
    END
  END la_output_core[14]
  PIN la_output_core[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1502.180 47.840 1502.460 50.240 ;
    END
  END la_output_core[15]
  PIN la_output_core[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.320 47.840 1506.600 50.240 ;
    END
  END la_output_core[16]
  PIN la_output_core[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.920 47.840 1511.200 50.240 ;
    END
  END la_output_core[17]
  PIN la_output_core[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1515.060 47.840 1515.340 50.240 ;
    END
  END la_output_core[18]
  PIN la_output_core[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1519.660 47.840 1519.940 50.240 ;
    END
  END la_output_core[19]
  PIN la_output_core[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1440.540 47.840 1440.820 50.240 ;
    END
  END la_output_core[1]
  PIN la_output_core[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1523.800 47.840 1524.080 50.240 ;
    END
  END la_output_core[20]
  PIN la_output_core[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1528.400 47.840 1528.680 50.240 ;
    END
  END la_output_core[21]
  PIN la_output_core[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1532.540 47.840 1532.820 50.240 ;
    END
  END la_output_core[22]
  PIN la_output_core[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1537.140 47.840 1537.420 50.240 ;
    END
  END la_output_core[23]
  PIN la_output_core[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1541.280 47.840 1541.560 50.240 ;
    END
  END la_output_core[24]
  PIN la_output_core[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.880 47.840 1546.160 50.240 ;
    END
  END la_output_core[25]
  PIN la_output_core[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1550.020 47.840 1550.300 50.240 ;
    END
  END la_output_core[26]
  PIN la_output_core[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.620 47.840 1554.900 50.240 ;
    END
  END la_output_core[27]
  PIN la_output_core[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1558.760 47.840 1559.040 50.240 ;
    END
  END la_output_core[28]
  PIN la_output_core[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1563.360 47.840 1563.640 50.240 ;
    END
  END la_output_core[29]
  PIN la_output_core[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1445.140 47.840 1445.420 50.240 ;
    END
  END la_output_core[2]
  PIN la_output_core[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1567.960 47.840 1568.240 50.240 ;
    END
  END la_output_core[30]
  PIN la_output_core[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.100 47.840 1572.380 50.240 ;
    END
  END la_output_core[31]
  PIN la_output_core[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.700 47.840 1576.980 50.240 ;
    END
  END la_output_core[32]
  PIN la_output_core[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1580.840 47.840 1581.120 50.240 ;
    END
  END la_output_core[33]
  PIN la_output_core[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1585.440 47.840 1585.720 50.240 ;
    END
  END la_output_core[34]
  PIN la_output_core[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.580 47.840 1589.860 50.240 ;
    END
  END la_output_core[35]
  PIN la_output_core[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1594.180 47.840 1594.460 50.240 ;
    END
  END la_output_core[36]
  PIN la_output_core[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1598.320 47.840 1598.600 50.240 ;
    END
  END la_output_core[37]
  PIN la_output_core[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1602.920 47.840 1603.200 50.240 ;
    END
  END la_output_core[38]
  PIN la_output_core[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1607.060 47.840 1607.340 50.240 ;
    END
  END la_output_core[39]
  PIN la_output_core[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1449.280 47.840 1449.560 50.240 ;
    END
  END la_output_core[3]
  PIN la_output_core[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1611.660 47.840 1611.940 50.240 ;
    END
  END la_output_core[40]
  PIN la_output_core[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1615.800 47.840 1616.080 50.240 ;
    END
  END la_output_core[41]
  PIN la_output_core[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1620.400 47.840 1620.680 50.240 ;
    END
  END la_output_core[42]
  PIN la_output_core[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1624.540 47.840 1624.820 50.240 ;
    END
  END la_output_core[43]
  PIN la_output_core[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1629.140 47.840 1629.420 50.240 ;
    END
  END la_output_core[44]
  PIN la_output_core[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.740 47.840 1634.020 50.240 ;
    END
  END la_output_core[45]
  PIN la_output_core[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.880 47.840 1638.160 50.240 ;
    END
  END la_output_core[46]
  PIN la_output_core[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1642.480 47.840 1642.760 50.240 ;
    END
  END la_output_core[47]
  PIN la_output_core[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1646.620 47.840 1646.900 50.240 ;
    END
  END la_output_core[48]
  PIN la_output_core[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1651.220 47.840 1651.500 50.240 ;
    END
  END la_output_core[49]
  PIN la_output_core[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.880 47.840 1454.160 50.240 ;
    END
  END la_output_core[4]
  PIN la_output_core[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1655.360 47.840 1655.640 50.240 ;
    END
  END la_output_core[50]
  PIN la_output_core[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1659.960 47.840 1660.240 50.240 ;
    END
  END la_output_core[51]
  PIN la_output_core[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1664.100 47.840 1664.380 50.240 ;
    END
  END la_output_core[52]
  PIN la_output_core[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1668.700 47.840 1668.980 50.240 ;
    END
  END la_output_core[53]
  PIN la_output_core[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1672.840 47.840 1673.120 50.240 ;
    END
  END la_output_core[54]
  PIN la_output_core[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1677.440 47.840 1677.720 50.240 ;
    END
  END la_output_core[55]
  PIN la_output_core[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1681.580 47.840 1681.860 50.240 ;
    END
  END la_output_core[56]
  PIN la_output_core[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1686.180 47.840 1686.460 50.240 ;
    END
  END la_output_core[57]
  PIN la_output_core[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1690.780 47.840 1691.060 50.240 ;
    END
  END la_output_core[58]
  PIN la_output_core[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1694.920 47.840 1695.200 50.240 ;
    END
  END la_output_core[59]
  PIN la_output_core[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1458.020 47.840 1458.300 50.240 ;
    END
  END la_output_core[5]
  PIN la_output_core[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1699.520 47.840 1699.800 50.240 ;
    END
  END la_output_core[60]
  PIN la_output_core[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.660 47.840 1703.940 50.240 ;
    END
  END la_output_core[61]
  PIN la_output_core[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1708.260 47.840 1708.540 50.240 ;
    END
  END la_output_core[62]
  PIN la_output_core[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1712.400 47.840 1712.680 50.240 ;
    END
  END la_output_core[63]
  PIN la_output_core[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1717.000 47.840 1717.280 50.240 ;
    END
  END la_output_core[64]
  PIN la_output_core[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.140 47.840 1721.420 50.240 ;
    END
  END la_output_core[65]
  PIN la_output_core[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1725.740 47.840 1726.020 50.240 ;
    END
  END la_output_core[66]
  PIN la_output_core[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1729.880 47.840 1730.160 50.240 ;
    END
  END la_output_core[67]
  PIN la_output_core[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1734.480 47.840 1734.760 50.240 ;
    END
  END la_output_core[68]
  PIN la_output_core[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.620 47.840 1738.900 50.240 ;
    END
  END la_output_core[69]
  PIN la_output_core[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1462.620 47.840 1462.900 50.240 ;
    END
  END la_output_core[6]
  PIN la_output_core[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1743.220 47.840 1743.500 50.240 ;
    END
  END la_output_core[70]
  PIN la_output_core[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.360 47.840 1747.640 50.240 ;
    END
  END la_output_core[71]
  PIN la_output_core[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.960 47.840 1752.240 50.240 ;
    END
  END la_output_core[72]
  PIN la_output_core[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.560 47.840 1756.840 50.240 ;
    END
  END la_output_core[73]
  PIN la_output_core[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1760.700 47.840 1760.980 50.240 ;
    END
  END la_output_core[74]
  PIN la_output_core[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1765.300 47.840 1765.580 50.240 ;
    END
  END la_output_core[75]
  PIN la_output_core[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1769.440 47.840 1769.720 50.240 ;
    END
  END la_output_core[76]
  PIN la_output_core[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.040 47.840 1774.320 50.240 ;
    END
  END la_output_core[77]
  PIN la_output_core[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1778.180 47.840 1778.460 50.240 ;
    END
  END la_output_core[78]
  PIN la_output_core[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1782.780 47.840 1783.060 50.240 ;
    END
  END la_output_core[79]
  PIN la_output_core[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1466.760 47.840 1467.040 50.240 ;
    END
  END la_output_core[7]
  PIN la_output_core[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.920 47.840 1787.200 50.240 ;
    END
  END la_output_core[80]
  PIN la_output_core[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1791.520 47.840 1791.800 50.240 ;
    END
  END la_output_core[81]
  PIN la_output_core[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1795.660 47.840 1795.940 50.240 ;
    END
  END la_output_core[82]
  PIN la_output_core[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1800.260 47.840 1800.540 50.240 ;
    END
  END la_output_core[83]
  PIN la_output_core[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.400 47.840 1804.680 50.240 ;
    END
  END la_output_core[84]
  PIN la_output_core[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1809.000 47.840 1809.280 50.240 ;
    END
  END la_output_core[85]
  PIN la_output_core[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1813.140 47.840 1813.420 50.240 ;
    END
  END la_output_core[86]
  PIN la_output_core[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1817.740 47.840 1818.020 50.240 ;
    END
  END la_output_core[87]
  PIN la_output_core[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.340 47.840 1822.620 50.240 ;
    END
  END la_output_core[88]
  PIN la_output_core[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1826.480 47.840 1826.760 50.240 ;
    END
  END la_output_core[89]
  PIN la_output_core[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.360 47.840 1471.640 50.240 ;
    END
  END la_output_core[8]
  PIN la_output_core[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1831.080 47.840 1831.360 50.240 ;
    END
  END la_output_core[90]
  PIN la_output_core[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1835.220 47.840 1835.500 50.240 ;
    END
  END la_output_core[91]
  PIN la_output_core[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.820 47.840 1840.100 50.240 ;
    END
  END la_output_core[92]
  PIN la_output_core[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1843.960 47.840 1844.240 50.240 ;
    END
  END la_output_core[93]
  PIN la_output_core[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1848.560 47.840 1848.840 50.240 ;
    END
  END la_output_core[94]
  PIN la_output_core[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1852.700 47.840 1852.980 50.240 ;
    END
  END la_output_core[95]
  PIN la_output_core[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.300 47.840 1857.580 50.240 ;
    END
  END la_output_core[96]
  PIN la_output_core[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1861.440 47.840 1861.720 50.240 ;
    END
  END la_output_core[97]
  PIN la_output_core[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1866.040 47.840 1866.320 50.240 ;
    END
  END la_output_core[98]
  PIN la_output_core[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1870.180 47.840 1870.460 50.240 ;
    END
  END la_output_core[99]
  PIN la_output_core[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1475.500 47.840 1475.780 50.240 ;
    END
  END la_output_core[9]
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.700 0.240 12.980 2.640 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.920 0.240 269.200 2.640 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.680 0.240 294.960 2.640 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.980 0.240 320.260 2.640 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.740 0.240 346.020 2.640 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.500 0.240 371.780 2.640 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.260 0.240 397.540 2.640 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.560 0.240 422.840 2.640 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.320 0.240 448.600 2.640 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.080 0.240 474.360 2.640 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.840 0.240 500.120 2.640 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.000 0.240 38.280 2.640 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.140 0.240 525.420 2.640 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.900 0.240 551.180 2.640 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.660 0.240 576.940 2.640 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.420 0.240 602.700 2.640 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.720 0.240 628.000 2.640 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.480 0.240 653.760 2.640 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.240 0.240 679.520 2.640 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.000 0.240 705.280 2.640 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.300 0.240 730.580 2.640 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.060 0.240 756.340 2.640 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.760 0.240 64.040 2.640 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.820 0.240 782.100 2.640 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.580 0.240 807.860 2.640 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.520 0.240 89.800 2.640 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.820 0.240 115.100 2.640 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.580 0.240 140.860 2.640 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.340 0.240 166.620 2.640 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.100 0.240 192.380 2.640 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.400 0.240 217.680 2.640 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.160 0.240 243.440 2.640 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.120 47.840 2.400 50.240 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.820 47.840 46.100 50.240 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.960 47.840 50.240 50.240 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.560 47.840 54.840 50.240 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.700 47.840 58.980 50.240 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.300 47.840 63.580 50.240 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.900 47.840 68.180 50.240 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.040 47.840 72.320 50.240 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.640 47.840 76.920 50.240 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.780 47.840 81.060 50.240 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.380 47.840 85.660 50.240 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.260 47.840 6.540 50.240 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.520 47.840 89.800 50.240 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.120 47.840 94.400 50.240 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.260 47.840 98.540 50.240 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.860 47.840 103.140 50.240 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.000 47.840 107.280 50.240 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.600 47.840 111.880 50.240 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.740 47.840 116.020 50.240 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.340 47.840 120.620 50.240 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.480 47.840 124.760 50.240 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.080 47.840 129.360 50.240 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.860 47.840 11.140 50.240 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.680 47.840 133.960 50.240 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.820 47.840 138.100 50.240 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.000 47.840 15.280 50.240 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.600 47.840 19.880 50.240 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.740 47.840 24.020 50.240 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.340 47.840 28.620 50.240 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.480 47.840 32.760 50.240 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.080 47.840 37.360 50.240 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.220 47.840 41.500 50.240 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 832.880 0.240 833.160 2.640 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.420 47.840 142.700 50.240 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.640 0.240 858.920 2.640 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.860 0.240 1115.140 2.640 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.620 0.240 1140.900 2.640 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1166.380 0.240 1166.660 2.640 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1192.140 0.240 1192.420 2.640 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1217.440 0.240 1217.720 2.640 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.200 0.240 1243.480 2.640 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.960 0.240 1269.240 2.640 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.720 0.240 1295.000 2.640 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.020 0.240 1320.300 2.640 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1345.780 0.240 1346.060 2.640 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.400 0.240 884.680 2.640 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1371.540 0.240 1371.820 2.640 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.300 0.240 1397.580 2.640 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1422.600 0.240 1422.880 2.640 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1448.360 0.240 1448.640 2.640 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1474.120 0.240 1474.400 2.640 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1499.880 0.240 1500.160 2.640 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1525.180 0.240 1525.460 2.640 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1550.940 0.240 1551.220 2.640 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.700 0.240 1576.980 2.640 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1602.460 0.240 1602.740 2.640 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.160 0.240 910.440 2.640 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.760 0.240 1628.040 2.640 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1653.520 0.240 1653.800 2.640 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.460 0.240 935.740 2.640 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.220 0.240 961.500 2.640 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.980 0.240 987.260 2.640 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.740 0.240 1013.020 2.640 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1038.040 0.240 1038.320 2.640 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.800 0.240 1064.080 2.640 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1089.560 0.240 1089.840 2.640 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.560 47.840 146.840 50.240 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.720 47.840 191.000 50.240 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.860 47.840 195.140 50.240 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.460 47.840 199.740 50.240 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.600 47.840 203.880 50.240 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.200 47.840 208.480 50.240 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.340 47.840 212.620 50.240 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.940 47.840 217.220 50.240 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.080 47.840 221.360 50.240 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.680 47.840 225.960 50.240 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.820 47.840 230.100 50.240 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.160 47.840 151.440 50.240 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.420 47.840 234.700 50.240 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 238.560 47.840 238.840 50.240 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.160 47.840 243.440 50.240 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.300 47.840 247.580 50.240 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 251.900 47.840 252.180 50.240 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.500 47.840 256.780 50.240 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.640 47.840 260.920 50.240 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.240 47.840 265.520 50.240 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.380 47.840 269.660 50.240 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.980 47.840 274.260 50.240 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.300 47.840 155.580 50.240 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.120 47.840 278.400 50.240 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 282.720 47.840 283.000 50.240 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.900 47.840 160.180 50.240 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.040 47.840 164.320 50.240 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.640 47.840 168.920 50.240 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.780 47.840 173.060 50.240 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.380 47.840 177.660 50.240 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.520 47.840 181.800 50.240 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.120 47.840 186.400 50.240 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.280 0.240 1679.560 2.640 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1705.040 0.240 1705.320 2.640 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1730.340 0.240 1730.620 2.640 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.100 0.240 1756.380 2.640 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.860 47.840 287.140 50.240 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.460 47.840 291.740 50.240 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.600 47.840 295.880 50.240 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.200 47.840 300.480 50.240 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1781.860 0.240 1782.140 2.640 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.340 47.840 304.620 50.240 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1807.620 0.240 1807.900 2.640 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.940 47.840 309.220 50.240 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1832.920 0.240 1833.200 2.640 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1858.680 0.240 1858.960 2.640 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1884.440 0.240 1884.720 2.640 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1910.200 0.240 1910.480 2.640 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.190 6.400 2.590 7.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1997.790 21.360 2000.190 21.960 ;
    END
  END user_clock2
  PIN user_resetn
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1997.790 28.160 2000.190 28.760 ;
    END
  END user_resetn
  PIN vccd
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1997.600 47.840 1997.880 50.240 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.190 18.640 2.590 19.240 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1935.500 0.240 1935.780 2.640 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1961.260 0.240 1961.540 2.640 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1987.020 0.240 1987.300 2.640 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 34.280 2000.190 34.880 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 40.400 2000.190 41.000 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.190 31.560 2.590 32.160 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1997.790 46.520 2000.190 47.120 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.190 43.800 2.590 44.400 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 0.190 0.155 8.470 3.045 ;
      LAYER met1 ;
        RECT 0.190 0.000 8.470 3.200 ;
  END
END mgmt_protect
END LIBRARY

