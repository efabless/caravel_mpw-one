magic
tech sky130A
magscale 1 2
timestamp 1624566096
<< obsli1 >>
rect 1104 2159 448868 167399
<< obsm1 >>
rect 78766 168008 78830 168020
rect 176102 168008 176166 168020
rect 78766 168000 176166 168008
rect 199838 168008 199902 168020
rect 276842 168008 276906 168020
rect 199838 168000 276906 168008
rect 14 1028 449498 168000
<< metal2 >>
rect 386 167200 442 168000
rect 1122 167200 1178 168000
rect 1858 167200 1914 168000
rect 2594 167200 2650 168000
rect 3330 167200 3386 168000
rect 4158 167200 4214 168000
rect 4894 167200 4950 168000
rect 5630 167200 5686 168000
rect 6366 167200 6422 168000
rect 7102 167200 7158 168000
rect 7930 167200 7986 168000
rect 8666 167200 8722 168000
rect 9402 167200 9458 168000
rect 10138 167200 10194 168000
rect 10874 167200 10930 168000
rect 11702 167200 11758 168000
rect 12438 167200 12494 168000
rect 13174 167200 13230 168000
rect 13910 167200 13966 168000
rect 14646 167200 14702 168000
rect 15474 167200 15530 168000
rect 16210 167200 16266 168000
rect 16946 167200 17002 168000
rect 17682 167200 17738 168000
rect 18418 167200 18474 168000
rect 19246 167200 19302 168000
rect 19982 167200 20038 168000
rect 20718 167200 20774 168000
rect 21454 167200 21510 168000
rect 22190 167200 22246 168000
rect 23018 167200 23074 168000
rect 23754 167200 23810 168000
rect 24490 167200 24546 168000
rect 25226 167200 25282 168000
rect 26054 167200 26110 168000
rect 26790 167200 26846 168000
rect 27526 167200 27582 168000
rect 28262 167200 28318 168000
rect 28998 167200 29054 168000
rect 29826 167200 29882 168000
rect 30562 167200 30618 168000
rect 31298 167200 31354 168000
rect 32034 167200 32090 168000
rect 32770 167200 32826 168000
rect 33598 167200 33654 168000
rect 34334 167200 34390 168000
rect 35070 167200 35126 168000
rect 35806 167200 35862 168000
rect 36542 167200 36598 168000
rect 37370 167200 37426 168000
rect 38106 167200 38162 168000
rect 38842 167200 38898 168000
rect 39578 167200 39634 168000
rect 40314 167200 40370 168000
rect 41142 167200 41198 168000
rect 41878 167200 41934 168000
rect 42614 167200 42670 168000
rect 43350 167200 43406 168000
rect 44086 167200 44142 168000
rect 44914 167200 44970 168000
rect 45650 167200 45706 168000
rect 46386 167200 46442 168000
rect 47122 167200 47178 168000
rect 47950 167200 48006 168000
rect 48686 167200 48742 168000
rect 49422 167200 49478 168000
rect 50158 167200 50214 168000
rect 50894 167200 50950 168000
rect 51722 167200 51778 168000
rect 52458 167200 52514 168000
rect 53194 167200 53250 168000
rect 53930 167200 53986 168000
rect 54666 167200 54722 168000
rect 55494 167200 55550 168000
rect 56230 167200 56286 168000
rect 56966 167200 57022 168000
rect 57702 167200 57758 168000
rect 58438 167200 58494 168000
rect 59266 167200 59322 168000
rect 60002 167200 60058 168000
rect 60738 167200 60794 168000
rect 61474 167200 61530 168000
rect 62210 167200 62266 168000
rect 63038 167200 63094 168000
rect 63774 167200 63830 168000
rect 64510 167200 64566 168000
rect 65246 167200 65302 168000
rect 65982 167200 66038 168000
rect 66810 167200 66866 168000
rect 67546 167200 67602 168000
rect 68282 167200 68338 168000
rect 69018 167200 69074 168000
rect 69754 167200 69810 168000
rect 70582 167200 70638 168000
rect 71318 167200 71374 168000
rect 72054 167200 72110 168000
rect 72790 167200 72846 168000
rect 73618 167200 73674 168000
rect 74354 167200 74410 168000
rect 75090 167200 75146 168000
rect 75826 167200 75882 168000
rect 76562 167200 76618 168000
rect 77390 167200 77446 168000
rect 78126 167200 78182 168000
rect 78862 167200 78918 168000
rect 79598 167200 79654 168000
rect 80334 167200 80390 168000
rect 81162 167200 81218 168000
rect 81898 167200 81954 168000
rect 82634 167200 82690 168000
rect 83370 167200 83426 168000
rect 84106 167200 84162 168000
rect 84934 167200 84990 168000
rect 85670 167200 85726 168000
rect 86406 167200 86462 168000
rect 87142 167200 87198 168000
rect 87878 167200 87934 168000
rect 88706 167200 88762 168000
rect 89442 167200 89498 168000
rect 90178 167200 90234 168000
rect 90914 167200 90970 168000
rect 91650 167200 91706 168000
rect 92478 167200 92534 168000
rect 93214 167200 93270 168000
rect 93950 167200 94006 168000
rect 94686 167200 94742 168000
rect 95514 167200 95570 168000
rect 96250 167200 96306 168000
rect 96986 167200 97042 168000
rect 97722 167200 97778 168000
rect 98458 167200 98514 168000
rect 99286 167200 99342 168000
rect 100022 167200 100078 168000
rect 100758 167200 100814 168000
rect 101494 167200 101550 168000
rect 102230 167200 102286 168000
rect 103058 167200 103114 168000
rect 103794 167200 103850 168000
rect 104530 167200 104586 168000
rect 105266 167200 105322 168000
rect 106002 167200 106058 168000
rect 106830 167200 106886 168000
rect 107566 167200 107622 168000
rect 108302 167200 108358 168000
rect 109038 167200 109094 168000
rect 109774 167200 109830 168000
rect 110602 167200 110658 168000
rect 111338 167200 111394 168000
rect 112074 167200 112130 168000
rect 112810 167200 112866 168000
rect 113546 167200 113602 168000
rect 114374 167200 114430 168000
rect 115110 167200 115166 168000
rect 115846 167200 115902 168000
rect 116582 167200 116638 168000
rect 117318 167200 117374 168000
rect 118146 167200 118202 168000
rect 118882 167200 118938 168000
rect 119618 167200 119674 168000
rect 120354 167200 120410 168000
rect 121182 167200 121238 168000
rect 121918 167200 121974 168000
rect 122654 167200 122710 168000
rect 123390 167200 123446 168000
rect 124126 167200 124182 168000
rect 124954 167200 125010 168000
rect 125690 167200 125746 168000
rect 126426 167200 126482 168000
rect 127162 167200 127218 168000
rect 127898 167200 127954 168000
rect 128726 167200 128782 168000
rect 129462 167200 129518 168000
rect 130198 167200 130254 168000
rect 130934 167200 130990 168000
rect 131670 167200 131726 168000
rect 132498 167200 132554 168000
rect 133234 167200 133290 168000
rect 133970 167200 134026 168000
rect 134706 167200 134762 168000
rect 135442 167200 135498 168000
rect 136270 167200 136326 168000
rect 137006 167200 137062 168000
rect 137742 167200 137798 168000
rect 138478 167200 138534 168000
rect 139214 167200 139270 168000
rect 140042 167200 140098 168000
rect 140778 167200 140834 168000
rect 141514 167200 141570 168000
rect 142250 167200 142306 168000
rect 143078 167200 143134 168000
rect 143814 167200 143870 168000
rect 144550 167200 144606 168000
rect 145286 167200 145342 168000
rect 146022 167200 146078 168000
rect 146850 167200 146906 168000
rect 147586 167200 147642 168000
rect 148322 167200 148378 168000
rect 149058 167200 149114 168000
rect 149794 167200 149850 168000
rect 150622 167200 150678 168000
rect 151358 167200 151414 168000
rect 152094 167200 152150 168000
rect 152830 167200 152886 168000
rect 153566 167200 153622 168000
rect 154394 167200 154450 168000
rect 155130 167200 155186 168000
rect 155866 167200 155922 168000
rect 156602 167200 156658 168000
rect 157338 167200 157394 168000
rect 158166 167200 158222 168000
rect 158902 167200 158958 168000
rect 159638 167200 159694 168000
rect 160374 167200 160430 168000
rect 161110 167200 161166 168000
rect 161938 167200 161994 168000
rect 162674 167200 162730 168000
rect 163410 167200 163466 168000
rect 164146 167200 164202 168000
rect 164882 167200 164938 168000
rect 165710 167200 165766 168000
rect 166446 167200 166502 168000
rect 167182 167200 167238 168000
rect 167918 167200 167974 168000
rect 168746 167200 168802 168000
rect 169482 167200 169538 168000
rect 170218 167200 170274 168000
rect 170954 167200 171010 168000
rect 171690 167200 171746 168000
rect 172518 167200 172574 168000
rect 173254 167200 173310 168000
rect 173990 167200 174046 168000
rect 174726 167200 174782 168000
rect 175462 167200 175518 168000
rect 176290 167200 176346 168000
rect 177026 167200 177082 168000
rect 177762 167200 177818 168000
rect 178498 167200 178554 168000
rect 179234 167200 179290 168000
rect 180062 167200 180118 168000
rect 180798 167200 180854 168000
rect 181534 167200 181590 168000
rect 182270 167200 182326 168000
rect 183006 167200 183062 168000
rect 183834 167200 183890 168000
rect 184570 167200 184626 168000
rect 185306 167200 185362 168000
rect 186042 167200 186098 168000
rect 186778 167200 186834 168000
rect 187606 167200 187662 168000
rect 188342 167200 188398 168000
rect 189078 167200 189134 168000
rect 189814 167200 189870 168000
rect 190642 167200 190698 168000
rect 191378 167200 191434 168000
rect 192114 167200 192170 168000
rect 192850 167200 192906 168000
rect 193586 167200 193642 168000
rect 194414 167200 194470 168000
rect 195150 167200 195206 168000
rect 195886 167200 195942 168000
rect 196622 167200 196678 168000
rect 197358 167200 197414 168000
rect 198186 167200 198242 168000
rect 198922 167200 198978 168000
rect 199658 167200 199714 168000
rect 200394 167200 200450 168000
rect 201130 167200 201186 168000
rect 201958 167200 202014 168000
rect 202694 167200 202750 168000
rect 203430 167200 203486 168000
rect 204166 167200 204222 168000
rect 204902 167200 204958 168000
rect 205730 167200 205786 168000
rect 206466 167200 206522 168000
rect 207202 167200 207258 168000
rect 207938 167200 207994 168000
rect 208674 167200 208730 168000
rect 209502 167200 209558 168000
rect 210238 167200 210294 168000
rect 210974 167200 211030 168000
rect 211710 167200 211766 168000
rect 212446 167200 212502 168000
rect 213274 167200 213330 168000
rect 214010 167200 214066 168000
rect 214746 167200 214802 168000
rect 215482 167200 215538 168000
rect 216310 167200 216366 168000
rect 217046 167200 217102 168000
rect 217782 167200 217838 168000
rect 218518 167200 218574 168000
rect 219254 167200 219310 168000
rect 220082 167200 220138 168000
rect 220818 167200 220874 168000
rect 221554 167200 221610 168000
rect 222290 167200 222346 168000
rect 223026 167200 223082 168000
rect 223854 167200 223910 168000
rect 224590 167200 224646 168000
rect 225326 167200 225382 168000
rect 226062 167200 226118 168000
rect 226798 167200 226854 168000
rect 227626 167200 227682 168000
rect 228362 167200 228418 168000
rect 229098 167200 229154 168000
rect 229834 167200 229890 168000
rect 230570 167200 230626 168000
rect 231398 167200 231454 168000
rect 232134 167200 232190 168000
rect 232870 167200 232926 168000
rect 233606 167200 233662 168000
rect 234342 167200 234398 168000
rect 235170 167200 235226 168000
rect 235906 167200 235962 168000
rect 236642 167200 236698 168000
rect 237378 167200 237434 168000
rect 238206 167200 238262 168000
rect 238942 167200 238998 168000
rect 239678 167200 239734 168000
rect 240414 167200 240470 168000
rect 241150 167200 241206 168000
rect 241978 167200 242034 168000
rect 242714 167200 242770 168000
rect 243450 167200 243506 168000
rect 244186 167200 244242 168000
rect 244922 167200 244978 168000
rect 245750 167200 245806 168000
rect 246486 167200 246542 168000
rect 247222 167200 247278 168000
rect 247958 167200 248014 168000
rect 248694 167200 248750 168000
rect 249522 167200 249578 168000
rect 250258 167200 250314 168000
rect 250994 167200 251050 168000
rect 251730 167200 251786 168000
rect 252466 167200 252522 168000
rect 253294 167200 253350 168000
rect 254030 167200 254086 168000
rect 254766 167200 254822 168000
rect 255502 167200 255558 168000
rect 256238 167200 256294 168000
rect 257066 167200 257122 168000
rect 257802 167200 257858 168000
rect 258538 167200 258594 168000
rect 259274 167200 259330 168000
rect 260010 167200 260066 168000
rect 260838 167200 260894 168000
rect 261574 167200 261630 168000
rect 262310 167200 262366 168000
rect 263046 167200 263102 168000
rect 263874 167200 263930 168000
rect 264610 167200 264666 168000
rect 265346 167200 265402 168000
rect 266082 167200 266138 168000
rect 266818 167200 266874 168000
rect 267646 167200 267702 168000
rect 268382 167200 268438 168000
rect 269118 167200 269174 168000
rect 269854 167200 269910 168000
rect 270590 167200 270646 168000
rect 271418 167200 271474 168000
rect 272154 167200 272210 168000
rect 272890 167200 272946 168000
rect 273626 167200 273682 168000
rect 274362 167200 274418 168000
rect 275190 167200 275246 168000
rect 275926 167200 275982 168000
rect 276662 167200 276718 168000
rect 277398 167200 277454 168000
rect 278134 167200 278190 168000
rect 278962 167200 279018 168000
rect 279698 167200 279754 168000
rect 280434 167200 280490 168000
rect 281170 167200 281226 168000
rect 281906 167200 281962 168000
rect 282734 167200 282790 168000
rect 283470 167200 283526 168000
rect 284206 167200 284262 168000
rect 284942 167200 284998 168000
rect 285770 167200 285826 168000
rect 286506 167200 286562 168000
rect 287242 167200 287298 168000
rect 287978 167200 288034 168000
rect 288714 167200 288770 168000
rect 289542 167200 289598 168000
rect 290278 167200 290334 168000
rect 291014 167200 291070 168000
rect 291750 167200 291806 168000
rect 292486 167200 292542 168000
rect 293314 167200 293370 168000
rect 294050 167200 294106 168000
rect 294786 167200 294842 168000
rect 295522 167200 295578 168000
rect 296258 167200 296314 168000
rect 297086 167200 297142 168000
rect 297822 167200 297878 168000
rect 298558 167200 298614 168000
rect 299294 167200 299350 168000
rect 300030 167200 300086 168000
rect 300858 167200 300914 168000
rect 301594 167200 301650 168000
rect 302330 167200 302386 168000
rect 303066 167200 303122 168000
rect 303802 167200 303858 168000
rect 304630 167200 304686 168000
rect 305366 167200 305422 168000
rect 306102 167200 306158 168000
rect 306838 167200 306894 168000
rect 307574 167200 307630 168000
rect 308402 167200 308458 168000
rect 309138 167200 309194 168000
rect 309874 167200 309930 168000
rect 310610 167200 310666 168000
rect 311438 167200 311494 168000
rect 312174 167200 312230 168000
rect 312910 167200 312966 168000
rect 313646 167200 313702 168000
rect 314382 167200 314438 168000
rect 315210 167200 315266 168000
rect 315946 167200 316002 168000
rect 316682 167200 316738 168000
rect 317418 167200 317474 168000
rect 318154 167200 318210 168000
rect 318982 167200 319038 168000
rect 319718 167200 319774 168000
rect 320454 167200 320510 168000
rect 321190 167200 321246 168000
rect 321926 167200 321982 168000
rect 322754 167200 322810 168000
rect 323490 167200 323546 168000
rect 324226 167200 324282 168000
rect 324962 167200 325018 168000
rect 325698 167200 325754 168000
rect 326526 167200 326582 168000
rect 327262 167200 327318 168000
rect 327998 167200 328054 168000
rect 328734 167200 328790 168000
rect 329470 167200 329526 168000
rect 330298 167200 330354 168000
rect 331034 167200 331090 168000
rect 331770 167200 331826 168000
rect 332506 167200 332562 168000
rect 333334 167200 333390 168000
rect 334070 167200 334126 168000
rect 334806 167200 334862 168000
rect 335542 167200 335598 168000
rect 336278 167200 336334 168000
rect 337106 167200 337162 168000
rect 337842 167200 337898 168000
rect 338578 167200 338634 168000
rect 339314 167200 339370 168000
rect 340050 167200 340106 168000
rect 340878 167200 340934 168000
rect 341614 167200 341670 168000
rect 342350 167200 342406 168000
rect 343086 167200 343142 168000
rect 343822 167200 343878 168000
rect 344650 167200 344706 168000
rect 345386 167200 345442 168000
rect 346122 167200 346178 168000
rect 346858 167200 346914 168000
rect 347594 167200 347650 168000
rect 348422 167200 348478 168000
rect 349158 167200 349214 168000
rect 349894 167200 349950 168000
rect 350630 167200 350686 168000
rect 351366 167200 351422 168000
rect 352194 167200 352250 168000
rect 352930 167200 352986 168000
rect 353666 167200 353722 168000
rect 354402 167200 354458 168000
rect 355138 167200 355194 168000
rect 355966 167200 356022 168000
rect 356702 167200 356758 168000
rect 357438 167200 357494 168000
rect 358174 167200 358230 168000
rect 359002 167200 359058 168000
rect 359738 167200 359794 168000
rect 360474 167200 360530 168000
rect 361210 167200 361266 168000
rect 361946 167200 362002 168000
rect 362774 167200 362830 168000
rect 363510 167200 363566 168000
rect 364246 167200 364302 168000
rect 364982 167200 365038 168000
rect 365718 167200 365774 168000
rect 366546 167200 366602 168000
rect 367282 167200 367338 168000
rect 368018 167200 368074 168000
rect 368754 167200 368810 168000
rect 369490 167200 369546 168000
rect 370318 167200 370374 168000
rect 371054 167200 371110 168000
rect 371790 167200 371846 168000
rect 372526 167200 372582 168000
rect 373262 167200 373318 168000
rect 374090 167200 374146 168000
rect 374826 167200 374882 168000
rect 375562 167200 375618 168000
rect 376298 167200 376354 168000
rect 377034 167200 377090 168000
rect 377862 167200 377918 168000
rect 378598 167200 378654 168000
rect 379334 167200 379390 168000
rect 380070 167200 380126 168000
rect 380898 167200 380954 168000
rect 381634 167200 381690 168000
rect 382370 167200 382426 168000
rect 383106 167200 383162 168000
rect 383842 167200 383898 168000
rect 384670 167200 384726 168000
rect 385406 167200 385462 168000
rect 386142 167200 386198 168000
rect 386878 167200 386934 168000
rect 387614 167200 387670 168000
rect 388442 167200 388498 168000
rect 389178 167200 389234 168000
rect 389914 167200 389970 168000
rect 390650 167200 390706 168000
rect 391386 167200 391442 168000
rect 392214 167200 392270 168000
rect 392950 167200 393006 168000
rect 393686 167200 393742 168000
rect 394422 167200 394478 168000
rect 395158 167200 395214 168000
rect 395986 167200 396042 168000
rect 396722 167200 396778 168000
rect 397458 167200 397514 168000
rect 398194 167200 398250 168000
rect 398930 167200 398986 168000
rect 399758 167200 399814 168000
rect 400494 167200 400550 168000
rect 401230 167200 401286 168000
rect 401966 167200 402022 168000
rect 402702 167200 402758 168000
rect 403530 167200 403586 168000
rect 404266 167200 404322 168000
rect 405002 167200 405058 168000
rect 405738 167200 405794 168000
rect 406566 167200 406622 168000
rect 407302 167200 407358 168000
rect 408038 167200 408094 168000
rect 408774 167200 408830 168000
rect 409510 167200 409566 168000
rect 410338 167200 410394 168000
rect 411074 167200 411130 168000
rect 411810 167200 411866 168000
rect 412546 167200 412602 168000
rect 413282 167200 413338 168000
rect 414110 167200 414166 168000
rect 414846 167200 414902 168000
rect 415582 167200 415638 168000
rect 416318 167200 416374 168000
rect 417054 167200 417110 168000
rect 417882 167200 417938 168000
rect 418618 167200 418674 168000
rect 419354 167200 419410 168000
rect 420090 167200 420146 168000
rect 420826 167200 420882 168000
rect 421654 167200 421710 168000
rect 422390 167200 422446 168000
rect 423126 167200 423182 168000
rect 423862 167200 423918 168000
rect 424598 167200 424654 168000
rect 425426 167200 425482 168000
rect 426162 167200 426218 168000
rect 426898 167200 426954 168000
rect 427634 167200 427690 168000
rect 428462 167200 428518 168000
rect 429198 167200 429254 168000
rect 429934 167200 429990 168000
rect 430670 167200 430726 168000
rect 431406 167200 431462 168000
rect 432234 167200 432290 168000
rect 432970 167200 433026 168000
rect 433706 167200 433762 168000
rect 434442 167200 434498 168000
rect 435178 167200 435234 168000
rect 436006 167200 436062 168000
rect 436742 167200 436798 168000
rect 437478 167200 437534 168000
rect 438214 167200 438270 168000
rect 438950 167200 439006 168000
rect 439778 167200 439834 168000
rect 440514 167200 440570 168000
rect 441250 167200 441306 168000
rect 441986 167200 442042 168000
rect 442722 167200 442778 168000
rect 443550 167200 443606 168000
rect 444286 167200 444342 168000
rect 445022 167200 445078 168000
rect 445758 167200 445814 168000
rect 446494 167200 446550 168000
rect 447322 167200 447378 168000
rect 448058 167200 448114 168000
rect 448794 167200 448850 168000
rect 449530 167200 449586 168000
rect 8666 0 8722 800
rect 25962 0 26018 800
rect 43258 0 43314 800
rect 60554 0 60610 800
rect 77850 0 77906 800
rect 95146 0 95202 800
rect 112442 0 112498 800
rect 129738 0 129794 800
rect 147034 0 147090 800
rect 164422 0 164478 800
rect 181718 0 181774 800
rect 199014 0 199070 800
rect 216310 0 216366 800
rect 233606 0 233662 800
rect 250902 0 250958 800
rect 268198 0 268254 800
rect 285494 0 285550 800
rect 302790 0 302846 800
rect 320178 0 320234 800
rect 337474 0 337530 800
rect 354770 0 354826 800
rect 372066 0 372122 800
rect 389362 0 389418 800
rect 406658 0 406714 800
rect 423954 0 424010 800
rect 441250 0 441306 800
<< obsm2 >>
rect 78772 168000 78824 168026
rect 176108 168000 176160 168026
rect 199844 168000 199896 168026
rect 276848 168000 276900 168026
rect 18 167144 330 168000
rect 498 167144 1066 168000
rect 1234 167144 1802 168000
rect 1970 167144 2538 168000
rect 2706 167144 3274 168000
rect 3442 167144 4102 168000
rect 4270 167144 4838 168000
rect 5006 167144 5574 168000
rect 5742 167144 6310 168000
rect 6478 167144 7046 168000
rect 7214 167144 7874 168000
rect 8042 167144 8610 168000
rect 8778 167144 9346 168000
rect 9514 167144 10082 168000
rect 10250 167144 10818 168000
rect 10986 167144 11646 168000
rect 11814 167144 12382 168000
rect 12550 167144 13118 168000
rect 13286 167144 13854 168000
rect 14022 167144 14590 168000
rect 14758 167144 15418 168000
rect 15586 167144 16154 168000
rect 16322 167144 16890 168000
rect 17058 167144 17626 168000
rect 17794 167144 18362 168000
rect 18530 167144 19190 168000
rect 19358 167144 19926 168000
rect 20094 167144 20662 168000
rect 20830 167144 21398 168000
rect 21566 167144 22134 168000
rect 22302 167144 22962 168000
rect 23130 167144 23698 168000
rect 23866 167144 24434 168000
rect 24602 167144 25170 168000
rect 25338 167144 25998 168000
rect 26166 167144 26734 168000
rect 26902 167144 27470 168000
rect 27638 167144 28206 168000
rect 28374 167144 28942 168000
rect 29110 167144 29770 168000
rect 29938 167144 30506 168000
rect 30674 167144 31242 168000
rect 31410 167144 31978 168000
rect 32146 167144 32714 168000
rect 32882 167144 33542 168000
rect 33710 167144 34278 168000
rect 34446 167144 35014 168000
rect 35182 167144 35750 168000
rect 35918 167144 36486 168000
rect 36654 167144 37314 168000
rect 37482 167144 38050 168000
rect 38218 167144 38786 168000
rect 38954 167144 39522 168000
rect 39690 167144 40258 168000
rect 40426 167144 41086 168000
rect 41254 167144 41822 168000
rect 41990 167144 42558 168000
rect 42726 167144 43294 168000
rect 43462 167144 44030 168000
rect 44198 167144 44858 168000
rect 45026 167144 45594 168000
rect 45762 167144 46330 168000
rect 46498 167144 47066 168000
rect 47234 167144 47894 168000
rect 48062 167144 48630 168000
rect 48798 167144 49366 168000
rect 49534 167144 50102 168000
rect 50270 167144 50838 168000
rect 51006 167144 51666 168000
rect 51834 167144 52402 168000
rect 52570 167144 53138 168000
rect 53306 167144 53874 168000
rect 54042 167144 54610 168000
rect 54778 167144 55438 168000
rect 55606 167144 56174 168000
rect 56342 167144 56910 168000
rect 57078 167144 57646 168000
rect 57814 167144 58382 168000
rect 58550 167144 59210 168000
rect 59378 167144 59946 168000
rect 60114 167144 60682 168000
rect 60850 167144 61418 168000
rect 61586 167144 62154 168000
rect 62322 167144 62982 168000
rect 63150 167144 63718 168000
rect 63886 167144 64454 168000
rect 64622 167144 65190 168000
rect 65358 167144 65926 168000
rect 66094 167144 66754 168000
rect 66922 167144 67490 168000
rect 67658 167144 68226 168000
rect 68394 167144 68962 168000
rect 69130 167144 69698 168000
rect 69866 167144 70526 168000
rect 70694 167144 71262 168000
rect 71430 167144 71998 168000
rect 72166 167144 72734 168000
rect 72902 167144 73562 168000
rect 73730 167144 74298 168000
rect 74466 167144 75034 168000
rect 75202 167144 75770 168000
rect 75938 167144 76506 168000
rect 76674 167144 77334 168000
rect 77502 167144 78070 168000
rect 78238 167968 78824 168000
rect 78238 167144 78806 167968
rect 78974 167144 79542 168000
rect 79710 167144 80278 168000
rect 80446 167144 81106 168000
rect 81274 167144 81842 168000
rect 82010 167144 82578 168000
rect 82746 167144 83314 168000
rect 83482 167144 84050 168000
rect 84218 167144 84878 168000
rect 85046 167144 85614 168000
rect 85782 167144 86350 168000
rect 86518 167144 87086 168000
rect 87254 167144 87822 168000
rect 87990 167144 88650 168000
rect 88818 167144 89386 168000
rect 89554 167144 90122 168000
rect 90290 167144 90858 168000
rect 91026 167144 91594 168000
rect 91762 167144 92422 168000
rect 92590 167144 93158 168000
rect 93326 167144 93894 168000
rect 94062 167144 94630 168000
rect 94798 167144 95458 168000
rect 95626 167144 96194 168000
rect 96362 167144 96930 168000
rect 97098 167144 97666 168000
rect 97834 167144 98402 168000
rect 98570 167144 99230 168000
rect 99398 167144 99966 168000
rect 100134 167144 100702 168000
rect 100870 167144 101438 168000
rect 101606 167144 102174 168000
rect 102342 167144 103002 168000
rect 103170 167144 103738 168000
rect 103906 167144 104474 168000
rect 104642 167144 105210 168000
rect 105378 167144 105946 168000
rect 106114 167144 106774 168000
rect 106942 167144 107510 168000
rect 107678 167144 108246 168000
rect 108414 167144 108982 168000
rect 109150 167144 109718 168000
rect 109886 167144 110546 168000
rect 110714 167144 111282 168000
rect 111450 167144 112018 168000
rect 112186 167144 112754 168000
rect 112922 167144 113490 168000
rect 113658 167144 114318 168000
rect 114486 167144 115054 168000
rect 115222 167144 115790 168000
rect 115958 167144 116526 168000
rect 116694 167144 117262 168000
rect 117430 167144 118090 168000
rect 118258 167144 118826 168000
rect 118994 167144 119562 168000
rect 119730 167144 120298 168000
rect 120466 167144 121126 168000
rect 121294 167144 121862 168000
rect 122030 167144 122598 168000
rect 122766 167144 123334 168000
rect 123502 167144 124070 168000
rect 124238 167144 124898 168000
rect 125066 167144 125634 168000
rect 125802 167144 126370 168000
rect 126538 167144 127106 168000
rect 127274 167144 127842 168000
rect 128010 167144 128670 168000
rect 128838 167144 129406 168000
rect 129574 167144 130142 168000
rect 130310 167144 130878 168000
rect 131046 167144 131614 168000
rect 131782 167144 132442 168000
rect 132610 167144 133178 168000
rect 133346 167144 133914 168000
rect 134082 167144 134650 168000
rect 134818 167144 135386 168000
rect 135554 167144 136214 168000
rect 136382 167144 136950 168000
rect 137118 167144 137686 168000
rect 137854 167144 138422 168000
rect 138590 167144 139158 168000
rect 139326 167144 139986 168000
rect 140154 167144 140722 168000
rect 140890 167144 141458 168000
rect 141626 167144 142194 168000
rect 142362 167144 143022 168000
rect 143190 167144 143758 168000
rect 143926 167144 144494 168000
rect 144662 167144 145230 168000
rect 145398 167144 145966 168000
rect 146134 167144 146794 168000
rect 146962 167144 147530 168000
rect 147698 167144 148266 168000
rect 148434 167144 149002 168000
rect 149170 167144 149738 168000
rect 149906 167144 150566 168000
rect 150734 167144 151302 168000
rect 151470 167144 152038 168000
rect 152206 167144 152774 168000
rect 152942 167144 153510 168000
rect 153678 167144 154338 168000
rect 154506 167144 155074 168000
rect 155242 167144 155810 168000
rect 155978 167144 156546 168000
rect 156714 167144 157282 168000
rect 157450 167144 158110 168000
rect 158278 167144 158846 168000
rect 159014 167144 159582 168000
rect 159750 167144 160318 168000
rect 160486 167144 161054 168000
rect 161222 167144 161882 168000
rect 162050 167144 162618 168000
rect 162786 167144 163354 168000
rect 163522 167144 164090 168000
rect 164258 167144 164826 168000
rect 164994 167144 165654 168000
rect 165822 167144 166390 168000
rect 166558 167144 167126 168000
rect 167294 167144 167862 168000
rect 168030 167144 168690 168000
rect 168858 167144 169426 168000
rect 169594 167144 170162 168000
rect 170330 167144 170898 168000
rect 171066 167144 171634 168000
rect 171802 167144 172462 168000
rect 172630 167144 173198 168000
rect 173366 167144 173934 168000
rect 174102 167144 174670 168000
rect 174838 167144 175406 168000
rect 175574 167144 176234 168000
rect 176402 167144 176970 168000
rect 177138 167144 177706 168000
rect 177874 167144 178442 168000
rect 178610 167144 179178 168000
rect 179346 167144 180006 168000
rect 180174 167144 180742 168000
rect 180910 167144 181478 168000
rect 181646 167144 182214 168000
rect 182382 167144 182950 168000
rect 183118 167144 183778 168000
rect 183946 167144 184514 168000
rect 184682 167144 185250 168000
rect 185418 167144 185986 168000
rect 186154 167144 186722 168000
rect 186890 167144 187550 168000
rect 187718 167144 188286 168000
rect 188454 167144 189022 168000
rect 189190 167144 189758 168000
rect 189926 167144 190586 168000
rect 190754 167144 191322 168000
rect 191490 167144 192058 168000
rect 192226 167144 192794 168000
rect 192962 167144 193530 168000
rect 193698 167144 194358 168000
rect 194526 167144 195094 168000
rect 195262 167144 195830 168000
rect 195998 167144 196566 168000
rect 196734 167144 197302 168000
rect 197470 167144 198130 168000
rect 198298 167144 198866 168000
rect 199034 167144 199602 168000
rect 199770 167144 200338 168000
rect 200506 167144 201074 168000
rect 201242 167144 201902 168000
rect 202070 167144 202638 168000
rect 202806 167144 203374 168000
rect 203542 167144 204110 168000
rect 204278 167144 204846 168000
rect 205014 167144 205674 168000
rect 205842 167144 206410 168000
rect 206578 167144 207146 168000
rect 207314 167144 207882 168000
rect 208050 167144 208618 168000
rect 208786 167144 209446 168000
rect 209614 167144 210182 168000
rect 210350 167144 210918 168000
rect 211086 167144 211654 168000
rect 211822 167144 212390 168000
rect 212558 167144 213218 168000
rect 213386 167144 213954 168000
rect 214122 167144 214690 168000
rect 214858 167144 215426 168000
rect 215594 167144 216254 168000
rect 216422 167144 216990 168000
rect 217158 167144 217726 168000
rect 217894 167144 218462 168000
rect 218630 167144 219198 168000
rect 219366 167144 220026 168000
rect 220194 167144 220762 168000
rect 220930 167144 221498 168000
rect 221666 167144 222234 168000
rect 222402 167144 222970 168000
rect 223138 167144 223798 168000
rect 223966 167144 224534 168000
rect 224702 167144 225270 168000
rect 225438 167144 226006 168000
rect 226174 167144 226742 168000
rect 226910 167144 227570 168000
rect 227738 167144 228306 168000
rect 228474 167144 229042 168000
rect 229210 167144 229778 168000
rect 229946 167144 230514 168000
rect 230682 167144 231342 168000
rect 231510 167144 232078 168000
rect 232246 167144 232814 168000
rect 232982 167144 233550 168000
rect 233718 167144 234286 168000
rect 234454 167144 235114 168000
rect 235282 167144 235850 168000
rect 236018 167144 236586 168000
rect 236754 167144 237322 168000
rect 237490 167144 238150 168000
rect 238318 167144 238886 168000
rect 239054 167144 239622 168000
rect 239790 167144 240358 168000
rect 240526 167144 241094 168000
rect 241262 167144 241922 168000
rect 242090 167144 242658 168000
rect 242826 167144 243394 168000
rect 243562 167144 244130 168000
rect 244298 167144 244866 168000
rect 245034 167144 245694 168000
rect 245862 167144 246430 168000
rect 246598 167144 247166 168000
rect 247334 167144 247902 168000
rect 248070 167144 248638 168000
rect 248806 167144 249466 168000
rect 249634 167144 250202 168000
rect 250370 167144 250938 168000
rect 251106 167144 251674 168000
rect 251842 167144 252410 168000
rect 252578 167144 253238 168000
rect 253406 167144 253974 168000
rect 254142 167144 254710 168000
rect 254878 167144 255446 168000
rect 255614 167144 256182 168000
rect 256350 167144 257010 168000
rect 257178 167144 257746 168000
rect 257914 167144 258482 168000
rect 258650 167144 259218 168000
rect 259386 167144 259954 168000
rect 260122 167144 260782 168000
rect 260950 167144 261518 168000
rect 261686 167144 262254 168000
rect 262422 167144 262990 168000
rect 263158 167144 263818 168000
rect 263986 167144 264554 168000
rect 264722 167144 265290 168000
rect 265458 167144 266026 168000
rect 266194 167144 266762 168000
rect 266930 167144 267590 168000
rect 267758 167144 268326 168000
rect 268494 167144 269062 168000
rect 269230 167144 269798 168000
rect 269966 167144 270534 168000
rect 270702 167144 271362 168000
rect 271530 167144 272098 168000
rect 272266 167144 272834 168000
rect 273002 167144 273570 168000
rect 273738 167144 274306 168000
rect 274474 167144 275134 168000
rect 275302 167144 275870 168000
rect 276038 167144 276606 168000
rect 276774 167144 277342 168000
rect 277510 167144 278078 168000
rect 278246 167144 278906 168000
rect 279074 167144 279642 168000
rect 279810 167144 280378 168000
rect 280546 167144 281114 168000
rect 281282 167144 281850 168000
rect 282018 167144 282678 168000
rect 282846 167144 283414 168000
rect 283582 167144 284150 168000
rect 284318 167144 284886 168000
rect 285054 167144 285714 168000
rect 285882 167144 286450 168000
rect 286618 167144 287186 168000
rect 287354 167144 287922 168000
rect 288090 167144 288658 168000
rect 288826 167144 289486 168000
rect 289654 167144 290222 168000
rect 290390 167144 290958 168000
rect 291126 167144 291694 168000
rect 291862 167144 292430 168000
rect 292598 167144 293258 168000
rect 293426 167144 293994 168000
rect 294162 167144 294730 168000
rect 294898 167144 295466 168000
rect 295634 167144 296202 168000
rect 296370 167144 297030 168000
rect 297198 167144 297766 168000
rect 297934 167144 298502 168000
rect 298670 167144 299238 168000
rect 299406 167144 299974 168000
rect 300142 167144 300802 168000
rect 300970 167144 301538 168000
rect 301706 167144 302274 168000
rect 302442 167144 303010 168000
rect 303178 167144 303746 168000
rect 303914 167144 304574 168000
rect 304742 167144 305310 168000
rect 305478 167144 306046 168000
rect 306214 167144 306782 168000
rect 306950 167144 307518 168000
rect 307686 167144 308346 168000
rect 308514 167144 309082 168000
rect 309250 167144 309818 168000
rect 309986 167144 310554 168000
rect 310722 167144 311382 168000
rect 311550 167144 312118 168000
rect 312286 167144 312854 168000
rect 313022 167144 313590 168000
rect 313758 167144 314326 168000
rect 314494 167144 315154 168000
rect 315322 167144 315890 168000
rect 316058 167144 316626 168000
rect 316794 167144 317362 168000
rect 317530 167144 318098 168000
rect 318266 167144 318926 168000
rect 319094 167144 319662 168000
rect 319830 167144 320398 168000
rect 320566 167144 321134 168000
rect 321302 167144 321870 168000
rect 322038 167144 322698 168000
rect 322866 167144 323434 168000
rect 323602 167144 324170 168000
rect 324338 167144 324906 168000
rect 325074 167144 325642 168000
rect 325810 167144 326470 168000
rect 326638 167144 327206 168000
rect 327374 167144 327942 168000
rect 328110 167144 328678 168000
rect 328846 167144 329414 168000
rect 329582 167144 330242 168000
rect 330410 167144 330978 168000
rect 331146 167144 331714 168000
rect 331882 167144 332450 168000
rect 332618 167144 333278 168000
rect 333446 167144 334014 168000
rect 334182 167144 334750 168000
rect 334918 167144 335486 168000
rect 335654 167144 336222 168000
rect 336390 167144 337050 168000
rect 337218 167144 337786 168000
rect 337954 167144 338522 168000
rect 338690 167144 339258 168000
rect 339426 167144 339994 168000
rect 340162 167144 340822 168000
rect 340990 167144 341558 168000
rect 341726 167144 342294 168000
rect 342462 167144 343030 168000
rect 343198 167144 343766 168000
rect 343934 167144 344594 168000
rect 344762 167144 345330 168000
rect 345498 167144 346066 168000
rect 346234 167144 346802 168000
rect 346970 167144 347538 168000
rect 347706 167144 348366 168000
rect 348534 167144 349102 168000
rect 349270 167144 349838 168000
rect 350006 167144 350574 168000
rect 350742 167144 351310 168000
rect 351478 167144 352138 168000
rect 352306 167144 352874 168000
rect 353042 167144 353610 168000
rect 353778 167144 354346 168000
rect 354514 167144 355082 168000
rect 355250 167144 355910 168000
rect 356078 167144 356646 168000
rect 356814 167144 357382 168000
rect 357550 167144 358118 168000
rect 358286 167144 358946 168000
rect 359114 167144 359682 168000
rect 359850 167144 360418 168000
rect 360586 167144 361154 168000
rect 361322 167144 361890 168000
rect 362058 167144 362718 168000
rect 362886 167144 363454 168000
rect 363622 167144 364190 168000
rect 364358 167144 364926 168000
rect 365094 167144 365662 168000
rect 365830 167144 366490 168000
rect 366658 167144 367226 168000
rect 367394 167144 367962 168000
rect 368130 167144 368698 168000
rect 368866 167144 369434 168000
rect 369602 167144 370262 168000
rect 370430 167144 370998 168000
rect 371166 167144 371734 168000
rect 371902 167144 372470 168000
rect 372638 167144 373206 168000
rect 373374 167144 374034 168000
rect 374202 167144 374770 168000
rect 374938 167144 375506 168000
rect 375674 167144 376242 168000
rect 376410 167144 376978 168000
rect 377146 167144 377806 168000
rect 377974 167144 378542 168000
rect 378710 167144 379278 168000
rect 379446 167144 380014 168000
rect 380182 167144 380842 168000
rect 381010 167144 381578 168000
rect 381746 167144 382314 168000
rect 382482 167144 383050 168000
rect 383218 167144 383786 168000
rect 383954 167144 384614 168000
rect 384782 167144 385350 168000
rect 385518 167144 386086 168000
rect 386254 167144 386822 168000
rect 386990 167144 387558 168000
rect 387726 167144 388386 168000
rect 388554 167144 389122 168000
rect 389290 167144 389858 168000
rect 390026 167144 390594 168000
rect 390762 167144 391330 168000
rect 391498 167144 392158 168000
rect 392326 167144 392894 168000
rect 393062 167144 393630 168000
rect 393798 167144 394366 168000
rect 394534 167144 395102 168000
rect 395270 167144 395930 168000
rect 396098 167144 396666 168000
rect 396834 167144 397402 168000
rect 397570 167144 398138 168000
rect 398306 167144 398874 168000
rect 399042 167144 399702 168000
rect 399870 167144 400438 168000
rect 400606 167144 401174 168000
rect 401342 167144 401910 168000
rect 402078 167144 402646 168000
rect 402814 167144 403474 168000
rect 403642 167144 404210 168000
rect 404378 167144 404946 168000
rect 405114 167144 405682 168000
rect 405850 167144 406510 168000
rect 406678 167144 407246 168000
rect 407414 167144 407982 168000
rect 408150 167144 408718 168000
rect 408886 167144 409454 168000
rect 409622 167144 410282 168000
rect 410450 167144 411018 168000
rect 411186 167144 411754 168000
rect 411922 167144 412490 168000
rect 412658 167144 413226 168000
rect 413394 167144 414054 168000
rect 414222 167144 414790 168000
rect 414958 167144 415526 168000
rect 415694 167144 416262 168000
rect 416430 167144 416998 168000
rect 417166 167144 417826 168000
rect 417994 167144 418562 168000
rect 418730 167144 419298 168000
rect 419466 167144 420034 168000
rect 420202 167144 420770 168000
rect 420938 167144 421598 168000
rect 421766 167144 422334 168000
rect 422502 167144 423070 168000
rect 423238 167144 423806 168000
rect 423974 167144 424542 168000
rect 424710 167144 425370 168000
rect 425538 167144 426106 168000
rect 426274 167144 426842 168000
rect 427010 167144 427578 168000
rect 427746 167144 428406 168000
rect 428574 167144 429142 168000
rect 429310 167144 429878 168000
rect 430046 167144 430614 168000
rect 430782 167144 431350 168000
rect 431518 167144 432178 168000
rect 432346 167144 432914 168000
rect 433082 167144 433650 168000
rect 433818 167144 434386 168000
rect 434554 167144 435122 168000
rect 435290 167144 435950 168000
rect 436118 167144 436686 168000
rect 436854 167144 437422 168000
rect 437590 167144 438158 168000
rect 438326 167144 438894 168000
rect 439062 167144 439722 168000
rect 439890 167144 440458 168000
rect 440626 167144 441194 168000
rect 441362 167144 441930 168000
rect 442098 167144 442666 168000
rect 442834 167144 443494 168000
rect 443662 167144 444230 168000
rect 444398 167144 444966 168000
rect 445134 167144 445702 168000
rect 445870 167144 446438 168000
rect 446606 167144 447266 168000
rect 447434 167144 448002 168000
rect 448170 167144 448738 168000
rect 448906 167144 449474 168000
rect 18 856 449572 167144
rect 18 800 8610 856
rect 8778 800 25906 856
rect 26074 800 43202 856
rect 43370 800 60498 856
rect 60666 800 77794 856
rect 77962 800 95090 856
rect 95258 800 112386 856
rect 112554 800 129682 856
rect 129850 800 146978 856
rect 147146 800 164366 856
rect 164534 800 181662 856
rect 181830 800 198958 856
rect 199126 800 216254 856
rect 216422 800 233550 856
rect 233718 800 250846 856
rect 251014 800 268142 856
rect 268310 800 285438 856
rect 285606 800 302734 856
rect 302902 800 320122 856
rect 320290 800 337418 856
rect 337586 800 354714 856
rect 354882 800 372010 856
rect 372178 800 389306 856
rect 389474 800 406602 856
rect 406770 800 423898 856
rect 424066 800 441194 856
rect 441362 800 449572 856
<< metal3 >>
rect 0 167424 800 167544
rect 449200 166880 450000 167000
rect 0 166608 800 166728
rect 0 165928 800 166048
rect 0 165112 800 165232
rect 449200 164976 450000 165096
rect 0 164432 800 164552
rect 0 163616 800 163736
rect 449200 163072 450000 163192
rect 0 162800 800 162920
rect 0 162120 800 162240
rect 0 161304 800 161424
rect 449200 161168 450000 161288
rect 0 160624 800 160744
rect 0 159808 800 159928
rect 449200 159264 450000 159384
rect 0 158992 800 159112
rect 0 158312 800 158432
rect 0 157496 800 157616
rect 449200 157360 450000 157480
rect 0 156816 800 156936
rect 0 156000 800 156120
rect 0 155320 800 155440
rect 449200 155456 450000 155576
rect 0 154504 800 154624
rect 0 153688 800 153808
rect 449200 153552 450000 153672
rect 0 153008 800 153128
rect 0 152192 800 152312
rect 0 151512 800 151632
rect 449200 151648 450000 151768
rect 0 150696 800 150816
rect 0 149880 800 150000
rect 449200 149744 450000 149864
rect 0 149200 800 149320
rect 0 148384 800 148504
rect 0 147704 800 147824
rect 449200 147840 450000 147960
rect 0 146888 800 147008
rect 0 146072 800 146192
rect 449200 145936 450000 146056
rect 0 145392 800 145512
rect 0 144576 800 144696
rect 0 143896 800 144016
rect 449200 144032 450000 144152
rect 0 143080 800 143200
rect 0 142400 800 142520
rect 449200 142128 450000 142248
rect 0 141584 800 141704
rect 0 140768 800 140888
rect 0 140088 800 140208
rect 449200 140224 450000 140344
rect 0 139272 800 139392
rect 0 138592 800 138712
rect 449200 138320 450000 138440
rect 0 137776 800 137896
rect 0 136960 800 137080
rect 0 136280 800 136400
rect 449200 136416 450000 136536
rect 0 135464 800 135584
rect 0 134784 800 134904
rect 449200 134512 450000 134632
rect 0 133968 800 134088
rect 0 133152 800 133272
rect 0 132472 800 132592
rect 449200 132608 450000 132728
rect 0 131656 800 131776
rect 0 130976 800 131096
rect 449200 130704 450000 130824
rect 0 130160 800 130280
rect 0 129480 800 129600
rect 0 128664 800 128784
rect 449200 128800 450000 128920
rect 0 127848 800 127968
rect 0 127168 800 127288
rect 449200 126896 450000 127016
rect 0 126352 800 126472
rect 0 125672 800 125792
rect 0 124856 800 124976
rect 449200 124992 450000 125112
rect 0 124040 800 124160
rect 0 123360 800 123480
rect 449200 123088 450000 123208
rect 0 122544 800 122664
rect 0 121864 800 121984
rect 0 121048 800 121168
rect 449200 121184 450000 121304
rect 0 120232 800 120352
rect 0 119552 800 119672
rect 449200 119280 450000 119400
rect 0 118736 800 118856
rect 0 118056 800 118176
rect 0 117240 800 117360
rect 449200 117376 450000 117496
rect 0 116560 800 116680
rect 0 115744 800 115864
rect 449200 115472 450000 115592
rect 0 114928 800 115048
rect 0 114248 800 114368
rect 0 113432 800 113552
rect 449200 113568 450000 113688
rect 0 112752 800 112872
rect 0 111936 800 112056
rect 449200 111528 450000 111648
rect 0 111120 800 111240
rect 0 110440 800 110560
rect 0 109624 800 109744
rect 449200 109624 450000 109744
rect 0 108944 800 109064
rect 0 108128 800 108248
rect 449200 107720 450000 107840
rect 0 107312 800 107432
rect 0 106632 800 106752
rect 0 105816 800 105936
rect 449200 105816 450000 105936
rect 0 105136 800 105256
rect 0 104320 800 104440
rect 449200 103912 450000 104032
rect 0 103640 800 103760
rect 0 102824 800 102944
rect 0 102008 800 102128
rect 449200 102008 450000 102128
rect 0 101328 800 101448
rect 0 100512 800 100632
rect 449200 100104 450000 100224
rect 0 99832 800 99952
rect 0 99016 800 99136
rect 0 98200 800 98320
rect 449200 98200 450000 98320
rect 0 97520 800 97640
rect 0 96704 800 96824
rect 449200 96296 450000 96416
rect 0 96024 800 96144
rect 0 95208 800 95328
rect 0 94392 800 94512
rect 449200 94392 450000 94512
rect 0 93712 800 93832
rect 0 92896 800 93016
rect 449200 92488 450000 92608
rect 0 92216 800 92336
rect 0 91400 800 91520
rect 0 90720 800 90840
rect 449200 90584 450000 90704
rect 0 89904 800 90024
rect 0 89088 800 89208
rect 449200 88680 450000 88800
rect 0 88408 800 88528
rect 0 87592 800 87712
rect 0 86912 800 87032
rect 449200 86776 450000 86896
rect 0 86096 800 86216
rect 0 85280 800 85400
rect 449200 84872 450000 84992
rect 0 84600 800 84720
rect 0 83784 800 83904
rect 0 83104 800 83224
rect 449200 82968 450000 83088
rect 0 82288 800 82408
rect 0 81472 800 81592
rect 449200 81064 450000 81184
rect 0 80792 800 80912
rect 0 79976 800 80096
rect 0 79296 800 79416
rect 449200 79160 450000 79280
rect 0 78480 800 78600
rect 0 77800 800 77920
rect 449200 77256 450000 77376
rect 0 76984 800 77104
rect 0 76168 800 76288
rect 0 75488 800 75608
rect 449200 75352 450000 75472
rect 0 74672 800 74792
rect 0 73992 800 74112
rect 449200 73448 450000 73568
rect 0 73176 800 73296
rect 0 72360 800 72480
rect 0 71680 800 71800
rect 449200 71544 450000 71664
rect 0 70864 800 70984
rect 0 70184 800 70304
rect 449200 69640 450000 69760
rect 0 69368 800 69488
rect 0 68552 800 68672
rect 0 67872 800 67992
rect 449200 67736 450000 67856
rect 0 67056 800 67176
rect 0 66376 800 66496
rect 449200 65832 450000 65952
rect 0 65560 800 65680
rect 0 64880 800 65000
rect 0 64064 800 64184
rect 449200 63928 450000 64048
rect 0 63248 800 63368
rect 0 62568 800 62688
rect 449200 62024 450000 62144
rect 0 61752 800 61872
rect 0 61072 800 61192
rect 0 60256 800 60376
rect 449200 60120 450000 60240
rect 0 59440 800 59560
rect 0 58760 800 58880
rect 449200 58216 450000 58336
rect 0 57944 800 58064
rect 0 57264 800 57384
rect 0 56448 800 56568
rect 449200 56176 450000 56296
rect 0 55632 800 55752
rect 0 54952 800 55072
rect 0 54136 800 54256
rect 449200 54272 450000 54392
rect 0 53456 800 53576
rect 0 52640 800 52760
rect 449200 52368 450000 52488
rect 0 51960 800 52080
rect 0 51144 800 51264
rect 0 50328 800 50448
rect 449200 50464 450000 50584
rect 0 49648 800 49768
rect 0 48832 800 48952
rect 449200 48560 450000 48680
rect 0 48152 800 48272
rect 0 47336 800 47456
rect 0 46520 800 46640
rect 449200 46656 450000 46776
rect 0 45840 800 45960
rect 0 45024 800 45144
rect 449200 44752 450000 44872
rect 0 44344 800 44464
rect 0 43528 800 43648
rect 0 42712 800 42832
rect 449200 42848 450000 42968
rect 0 42032 800 42152
rect 0 41216 800 41336
rect 449200 40944 450000 41064
rect 0 40536 800 40656
rect 0 39720 800 39840
rect 0 39040 800 39160
rect 449200 39040 450000 39160
rect 0 38224 800 38344
rect 0 37408 800 37528
rect 449200 37136 450000 37256
rect 0 36728 800 36848
rect 0 35912 800 36032
rect 0 35232 800 35352
rect 449200 35232 450000 35352
rect 0 34416 800 34536
rect 0 33600 800 33720
rect 449200 33328 450000 33448
rect 0 32920 800 33040
rect 0 32104 800 32224
rect 0 31424 800 31544
rect 449200 31424 450000 31544
rect 0 30608 800 30728
rect 0 29792 800 29912
rect 449200 29520 450000 29640
rect 0 29112 800 29232
rect 0 28296 800 28416
rect 0 27616 800 27736
rect 449200 27616 450000 27736
rect 0 26800 800 26920
rect 0 26120 800 26240
rect 449200 25712 450000 25832
rect 0 25304 800 25424
rect 0 24488 800 24608
rect 0 23808 800 23928
rect 449200 23808 450000 23928
rect 0 22992 800 23112
rect 0 22312 800 22432
rect 449200 21904 450000 22024
rect 0 21496 800 21616
rect 0 20680 800 20800
rect 0 20000 800 20120
rect 449200 20000 450000 20120
rect 0 19184 800 19304
rect 0 18504 800 18624
rect 449200 18096 450000 18216
rect 0 17688 800 17808
rect 0 16872 800 16992
rect 0 16192 800 16312
rect 449200 16192 450000 16312
rect 0 15376 800 15496
rect 0 14696 800 14816
rect 449200 14288 450000 14408
rect 0 13880 800 14000
rect 0 13200 800 13320
rect 0 12384 800 12504
rect 449200 12384 450000 12504
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 449200 10480 450000 10600
rect 0 10072 800 10192
rect 0 9392 800 9512
rect 0 8576 800 8696
rect 449200 8576 450000 8696
rect 0 7760 800 7880
rect 0 7080 800 7200
rect 449200 6672 450000 6792
rect 0 6264 800 6384
rect 0 5584 800 5704
rect 0 4768 800 4888
rect 449200 4768 450000 4888
rect 0 3952 800 4072
rect 0 3272 800 3392
rect 449200 2864 450000 2984
rect 0 2456 800 2576
rect 0 1776 800 1896
rect 0 960 800 1080
rect 449200 960 450000 1080
rect 0 280 800 400
<< obsm3 >>
rect 880 167344 449200 167517
rect 13 167080 449200 167344
rect 13 166808 449120 167080
rect 880 166800 449120 166808
rect 880 166528 449200 166800
rect 13 166128 449200 166528
rect 880 165848 449200 166128
rect 13 165312 449200 165848
rect 880 165176 449200 165312
rect 880 165032 449120 165176
rect 13 164896 449120 165032
rect 13 164632 449200 164896
rect 880 164352 449200 164632
rect 13 163816 449200 164352
rect 880 163536 449200 163816
rect 13 163272 449200 163536
rect 13 163000 449120 163272
rect 880 162992 449120 163000
rect 880 162720 449200 162992
rect 13 162320 449200 162720
rect 880 162040 449200 162320
rect 13 161504 449200 162040
rect 880 161368 449200 161504
rect 880 161224 449120 161368
rect 13 161088 449120 161224
rect 13 160824 449200 161088
rect 880 160544 449200 160824
rect 13 160008 449200 160544
rect 880 159728 449200 160008
rect 13 159464 449200 159728
rect 13 159192 449120 159464
rect 880 159184 449120 159192
rect 880 158912 449200 159184
rect 13 158512 449200 158912
rect 880 158232 449200 158512
rect 13 157696 449200 158232
rect 880 157560 449200 157696
rect 880 157416 449120 157560
rect 13 157280 449120 157416
rect 13 157016 449200 157280
rect 880 156736 449200 157016
rect 13 156200 449200 156736
rect 880 155920 449200 156200
rect 13 155656 449200 155920
rect 13 155520 449120 155656
rect 880 155376 449120 155520
rect 880 155240 449200 155376
rect 13 154704 449200 155240
rect 880 154424 449200 154704
rect 13 153888 449200 154424
rect 880 153752 449200 153888
rect 880 153608 449120 153752
rect 13 153472 449120 153608
rect 13 153208 449200 153472
rect 880 152928 449200 153208
rect 13 152392 449200 152928
rect 880 152112 449200 152392
rect 13 151848 449200 152112
rect 13 151712 449120 151848
rect 880 151568 449120 151712
rect 880 151432 449200 151568
rect 13 150896 449200 151432
rect 880 150616 449200 150896
rect 13 150080 449200 150616
rect 880 149944 449200 150080
rect 880 149800 449120 149944
rect 13 149664 449120 149800
rect 13 149400 449200 149664
rect 880 149120 449200 149400
rect 13 148584 449200 149120
rect 880 148304 449200 148584
rect 13 148040 449200 148304
rect 13 147904 449120 148040
rect 880 147760 449120 147904
rect 880 147624 449200 147760
rect 13 147088 449200 147624
rect 880 146808 449200 147088
rect 13 146272 449200 146808
rect 880 146136 449200 146272
rect 880 145992 449120 146136
rect 13 145856 449120 145992
rect 13 145592 449200 145856
rect 880 145312 449200 145592
rect 13 144776 449200 145312
rect 880 144496 449200 144776
rect 13 144232 449200 144496
rect 13 144096 449120 144232
rect 880 143952 449120 144096
rect 880 143816 449200 143952
rect 13 143280 449200 143816
rect 880 143000 449200 143280
rect 13 142600 449200 143000
rect 880 142328 449200 142600
rect 880 142320 449120 142328
rect 13 142048 449120 142320
rect 13 141784 449200 142048
rect 880 141504 449200 141784
rect 13 140968 449200 141504
rect 880 140688 449200 140968
rect 13 140424 449200 140688
rect 13 140288 449120 140424
rect 880 140144 449120 140288
rect 880 140008 449200 140144
rect 13 139472 449200 140008
rect 880 139192 449200 139472
rect 13 138792 449200 139192
rect 880 138520 449200 138792
rect 880 138512 449120 138520
rect 13 138240 449120 138512
rect 13 137976 449200 138240
rect 880 137696 449200 137976
rect 13 137160 449200 137696
rect 880 136880 449200 137160
rect 13 136616 449200 136880
rect 13 136480 449120 136616
rect 880 136336 449120 136480
rect 880 136200 449200 136336
rect 13 135664 449200 136200
rect 880 135384 449200 135664
rect 13 134984 449200 135384
rect 880 134712 449200 134984
rect 880 134704 449120 134712
rect 13 134432 449120 134704
rect 13 134168 449200 134432
rect 880 133888 449200 134168
rect 13 133352 449200 133888
rect 880 133072 449200 133352
rect 13 132808 449200 133072
rect 13 132672 449120 132808
rect 880 132528 449120 132672
rect 880 132392 449200 132528
rect 13 131856 449200 132392
rect 880 131576 449200 131856
rect 13 131176 449200 131576
rect 880 130904 449200 131176
rect 880 130896 449120 130904
rect 13 130624 449120 130896
rect 13 130360 449200 130624
rect 880 130080 449200 130360
rect 13 129680 449200 130080
rect 880 129400 449200 129680
rect 13 129000 449200 129400
rect 13 128864 449120 129000
rect 880 128720 449120 128864
rect 880 128584 449200 128720
rect 13 128048 449200 128584
rect 880 127768 449200 128048
rect 13 127368 449200 127768
rect 880 127096 449200 127368
rect 880 127088 449120 127096
rect 13 126816 449120 127088
rect 13 126552 449200 126816
rect 880 126272 449200 126552
rect 13 125872 449200 126272
rect 880 125592 449200 125872
rect 13 125192 449200 125592
rect 13 125056 449120 125192
rect 880 124912 449120 125056
rect 880 124776 449200 124912
rect 13 124240 449200 124776
rect 880 123960 449200 124240
rect 13 123560 449200 123960
rect 880 123288 449200 123560
rect 880 123280 449120 123288
rect 13 123008 449120 123280
rect 13 122744 449200 123008
rect 880 122464 449200 122744
rect 13 122064 449200 122464
rect 880 121784 449200 122064
rect 13 121384 449200 121784
rect 13 121248 449120 121384
rect 880 121104 449120 121248
rect 880 120968 449200 121104
rect 13 120432 449200 120968
rect 880 120152 449200 120432
rect 13 119752 449200 120152
rect 880 119480 449200 119752
rect 880 119472 449120 119480
rect 13 119200 449120 119472
rect 13 118936 449200 119200
rect 880 118656 449200 118936
rect 13 118256 449200 118656
rect 880 117976 449200 118256
rect 13 117576 449200 117976
rect 13 117440 449120 117576
rect 880 117296 449120 117440
rect 880 117160 449200 117296
rect 13 116760 449200 117160
rect 880 116480 449200 116760
rect 13 115944 449200 116480
rect 880 115672 449200 115944
rect 880 115664 449120 115672
rect 13 115392 449120 115664
rect 13 115128 449200 115392
rect 880 114848 449200 115128
rect 13 114448 449200 114848
rect 880 114168 449200 114448
rect 13 113768 449200 114168
rect 13 113632 449120 113768
rect 880 113488 449120 113632
rect 880 113352 449200 113488
rect 13 112952 449200 113352
rect 880 112672 449200 112952
rect 13 112136 449200 112672
rect 880 111856 449200 112136
rect 13 111728 449200 111856
rect 13 111448 449120 111728
rect 13 111320 449200 111448
rect 880 111040 449200 111320
rect 13 110640 449200 111040
rect 880 110360 449200 110640
rect 13 109824 449200 110360
rect 880 109544 449120 109824
rect 13 109144 449200 109544
rect 880 108864 449200 109144
rect 13 108328 449200 108864
rect 880 108048 449200 108328
rect 13 107920 449200 108048
rect 13 107640 449120 107920
rect 13 107512 449200 107640
rect 880 107232 449200 107512
rect 13 106832 449200 107232
rect 880 106552 449200 106832
rect 13 106016 449200 106552
rect 880 105736 449120 106016
rect 13 105336 449200 105736
rect 880 105056 449200 105336
rect 13 104520 449200 105056
rect 880 104240 449200 104520
rect 13 104112 449200 104240
rect 13 103840 449120 104112
rect 880 103832 449120 103840
rect 880 103560 449200 103832
rect 13 103024 449200 103560
rect 880 102744 449200 103024
rect 13 102208 449200 102744
rect 880 101928 449120 102208
rect 13 101528 449200 101928
rect 880 101248 449200 101528
rect 13 100712 449200 101248
rect 880 100432 449200 100712
rect 13 100304 449200 100432
rect 13 100032 449120 100304
rect 880 100024 449120 100032
rect 880 99752 449200 100024
rect 13 99216 449200 99752
rect 880 98936 449200 99216
rect 13 98400 449200 98936
rect 880 98120 449120 98400
rect 13 97720 449200 98120
rect 880 97440 449200 97720
rect 13 96904 449200 97440
rect 880 96624 449200 96904
rect 13 96496 449200 96624
rect 13 96224 449120 96496
rect 880 96216 449120 96224
rect 880 95944 449200 96216
rect 13 95408 449200 95944
rect 880 95128 449200 95408
rect 13 94592 449200 95128
rect 880 94312 449120 94592
rect 13 93912 449200 94312
rect 880 93632 449200 93912
rect 13 93096 449200 93632
rect 880 92816 449200 93096
rect 13 92688 449200 92816
rect 13 92416 449120 92688
rect 880 92408 449120 92416
rect 880 92136 449200 92408
rect 13 91600 449200 92136
rect 880 91320 449200 91600
rect 13 90920 449200 91320
rect 880 90784 449200 90920
rect 880 90640 449120 90784
rect 13 90504 449120 90640
rect 13 90104 449200 90504
rect 880 89824 449200 90104
rect 13 89288 449200 89824
rect 880 89008 449200 89288
rect 13 88880 449200 89008
rect 13 88608 449120 88880
rect 880 88600 449120 88608
rect 880 88328 449200 88600
rect 13 87792 449200 88328
rect 880 87512 449200 87792
rect 13 87112 449200 87512
rect 880 86976 449200 87112
rect 880 86832 449120 86976
rect 13 86696 449120 86832
rect 13 86296 449200 86696
rect 880 86016 449200 86296
rect 13 85480 449200 86016
rect 880 85200 449200 85480
rect 13 85072 449200 85200
rect 13 84800 449120 85072
rect 880 84792 449120 84800
rect 880 84520 449200 84792
rect 13 83984 449200 84520
rect 880 83704 449200 83984
rect 13 83304 449200 83704
rect 880 83168 449200 83304
rect 880 83024 449120 83168
rect 13 82888 449120 83024
rect 13 82488 449200 82888
rect 880 82208 449200 82488
rect 13 81672 449200 82208
rect 880 81392 449200 81672
rect 13 81264 449200 81392
rect 13 80992 449120 81264
rect 880 80984 449120 80992
rect 880 80712 449200 80984
rect 13 80176 449200 80712
rect 880 79896 449200 80176
rect 13 79496 449200 79896
rect 880 79360 449200 79496
rect 880 79216 449120 79360
rect 13 79080 449120 79216
rect 13 78680 449200 79080
rect 880 78400 449200 78680
rect 13 78000 449200 78400
rect 880 77720 449200 78000
rect 13 77456 449200 77720
rect 13 77184 449120 77456
rect 880 77176 449120 77184
rect 880 76904 449200 77176
rect 13 76368 449200 76904
rect 880 76088 449200 76368
rect 13 75688 449200 76088
rect 880 75552 449200 75688
rect 880 75408 449120 75552
rect 13 75272 449120 75408
rect 13 74872 449200 75272
rect 880 74592 449200 74872
rect 13 74192 449200 74592
rect 880 73912 449200 74192
rect 13 73648 449200 73912
rect 13 73376 449120 73648
rect 880 73368 449120 73376
rect 880 73096 449200 73368
rect 13 72560 449200 73096
rect 880 72280 449200 72560
rect 13 71880 449200 72280
rect 880 71744 449200 71880
rect 880 71600 449120 71744
rect 13 71464 449120 71600
rect 13 71064 449200 71464
rect 880 70784 449200 71064
rect 13 70384 449200 70784
rect 880 70104 449200 70384
rect 13 69840 449200 70104
rect 13 69568 449120 69840
rect 880 69560 449120 69568
rect 880 69288 449200 69560
rect 13 68752 449200 69288
rect 880 68472 449200 68752
rect 13 68072 449200 68472
rect 880 67936 449200 68072
rect 880 67792 449120 67936
rect 13 67656 449120 67792
rect 13 67256 449200 67656
rect 880 66976 449200 67256
rect 13 66576 449200 66976
rect 880 66296 449200 66576
rect 13 66032 449200 66296
rect 13 65760 449120 66032
rect 880 65752 449120 65760
rect 880 65480 449200 65752
rect 13 65080 449200 65480
rect 880 64800 449200 65080
rect 13 64264 449200 64800
rect 880 64128 449200 64264
rect 880 63984 449120 64128
rect 13 63848 449120 63984
rect 13 63448 449200 63848
rect 880 63168 449200 63448
rect 13 62768 449200 63168
rect 880 62488 449200 62768
rect 13 62224 449200 62488
rect 13 61952 449120 62224
rect 880 61944 449120 61952
rect 880 61672 449200 61944
rect 13 61272 449200 61672
rect 880 60992 449200 61272
rect 13 60456 449200 60992
rect 880 60320 449200 60456
rect 880 60176 449120 60320
rect 13 60040 449120 60176
rect 13 59640 449200 60040
rect 880 59360 449200 59640
rect 13 58960 449200 59360
rect 880 58680 449200 58960
rect 13 58416 449200 58680
rect 13 58144 449120 58416
rect 880 58136 449120 58144
rect 880 57864 449200 58136
rect 13 57464 449200 57864
rect 880 57184 449200 57464
rect 13 56648 449200 57184
rect 880 56376 449200 56648
rect 880 56368 449120 56376
rect 13 56096 449120 56368
rect 13 55832 449200 56096
rect 880 55552 449200 55832
rect 13 55152 449200 55552
rect 880 54872 449200 55152
rect 13 54472 449200 54872
rect 13 54336 449120 54472
rect 880 54192 449120 54336
rect 880 54056 449200 54192
rect 13 53656 449200 54056
rect 880 53376 449200 53656
rect 13 52840 449200 53376
rect 880 52568 449200 52840
rect 880 52560 449120 52568
rect 13 52288 449120 52560
rect 13 52160 449200 52288
rect 880 51880 449200 52160
rect 13 51344 449200 51880
rect 880 51064 449200 51344
rect 13 50664 449200 51064
rect 13 50528 449120 50664
rect 880 50384 449120 50528
rect 880 50248 449200 50384
rect 13 49848 449200 50248
rect 880 49568 449200 49848
rect 13 49032 449200 49568
rect 880 48760 449200 49032
rect 880 48752 449120 48760
rect 13 48480 449120 48752
rect 13 48352 449200 48480
rect 880 48072 449200 48352
rect 13 47536 449200 48072
rect 880 47256 449200 47536
rect 13 46856 449200 47256
rect 13 46720 449120 46856
rect 880 46576 449120 46720
rect 880 46440 449200 46576
rect 13 46040 449200 46440
rect 880 45760 449200 46040
rect 13 45224 449200 45760
rect 880 44952 449200 45224
rect 880 44944 449120 44952
rect 13 44672 449120 44944
rect 13 44544 449200 44672
rect 880 44264 449200 44544
rect 13 43728 449200 44264
rect 880 43448 449200 43728
rect 13 43048 449200 43448
rect 13 42912 449120 43048
rect 880 42768 449120 42912
rect 880 42632 449200 42768
rect 13 42232 449200 42632
rect 880 41952 449200 42232
rect 13 41416 449200 41952
rect 880 41144 449200 41416
rect 880 41136 449120 41144
rect 13 40864 449120 41136
rect 13 40736 449200 40864
rect 880 40456 449200 40736
rect 13 39920 449200 40456
rect 880 39640 449200 39920
rect 13 39240 449200 39640
rect 880 38960 449120 39240
rect 13 38424 449200 38960
rect 880 38144 449200 38424
rect 13 37608 449200 38144
rect 880 37336 449200 37608
rect 880 37328 449120 37336
rect 13 37056 449120 37328
rect 13 36928 449200 37056
rect 880 36648 449200 36928
rect 13 36112 449200 36648
rect 880 35832 449200 36112
rect 13 35432 449200 35832
rect 880 35152 449120 35432
rect 13 34616 449200 35152
rect 880 34336 449200 34616
rect 13 33800 449200 34336
rect 880 33528 449200 33800
rect 880 33520 449120 33528
rect 13 33248 449120 33520
rect 13 33120 449200 33248
rect 880 32840 449200 33120
rect 13 32304 449200 32840
rect 880 32024 449200 32304
rect 13 31624 449200 32024
rect 880 31344 449120 31624
rect 13 30808 449200 31344
rect 880 30528 449200 30808
rect 13 29992 449200 30528
rect 880 29720 449200 29992
rect 880 29712 449120 29720
rect 13 29440 449120 29712
rect 13 29312 449200 29440
rect 880 29032 449200 29312
rect 13 28496 449200 29032
rect 880 28216 449200 28496
rect 13 27816 449200 28216
rect 880 27536 449120 27816
rect 13 27000 449200 27536
rect 880 26720 449200 27000
rect 13 26320 449200 26720
rect 880 26040 449200 26320
rect 13 25912 449200 26040
rect 13 25632 449120 25912
rect 13 25504 449200 25632
rect 880 25224 449200 25504
rect 13 24688 449200 25224
rect 880 24408 449200 24688
rect 13 24008 449200 24408
rect 880 23728 449120 24008
rect 13 23192 449200 23728
rect 880 22912 449200 23192
rect 13 22512 449200 22912
rect 880 22232 449200 22512
rect 13 22104 449200 22232
rect 13 21824 449120 22104
rect 13 21696 449200 21824
rect 880 21416 449200 21696
rect 13 20880 449200 21416
rect 880 20600 449200 20880
rect 13 20200 449200 20600
rect 880 19920 449120 20200
rect 13 19384 449200 19920
rect 880 19104 449200 19384
rect 13 18704 449200 19104
rect 880 18424 449200 18704
rect 13 18296 449200 18424
rect 13 18016 449120 18296
rect 13 17888 449200 18016
rect 880 17608 449200 17888
rect 13 17072 449200 17608
rect 880 16792 449200 17072
rect 13 16392 449200 16792
rect 880 16112 449120 16392
rect 13 15576 449200 16112
rect 880 15296 449200 15576
rect 13 14896 449200 15296
rect 880 14616 449200 14896
rect 13 14488 449200 14616
rect 13 14208 449120 14488
rect 13 14080 449200 14208
rect 880 13800 449200 14080
rect 13 13400 449200 13800
rect 880 13120 449200 13400
rect 13 12584 449200 13120
rect 880 12304 449120 12584
rect 13 11768 449200 12304
rect 880 11488 449200 11768
rect 13 11088 449200 11488
rect 880 10808 449200 11088
rect 13 10680 449200 10808
rect 13 10400 449120 10680
rect 13 10272 449200 10400
rect 880 9992 449200 10272
rect 13 9592 449200 9992
rect 880 9312 449200 9592
rect 13 8776 449200 9312
rect 880 8496 449120 8776
rect 13 7960 449200 8496
rect 880 7680 449200 7960
rect 13 7280 449200 7680
rect 880 7000 449200 7280
rect 13 6872 449200 7000
rect 13 6592 449120 6872
rect 13 6464 449200 6592
rect 880 6184 449200 6464
rect 13 5784 449200 6184
rect 880 5504 449200 5784
rect 13 4968 449200 5504
rect 880 4688 449120 4968
rect 13 4152 449200 4688
rect 880 3872 449200 4152
rect 13 3472 449200 3872
rect 880 3192 449200 3472
rect 13 3064 449200 3192
rect 13 2784 449120 3064
rect 13 2656 449200 2784
rect 880 2376 449200 2656
rect 13 1976 449200 2376
rect 880 1696 449200 1976
rect 13 1160 449200 1696
rect 880 880 449120 1160
rect 13 480 449200 880
rect 880 308 449200 480
<< metal4 >>
rect 4208 2128 4528 165424
rect 9208 2128 9528 165424
rect 14208 2128 14528 165424
rect 19208 2128 19528 165424
rect 24208 128152 24528 165424
rect 29208 128152 29528 165424
rect 34208 128152 34528 165424
rect 39208 128152 39528 165424
rect 44208 128152 44528 165424
rect 49208 128152 49528 165424
rect 54208 128152 54528 165424
rect 59208 128152 59528 165424
rect 64208 128152 64528 165424
rect 69208 128152 69528 165424
rect 74208 128152 74528 165424
rect 79208 128152 79528 165424
rect 84208 128152 84528 165424
rect 89208 128152 89528 165424
rect 94208 128152 94528 165424
rect 99208 128152 99528 165424
rect 104208 128152 104528 165424
rect 109208 128152 109528 165424
rect 114208 128152 114528 165424
rect 119208 128152 119528 165424
rect 124208 128152 124528 165424
rect 129208 128152 129528 165424
rect 134208 128152 134528 165424
rect 139208 128152 139528 165424
rect 144208 128152 144528 165424
rect 149208 128152 149528 165424
rect 154208 128152 154528 165424
rect 159208 128152 159528 165424
rect 164208 128152 164528 165424
rect 169208 128152 169528 165424
rect 174208 128152 174528 165424
rect 24208 2128 24528 21248
rect 29208 2128 29528 21248
rect 34208 2128 34528 21248
rect 39208 2128 39528 21248
rect 44208 2128 44528 21248
rect 49208 2128 49528 21248
rect 54208 2128 54528 21248
rect 59208 2128 59528 21248
rect 64208 2128 64528 21248
rect 69208 2128 69528 21248
rect 74208 2128 74528 21248
rect 79208 2128 79528 21248
rect 84208 2128 84528 21248
rect 89208 2128 89528 21248
rect 94208 2128 94528 21248
rect 99208 2128 99528 21248
rect 104208 2128 104528 21248
rect 109208 2128 109528 21248
rect 114208 2128 114528 21248
rect 119208 2128 119528 21248
rect 124208 2128 124528 21248
rect 129208 2128 129528 21248
rect 134208 2128 134528 21248
rect 139208 2128 139528 21248
rect 144208 2128 144528 21248
rect 149208 2128 149528 21248
rect 154208 2128 154528 21248
rect 159208 2128 159528 21248
rect 164208 2128 164528 21248
rect 169208 2128 169528 21248
rect 174208 2128 174528 21248
rect 179208 2128 179528 165424
rect 184208 2128 184528 165424
rect 189208 2128 189528 165424
rect 194208 2128 194528 165424
rect 199208 2128 199528 165424
rect 204208 2128 204528 165424
rect 209208 2128 209528 165424
rect 214208 2128 214528 165424
rect 219208 2128 219528 165424
rect 224208 2128 224528 165424
rect 229208 2128 229528 165424
rect 234208 2128 234528 165424
rect 239208 2128 239528 165424
rect 244208 2128 244528 165424
rect 249208 2128 249528 165424
rect 254208 2128 254528 165424
rect 259208 2128 259528 165424
rect 264208 2128 264528 165424
rect 269208 2128 269528 165424
rect 274208 2128 274528 165424
rect 279208 2128 279528 165424
rect 284208 2128 284528 165424
rect 289208 2128 289528 165424
rect 294208 2128 294528 165424
rect 299208 2128 299528 165424
rect 304208 2128 304528 165424
rect 309208 2128 309528 165424
rect 314208 2128 314528 165424
rect 319208 2128 319528 165424
rect 324208 2128 324528 165424
rect 329208 2128 329528 165424
rect 334208 2128 334528 165424
rect 339208 2128 339528 165424
rect 344208 2128 344528 165424
rect 349208 2128 349528 165424
rect 354208 2128 354528 165424
rect 359208 2128 359528 165424
rect 364208 2128 364528 165424
rect 369208 2128 369528 165424
rect 374208 2128 374528 165424
rect 379208 2128 379528 165424
rect 384208 2128 384528 165424
rect 389208 164296 389528 165424
rect 394208 164296 394528 165424
rect 399208 164296 399528 165424
rect 389208 2128 389528 145392
rect 394208 2128 394528 145392
rect 399208 2128 399528 145392
rect 404208 2128 404528 165424
rect 409208 2128 409528 165424
rect 414208 2128 414528 165424
rect 419208 2128 419528 165424
rect 424208 2128 424528 165424
rect 429208 2128 429528 165424
rect 434208 2128 434528 165424
rect 439208 2128 439528 165424
rect 444208 2128 444528 165424
<< obsm4 >>
rect 1899 165504 446877 166701
rect 1899 2048 4128 165504
rect 4608 2048 9128 165504
rect 9608 2048 14128 165504
rect 14608 2048 19128 165504
rect 19608 128072 24128 165504
rect 24608 128072 29128 165504
rect 29608 128072 34128 165504
rect 34608 128072 39128 165504
rect 39608 128072 44128 165504
rect 44608 128072 49128 165504
rect 49608 128072 54128 165504
rect 54608 128072 59128 165504
rect 59608 128072 64128 165504
rect 64608 128072 69128 165504
rect 69608 128072 74128 165504
rect 74608 128072 79128 165504
rect 79608 128072 84128 165504
rect 84608 128072 89128 165504
rect 89608 128072 94128 165504
rect 94608 128072 99128 165504
rect 99608 128072 104128 165504
rect 104608 128072 109128 165504
rect 109608 128072 114128 165504
rect 114608 128072 119128 165504
rect 119608 128072 124128 165504
rect 124608 128072 129128 165504
rect 129608 128072 134128 165504
rect 134608 128072 139128 165504
rect 139608 128072 144128 165504
rect 144608 128072 149128 165504
rect 149608 128072 154128 165504
rect 154608 128072 159128 165504
rect 159608 128072 164128 165504
rect 164608 128072 169128 165504
rect 169608 128072 174128 165504
rect 174608 128072 179128 165504
rect 19608 21328 179128 128072
rect 19608 2048 24128 21328
rect 24608 2048 29128 21328
rect 29608 2048 34128 21328
rect 34608 2048 39128 21328
rect 39608 2048 44128 21328
rect 44608 2048 49128 21328
rect 49608 2048 54128 21328
rect 54608 2048 59128 21328
rect 59608 2048 64128 21328
rect 64608 2048 69128 21328
rect 69608 2048 74128 21328
rect 74608 2048 79128 21328
rect 79608 2048 84128 21328
rect 84608 2048 89128 21328
rect 89608 2048 94128 21328
rect 94608 2048 99128 21328
rect 99608 2048 104128 21328
rect 104608 2048 109128 21328
rect 109608 2048 114128 21328
rect 114608 2048 119128 21328
rect 119608 2048 124128 21328
rect 124608 2048 129128 21328
rect 129608 2048 134128 21328
rect 134608 2048 139128 21328
rect 139608 2048 144128 21328
rect 144608 2048 149128 21328
rect 149608 2048 154128 21328
rect 154608 2048 159128 21328
rect 159608 2048 164128 21328
rect 164608 2048 169128 21328
rect 169608 2048 174128 21328
rect 174608 2048 179128 21328
rect 179608 2048 184128 165504
rect 184608 2048 189128 165504
rect 189608 2048 194128 165504
rect 194608 2048 199128 165504
rect 199608 2048 204128 165504
rect 204608 2048 209128 165504
rect 209608 2048 214128 165504
rect 214608 2048 219128 165504
rect 219608 2048 224128 165504
rect 224608 2048 229128 165504
rect 229608 2048 234128 165504
rect 234608 2048 239128 165504
rect 239608 2048 244128 165504
rect 244608 2048 249128 165504
rect 249608 2048 254128 165504
rect 254608 2048 259128 165504
rect 259608 2048 264128 165504
rect 264608 2048 269128 165504
rect 269608 2048 274128 165504
rect 274608 2048 279128 165504
rect 279608 2048 284128 165504
rect 284608 2048 289128 165504
rect 289608 2048 294128 165504
rect 294608 2048 299128 165504
rect 299608 2048 304128 165504
rect 304608 2048 309128 165504
rect 309608 2048 314128 165504
rect 314608 2048 319128 165504
rect 319608 2048 324128 165504
rect 324608 2048 329128 165504
rect 329608 2048 334128 165504
rect 334608 2048 339128 165504
rect 339608 2048 344128 165504
rect 344608 2048 349128 165504
rect 349608 2048 354128 165504
rect 354608 2048 359128 165504
rect 359608 2048 364128 165504
rect 364608 2048 369128 165504
rect 369608 2048 374128 165504
rect 374608 2048 379128 165504
rect 379608 2048 384128 165504
rect 384608 164216 389128 165504
rect 389608 164216 394128 165504
rect 394608 164216 399128 165504
rect 399608 164216 404128 165504
rect 384608 145472 404128 164216
rect 384608 2048 389128 145472
rect 389608 2048 394128 145472
rect 394608 2048 399128 145472
rect 399608 2048 404128 145472
rect 404608 2048 409128 165504
rect 409608 2048 414128 165504
rect 414608 2048 419128 165504
rect 419608 2048 424128 165504
rect 424608 2048 429128 165504
rect 429608 2048 434128 165504
rect 434608 2048 439128 165504
rect 439608 2048 444128 165504
rect 444608 2048 446877 165504
rect 1899 307 446877 2048
<< metal5 >>
rect 1104 161298 448868 161618
rect 1104 148298 448868 148618
rect 1104 135298 448868 135618
rect 1104 122298 448868 122618
rect 1104 109298 448868 109618
rect 1104 96298 448868 96618
rect 1104 83298 448868 83618
rect 1104 70298 448868 70618
rect 1104 57298 448868 57618
rect 1104 44298 448868 44618
rect 1104 31298 448868 31618
rect 1104 18298 448868 18618
rect 1104 5298 448868 5618
<< labels >>
rlabel metal2 s 25962 0 26018 800 6 clock
port 1 nsew signal input
rlabel metal2 s 386 167200 442 168000 6 core_clk
port 2 nsew signal output
rlabel metal2 s 1122 167200 1178 168000 6 core_rstn
port 3 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 216310 0 216366 800 6 flash_clk_ieb
port 5 nsew signal output
rlabel metal2 s 233606 0 233662 800 6 flash_clk_oeb
port 6 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 flash_csb
port 7 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 flash_csb_ieb
port 8 nsew signal output
rlabel metal2 s 181718 0 181774 800 6 flash_csb_oeb
port 9 nsew signal output
rlabel metal2 s 250902 0 250958 800 6 flash_io0_di
port 10 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 flash_io0_do
port 11 nsew signal output
rlabel metal2 s 285494 0 285550 800 6 flash_io0_ieb
port 12 nsew signal output
rlabel metal2 s 302790 0 302846 800 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal2 s 320178 0 320234 800 6 flash_io1_di
port 14 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 flash_io1_do
port 15 nsew signal output
rlabel metal2 s 354770 0 354826 800 6 flash_io1_ieb
port 16 nsew signal output
rlabel metal2 s 372066 0 372122 800 6 flash_io1_oeb
port 17 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 flash_io2_oeb
port 18 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 flash_io3_oeb
port 19 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 gpio_in_pad
port 20 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 gpio_inenb_pad
port 21 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 gpio_mode0_pad
port 22 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 gpio_mode1_pad
port 23 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 gpio_out_pad
port 24 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 gpio_outenb_pad
port 25 nsew signal output
rlabel metal3 s 449200 63928 450000 64048 6 jtag_out
port 26 nsew signal output
rlabel metal3 s 449200 65832 450000 65952 6 jtag_outenb
port 27 nsew signal output
rlabel metal2 s 2594 167200 2650 168000 6 la_iena[0]
port 28 nsew signal output
rlabel metal2 s 304630 167200 304686 168000 6 la_iena[100]
port 29 nsew signal output
rlabel metal2 s 307574 167200 307630 168000 6 la_iena[101]
port 30 nsew signal output
rlabel metal2 s 310610 167200 310666 168000 6 la_iena[102]
port 31 nsew signal output
rlabel metal2 s 313646 167200 313702 168000 6 la_iena[103]
port 32 nsew signal output
rlabel metal2 s 316682 167200 316738 168000 6 la_iena[104]
port 33 nsew signal output
rlabel metal2 s 319718 167200 319774 168000 6 la_iena[105]
port 34 nsew signal output
rlabel metal2 s 322754 167200 322810 168000 6 la_iena[106]
port 35 nsew signal output
rlabel metal2 s 325698 167200 325754 168000 6 la_iena[107]
port 36 nsew signal output
rlabel metal2 s 328734 167200 328790 168000 6 la_iena[108]
port 37 nsew signal output
rlabel metal2 s 331770 167200 331826 168000 6 la_iena[109]
port 38 nsew signal output
rlabel metal2 s 32770 167200 32826 168000 6 la_iena[10]
port 39 nsew signal output
rlabel metal2 s 334806 167200 334862 168000 6 la_iena[110]
port 40 nsew signal output
rlabel metal2 s 337842 167200 337898 168000 6 la_iena[111]
port 41 nsew signal output
rlabel metal2 s 340878 167200 340934 168000 6 la_iena[112]
port 42 nsew signal output
rlabel metal2 s 343822 167200 343878 168000 6 la_iena[113]
port 43 nsew signal output
rlabel metal2 s 346858 167200 346914 168000 6 la_iena[114]
port 44 nsew signal output
rlabel metal2 s 349894 167200 349950 168000 6 la_iena[115]
port 45 nsew signal output
rlabel metal2 s 352930 167200 352986 168000 6 la_iena[116]
port 46 nsew signal output
rlabel metal2 s 355966 167200 356022 168000 6 la_iena[117]
port 47 nsew signal output
rlabel metal2 s 359002 167200 359058 168000 6 la_iena[118]
port 48 nsew signal output
rlabel metal2 s 361946 167200 362002 168000 6 la_iena[119]
port 49 nsew signal output
rlabel metal2 s 35806 167200 35862 168000 6 la_iena[11]
port 50 nsew signal output
rlabel metal2 s 364982 167200 365038 168000 6 la_iena[120]
port 51 nsew signal output
rlabel metal2 s 368018 167200 368074 168000 6 la_iena[121]
port 52 nsew signal output
rlabel metal2 s 371054 167200 371110 168000 6 la_iena[122]
port 53 nsew signal output
rlabel metal2 s 374090 167200 374146 168000 6 la_iena[123]
port 54 nsew signal output
rlabel metal2 s 377034 167200 377090 168000 6 la_iena[124]
port 55 nsew signal output
rlabel metal2 s 380070 167200 380126 168000 6 la_iena[125]
port 56 nsew signal output
rlabel metal2 s 383106 167200 383162 168000 6 la_iena[126]
port 57 nsew signal output
rlabel metal2 s 386142 167200 386198 168000 6 la_iena[127]
port 58 nsew signal output
rlabel metal2 s 38842 167200 38898 168000 6 la_iena[12]
port 59 nsew signal output
rlabel metal2 s 41878 167200 41934 168000 6 la_iena[13]
port 60 nsew signal output
rlabel metal2 s 44914 167200 44970 168000 6 la_iena[14]
port 61 nsew signal output
rlabel metal2 s 47950 167200 48006 168000 6 la_iena[15]
port 62 nsew signal output
rlabel metal2 s 50894 167200 50950 168000 6 la_iena[16]
port 63 nsew signal output
rlabel metal2 s 53930 167200 53986 168000 6 la_iena[17]
port 64 nsew signal output
rlabel metal2 s 56966 167200 57022 168000 6 la_iena[18]
port 65 nsew signal output
rlabel metal2 s 60002 167200 60058 168000 6 la_iena[19]
port 66 nsew signal output
rlabel metal2 s 5630 167200 5686 168000 6 la_iena[1]
port 67 nsew signal output
rlabel metal2 s 63038 167200 63094 168000 6 la_iena[20]
port 68 nsew signal output
rlabel metal2 s 65982 167200 66038 168000 6 la_iena[21]
port 69 nsew signal output
rlabel metal2 s 69018 167200 69074 168000 6 la_iena[22]
port 70 nsew signal output
rlabel metal2 s 72054 167200 72110 168000 6 la_iena[23]
port 71 nsew signal output
rlabel metal2 s 75090 167200 75146 168000 6 la_iena[24]
port 72 nsew signal output
rlabel metal2 s 78126 167200 78182 168000 6 la_iena[25]
port 73 nsew signal output
rlabel metal2 s 81162 167200 81218 168000 6 la_iena[26]
port 74 nsew signal output
rlabel metal2 s 84106 167200 84162 168000 6 la_iena[27]
port 75 nsew signal output
rlabel metal2 s 87142 167200 87198 168000 6 la_iena[28]
port 76 nsew signal output
rlabel metal2 s 90178 167200 90234 168000 6 la_iena[29]
port 77 nsew signal output
rlabel metal2 s 8666 167200 8722 168000 6 la_iena[2]
port 78 nsew signal output
rlabel metal2 s 93214 167200 93270 168000 6 la_iena[30]
port 79 nsew signal output
rlabel metal2 s 96250 167200 96306 168000 6 la_iena[31]
port 80 nsew signal output
rlabel metal2 s 99286 167200 99342 168000 6 la_iena[32]
port 81 nsew signal output
rlabel metal2 s 102230 167200 102286 168000 6 la_iena[33]
port 82 nsew signal output
rlabel metal2 s 105266 167200 105322 168000 6 la_iena[34]
port 83 nsew signal output
rlabel metal2 s 108302 167200 108358 168000 6 la_iena[35]
port 84 nsew signal output
rlabel metal2 s 111338 167200 111394 168000 6 la_iena[36]
port 85 nsew signal output
rlabel metal2 s 114374 167200 114430 168000 6 la_iena[37]
port 86 nsew signal output
rlabel metal2 s 117318 167200 117374 168000 6 la_iena[38]
port 87 nsew signal output
rlabel metal2 s 120354 167200 120410 168000 6 la_iena[39]
port 88 nsew signal output
rlabel metal2 s 11702 167200 11758 168000 6 la_iena[3]
port 89 nsew signal output
rlabel metal2 s 123390 167200 123446 168000 6 la_iena[40]
port 90 nsew signal output
rlabel metal2 s 126426 167200 126482 168000 6 la_iena[41]
port 91 nsew signal output
rlabel metal2 s 129462 167200 129518 168000 6 la_iena[42]
port 92 nsew signal output
rlabel metal2 s 132498 167200 132554 168000 6 la_iena[43]
port 93 nsew signal output
rlabel metal2 s 135442 167200 135498 168000 6 la_iena[44]
port 94 nsew signal output
rlabel metal2 s 138478 167200 138534 168000 6 la_iena[45]
port 95 nsew signal output
rlabel metal2 s 141514 167200 141570 168000 6 la_iena[46]
port 96 nsew signal output
rlabel metal2 s 144550 167200 144606 168000 6 la_iena[47]
port 97 nsew signal output
rlabel metal2 s 147586 167200 147642 168000 6 la_iena[48]
port 98 nsew signal output
rlabel metal2 s 150622 167200 150678 168000 6 la_iena[49]
port 99 nsew signal output
rlabel metal2 s 14646 167200 14702 168000 6 la_iena[4]
port 100 nsew signal output
rlabel metal2 s 153566 167200 153622 168000 6 la_iena[50]
port 101 nsew signal output
rlabel metal2 s 156602 167200 156658 168000 6 la_iena[51]
port 102 nsew signal output
rlabel metal2 s 159638 167200 159694 168000 6 la_iena[52]
port 103 nsew signal output
rlabel metal2 s 162674 167200 162730 168000 6 la_iena[53]
port 104 nsew signal output
rlabel metal2 s 165710 167200 165766 168000 6 la_iena[54]
port 105 nsew signal output
rlabel metal2 s 168746 167200 168802 168000 6 la_iena[55]
port 106 nsew signal output
rlabel metal2 s 171690 167200 171746 168000 6 la_iena[56]
port 107 nsew signal output
rlabel metal2 s 174726 167200 174782 168000 6 la_iena[57]
port 108 nsew signal output
rlabel metal2 s 177762 167200 177818 168000 6 la_iena[58]
port 109 nsew signal output
rlabel metal2 s 180798 167200 180854 168000 6 la_iena[59]
port 110 nsew signal output
rlabel metal2 s 17682 167200 17738 168000 6 la_iena[5]
port 111 nsew signal output
rlabel metal2 s 183834 167200 183890 168000 6 la_iena[60]
port 112 nsew signal output
rlabel metal2 s 186778 167200 186834 168000 6 la_iena[61]
port 113 nsew signal output
rlabel metal2 s 189814 167200 189870 168000 6 la_iena[62]
port 114 nsew signal output
rlabel metal2 s 192850 167200 192906 168000 6 la_iena[63]
port 115 nsew signal output
rlabel metal2 s 195886 167200 195942 168000 6 la_iena[64]
port 116 nsew signal output
rlabel metal2 s 198922 167200 198978 168000 6 la_iena[65]
port 117 nsew signal output
rlabel metal2 s 201958 167200 202014 168000 6 la_iena[66]
port 118 nsew signal output
rlabel metal2 s 204902 167200 204958 168000 6 la_iena[67]
port 119 nsew signal output
rlabel metal2 s 207938 167200 207994 168000 6 la_iena[68]
port 120 nsew signal output
rlabel metal2 s 210974 167200 211030 168000 6 la_iena[69]
port 121 nsew signal output
rlabel metal2 s 20718 167200 20774 168000 6 la_iena[6]
port 122 nsew signal output
rlabel metal2 s 214010 167200 214066 168000 6 la_iena[70]
port 123 nsew signal output
rlabel metal2 s 217046 167200 217102 168000 6 la_iena[71]
port 124 nsew signal output
rlabel metal2 s 220082 167200 220138 168000 6 la_iena[72]
port 125 nsew signal output
rlabel metal2 s 223026 167200 223082 168000 6 la_iena[73]
port 126 nsew signal output
rlabel metal2 s 226062 167200 226118 168000 6 la_iena[74]
port 127 nsew signal output
rlabel metal2 s 229098 167200 229154 168000 6 la_iena[75]
port 128 nsew signal output
rlabel metal2 s 232134 167200 232190 168000 6 la_iena[76]
port 129 nsew signal output
rlabel metal2 s 235170 167200 235226 168000 6 la_iena[77]
port 130 nsew signal output
rlabel metal2 s 238206 167200 238262 168000 6 la_iena[78]
port 131 nsew signal output
rlabel metal2 s 241150 167200 241206 168000 6 la_iena[79]
port 132 nsew signal output
rlabel metal2 s 23754 167200 23810 168000 6 la_iena[7]
port 133 nsew signal output
rlabel metal2 s 244186 167200 244242 168000 6 la_iena[80]
port 134 nsew signal output
rlabel metal2 s 247222 167200 247278 168000 6 la_iena[81]
port 135 nsew signal output
rlabel metal2 s 250258 167200 250314 168000 6 la_iena[82]
port 136 nsew signal output
rlabel metal2 s 253294 167200 253350 168000 6 la_iena[83]
port 137 nsew signal output
rlabel metal2 s 256238 167200 256294 168000 6 la_iena[84]
port 138 nsew signal output
rlabel metal2 s 259274 167200 259330 168000 6 la_iena[85]
port 139 nsew signal output
rlabel metal2 s 262310 167200 262366 168000 6 la_iena[86]
port 140 nsew signal output
rlabel metal2 s 265346 167200 265402 168000 6 la_iena[87]
port 141 nsew signal output
rlabel metal2 s 268382 167200 268438 168000 6 la_iena[88]
port 142 nsew signal output
rlabel metal2 s 271418 167200 271474 168000 6 la_iena[89]
port 143 nsew signal output
rlabel metal2 s 26790 167200 26846 168000 6 la_iena[8]
port 144 nsew signal output
rlabel metal2 s 274362 167200 274418 168000 6 la_iena[90]
port 145 nsew signal output
rlabel metal2 s 277398 167200 277454 168000 6 la_iena[91]
port 146 nsew signal output
rlabel metal2 s 280434 167200 280490 168000 6 la_iena[92]
port 147 nsew signal output
rlabel metal2 s 283470 167200 283526 168000 6 la_iena[93]
port 148 nsew signal output
rlabel metal2 s 286506 167200 286562 168000 6 la_iena[94]
port 149 nsew signal output
rlabel metal2 s 289542 167200 289598 168000 6 la_iena[95]
port 150 nsew signal output
rlabel metal2 s 292486 167200 292542 168000 6 la_iena[96]
port 151 nsew signal output
rlabel metal2 s 295522 167200 295578 168000 6 la_iena[97]
port 152 nsew signal output
rlabel metal2 s 298558 167200 298614 168000 6 la_iena[98]
port 153 nsew signal output
rlabel metal2 s 301594 167200 301650 168000 6 la_iena[99]
port 154 nsew signal output
rlabel metal2 s 29826 167200 29882 168000 6 la_iena[9]
port 155 nsew signal output
rlabel metal2 s 3330 167200 3386 168000 6 la_input[0]
port 156 nsew signal input
rlabel metal2 s 305366 167200 305422 168000 6 la_input[100]
port 157 nsew signal input
rlabel metal2 s 308402 167200 308458 168000 6 la_input[101]
port 158 nsew signal input
rlabel metal2 s 311438 167200 311494 168000 6 la_input[102]
port 159 nsew signal input
rlabel metal2 s 314382 167200 314438 168000 6 la_input[103]
port 160 nsew signal input
rlabel metal2 s 317418 167200 317474 168000 6 la_input[104]
port 161 nsew signal input
rlabel metal2 s 320454 167200 320510 168000 6 la_input[105]
port 162 nsew signal input
rlabel metal2 s 323490 167200 323546 168000 6 la_input[106]
port 163 nsew signal input
rlabel metal2 s 326526 167200 326582 168000 6 la_input[107]
port 164 nsew signal input
rlabel metal2 s 329470 167200 329526 168000 6 la_input[108]
port 165 nsew signal input
rlabel metal2 s 332506 167200 332562 168000 6 la_input[109]
port 166 nsew signal input
rlabel metal2 s 33598 167200 33654 168000 6 la_input[10]
port 167 nsew signal input
rlabel metal2 s 335542 167200 335598 168000 6 la_input[110]
port 168 nsew signal input
rlabel metal2 s 338578 167200 338634 168000 6 la_input[111]
port 169 nsew signal input
rlabel metal2 s 341614 167200 341670 168000 6 la_input[112]
port 170 nsew signal input
rlabel metal2 s 344650 167200 344706 168000 6 la_input[113]
port 171 nsew signal input
rlabel metal2 s 347594 167200 347650 168000 6 la_input[114]
port 172 nsew signal input
rlabel metal2 s 350630 167200 350686 168000 6 la_input[115]
port 173 nsew signal input
rlabel metal2 s 353666 167200 353722 168000 6 la_input[116]
port 174 nsew signal input
rlabel metal2 s 356702 167200 356758 168000 6 la_input[117]
port 175 nsew signal input
rlabel metal2 s 359738 167200 359794 168000 6 la_input[118]
port 176 nsew signal input
rlabel metal2 s 362774 167200 362830 168000 6 la_input[119]
port 177 nsew signal input
rlabel metal2 s 36542 167200 36598 168000 6 la_input[11]
port 178 nsew signal input
rlabel metal2 s 365718 167200 365774 168000 6 la_input[120]
port 179 nsew signal input
rlabel metal2 s 368754 167200 368810 168000 6 la_input[121]
port 180 nsew signal input
rlabel metal2 s 371790 167200 371846 168000 6 la_input[122]
port 181 nsew signal input
rlabel metal2 s 374826 167200 374882 168000 6 la_input[123]
port 182 nsew signal input
rlabel metal2 s 377862 167200 377918 168000 6 la_input[124]
port 183 nsew signal input
rlabel metal2 s 380898 167200 380954 168000 6 la_input[125]
port 184 nsew signal input
rlabel metal2 s 383842 167200 383898 168000 6 la_input[126]
port 185 nsew signal input
rlabel metal2 s 386878 167200 386934 168000 6 la_input[127]
port 186 nsew signal input
rlabel metal2 s 39578 167200 39634 168000 6 la_input[12]
port 187 nsew signal input
rlabel metal2 s 42614 167200 42670 168000 6 la_input[13]
port 188 nsew signal input
rlabel metal2 s 45650 167200 45706 168000 6 la_input[14]
port 189 nsew signal input
rlabel metal2 s 48686 167200 48742 168000 6 la_input[15]
port 190 nsew signal input
rlabel metal2 s 51722 167200 51778 168000 6 la_input[16]
port 191 nsew signal input
rlabel metal2 s 54666 167200 54722 168000 6 la_input[17]
port 192 nsew signal input
rlabel metal2 s 57702 167200 57758 168000 6 la_input[18]
port 193 nsew signal input
rlabel metal2 s 60738 167200 60794 168000 6 la_input[19]
port 194 nsew signal input
rlabel metal2 s 6366 167200 6422 168000 6 la_input[1]
port 195 nsew signal input
rlabel metal2 s 63774 167200 63830 168000 6 la_input[20]
port 196 nsew signal input
rlabel metal2 s 66810 167200 66866 168000 6 la_input[21]
port 197 nsew signal input
rlabel metal2 s 69754 167200 69810 168000 6 la_input[22]
port 198 nsew signal input
rlabel metal2 s 72790 167200 72846 168000 6 la_input[23]
port 199 nsew signal input
rlabel metal2 s 75826 167200 75882 168000 6 la_input[24]
port 200 nsew signal input
rlabel metal2 s 78862 167200 78918 168000 6 la_input[25]
port 201 nsew signal input
rlabel metal2 s 81898 167200 81954 168000 6 la_input[26]
port 202 nsew signal input
rlabel metal2 s 84934 167200 84990 168000 6 la_input[27]
port 203 nsew signal input
rlabel metal2 s 87878 167200 87934 168000 6 la_input[28]
port 204 nsew signal input
rlabel metal2 s 90914 167200 90970 168000 6 la_input[29]
port 205 nsew signal input
rlabel metal2 s 9402 167200 9458 168000 6 la_input[2]
port 206 nsew signal input
rlabel metal2 s 93950 167200 94006 168000 6 la_input[30]
port 207 nsew signal input
rlabel metal2 s 96986 167200 97042 168000 6 la_input[31]
port 208 nsew signal input
rlabel metal2 s 100022 167200 100078 168000 6 la_input[32]
port 209 nsew signal input
rlabel metal2 s 103058 167200 103114 168000 6 la_input[33]
port 210 nsew signal input
rlabel metal2 s 106002 167200 106058 168000 6 la_input[34]
port 211 nsew signal input
rlabel metal2 s 109038 167200 109094 168000 6 la_input[35]
port 212 nsew signal input
rlabel metal2 s 112074 167200 112130 168000 6 la_input[36]
port 213 nsew signal input
rlabel metal2 s 115110 167200 115166 168000 6 la_input[37]
port 214 nsew signal input
rlabel metal2 s 118146 167200 118202 168000 6 la_input[38]
port 215 nsew signal input
rlabel metal2 s 121182 167200 121238 168000 6 la_input[39]
port 216 nsew signal input
rlabel metal2 s 12438 167200 12494 168000 6 la_input[3]
port 217 nsew signal input
rlabel metal2 s 124126 167200 124182 168000 6 la_input[40]
port 218 nsew signal input
rlabel metal2 s 127162 167200 127218 168000 6 la_input[41]
port 219 nsew signal input
rlabel metal2 s 130198 167200 130254 168000 6 la_input[42]
port 220 nsew signal input
rlabel metal2 s 133234 167200 133290 168000 6 la_input[43]
port 221 nsew signal input
rlabel metal2 s 136270 167200 136326 168000 6 la_input[44]
port 222 nsew signal input
rlabel metal2 s 139214 167200 139270 168000 6 la_input[45]
port 223 nsew signal input
rlabel metal2 s 142250 167200 142306 168000 6 la_input[46]
port 224 nsew signal input
rlabel metal2 s 145286 167200 145342 168000 6 la_input[47]
port 225 nsew signal input
rlabel metal2 s 148322 167200 148378 168000 6 la_input[48]
port 226 nsew signal input
rlabel metal2 s 151358 167200 151414 168000 6 la_input[49]
port 227 nsew signal input
rlabel metal2 s 15474 167200 15530 168000 6 la_input[4]
port 228 nsew signal input
rlabel metal2 s 154394 167200 154450 168000 6 la_input[50]
port 229 nsew signal input
rlabel metal2 s 157338 167200 157394 168000 6 la_input[51]
port 230 nsew signal input
rlabel metal2 s 160374 167200 160430 168000 6 la_input[52]
port 231 nsew signal input
rlabel metal2 s 163410 167200 163466 168000 6 la_input[53]
port 232 nsew signal input
rlabel metal2 s 166446 167200 166502 168000 6 la_input[54]
port 233 nsew signal input
rlabel metal2 s 169482 167200 169538 168000 6 la_input[55]
port 234 nsew signal input
rlabel metal2 s 172518 167200 172574 168000 6 la_input[56]
port 235 nsew signal input
rlabel metal2 s 175462 167200 175518 168000 6 la_input[57]
port 236 nsew signal input
rlabel metal2 s 178498 167200 178554 168000 6 la_input[58]
port 237 nsew signal input
rlabel metal2 s 181534 167200 181590 168000 6 la_input[59]
port 238 nsew signal input
rlabel metal2 s 18418 167200 18474 168000 6 la_input[5]
port 239 nsew signal input
rlabel metal2 s 184570 167200 184626 168000 6 la_input[60]
port 240 nsew signal input
rlabel metal2 s 187606 167200 187662 168000 6 la_input[61]
port 241 nsew signal input
rlabel metal2 s 190642 167200 190698 168000 6 la_input[62]
port 242 nsew signal input
rlabel metal2 s 193586 167200 193642 168000 6 la_input[63]
port 243 nsew signal input
rlabel metal2 s 196622 167200 196678 168000 6 la_input[64]
port 244 nsew signal input
rlabel metal2 s 199658 167200 199714 168000 6 la_input[65]
port 245 nsew signal input
rlabel metal2 s 202694 167200 202750 168000 6 la_input[66]
port 246 nsew signal input
rlabel metal2 s 205730 167200 205786 168000 6 la_input[67]
port 247 nsew signal input
rlabel metal2 s 208674 167200 208730 168000 6 la_input[68]
port 248 nsew signal input
rlabel metal2 s 211710 167200 211766 168000 6 la_input[69]
port 249 nsew signal input
rlabel metal2 s 21454 167200 21510 168000 6 la_input[6]
port 250 nsew signal input
rlabel metal2 s 214746 167200 214802 168000 6 la_input[70]
port 251 nsew signal input
rlabel metal2 s 217782 167200 217838 168000 6 la_input[71]
port 252 nsew signal input
rlabel metal2 s 220818 167200 220874 168000 6 la_input[72]
port 253 nsew signal input
rlabel metal2 s 223854 167200 223910 168000 6 la_input[73]
port 254 nsew signal input
rlabel metal2 s 226798 167200 226854 168000 6 la_input[74]
port 255 nsew signal input
rlabel metal2 s 229834 167200 229890 168000 6 la_input[75]
port 256 nsew signal input
rlabel metal2 s 232870 167200 232926 168000 6 la_input[76]
port 257 nsew signal input
rlabel metal2 s 235906 167200 235962 168000 6 la_input[77]
port 258 nsew signal input
rlabel metal2 s 238942 167200 238998 168000 6 la_input[78]
port 259 nsew signal input
rlabel metal2 s 241978 167200 242034 168000 6 la_input[79]
port 260 nsew signal input
rlabel metal2 s 24490 167200 24546 168000 6 la_input[7]
port 261 nsew signal input
rlabel metal2 s 244922 167200 244978 168000 6 la_input[80]
port 262 nsew signal input
rlabel metal2 s 247958 167200 248014 168000 6 la_input[81]
port 263 nsew signal input
rlabel metal2 s 250994 167200 251050 168000 6 la_input[82]
port 264 nsew signal input
rlabel metal2 s 254030 167200 254086 168000 6 la_input[83]
port 265 nsew signal input
rlabel metal2 s 257066 167200 257122 168000 6 la_input[84]
port 266 nsew signal input
rlabel metal2 s 260010 167200 260066 168000 6 la_input[85]
port 267 nsew signal input
rlabel metal2 s 263046 167200 263102 168000 6 la_input[86]
port 268 nsew signal input
rlabel metal2 s 266082 167200 266138 168000 6 la_input[87]
port 269 nsew signal input
rlabel metal2 s 269118 167200 269174 168000 6 la_input[88]
port 270 nsew signal input
rlabel metal2 s 272154 167200 272210 168000 6 la_input[89]
port 271 nsew signal input
rlabel metal2 s 27526 167200 27582 168000 6 la_input[8]
port 272 nsew signal input
rlabel metal2 s 275190 167200 275246 168000 6 la_input[90]
port 273 nsew signal input
rlabel metal2 s 278134 167200 278190 168000 6 la_input[91]
port 274 nsew signal input
rlabel metal2 s 281170 167200 281226 168000 6 la_input[92]
port 275 nsew signal input
rlabel metal2 s 284206 167200 284262 168000 6 la_input[93]
port 276 nsew signal input
rlabel metal2 s 287242 167200 287298 168000 6 la_input[94]
port 277 nsew signal input
rlabel metal2 s 290278 167200 290334 168000 6 la_input[95]
port 278 nsew signal input
rlabel metal2 s 293314 167200 293370 168000 6 la_input[96]
port 279 nsew signal input
rlabel metal2 s 296258 167200 296314 168000 6 la_input[97]
port 280 nsew signal input
rlabel metal2 s 299294 167200 299350 168000 6 la_input[98]
port 281 nsew signal input
rlabel metal2 s 302330 167200 302386 168000 6 la_input[99]
port 282 nsew signal input
rlabel metal2 s 30562 167200 30618 168000 6 la_input[9]
port 283 nsew signal input
rlabel metal2 s 4158 167200 4214 168000 6 la_oenb[0]
port 284 nsew signal output
rlabel metal2 s 306102 167200 306158 168000 6 la_oenb[100]
port 285 nsew signal output
rlabel metal2 s 309138 167200 309194 168000 6 la_oenb[101]
port 286 nsew signal output
rlabel metal2 s 312174 167200 312230 168000 6 la_oenb[102]
port 287 nsew signal output
rlabel metal2 s 315210 167200 315266 168000 6 la_oenb[103]
port 288 nsew signal output
rlabel metal2 s 318154 167200 318210 168000 6 la_oenb[104]
port 289 nsew signal output
rlabel metal2 s 321190 167200 321246 168000 6 la_oenb[105]
port 290 nsew signal output
rlabel metal2 s 324226 167200 324282 168000 6 la_oenb[106]
port 291 nsew signal output
rlabel metal2 s 327262 167200 327318 168000 6 la_oenb[107]
port 292 nsew signal output
rlabel metal2 s 330298 167200 330354 168000 6 la_oenb[108]
port 293 nsew signal output
rlabel metal2 s 333334 167200 333390 168000 6 la_oenb[109]
port 294 nsew signal output
rlabel metal2 s 34334 167200 34390 168000 6 la_oenb[10]
port 295 nsew signal output
rlabel metal2 s 336278 167200 336334 168000 6 la_oenb[110]
port 296 nsew signal output
rlabel metal2 s 339314 167200 339370 168000 6 la_oenb[111]
port 297 nsew signal output
rlabel metal2 s 342350 167200 342406 168000 6 la_oenb[112]
port 298 nsew signal output
rlabel metal2 s 345386 167200 345442 168000 6 la_oenb[113]
port 299 nsew signal output
rlabel metal2 s 348422 167200 348478 168000 6 la_oenb[114]
port 300 nsew signal output
rlabel metal2 s 351366 167200 351422 168000 6 la_oenb[115]
port 301 nsew signal output
rlabel metal2 s 354402 167200 354458 168000 6 la_oenb[116]
port 302 nsew signal output
rlabel metal2 s 357438 167200 357494 168000 6 la_oenb[117]
port 303 nsew signal output
rlabel metal2 s 360474 167200 360530 168000 6 la_oenb[118]
port 304 nsew signal output
rlabel metal2 s 363510 167200 363566 168000 6 la_oenb[119]
port 305 nsew signal output
rlabel metal2 s 37370 167200 37426 168000 6 la_oenb[11]
port 306 nsew signal output
rlabel metal2 s 366546 167200 366602 168000 6 la_oenb[120]
port 307 nsew signal output
rlabel metal2 s 369490 167200 369546 168000 6 la_oenb[121]
port 308 nsew signal output
rlabel metal2 s 372526 167200 372582 168000 6 la_oenb[122]
port 309 nsew signal output
rlabel metal2 s 375562 167200 375618 168000 6 la_oenb[123]
port 310 nsew signal output
rlabel metal2 s 378598 167200 378654 168000 6 la_oenb[124]
port 311 nsew signal output
rlabel metal2 s 381634 167200 381690 168000 6 la_oenb[125]
port 312 nsew signal output
rlabel metal2 s 384670 167200 384726 168000 6 la_oenb[126]
port 313 nsew signal output
rlabel metal2 s 387614 167200 387670 168000 6 la_oenb[127]
port 314 nsew signal output
rlabel metal2 s 40314 167200 40370 168000 6 la_oenb[12]
port 315 nsew signal output
rlabel metal2 s 43350 167200 43406 168000 6 la_oenb[13]
port 316 nsew signal output
rlabel metal2 s 46386 167200 46442 168000 6 la_oenb[14]
port 317 nsew signal output
rlabel metal2 s 49422 167200 49478 168000 6 la_oenb[15]
port 318 nsew signal output
rlabel metal2 s 52458 167200 52514 168000 6 la_oenb[16]
port 319 nsew signal output
rlabel metal2 s 55494 167200 55550 168000 6 la_oenb[17]
port 320 nsew signal output
rlabel metal2 s 58438 167200 58494 168000 6 la_oenb[18]
port 321 nsew signal output
rlabel metal2 s 61474 167200 61530 168000 6 la_oenb[19]
port 322 nsew signal output
rlabel metal2 s 7102 167200 7158 168000 6 la_oenb[1]
port 323 nsew signal output
rlabel metal2 s 64510 167200 64566 168000 6 la_oenb[20]
port 324 nsew signal output
rlabel metal2 s 67546 167200 67602 168000 6 la_oenb[21]
port 325 nsew signal output
rlabel metal2 s 70582 167200 70638 168000 6 la_oenb[22]
port 326 nsew signal output
rlabel metal2 s 73618 167200 73674 168000 6 la_oenb[23]
port 327 nsew signal output
rlabel metal2 s 76562 167200 76618 168000 6 la_oenb[24]
port 328 nsew signal output
rlabel metal2 s 79598 167200 79654 168000 6 la_oenb[25]
port 329 nsew signal output
rlabel metal2 s 82634 167200 82690 168000 6 la_oenb[26]
port 330 nsew signal output
rlabel metal2 s 85670 167200 85726 168000 6 la_oenb[27]
port 331 nsew signal output
rlabel metal2 s 88706 167200 88762 168000 6 la_oenb[28]
port 332 nsew signal output
rlabel metal2 s 91650 167200 91706 168000 6 la_oenb[29]
port 333 nsew signal output
rlabel metal2 s 10138 167200 10194 168000 6 la_oenb[2]
port 334 nsew signal output
rlabel metal2 s 94686 167200 94742 168000 6 la_oenb[30]
port 335 nsew signal output
rlabel metal2 s 97722 167200 97778 168000 6 la_oenb[31]
port 336 nsew signal output
rlabel metal2 s 100758 167200 100814 168000 6 la_oenb[32]
port 337 nsew signal output
rlabel metal2 s 103794 167200 103850 168000 6 la_oenb[33]
port 338 nsew signal output
rlabel metal2 s 106830 167200 106886 168000 6 la_oenb[34]
port 339 nsew signal output
rlabel metal2 s 109774 167200 109830 168000 6 la_oenb[35]
port 340 nsew signal output
rlabel metal2 s 112810 167200 112866 168000 6 la_oenb[36]
port 341 nsew signal output
rlabel metal2 s 115846 167200 115902 168000 6 la_oenb[37]
port 342 nsew signal output
rlabel metal2 s 118882 167200 118938 168000 6 la_oenb[38]
port 343 nsew signal output
rlabel metal2 s 121918 167200 121974 168000 6 la_oenb[39]
port 344 nsew signal output
rlabel metal2 s 13174 167200 13230 168000 6 la_oenb[3]
port 345 nsew signal output
rlabel metal2 s 124954 167200 125010 168000 6 la_oenb[40]
port 346 nsew signal output
rlabel metal2 s 127898 167200 127954 168000 6 la_oenb[41]
port 347 nsew signal output
rlabel metal2 s 130934 167200 130990 168000 6 la_oenb[42]
port 348 nsew signal output
rlabel metal2 s 133970 167200 134026 168000 6 la_oenb[43]
port 349 nsew signal output
rlabel metal2 s 137006 167200 137062 168000 6 la_oenb[44]
port 350 nsew signal output
rlabel metal2 s 140042 167200 140098 168000 6 la_oenb[45]
port 351 nsew signal output
rlabel metal2 s 143078 167200 143134 168000 6 la_oenb[46]
port 352 nsew signal output
rlabel metal2 s 146022 167200 146078 168000 6 la_oenb[47]
port 353 nsew signal output
rlabel metal2 s 149058 167200 149114 168000 6 la_oenb[48]
port 354 nsew signal output
rlabel metal2 s 152094 167200 152150 168000 6 la_oenb[49]
port 355 nsew signal output
rlabel metal2 s 16210 167200 16266 168000 6 la_oenb[4]
port 356 nsew signal output
rlabel metal2 s 155130 167200 155186 168000 6 la_oenb[50]
port 357 nsew signal output
rlabel metal2 s 158166 167200 158222 168000 6 la_oenb[51]
port 358 nsew signal output
rlabel metal2 s 161110 167200 161166 168000 6 la_oenb[52]
port 359 nsew signal output
rlabel metal2 s 164146 167200 164202 168000 6 la_oenb[53]
port 360 nsew signal output
rlabel metal2 s 167182 167200 167238 168000 6 la_oenb[54]
port 361 nsew signal output
rlabel metal2 s 170218 167200 170274 168000 6 la_oenb[55]
port 362 nsew signal output
rlabel metal2 s 173254 167200 173310 168000 6 la_oenb[56]
port 363 nsew signal output
rlabel metal2 s 176290 167200 176346 168000 6 la_oenb[57]
port 364 nsew signal output
rlabel metal2 s 179234 167200 179290 168000 6 la_oenb[58]
port 365 nsew signal output
rlabel metal2 s 182270 167200 182326 168000 6 la_oenb[59]
port 366 nsew signal output
rlabel metal2 s 19246 167200 19302 168000 6 la_oenb[5]
port 367 nsew signal output
rlabel metal2 s 185306 167200 185362 168000 6 la_oenb[60]
port 368 nsew signal output
rlabel metal2 s 188342 167200 188398 168000 6 la_oenb[61]
port 369 nsew signal output
rlabel metal2 s 191378 167200 191434 168000 6 la_oenb[62]
port 370 nsew signal output
rlabel metal2 s 194414 167200 194470 168000 6 la_oenb[63]
port 371 nsew signal output
rlabel metal2 s 197358 167200 197414 168000 6 la_oenb[64]
port 372 nsew signal output
rlabel metal2 s 200394 167200 200450 168000 6 la_oenb[65]
port 373 nsew signal output
rlabel metal2 s 203430 167200 203486 168000 6 la_oenb[66]
port 374 nsew signal output
rlabel metal2 s 206466 167200 206522 168000 6 la_oenb[67]
port 375 nsew signal output
rlabel metal2 s 209502 167200 209558 168000 6 la_oenb[68]
port 376 nsew signal output
rlabel metal2 s 212446 167200 212502 168000 6 la_oenb[69]
port 377 nsew signal output
rlabel metal2 s 22190 167200 22246 168000 6 la_oenb[6]
port 378 nsew signal output
rlabel metal2 s 215482 167200 215538 168000 6 la_oenb[70]
port 379 nsew signal output
rlabel metal2 s 218518 167200 218574 168000 6 la_oenb[71]
port 380 nsew signal output
rlabel metal2 s 221554 167200 221610 168000 6 la_oenb[72]
port 381 nsew signal output
rlabel metal2 s 224590 167200 224646 168000 6 la_oenb[73]
port 382 nsew signal output
rlabel metal2 s 227626 167200 227682 168000 6 la_oenb[74]
port 383 nsew signal output
rlabel metal2 s 230570 167200 230626 168000 6 la_oenb[75]
port 384 nsew signal output
rlabel metal2 s 233606 167200 233662 168000 6 la_oenb[76]
port 385 nsew signal output
rlabel metal2 s 236642 167200 236698 168000 6 la_oenb[77]
port 386 nsew signal output
rlabel metal2 s 239678 167200 239734 168000 6 la_oenb[78]
port 387 nsew signal output
rlabel metal2 s 242714 167200 242770 168000 6 la_oenb[79]
port 388 nsew signal output
rlabel metal2 s 25226 167200 25282 168000 6 la_oenb[7]
port 389 nsew signal output
rlabel metal2 s 245750 167200 245806 168000 6 la_oenb[80]
port 390 nsew signal output
rlabel metal2 s 248694 167200 248750 168000 6 la_oenb[81]
port 391 nsew signal output
rlabel metal2 s 251730 167200 251786 168000 6 la_oenb[82]
port 392 nsew signal output
rlabel metal2 s 254766 167200 254822 168000 6 la_oenb[83]
port 393 nsew signal output
rlabel metal2 s 257802 167200 257858 168000 6 la_oenb[84]
port 394 nsew signal output
rlabel metal2 s 260838 167200 260894 168000 6 la_oenb[85]
port 395 nsew signal output
rlabel metal2 s 263874 167200 263930 168000 6 la_oenb[86]
port 396 nsew signal output
rlabel metal2 s 266818 167200 266874 168000 6 la_oenb[87]
port 397 nsew signal output
rlabel metal2 s 269854 167200 269910 168000 6 la_oenb[88]
port 398 nsew signal output
rlabel metal2 s 272890 167200 272946 168000 6 la_oenb[89]
port 399 nsew signal output
rlabel metal2 s 28262 167200 28318 168000 6 la_oenb[8]
port 400 nsew signal output
rlabel metal2 s 275926 167200 275982 168000 6 la_oenb[90]
port 401 nsew signal output
rlabel metal2 s 278962 167200 279018 168000 6 la_oenb[91]
port 402 nsew signal output
rlabel metal2 s 281906 167200 281962 168000 6 la_oenb[92]
port 403 nsew signal output
rlabel metal2 s 284942 167200 284998 168000 6 la_oenb[93]
port 404 nsew signal output
rlabel metal2 s 287978 167200 288034 168000 6 la_oenb[94]
port 405 nsew signal output
rlabel metal2 s 291014 167200 291070 168000 6 la_oenb[95]
port 406 nsew signal output
rlabel metal2 s 294050 167200 294106 168000 6 la_oenb[96]
port 407 nsew signal output
rlabel metal2 s 297086 167200 297142 168000 6 la_oenb[97]
port 408 nsew signal output
rlabel metal2 s 300030 167200 300086 168000 6 la_oenb[98]
port 409 nsew signal output
rlabel metal2 s 303066 167200 303122 168000 6 la_oenb[99]
port 410 nsew signal output
rlabel metal2 s 31298 167200 31354 168000 6 la_oenb[9]
port 411 nsew signal output
rlabel metal2 s 4894 167200 4950 168000 6 la_output[0]
port 412 nsew signal output
rlabel metal2 s 306838 167200 306894 168000 6 la_output[100]
port 413 nsew signal output
rlabel metal2 s 309874 167200 309930 168000 6 la_output[101]
port 414 nsew signal output
rlabel metal2 s 312910 167200 312966 168000 6 la_output[102]
port 415 nsew signal output
rlabel metal2 s 315946 167200 316002 168000 6 la_output[103]
port 416 nsew signal output
rlabel metal2 s 318982 167200 319038 168000 6 la_output[104]
port 417 nsew signal output
rlabel metal2 s 321926 167200 321982 168000 6 la_output[105]
port 418 nsew signal output
rlabel metal2 s 324962 167200 325018 168000 6 la_output[106]
port 419 nsew signal output
rlabel metal2 s 327998 167200 328054 168000 6 la_output[107]
port 420 nsew signal output
rlabel metal2 s 331034 167200 331090 168000 6 la_output[108]
port 421 nsew signal output
rlabel metal2 s 334070 167200 334126 168000 6 la_output[109]
port 422 nsew signal output
rlabel metal2 s 35070 167200 35126 168000 6 la_output[10]
port 423 nsew signal output
rlabel metal2 s 337106 167200 337162 168000 6 la_output[110]
port 424 nsew signal output
rlabel metal2 s 340050 167200 340106 168000 6 la_output[111]
port 425 nsew signal output
rlabel metal2 s 343086 167200 343142 168000 6 la_output[112]
port 426 nsew signal output
rlabel metal2 s 346122 167200 346178 168000 6 la_output[113]
port 427 nsew signal output
rlabel metal2 s 349158 167200 349214 168000 6 la_output[114]
port 428 nsew signal output
rlabel metal2 s 352194 167200 352250 168000 6 la_output[115]
port 429 nsew signal output
rlabel metal2 s 355138 167200 355194 168000 6 la_output[116]
port 430 nsew signal output
rlabel metal2 s 358174 167200 358230 168000 6 la_output[117]
port 431 nsew signal output
rlabel metal2 s 361210 167200 361266 168000 6 la_output[118]
port 432 nsew signal output
rlabel metal2 s 364246 167200 364302 168000 6 la_output[119]
port 433 nsew signal output
rlabel metal2 s 38106 167200 38162 168000 6 la_output[11]
port 434 nsew signal output
rlabel metal2 s 367282 167200 367338 168000 6 la_output[120]
port 435 nsew signal output
rlabel metal2 s 370318 167200 370374 168000 6 la_output[121]
port 436 nsew signal output
rlabel metal2 s 373262 167200 373318 168000 6 la_output[122]
port 437 nsew signal output
rlabel metal2 s 376298 167200 376354 168000 6 la_output[123]
port 438 nsew signal output
rlabel metal2 s 379334 167200 379390 168000 6 la_output[124]
port 439 nsew signal output
rlabel metal2 s 382370 167200 382426 168000 6 la_output[125]
port 440 nsew signal output
rlabel metal2 s 385406 167200 385462 168000 6 la_output[126]
port 441 nsew signal output
rlabel metal2 s 388442 167200 388498 168000 6 la_output[127]
port 442 nsew signal output
rlabel metal2 s 41142 167200 41198 168000 6 la_output[12]
port 443 nsew signal output
rlabel metal2 s 44086 167200 44142 168000 6 la_output[13]
port 444 nsew signal output
rlabel metal2 s 47122 167200 47178 168000 6 la_output[14]
port 445 nsew signal output
rlabel metal2 s 50158 167200 50214 168000 6 la_output[15]
port 446 nsew signal output
rlabel metal2 s 53194 167200 53250 168000 6 la_output[16]
port 447 nsew signal output
rlabel metal2 s 56230 167200 56286 168000 6 la_output[17]
port 448 nsew signal output
rlabel metal2 s 59266 167200 59322 168000 6 la_output[18]
port 449 nsew signal output
rlabel metal2 s 62210 167200 62266 168000 6 la_output[19]
port 450 nsew signal output
rlabel metal2 s 7930 167200 7986 168000 6 la_output[1]
port 451 nsew signal output
rlabel metal2 s 65246 167200 65302 168000 6 la_output[20]
port 452 nsew signal output
rlabel metal2 s 68282 167200 68338 168000 6 la_output[21]
port 453 nsew signal output
rlabel metal2 s 71318 167200 71374 168000 6 la_output[22]
port 454 nsew signal output
rlabel metal2 s 74354 167200 74410 168000 6 la_output[23]
port 455 nsew signal output
rlabel metal2 s 77390 167200 77446 168000 6 la_output[24]
port 456 nsew signal output
rlabel metal2 s 80334 167200 80390 168000 6 la_output[25]
port 457 nsew signal output
rlabel metal2 s 83370 167200 83426 168000 6 la_output[26]
port 458 nsew signal output
rlabel metal2 s 86406 167200 86462 168000 6 la_output[27]
port 459 nsew signal output
rlabel metal2 s 89442 167200 89498 168000 6 la_output[28]
port 460 nsew signal output
rlabel metal2 s 92478 167200 92534 168000 6 la_output[29]
port 461 nsew signal output
rlabel metal2 s 10874 167200 10930 168000 6 la_output[2]
port 462 nsew signal output
rlabel metal2 s 95514 167200 95570 168000 6 la_output[30]
port 463 nsew signal output
rlabel metal2 s 98458 167200 98514 168000 6 la_output[31]
port 464 nsew signal output
rlabel metal2 s 101494 167200 101550 168000 6 la_output[32]
port 465 nsew signal output
rlabel metal2 s 104530 167200 104586 168000 6 la_output[33]
port 466 nsew signal output
rlabel metal2 s 107566 167200 107622 168000 6 la_output[34]
port 467 nsew signal output
rlabel metal2 s 110602 167200 110658 168000 6 la_output[35]
port 468 nsew signal output
rlabel metal2 s 113546 167200 113602 168000 6 la_output[36]
port 469 nsew signal output
rlabel metal2 s 116582 167200 116638 168000 6 la_output[37]
port 470 nsew signal output
rlabel metal2 s 119618 167200 119674 168000 6 la_output[38]
port 471 nsew signal output
rlabel metal2 s 122654 167200 122710 168000 6 la_output[39]
port 472 nsew signal output
rlabel metal2 s 13910 167200 13966 168000 6 la_output[3]
port 473 nsew signal output
rlabel metal2 s 125690 167200 125746 168000 6 la_output[40]
port 474 nsew signal output
rlabel metal2 s 128726 167200 128782 168000 6 la_output[41]
port 475 nsew signal output
rlabel metal2 s 131670 167200 131726 168000 6 la_output[42]
port 476 nsew signal output
rlabel metal2 s 134706 167200 134762 168000 6 la_output[43]
port 477 nsew signal output
rlabel metal2 s 137742 167200 137798 168000 6 la_output[44]
port 478 nsew signal output
rlabel metal2 s 140778 167200 140834 168000 6 la_output[45]
port 479 nsew signal output
rlabel metal2 s 143814 167200 143870 168000 6 la_output[46]
port 480 nsew signal output
rlabel metal2 s 146850 167200 146906 168000 6 la_output[47]
port 481 nsew signal output
rlabel metal2 s 149794 167200 149850 168000 6 la_output[48]
port 482 nsew signal output
rlabel metal2 s 152830 167200 152886 168000 6 la_output[49]
port 483 nsew signal output
rlabel metal2 s 16946 167200 17002 168000 6 la_output[4]
port 484 nsew signal output
rlabel metal2 s 155866 167200 155922 168000 6 la_output[50]
port 485 nsew signal output
rlabel metal2 s 158902 167200 158958 168000 6 la_output[51]
port 486 nsew signal output
rlabel metal2 s 161938 167200 161994 168000 6 la_output[52]
port 487 nsew signal output
rlabel metal2 s 164882 167200 164938 168000 6 la_output[53]
port 488 nsew signal output
rlabel metal2 s 167918 167200 167974 168000 6 la_output[54]
port 489 nsew signal output
rlabel metal2 s 170954 167200 171010 168000 6 la_output[55]
port 490 nsew signal output
rlabel metal2 s 173990 167200 174046 168000 6 la_output[56]
port 491 nsew signal output
rlabel metal2 s 177026 167200 177082 168000 6 la_output[57]
port 492 nsew signal output
rlabel metal2 s 180062 167200 180118 168000 6 la_output[58]
port 493 nsew signal output
rlabel metal2 s 183006 167200 183062 168000 6 la_output[59]
port 494 nsew signal output
rlabel metal2 s 19982 167200 20038 168000 6 la_output[5]
port 495 nsew signal output
rlabel metal2 s 186042 167200 186098 168000 6 la_output[60]
port 496 nsew signal output
rlabel metal2 s 189078 167200 189134 168000 6 la_output[61]
port 497 nsew signal output
rlabel metal2 s 192114 167200 192170 168000 6 la_output[62]
port 498 nsew signal output
rlabel metal2 s 195150 167200 195206 168000 6 la_output[63]
port 499 nsew signal output
rlabel metal2 s 198186 167200 198242 168000 6 la_output[64]
port 500 nsew signal output
rlabel metal2 s 201130 167200 201186 168000 6 la_output[65]
port 501 nsew signal output
rlabel metal2 s 204166 167200 204222 168000 6 la_output[66]
port 502 nsew signal output
rlabel metal2 s 207202 167200 207258 168000 6 la_output[67]
port 503 nsew signal output
rlabel metal2 s 210238 167200 210294 168000 6 la_output[68]
port 504 nsew signal output
rlabel metal2 s 213274 167200 213330 168000 6 la_output[69]
port 505 nsew signal output
rlabel metal2 s 23018 167200 23074 168000 6 la_output[6]
port 506 nsew signal output
rlabel metal2 s 216310 167200 216366 168000 6 la_output[70]
port 507 nsew signal output
rlabel metal2 s 219254 167200 219310 168000 6 la_output[71]
port 508 nsew signal output
rlabel metal2 s 222290 167200 222346 168000 6 la_output[72]
port 509 nsew signal output
rlabel metal2 s 225326 167200 225382 168000 6 la_output[73]
port 510 nsew signal output
rlabel metal2 s 228362 167200 228418 168000 6 la_output[74]
port 511 nsew signal output
rlabel metal2 s 231398 167200 231454 168000 6 la_output[75]
port 512 nsew signal output
rlabel metal2 s 234342 167200 234398 168000 6 la_output[76]
port 513 nsew signal output
rlabel metal2 s 237378 167200 237434 168000 6 la_output[77]
port 514 nsew signal output
rlabel metal2 s 240414 167200 240470 168000 6 la_output[78]
port 515 nsew signal output
rlabel metal2 s 243450 167200 243506 168000 6 la_output[79]
port 516 nsew signal output
rlabel metal2 s 26054 167200 26110 168000 6 la_output[7]
port 517 nsew signal output
rlabel metal2 s 246486 167200 246542 168000 6 la_output[80]
port 518 nsew signal output
rlabel metal2 s 249522 167200 249578 168000 6 la_output[81]
port 519 nsew signal output
rlabel metal2 s 252466 167200 252522 168000 6 la_output[82]
port 520 nsew signal output
rlabel metal2 s 255502 167200 255558 168000 6 la_output[83]
port 521 nsew signal output
rlabel metal2 s 258538 167200 258594 168000 6 la_output[84]
port 522 nsew signal output
rlabel metal2 s 261574 167200 261630 168000 6 la_output[85]
port 523 nsew signal output
rlabel metal2 s 264610 167200 264666 168000 6 la_output[86]
port 524 nsew signal output
rlabel metal2 s 267646 167200 267702 168000 6 la_output[87]
port 525 nsew signal output
rlabel metal2 s 270590 167200 270646 168000 6 la_output[88]
port 526 nsew signal output
rlabel metal2 s 273626 167200 273682 168000 6 la_output[89]
port 527 nsew signal output
rlabel metal2 s 28998 167200 29054 168000 6 la_output[8]
port 528 nsew signal output
rlabel metal2 s 276662 167200 276718 168000 6 la_output[90]
port 529 nsew signal output
rlabel metal2 s 279698 167200 279754 168000 6 la_output[91]
port 530 nsew signal output
rlabel metal2 s 282734 167200 282790 168000 6 la_output[92]
port 531 nsew signal output
rlabel metal2 s 285770 167200 285826 168000 6 la_output[93]
port 532 nsew signal output
rlabel metal2 s 288714 167200 288770 168000 6 la_output[94]
port 533 nsew signal output
rlabel metal2 s 291750 167200 291806 168000 6 la_output[95]
port 534 nsew signal output
rlabel metal2 s 294786 167200 294842 168000 6 la_output[96]
port 535 nsew signal output
rlabel metal2 s 297822 167200 297878 168000 6 la_output[97]
port 536 nsew signal output
rlabel metal2 s 300858 167200 300914 168000 6 la_output[98]
port 537 nsew signal output
rlabel metal2 s 303802 167200 303858 168000 6 la_output[99]
port 538 nsew signal output
rlabel metal2 s 32034 167200 32090 168000 6 la_output[9]
port 539 nsew signal output
rlabel metal3 s 449200 960 450000 1080 6 mask_rev[0]
port 540 nsew signal input
rlabel metal3 s 449200 20000 450000 20120 6 mask_rev[10]
port 541 nsew signal input
rlabel metal3 s 449200 21904 450000 22024 6 mask_rev[11]
port 542 nsew signal input
rlabel metal3 s 449200 23808 450000 23928 6 mask_rev[12]
port 543 nsew signal input
rlabel metal3 s 449200 25712 450000 25832 6 mask_rev[13]
port 544 nsew signal input
rlabel metal3 s 449200 27616 450000 27736 6 mask_rev[14]
port 545 nsew signal input
rlabel metal3 s 449200 29520 450000 29640 6 mask_rev[15]
port 546 nsew signal input
rlabel metal3 s 449200 31424 450000 31544 6 mask_rev[16]
port 547 nsew signal input
rlabel metal3 s 449200 33328 450000 33448 6 mask_rev[17]
port 548 nsew signal input
rlabel metal3 s 449200 35232 450000 35352 6 mask_rev[18]
port 549 nsew signal input
rlabel metal3 s 449200 37136 450000 37256 6 mask_rev[19]
port 550 nsew signal input
rlabel metal3 s 449200 2864 450000 2984 6 mask_rev[1]
port 551 nsew signal input
rlabel metal3 s 449200 39040 450000 39160 6 mask_rev[20]
port 552 nsew signal input
rlabel metal3 s 449200 40944 450000 41064 6 mask_rev[21]
port 553 nsew signal input
rlabel metal3 s 449200 42848 450000 42968 6 mask_rev[22]
port 554 nsew signal input
rlabel metal3 s 449200 44752 450000 44872 6 mask_rev[23]
port 555 nsew signal input
rlabel metal3 s 449200 46656 450000 46776 6 mask_rev[24]
port 556 nsew signal input
rlabel metal3 s 449200 48560 450000 48680 6 mask_rev[25]
port 557 nsew signal input
rlabel metal3 s 449200 50464 450000 50584 6 mask_rev[26]
port 558 nsew signal input
rlabel metal3 s 449200 52368 450000 52488 6 mask_rev[27]
port 559 nsew signal input
rlabel metal3 s 449200 54272 450000 54392 6 mask_rev[28]
port 560 nsew signal input
rlabel metal3 s 449200 56176 450000 56296 6 mask_rev[29]
port 561 nsew signal input
rlabel metal3 s 449200 4768 450000 4888 6 mask_rev[2]
port 562 nsew signal input
rlabel metal3 s 449200 58216 450000 58336 6 mask_rev[30]
port 563 nsew signal input
rlabel metal3 s 449200 60120 450000 60240 6 mask_rev[31]
port 564 nsew signal input
rlabel metal3 s 449200 6672 450000 6792 6 mask_rev[3]
port 565 nsew signal input
rlabel metal3 s 449200 8576 450000 8696 6 mask_rev[4]
port 566 nsew signal input
rlabel metal3 s 449200 10480 450000 10600 6 mask_rev[5]
port 567 nsew signal input
rlabel metal3 s 449200 12384 450000 12504 6 mask_rev[6]
port 568 nsew signal input
rlabel metal3 s 449200 14288 450000 14408 6 mask_rev[7]
port 569 nsew signal input
rlabel metal3 s 449200 16192 450000 16312 6 mask_rev[8]
port 570 nsew signal input
rlabel metal3 s 449200 18096 450000 18216 6 mask_rev[9]
port 571 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 mgmt_addr[0]
port 572 nsew signal output
rlabel metal3 s 0 61072 800 61192 6 mgmt_addr[1]
port 573 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 mgmt_addr[2]
port 574 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 mgmt_addr[3]
port 575 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 mgmt_addr[4]
port 576 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 mgmt_addr[5]
port 577 nsew signal output
rlabel metal3 s 0 64880 800 65000 6 mgmt_addr[6]
port 578 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 mgmt_addr[7]
port 579 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 mgmt_addr_ro[0]
port 580 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 mgmt_addr_ro[1]
port 581 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 mgmt_addr_ro[2]
port 582 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 mgmt_addr_ro[3]
port 583 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 mgmt_addr_ro[4]
port 584 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 mgmt_addr_ro[5]
port 585 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 mgmt_addr_ro[6]
port 586 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 mgmt_addr_ro[7]
port 587 nsew signal output
rlabel metal3 s 0 280 800 400 6 mgmt_ena[0]
port 588 nsew signal output
rlabel metal3 s 0 90720 800 90840 6 mgmt_ena[1]
port 589 nsew signal output
rlabel metal3 s 0 960 800 1080 6 mgmt_ena_ro
port 590 nsew signal output
rlabel metal3 s 449200 77256 450000 77376 6 mgmt_in_data[0]
port 591 nsew signal input
rlabel metal3 s 449200 115472 450000 115592 6 mgmt_in_data[10]
port 592 nsew signal input
rlabel metal3 s 449200 119280 450000 119400 6 mgmt_in_data[11]
port 593 nsew signal input
rlabel metal3 s 449200 123088 450000 123208 6 mgmt_in_data[12]
port 594 nsew signal input
rlabel metal3 s 449200 126896 450000 127016 6 mgmt_in_data[13]
port 595 nsew signal input
rlabel metal3 s 449200 130704 450000 130824 6 mgmt_in_data[14]
port 596 nsew signal input
rlabel metal3 s 449200 134512 450000 134632 6 mgmt_in_data[15]
port 597 nsew signal input
rlabel metal3 s 449200 138320 450000 138440 6 mgmt_in_data[16]
port 598 nsew signal input
rlabel metal3 s 449200 142128 450000 142248 6 mgmt_in_data[17]
port 599 nsew signal input
rlabel metal3 s 449200 145936 450000 146056 6 mgmt_in_data[18]
port 600 nsew signal input
rlabel metal3 s 449200 149744 450000 149864 6 mgmt_in_data[19]
port 601 nsew signal input
rlabel metal3 s 449200 81064 450000 81184 6 mgmt_in_data[1]
port 602 nsew signal input
rlabel metal3 s 449200 153552 450000 153672 6 mgmt_in_data[20]
port 603 nsew signal input
rlabel metal3 s 449200 157360 450000 157480 6 mgmt_in_data[21]
port 604 nsew signal input
rlabel metal3 s 449200 161168 450000 161288 6 mgmt_in_data[22]
port 605 nsew signal input
rlabel metal3 s 449200 164976 450000 165096 6 mgmt_in_data[23]
port 606 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 mgmt_in_data[24]
port 607 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 mgmt_in_data[25]
port 608 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 mgmt_in_data[26]
port 609 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 mgmt_in_data[27]
port 610 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 mgmt_in_data[28]
port 611 nsew signal input
rlabel metal3 s 0 154504 800 154624 6 mgmt_in_data[29]
port 612 nsew signal input
rlabel metal3 s 449200 84872 450000 84992 6 mgmt_in_data[2]
port 613 nsew signal input
rlabel metal3 s 0 156000 800 156120 6 mgmt_in_data[30]
port 614 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 mgmt_in_data[31]
port 615 nsew signal input
rlabel metal3 s 0 158992 800 159112 6 mgmt_in_data[32]
port 616 nsew signal input
rlabel metal3 s 0 160624 800 160744 6 mgmt_in_data[33]
port 617 nsew signal input
rlabel metal3 s 0 162120 800 162240 6 mgmt_in_data[34]
port 618 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 mgmt_in_data[35]
port 619 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 mgmt_in_data[36]
port 620 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 mgmt_in_data[37]
port 621 nsew signal input
rlabel metal3 s 449200 88680 450000 88800 6 mgmt_in_data[3]
port 622 nsew signal input
rlabel metal3 s 449200 92488 450000 92608 6 mgmt_in_data[4]
port 623 nsew signal input
rlabel metal3 s 449200 96296 450000 96416 6 mgmt_in_data[5]
port 624 nsew signal input
rlabel metal3 s 449200 100104 450000 100224 6 mgmt_in_data[6]
port 625 nsew signal input
rlabel metal3 s 449200 103912 450000 104032 6 mgmt_in_data[7]
port 626 nsew signal input
rlabel metal3 s 449200 107720 450000 107840 6 mgmt_in_data[8]
port 627 nsew signal input
rlabel metal3 s 449200 111528 450000 111648 6 mgmt_in_data[9]
port 628 nsew signal input
rlabel metal3 s 449200 79160 450000 79280 6 mgmt_out_data[0]
port 629 nsew signal output
rlabel metal3 s 449200 117376 450000 117496 6 mgmt_out_data[10]
port 630 nsew signal output
rlabel metal3 s 449200 121184 450000 121304 6 mgmt_out_data[11]
port 631 nsew signal output
rlabel metal3 s 449200 124992 450000 125112 6 mgmt_out_data[12]
port 632 nsew signal output
rlabel metal3 s 449200 128800 450000 128920 6 mgmt_out_data[13]
port 633 nsew signal output
rlabel metal3 s 449200 132608 450000 132728 6 mgmt_out_data[14]
port 634 nsew signal output
rlabel metal3 s 449200 136416 450000 136536 6 mgmt_out_data[15]
port 635 nsew signal output
rlabel metal3 s 449200 140224 450000 140344 6 mgmt_out_data[16]
port 636 nsew signal output
rlabel metal3 s 449200 144032 450000 144152 6 mgmt_out_data[17]
port 637 nsew signal output
rlabel metal3 s 449200 147840 450000 147960 6 mgmt_out_data[18]
port 638 nsew signal output
rlabel metal3 s 449200 151648 450000 151768 6 mgmt_out_data[19]
port 639 nsew signal output
rlabel metal3 s 449200 82968 450000 83088 6 mgmt_out_data[1]
port 640 nsew signal output
rlabel metal3 s 449200 155456 450000 155576 6 mgmt_out_data[20]
port 641 nsew signal output
rlabel metal3 s 449200 159264 450000 159384 6 mgmt_out_data[21]
port 642 nsew signal output
rlabel metal3 s 449200 163072 450000 163192 6 mgmt_out_data[22]
port 643 nsew signal output
rlabel metal3 s 449200 166880 450000 167000 6 mgmt_out_data[23]
port 644 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 mgmt_out_data[24]
port 645 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 mgmt_out_data[25]
port 646 nsew signal output
rlabel metal3 s 0 150696 800 150816 6 mgmt_out_data[26]
port 647 nsew signal output
rlabel metal3 s 0 152192 800 152312 6 mgmt_out_data[27]
port 648 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 mgmt_out_data[28]
port 649 nsew signal output
rlabel metal3 s 0 155320 800 155440 6 mgmt_out_data[29]
port 650 nsew signal output
rlabel metal3 s 449200 86776 450000 86896 6 mgmt_out_data[2]
port 651 nsew signal output
rlabel metal3 s 0 156816 800 156936 6 mgmt_out_data[30]
port 652 nsew signal output
rlabel metal3 s 0 158312 800 158432 6 mgmt_out_data[31]
port 653 nsew signal output
rlabel metal3 s 0 159808 800 159928 6 mgmt_out_data[32]
port 654 nsew signal output
rlabel metal3 s 0 161304 800 161424 6 mgmt_out_data[33]
port 655 nsew signal output
rlabel metal3 s 0 162800 800 162920 6 mgmt_out_data[34]
port 656 nsew signal output
rlabel metal3 s 0 164432 800 164552 6 mgmt_out_data[35]
port 657 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 mgmt_out_data[36]
port 658 nsew signal output
rlabel metal3 s 0 167424 800 167544 6 mgmt_out_data[37]
port 659 nsew signal output
rlabel metal3 s 449200 90584 450000 90704 6 mgmt_out_data[3]
port 660 nsew signal output
rlabel metal3 s 449200 94392 450000 94512 6 mgmt_out_data[4]
port 661 nsew signal output
rlabel metal3 s 449200 98200 450000 98320 6 mgmt_out_data[5]
port 662 nsew signal output
rlabel metal3 s 449200 102008 450000 102128 6 mgmt_out_data[6]
port 663 nsew signal output
rlabel metal3 s 449200 105816 450000 105936 6 mgmt_out_data[7]
port 664 nsew signal output
rlabel metal3 s 449200 109624 450000 109744 6 mgmt_out_data[8]
port 665 nsew signal output
rlabel metal3 s 449200 113568 450000 113688 6 mgmt_out_data[9]
port 666 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 mgmt_rdata[0]
port 667 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 mgmt_rdata[10]
port 668 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 mgmt_rdata[11]
port 669 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 mgmt_rdata[12]
port 670 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 mgmt_rdata[13]
port 671 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 mgmt_rdata[14]
port 672 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 mgmt_rdata[15]
port 673 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 mgmt_rdata[16]
port 674 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 mgmt_rdata[17]
port 675 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 mgmt_rdata[18]
port 676 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 mgmt_rdata[19]
port 677 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 mgmt_rdata[1]
port 678 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 mgmt_rdata[20]
port 679 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 mgmt_rdata[21]
port 680 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 mgmt_rdata[22]
port 681 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 mgmt_rdata[23]
port 682 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 mgmt_rdata[24]
port 683 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 mgmt_rdata[25]
port 684 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 mgmt_rdata[26]
port 685 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 mgmt_rdata[27]
port 686 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 mgmt_rdata[28]
port 687 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 mgmt_rdata[29]
port 688 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 mgmt_rdata[2]
port 689 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 mgmt_rdata[30]
port 690 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 mgmt_rdata[31]
port 691 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 mgmt_rdata[32]
port 692 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 mgmt_rdata[33]
port 693 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 mgmt_rdata[34]
port 694 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 mgmt_rdata[35]
port 695 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 mgmt_rdata[36]
port 696 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 mgmt_rdata[37]
port 697 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 mgmt_rdata[38]
port 698 nsew signal input
rlabel metal3 s 0 100512 800 100632 6 mgmt_rdata[39]
port 699 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 mgmt_rdata[3]
port 700 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 mgmt_rdata[40]
port 701 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 mgmt_rdata[41]
port 702 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 mgmt_rdata[42]
port 703 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 mgmt_rdata[43]
port 704 nsew signal input
rlabel metal3 s 0 104320 800 104440 6 mgmt_rdata[44]
port 705 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 mgmt_rdata[45]
port 706 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 mgmt_rdata[46]
port 707 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 mgmt_rdata[47]
port 708 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 mgmt_rdata[48]
port 709 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 mgmt_rdata[49]
port 710 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 mgmt_rdata[4]
port 711 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 mgmt_rdata[50]
port 712 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 mgmt_rdata[51]
port 713 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 mgmt_rdata[52]
port 714 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 mgmt_rdata[53]
port 715 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 mgmt_rdata[54]
port 716 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 mgmt_rdata[55]
port 717 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 mgmt_rdata[56]
port 718 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 mgmt_rdata[57]
port 719 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 mgmt_rdata[58]
port 720 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 mgmt_rdata[59]
port 721 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 mgmt_rdata[5]
port 722 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 mgmt_rdata[60]
port 723 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 mgmt_rdata[61]
port 724 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 mgmt_rdata[62]
port 725 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 mgmt_rdata[63]
port 726 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 mgmt_rdata[6]
port 727 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 mgmt_rdata[7]
port 728 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 mgmt_rdata[8]
port 729 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 mgmt_rdata[9]
port 730 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 mgmt_rdata_ro[0]
port 731 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 mgmt_rdata_ro[10]
port 732 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 mgmt_rdata_ro[11]
port 733 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 mgmt_rdata_ro[12]
port 734 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 mgmt_rdata_ro[13]
port 735 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 mgmt_rdata_ro[14]
port 736 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 mgmt_rdata_ro[15]
port 737 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 mgmt_rdata_ro[16]
port 738 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 mgmt_rdata_ro[17]
port 739 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 mgmt_rdata_ro[18]
port 740 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 mgmt_rdata_ro[19]
port 741 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 mgmt_rdata_ro[1]
port 742 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 mgmt_rdata_ro[20]
port 743 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 mgmt_rdata_ro[21]
port 744 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 mgmt_rdata_ro[22]
port 745 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 mgmt_rdata_ro[23]
port 746 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 mgmt_rdata_ro[24]
port 747 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 mgmt_rdata_ro[25]
port 748 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 mgmt_rdata_ro[26]
port 749 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 mgmt_rdata_ro[27]
port 750 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 mgmt_rdata_ro[28]
port 751 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 mgmt_rdata_ro[29]
port 752 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 mgmt_rdata_ro[2]
port 753 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 mgmt_rdata_ro[30]
port 754 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 mgmt_rdata_ro[31]
port 755 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 mgmt_rdata_ro[3]
port 756 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 mgmt_rdata_ro[4]
port 757 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 mgmt_rdata_ro[5]
port 758 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 mgmt_rdata_ro[6]
port 759 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 mgmt_rdata_ro[7]
port 760 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 mgmt_rdata_ro[8]
port 761 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 mgmt_rdata_ro[9]
port 762 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 mgmt_wdata[0]
port 763 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 mgmt_wdata[10]
port 764 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 mgmt_wdata[11]
port 765 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 mgmt_wdata[12]
port 766 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 mgmt_wdata[13]
port 767 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 mgmt_wdata[14]
port 768 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 mgmt_wdata[15]
port 769 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 mgmt_wdata[16]
port 770 nsew signal output
rlabel metal3 s 0 79296 800 79416 6 mgmt_wdata[17]
port 771 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 mgmt_wdata[18]
port 772 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 mgmt_wdata[19]
port 773 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 mgmt_wdata[1]
port 774 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 mgmt_wdata[20]
port 775 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 mgmt_wdata[21]
port 776 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 mgmt_wdata[22]
port 777 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 mgmt_wdata[23]
port 778 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 mgmt_wdata[24]
port 779 nsew signal output
rlabel metal3 s 0 85280 800 85400 6 mgmt_wdata[25]
port 780 nsew signal output
rlabel metal3 s 0 86096 800 86216 6 mgmt_wdata[26]
port 781 nsew signal output
rlabel metal3 s 0 86912 800 87032 6 mgmt_wdata[27]
port 782 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 mgmt_wdata[28]
port 783 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 mgmt_wdata[29]
port 784 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 mgmt_wdata[2]
port 785 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 mgmt_wdata[30]
port 786 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 mgmt_wdata[31]
port 787 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 mgmt_wdata[3]
port 788 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 mgmt_wdata[4]
port 789 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 mgmt_wdata[5]
port 790 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 mgmt_wdata[6]
port 791 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 mgmt_wdata[7]
port 792 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 mgmt_wdata[8]
port 793 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 mgmt_wdata[9]
port 794 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 mgmt_wen[0]
port 795 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 mgmt_wen[1]
port 796 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 mgmt_wen_mask[0]
port 797 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 mgmt_wen_mask[1]
port 798 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 mgmt_wen_mask[2]
port 799 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 mgmt_wen_mask[3]
port 800 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 mgmt_wen_mask[4]
port 801 nsew signal output
rlabel metal3 s 0 92896 800 93016 6 mgmt_wen_mask[5]
port 802 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 mgmt_wen_mask[6]
port 803 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 mgmt_wen_mask[7]
port 804 nsew signal output
rlabel metal2 s 443550 167200 443606 168000 6 mprj2_vcc_pwrgood
port 805 nsew signal input
rlabel metal2 s 445022 167200 445078 168000 6 mprj2_vdd_pwrgood
port 806 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 mprj_ack_i
port 807 nsew signal input
rlabel metal2 s 391386 167200 391442 168000 6 mprj_adr_o[0]
port 808 nsew signal output
rlabel metal2 s 409510 167200 409566 168000 6 mprj_adr_o[10]
port 809 nsew signal output
rlabel metal2 s 411074 167200 411130 168000 6 mprj_adr_o[11]
port 810 nsew signal output
rlabel metal2 s 412546 167200 412602 168000 6 mprj_adr_o[12]
port 811 nsew signal output
rlabel metal2 s 414110 167200 414166 168000 6 mprj_adr_o[13]
port 812 nsew signal output
rlabel metal2 s 415582 167200 415638 168000 6 mprj_adr_o[14]
port 813 nsew signal output
rlabel metal2 s 417054 167200 417110 168000 6 mprj_adr_o[15]
port 814 nsew signal output
rlabel metal2 s 418618 167200 418674 168000 6 mprj_adr_o[16]
port 815 nsew signal output
rlabel metal2 s 420090 167200 420146 168000 6 mprj_adr_o[17]
port 816 nsew signal output
rlabel metal2 s 421654 167200 421710 168000 6 mprj_adr_o[18]
port 817 nsew signal output
rlabel metal2 s 423126 167200 423182 168000 6 mprj_adr_o[19]
port 818 nsew signal output
rlabel metal2 s 393686 167200 393742 168000 6 mprj_adr_o[1]
port 819 nsew signal output
rlabel metal2 s 424598 167200 424654 168000 6 mprj_adr_o[20]
port 820 nsew signal output
rlabel metal2 s 426162 167200 426218 168000 6 mprj_adr_o[21]
port 821 nsew signal output
rlabel metal2 s 427634 167200 427690 168000 6 mprj_adr_o[22]
port 822 nsew signal output
rlabel metal2 s 429198 167200 429254 168000 6 mprj_adr_o[23]
port 823 nsew signal output
rlabel metal2 s 430670 167200 430726 168000 6 mprj_adr_o[24]
port 824 nsew signal output
rlabel metal2 s 432234 167200 432290 168000 6 mprj_adr_o[25]
port 825 nsew signal output
rlabel metal2 s 433706 167200 433762 168000 6 mprj_adr_o[26]
port 826 nsew signal output
rlabel metal2 s 435178 167200 435234 168000 6 mprj_adr_o[27]
port 827 nsew signal output
rlabel metal2 s 436742 167200 436798 168000 6 mprj_adr_o[28]
port 828 nsew signal output
rlabel metal2 s 438214 167200 438270 168000 6 mprj_adr_o[29]
port 829 nsew signal output
rlabel metal2 s 395986 167200 396042 168000 6 mprj_adr_o[2]
port 830 nsew signal output
rlabel metal2 s 439778 167200 439834 168000 6 mprj_adr_o[30]
port 831 nsew signal output
rlabel metal2 s 441250 167200 441306 168000 6 mprj_adr_o[31]
port 832 nsew signal output
rlabel metal2 s 398194 167200 398250 168000 6 mprj_adr_o[3]
port 833 nsew signal output
rlabel metal2 s 400494 167200 400550 168000 6 mprj_adr_o[4]
port 834 nsew signal output
rlabel metal2 s 401966 167200 402022 168000 6 mprj_adr_o[5]
port 835 nsew signal output
rlabel metal2 s 403530 167200 403586 168000 6 mprj_adr_o[6]
port 836 nsew signal output
rlabel metal2 s 405002 167200 405058 168000 6 mprj_adr_o[7]
port 837 nsew signal output
rlabel metal2 s 406566 167200 406622 168000 6 mprj_adr_o[8]
port 838 nsew signal output
rlabel metal2 s 408038 167200 408094 168000 6 mprj_adr_o[9]
port 839 nsew signal output
rlabel metal2 s 389178 167200 389234 168000 6 mprj_cyc_o
port 840 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 mprj_dat_i[0]
port 841 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 mprj_dat_i[10]
port 842 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 mprj_dat_i[11]
port 843 nsew signal input
rlabel metal3 s 0 130976 800 131096 6 mprj_dat_i[12]
port 844 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 mprj_dat_i[13]
port 845 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 mprj_dat_i[14]
port 846 nsew signal input
rlabel metal3 s 0 133152 800 133272 6 mprj_dat_i[15]
port 847 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 mprj_dat_i[16]
port 848 nsew signal input
rlabel metal3 s 0 134784 800 134904 6 mprj_dat_i[17]
port 849 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 mprj_dat_i[18]
port 850 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 mprj_dat_i[19]
port 851 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 mprj_dat_i[1]
port 852 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 mprj_dat_i[20]
port 853 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 mprj_dat_i[21]
port 854 nsew signal input
rlabel metal3 s 0 138592 800 138712 6 mprj_dat_i[22]
port 855 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 mprj_dat_i[23]
port 856 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 mprj_dat_i[24]
port 857 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 mprj_dat_i[25]
port 858 nsew signal input
rlabel metal3 s 0 141584 800 141704 6 mprj_dat_i[26]
port 859 nsew signal input
rlabel metal3 s 0 142400 800 142520 6 mprj_dat_i[27]
port 860 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 mprj_dat_i[28]
port 861 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 mprj_dat_i[29]
port 862 nsew signal input
rlabel metal3 s 0 123360 800 123480 6 mprj_dat_i[2]
port 863 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 mprj_dat_i[30]
port 864 nsew signal input
rlabel metal3 s 0 145392 800 145512 6 mprj_dat_i[31]
port 865 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 mprj_dat_i[3]
port 866 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 mprj_dat_i[4]
port 867 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 mprj_dat_i[5]
port 868 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 mprj_dat_i[6]
port 869 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 mprj_dat_i[7]
port 870 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 mprj_dat_i[8]
port 871 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 mprj_dat_i[9]
port 872 nsew signal input
rlabel metal2 s 392214 167200 392270 168000 6 mprj_dat_o[0]
port 873 nsew signal output
rlabel metal2 s 410338 167200 410394 168000 6 mprj_dat_o[10]
port 874 nsew signal output
rlabel metal2 s 411810 167200 411866 168000 6 mprj_dat_o[11]
port 875 nsew signal output
rlabel metal2 s 413282 167200 413338 168000 6 mprj_dat_o[12]
port 876 nsew signal output
rlabel metal2 s 414846 167200 414902 168000 6 mprj_dat_o[13]
port 877 nsew signal output
rlabel metal2 s 416318 167200 416374 168000 6 mprj_dat_o[14]
port 878 nsew signal output
rlabel metal2 s 417882 167200 417938 168000 6 mprj_dat_o[15]
port 879 nsew signal output
rlabel metal2 s 419354 167200 419410 168000 6 mprj_dat_o[16]
port 880 nsew signal output
rlabel metal2 s 420826 167200 420882 168000 6 mprj_dat_o[17]
port 881 nsew signal output
rlabel metal2 s 422390 167200 422446 168000 6 mprj_dat_o[18]
port 882 nsew signal output
rlabel metal2 s 423862 167200 423918 168000 6 mprj_dat_o[19]
port 883 nsew signal output
rlabel metal2 s 394422 167200 394478 168000 6 mprj_dat_o[1]
port 884 nsew signal output
rlabel metal2 s 425426 167200 425482 168000 6 mprj_dat_o[20]
port 885 nsew signal output
rlabel metal2 s 426898 167200 426954 168000 6 mprj_dat_o[21]
port 886 nsew signal output
rlabel metal2 s 428462 167200 428518 168000 6 mprj_dat_o[22]
port 887 nsew signal output
rlabel metal2 s 429934 167200 429990 168000 6 mprj_dat_o[23]
port 888 nsew signal output
rlabel metal2 s 431406 167200 431462 168000 6 mprj_dat_o[24]
port 889 nsew signal output
rlabel metal2 s 432970 167200 433026 168000 6 mprj_dat_o[25]
port 890 nsew signal output
rlabel metal2 s 434442 167200 434498 168000 6 mprj_dat_o[26]
port 891 nsew signal output
rlabel metal2 s 436006 167200 436062 168000 6 mprj_dat_o[27]
port 892 nsew signal output
rlabel metal2 s 437478 167200 437534 168000 6 mprj_dat_o[28]
port 893 nsew signal output
rlabel metal2 s 438950 167200 439006 168000 6 mprj_dat_o[29]
port 894 nsew signal output
rlabel metal2 s 396722 167200 396778 168000 6 mprj_dat_o[2]
port 895 nsew signal output
rlabel metal2 s 440514 167200 440570 168000 6 mprj_dat_o[30]
port 896 nsew signal output
rlabel metal2 s 441986 167200 442042 168000 6 mprj_dat_o[31]
port 897 nsew signal output
rlabel metal2 s 398930 167200 398986 168000 6 mprj_dat_o[3]
port 898 nsew signal output
rlabel metal2 s 401230 167200 401286 168000 6 mprj_dat_o[4]
port 899 nsew signal output
rlabel metal2 s 402702 167200 402758 168000 6 mprj_dat_o[5]
port 900 nsew signal output
rlabel metal2 s 404266 167200 404322 168000 6 mprj_dat_o[6]
port 901 nsew signal output
rlabel metal2 s 405738 167200 405794 168000 6 mprj_dat_o[7]
port 902 nsew signal output
rlabel metal2 s 407302 167200 407358 168000 6 mprj_dat_o[8]
port 903 nsew signal output
rlabel metal2 s 408774 167200 408830 168000 6 mprj_dat_o[9]
port 904 nsew signal output
rlabel metal3 s 449200 69640 450000 69760 6 mprj_io_loader_clock
port 905 nsew signal output
rlabel metal3 s 449200 75352 450000 75472 6 mprj_io_loader_data_1
port 906 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 mprj_io_loader_data_2
port 907 nsew signal output
rlabel metal3 s 449200 67736 450000 67856 6 mprj_io_loader_resetn
port 908 nsew signal output
rlabel metal2 s 392950 167200 393006 168000 6 mprj_sel_o[0]
port 909 nsew signal output
rlabel metal2 s 395158 167200 395214 168000 6 mprj_sel_o[1]
port 910 nsew signal output
rlabel metal2 s 397458 167200 397514 168000 6 mprj_sel_o[2]
port 911 nsew signal output
rlabel metal2 s 399758 167200 399814 168000 6 mprj_sel_o[3]
port 912 nsew signal output
rlabel metal2 s 389914 167200 389970 168000 6 mprj_stb_o
port 913 nsew signal output
rlabel metal2 s 442722 167200 442778 168000 6 mprj_vcc_pwrgood
port 914 nsew signal input
rlabel metal2 s 444286 167200 444342 168000 6 mprj_vdd_pwrgood
port 915 nsew signal input
rlabel metal2 s 390650 167200 390706 168000 6 mprj_we_o
port 916 nsew signal output
rlabel metal3 s 449200 62024 450000 62144 6 porb
port 917 nsew signal input
rlabel metal2 s 389362 0 389418 800 6 pwr_ctrl_out[0]
port 918 nsew signal output
rlabel metal2 s 406658 0 406714 800 6 pwr_ctrl_out[1]
port 919 nsew signal output
rlabel metal2 s 423954 0 424010 800 6 pwr_ctrl_out[2]
port 920 nsew signal output
rlabel metal2 s 441250 0 441306 800 6 pwr_ctrl_out[3]
port 921 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 resetb
port 922 nsew signal input
rlabel metal3 s 449200 71544 450000 71664 6 sdo_out
port 923 nsew signal output
rlabel metal3 s 449200 73448 450000 73568 6 sdo_outenb
port 924 nsew signal output
rlabel metal2 s 1858 167200 1914 168000 6 user_clk
port 925 nsew signal output
rlabel metal2 s 445758 167200 445814 168000 6 user_irq[0]
port 926 nsew signal input
rlabel metal2 s 446494 167200 446550 168000 6 user_irq[1]
port 927 nsew signal input
rlabel metal2 s 447322 167200 447378 168000 6 user_irq[2]
port 928 nsew signal input
rlabel metal2 s 448058 167200 448114 168000 6 user_irq_ena[0]
port 929 nsew signal output
rlabel metal2 s 448794 167200 448850 168000 6 user_irq_ena[1]
port 930 nsew signal output
rlabel metal2 s 449530 167200 449586 168000 6 user_irq_ena[2]
port 931 nsew signal output
rlabel metal4 s 444208 2128 444528 165424 6 VPWR
port 932 nsew power bidirectional
rlabel metal4 s 434208 2128 434528 165424 6 VPWR
port 933 nsew power bidirectional
rlabel metal4 s 424208 2128 424528 165424 6 VPWR
port 934 nsew power bidirectional
rlabel metal4 s 414208 2128 414528 165424 6 VPWR
port 935 nsew power bidirectional
rlabel metal4 s 404208 2128 404528 165424 6 VPWR
port 936 nsew power bidirectional
rlabel metal4 s 394208 164296 394528 165424 6 VPWR
port 937 nsew power bidirectional
rlabel metal4 s 384208 2128 384528 165424 6 VPWR
port 938 nsew power bidirectional
rlabel metal4 s 374208 2128 374528 165424 6 VPWR
port 939 nsew power bidirectional
rlabel metal4 s 364208 2128 364528 165424 6 VPWR
port 940 nsew power bidirectional
rlabel metal4 s 354208 2128 354528 165424 6 VPWR
port 941 nsew power bidirectional
rlabel metal4 s 344208 2128 344528 165424 6 VPWR
port 942 nsew power bidirectional
rlabel metal4 s 334208 2128 334528 165424 6 VPWR
port 943 nsew power bidirectional
rlabel metal4 s 324208 2128 324528 165424 6 VPWR
port 944 nsew power bidirectional
rlabel metal4 s 314208 2128 314528 165424 6 VPWR
port 945 nsew power bidirectional
rlabel metal4 s 304208 2128 304528 165424 6 VPWR
port 946 nsew power bidirectional
rlabel metal4 s 294208 2128 294528 165424 6 VPWR
port 947 nsew power bidirectional
rlabel metal4 s 284208 2128 284528 165424 6 VPWR
port 948 nsew power bidirectional
rlabel metal4 s 274208 2128 274528 165424 6 VPWR
port 949 nsew power bidirectional
rlabel metal4 s 264208 2128 264528 165424 6 VPWR
port 950 nsew power bidirectional
rlabel metal4 s 254208 2128 254528 165424 6 VPWR
port 951 nsew power bidirectional
rlabel metal4 s 244208 2128 244528 165424 6 VPWR
port 952 nsew power bidirectional
rlabel metal4 s 234208 2128 234528 165424 6 VPWR
port 953 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 165424 6 VPWR
port 954 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 165424 6 VPWR
port 955 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 165424 6 VPWR
port 956 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 165424 6 VPWR
port 957 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 165424 6 VPWR
port 958 nsew power bidirectional
rlabel metal4 s 174208 128152 174528 165424 6 VPWR
port 959 nsew power bidirectional
rlabel metal4 s 164208 128152 164528 165424 6 VPWR
port 960 nsew power bidirectional
rlabel metal4 s 154208 128152 154528 165424 6 VPWR
port 961 nsew power bidirectional
rlabel metal4 s 144208 128152 144528 165424 6 VPWR
port 962 nsew power bidirectional
rlabel metal4 s 134208 128152 134528 165424 6 VPWR
port 963 nsew power bidirectional
rlabel metal4 s 124208 128152 124528 165424 6 VPWR
port 964 nsew power bidirectional
rlabel metal4 s 114208 128152 114528 165424 6 VPWR
port 965 nsew power bidirectional
rlabel metal4 s 104208 128152 104528 165424 6 VPWR
port 966 nsew power bidirectional
rlabel metal4 s 94208 128152 94528 165424 6 VPWR
port 967 nsew power bidirectional
rlabel metal4 s 84208 128152 84528 165424 6 VPWR
port 968 nsew power bidirectional
rlabel metal4 s 74208 128152 74528 165424 6 VPWR
port 969 nsew power bidirectional
rlabel metal4 s 64208 128152 64528 165424 6 VPWR
port 970 nsew power bidirectional
rlabel metal4 s 54208 128152 54528 165424 6 VPWR
port 971 nsew power bidirectional
rlabel metal4 s 44208 128152 44528 165424 6 VPWR
port 972 nsew power bidirectional
rlabel metal4 s 34208 128152 34528 165424 6 VPWR
port 973 nsew power bidirectional
rlabel metal4 s 24208 128152 24528 165424 6 VPWR
port 974 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 165424 6 VPWR
port 975 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 165424 6 VPWR
port 976 nsew power bidirectional
rlabel metal4 s 394208 2128 394528 145392 6 VPWR
port 977 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 21248 6 VPWR
port 978 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 21248 6 VPWR
port 979 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 21248 6 VPWR
port 980 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 21248 6 VPWR
port 981 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 21248 6 VPWR
port 982 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 21248 6 VPWR
port 983 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 21248 6 VPWR
port 984 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 21248 6 VPWR
port 985 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 21248 6 VPWR
port 986 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 21248 6 VPWR
port 987 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 21248 6 VPWR
port 988 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 21248 6 VPWR
port 989 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 21248 6 VPWR
port 990 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 21248 6 VPWR
port 991 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 21248 6 VPWR
port 992 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 21248 6 VPWR
port 993 nsew power bidirectional
rlabel metal5 s 1104 161298 448868 161618 6 VPWR
port 994 nsew power bidirectional
rlabel metal5 s 1104 135298 448868 135618 6 VPWR
port 995 nsew power bidirectional
rlabel metal5 s 1104 109298 448868 109618 6 VPWR
port 996 nsew power bidirectional
rlabel metal5 s 1104 83298 448868 83618 6 VPWR
port 997 nsew power bidirectional
rlabel metal5 s 1104 57298 448868 57618 6 VPWR
port 998 nsew power bidirectional
rlabel metal5 s 1104 31298 448868 31618 6 VPWR
port 999 nsew power bidirectional
rlabel metal5 s 1104 5298 448868 5618 6 VPWR
port 1000 nsew power bidirectional
rlabel metal4 s 439208 2128 439528 165424 6 VGND
port 1001 nsew ground bidirectional
rlabel metal4 s 429208 2128 429528 165424 6 VGND
port 1002 nsew ground bidirectional
rlabel metal4 s 419208 2128 419528 165424 6 VGND
port 1003 nsew ground bidirectional
rlabel metal4 s 409208 2128 409528 165424 6 VGND
port 1004 nsew ground bidirectional
rlabel metal4 s 399208 164296 399528 165424 6 VGND
port 1005 nsew ground bidirectional
rlabel metal4 s 389208 164296 389528 165424 6 VGND
port 1006 nsew ground bidirectional
rlabel metal4 s 379208 2128 379528 165424 6 VGND
port 1007 nsew ground bidirectional
rlabel metal4 s 369208 2128 369528 165424 6 VGND
port 1008 nsew ground bidirectional
rlabel metal4 s 359208 2128 359528 165424 6 VGND
port 1009 nsew ground bidirectional
rlabel metal4 s 349208 2128 349528 165424 6 VGND
port 1010 nsew ground bidirectional
rlabel metal4 s 339208 2128 339528 165424 6 VGND
port 1011 nsew ground bidirectional
rlabel metal4 s 329208 2128 329528 165424 6 VGND
port 1012 nsew ground bidirectional
rlabel metal4 s 319208 2128 319528 165424 6 VGND
port 1013 nsew ground bidirectional
rlabel metal4 s 309208 2128 309528 165424 6 VGND
port 1014 nsew ground bidirectional
rlabel metal4 s 299208 2128 299528 165424 6 VGND
port 1015 nsew ground bidirectional
rlabel metal4 s 289208 2128 289528 165424 6 VGND
port 1016 nsew ground bidirectional
rlabel metal4 s 279208 2128 279528 165424 6 VGND
port 1017 nsew ground bidirectional
rlabel metal4 s 269208 2128 269528 165424 6 VGND
port 1018 nsew ground bidirectional
rlabel metal4 s 259208 2128 259528 165424 6 VGND
port 1019 nsew ground bidirectional
rlabel metal4 s 249208 2128 249528 165424 6 VGND
port 1020 nsew ground bidirectional
rlabel metal4 s 239208 2128 239528 165424 6 VGND
port 1021 nsew ground bidirectional
rlabel metal4 s 229208 2128 229528 165424 6 VGND
port 1022 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 165424 6 VGND
port 1023 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 165424 6 VGND
port 1024 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 165424 6 VGND
port 1025 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 165424 6 VGND
port 1026 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 165424 6 VGND
port 1027 nsew ground bidirectional
rlabel metal4 s 169208 128152 169528 165424 6 VGND
port 1028 nsew ground bidirectional
rlabel metal4 s 159208 128152 159528 165424 6 VGND
port 1029 nsew ground bidirectional
rlabel metal4 s 149208 128152 149528 165424 6 VGND
port 1030 nsew ground bidirectional
rlabel metal4 s 139208 128152 139528 165424 6 VGND
port 1031 nsew ground bidirectional
rlabel metal4 s 129208 128152 129528 165424 6 VGND
port 1032 nsew ground bidirectional
rlabel metal4 s 119208 128152 119528 165424 6 VGND
port 1033 nsew ground bidirectional
rlabel metal4 s 109208 128152 109528 165424 6 VGND
port 1034 nsew ground bidirectional
rlabel metal4 s 99208 128152 99528 165424 6 VGND
port 1035 nsew ground bidirectional
rlabel metal4 s 89208 128152 89528 165424 6 VGND
port 1036 nsew ground bidirectional
rlabel metal4 s 79208 128152 79528 165424 6 VGND
port 1037 nsew ground bidirectional
rlabel metal4 s 69208 128152 69528 165424 6 VGND
port 1038 nsew ground bidirectional
rlabel metal4 s 59208 128152 59528 165424 6 VGND
port 1039 nsew ground bidirectional
rlabel metal4 s 49208 128152 49528 165424 6 VGND
port 1040 nsew ground bidirectional
rlabel metal4 s 39208 128152 39528 165424 6 VGND
port 1041 nsew ground bidirectional
rlabel metal4 s 29208 128152 29528 165424 6 VGND
port 1042 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 165424 6 VGND
port 1043 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 165424 6 VGND
port 1044 nsew ground bidirectional
rlabel metal4 s 399208 2128 399528 145392 6 VGND
port 1045 nsew ground bidirectional
rlabel metal4 s 389208 2128 389528 145392 6 VGND
port 1046 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 21248 6 VGND
port 1047 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 21248 6 VGND
port 1048 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 21248 6 VGND
port 1049 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 21248 6 VGND
port 1050 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 21248 6 VGND
port 1051 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 21248 6 VGND
port 1052 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 21248 6 VGND
port 1053 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 21248 6 VGND
port 1054 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 21248 6 VGND
port 1055 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 21248 6 VGND
port 1056 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 21248 6 VGND
port 1057 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 21248 6 VGND
port 1058 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 21248 6 VGND
port 1059 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 21248 6 VGND
port 1060 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 21248 6 VGND
port 1061 nsew ground bidirectional
rlabel metal5 s 1104 148298 448868 148618 6 VGND
port 1062 nsew ground bidirectional
rlabel metal5 s 1104 122298 448868 122618 6 VGND
port 1063 nsew ground bidirectional
rlabel metal5 s 1104 96298 448868 96618 6 VGND
port 1064 nsew ground bidirectional
rlabel metal5 s 1104 70298 448868 70618 6 VGND
port 1065 nsew ground bidirectional
rlabel metal5 s 1104 44298 448868 44618 6 VGND
port 1066 nsew ground bidirectional
rlabel metal5 s 1104 18298 448868 18618 6 VGND
port 1067 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 450000 168000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core/runs/mgmt_core/results/magic/mgmt_core.gds
string GDS_END 175437274
string GDS_START 62915804
<< end >>

