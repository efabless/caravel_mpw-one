magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 2168 2245
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_0
timestamp 1623348570
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_1
timestamp 1623348570
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_2
timestamp 1623348570
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_3
timestamp 1623348570
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_4
timestamp 1623348570
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_1
timestamp 1623348570
transform 1 0 880 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 908 985 908 985 0 FreeSans 300 0 0 0 S
flabel comment s 752 985 752 985 0 FreeSans 300 0 0 0 D
flabel comment s 596 985 596 985 0 FreeSans 300 0 0 0 S
flabel comment s 440 985 440 985 0 FreeSans 300 0 0 0 D
flabel comment s 284 985 284 985 0 FreeSans 300 0 0 0 S
flabel comment s 128 985 128 985 0 FreeSans 300 0 0 0 D
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 43805558
string GDS_START 43801924
<< end >>
