// Copyright 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module caravel(vddio, vssio, vdda, vssa, vccd, vssd, vdda1, vdda2, vssa1, vssa2, vccd1, vccd2, vssd1, vssd2, gpio, mprj_io, pwr_ctrl_out, clock, resetb, flash_csb, flash_clk, flash_io0, flash_io1);
  wire caravel_clk;
  wire caravel_clk2;
  wire caravel_rstn;
  input clock;
  wire clock_core;
  output flash_clk;
  wire flash_clk_core;
  wire flash_clk_ieb_core;
  wire flash_clk_oeb_core;
  output flash_csb;
  wire flash_csb_core;
  wire flash_csb_ieb_core;
  wire flash_csb_oeb_core;
  output flash_io0;
  wire flash_io0_di_core;
  wire flash_io0_do_core;
  wire flash_io0_ieb_core;
  wire flash_io0_oeb_core;
  output flash_io1;
  wire flash_io1_di_core;
  wire flash_io1_do_core;
  wire flash_io1_ieb_core;
  wire flash_io1_oeb_core;
  wire flash_io2_di_core;
  wire flash_io2_do_core;
  wire flash_io2_ieb_core;
  wire flash_io2_oeb_core;
  wire flash_io3_di_core;
  wire flash_io3_do_core;
  wire flash_io3_ieb_core;
  wire flash_io3_oeb_core;
  inout gpio;
  wire gpio_in_core;
  wire gpio_inenb_core;
  wire gpio_mode0_core;
  wire gpio_mode1_core;
  wire gpio_out_core;
  wire gpio_outenb_core;
  wire \gpio_serial_link[0] ;
  wire \gpio_serial_link[10] ;
  wire \gpio_serial_link[11] ;
  wire \gpio_serial_link[12] ;
  wire \gpio_serial_link[13] ;
  wire \gpio_serial_link[14] ;
  wire \gpio_serial_link[15] ;
  wire \gpio_serial_link[16] ;
  wire \gpio_serial_link[17] ;
  wire \gpio_serial_link[18] ;
  wire \gpio_serial_link[19] ;
  wire \gpio_serial_link[1] ;
  wire \gpio_serial_link[20] ;
  wire \gpio_serial_link[21] ;
  wire \gpio_serial_link[22] ;
  wire \gpio_serial_link[23] ;
  wire \gpio_serial_link[24] ;
  wire \gpio_serial_link[25] ;
  wire \gpio_serial_link[26] ;
  wire \gpio_serial_link[27] ;
  wire \gpio_serial_link[28] ;
  wire \gpio_serial_link[29] ;
  wire \gpio_serial_link[2] ;
  wire \gpio_serial_link[30] ;
  wire \gpio_serial_link[31] ;
  wire \gpio_serial_link[32] ;
  wire \gpio_serial_link[33] ;
  wire \gpio_serial_link[34] ;
  wire \gpio_serial_link[35] ;
  wire \gpio_serial_link[36] ;
  wire \gpio_serial_link[37] ;
  wire \gpio_serial_link[3] ;
  wire \gpio_serial_link[4] ;
  wire \gpio_serial_link[5] ;
  wire \gpio_serial_link[6] ;
  wire \gpio_serial_link[7] ;
  wire \gpio_serial_link[8] ;
  wire \gpio_serial_link[9] ;
  wire \gpio_serial_link_shifted[0] ;
  wire \gpio_serial_link_shifted[10] ;
  wire \gpio_serial_link_shifted[11] ;
  wire \gpio_serial_link_shifted[12] ;
  wire \gpio_serial_link_shifted[13] ;
  wire \gpio_serial_link_shifted[14] ;
  wire \gpio_serial_link_shifted[15] ;
  wire \gpio_serial_link_shifted[16] ;
  wire \gpio_serial_link_shifted[17] ;
  wire \gpio_serial_link_shifted[18] ;
  wire \gpio_serial_link_shifted[19] ;
  wire \gpio_serial_link_shifted[1] ;
  wire \gpio_serial_link_shifted[20] ;
  wire \gpio_serial_link_shifted[21] ;
  wire \gpio_serial_link_shifted[22] ;
  wire \gpio_serial_link_shifted[23] ;
  wire \gpio_serial_link_shifted[24] ;
  wire \gpio_serial_link_shifted[25] ;
  wire \gpio_serial_link_shifted[26] ;
  wire \gpio_serial_link_shifted[27] ;
  wire \gpio_serial_link_shifted[28] ;
  wire \gpio_serial_link_shifted[29] ;
  wire \gpio_serial_link_shifted[2] ;
  wire \gpio_serial_link_shifted[30] ;
  wire \gpio_serial_link_shifted[31] ;
  wire \gpio_serial_link_shifted[32] ;
  wire \gpio_serial_link_shifted[33] ;
  wire \gpio_serial_link_shifted[34] ;
  wire \gpio_serial_link_shifted[35] ;
  wire \gpio_serial_link_shifted[36] ;
  wire \gpio_serial_link_shifted[37] ;
  wire \gpio_serial_link_shifted[3] ;
  wire \gpio_serial_link_shifted[4] ;
  wire \gpio_serial_link_shifted[5] ;
  wire \gpio_serial_link_shifted[6] ;
  wire \gpio_serial_link_shifted[7] ;
  wire \gpio_serial_link_shifted[8] ;
  wire \gpio_serial_link_shifted[9] ;
  wire jtag_out;
  wire jtag_outenb;
  wire \la_data_in_mprj[0] ;
  wire \la_data_in_mprj[100] ;
  wire \la_data_in_mprj[101] ;
  wire \la_data_in_mprj[102] ;
  wire \la_data_in_mprj[103] ;
  wire \la_data_in_mprj[104] ;
  wire \la_data_in_mprj[105] ;
  wire \la_data_in_mprj[106] ;
  wire \la_data_in_mprj[107] ;
  wire \la_data_in_mprj[108] ;
  wire \la_data_in_mprj[109] ;
  wire \la_data_in_mprj[10] ;
  wire \la_data_in_mprj[110] ;
  wire \la_data_in_mprj[111] ;
  wire \la_data_in_mprj[112] ;
  wire \la_data_in_mprj[113] ;
  wire \la_data_in_mprj[114] ;
  wire \la_data_in_mprj[115] ;
  wire \la_data_in_mprj[116] ;
  wire \la_data_in_mprj[117] ;
  wire \la_data_in_mprj[118] ;
  wire \la_data_in_mprj[119] ;
  wire \la_data_in_mprj[11] ;
  wire \la_data_in_mprj[120] ;
  wire \la_data_in_mprj[121] ;
  wire \la_data_in_mprj[122] ;
  wire \la_data_in_mprj[123] ;
  wire \la_data_in_mprj[124] ;
  wire \la_data_in_mprj[125] ;
  wire \la_data_in_mprj[126] ;
  wire \la_data_in_mprj[127] ;
  wire \la_data_in_mprj[12] ;
  wire \la_data_in_mprj[13] ;
  wire \la_data_in_mprj[14] ;
  wire \la_data_in_mprj[15] ;
  wire \la_data_in_mprj[16] ;
  wire \la_data_in_mprj[17] ;
  wire \la_data_in_mprj[18] ;
  wire \la_data_in_mprj[19] ;
  wire \la_data_in_mprj[1] ;
  wire \la_data_in_mprj[20] ;
  wire \la_data_in_mprj[21] ;
  wire \la_data_in_mprj[22] ;
  wire \la_data_in_mprj[23] ;
  wire \la_data_in_mprj[24] ;
  wire \la_data_in_mprj[25] ;
  wire \la_data_in_mprj[26] ;
  wire \la_data_in_mprj[27] ;
  wire \la_data_in_mprj[28] ;
  wire \la_data_in_mprj[29] ;
  wire \la_data_in_mprj[2] ;
  wire \la_data_in_mprj[30] ;
  wire \la_data_in_mprj[31] ;
  wire \la_data_in_mprj[32] ;
  wire \la_data_in_mprj[33] ;
  wire \la_data_in_mprj[34] ;
  wire \la_data_in_mprj[35] ;
  wire \la_data_in_mprj[36] ;
  wire \la_data_in_mprj[37] ;
  wire \la_data_in_mprj[38] ;
  wire \la_data_in_mprj[39] ;
  wire \la_data_in_mprj[3] ;
  wire \la_data_in_mprj[40] ;
  wire \la_data_in_mprj[41] ;
  wire \la_data_in_mprj[42] ;
  wire \la_data_in_mprj[43] ;
  wire \la_data_in_mprj[44] ;
  wire \la_data_in_mprj[45] ;
  wire \la_data_in_mprj[46] ;
  wire \la_data_in_mprj[47] ;
  wire \la_data_in_mprj[48] ;
  wire \la_data_in_mprj[49] ;
  wire \la_data_in_mprj[4] ;
  wire \la_data_in_mprj[50] ;
  wire \la_data_in_mprj[51] ;
  wire \la_data_in_mprj[52] ;
  wire \la_data_in_mprj[53] ;
  wire \la_data_in_mprj[54] ;
  wire \la_data_in_mprj[55] ;
  wire \la_data_in_mprj[56] ;
  wire \la_data_in_mprj[57] ;
  wire \la_data_in_mprj[58] ;
  wire \la_data_in_mprj[59] ;
  wire \la_data_in_mprj[5] ;
  wire \la_data_in_mprj[60] ;
  wire \la_data_in_mprj[61] ;
  wire \la_data_in_mprj[62] ;
  wire \la_data_in_mprj[63] ;
  wire \la_data_in_mprj[64] ;
  wire \la_data_in_mprj[65] ;
  wire \la_data_in_mprj[66] ;
  wire \la_data_in_mprj[67] ;
  wire \la_data_in_mprj[68] ;
  wire \la_data_in_mprj[69] ;
  wire \la_data_in_mprj[6] ;
  wire \la_data_in_mprj[70] ;
  wire \la_data_in_mprj[71] ;
  wire \la_data_in_mprj[72] ;
  wire \la_data_in_mprj[73] ;
  wire \la_data_in_mprj[74] ;
  wire \la_data_in_mprj[75] ;
  wire \la_data_in_mprj[76] ;
  wire \la_data_in_mprj[77] ;
  wire \la_data_in_mprj[78] ;
  wire \la_data_in_mprj[79] ;
  wire \la_data_in_mprj[7] ;
  wire \la_data_in_mprj[80] ;
  wire \la_data_in_mprj[81] ;
  wire \la_data_in_mprj[82] ;
  wire \la_data_in_mprj[83] ;
  wire \la_data_in_mprj[84] ;
  wire \la_data_in_mprj[85] ;
  wire \la_data_in_mprj[86] ;
  wire \la_data_in_mprj[87] ;
  wire \la_data_in_mprj[88] ;
  wire \la_data_in_mprj[89] ;
  wire \la_data_in_mprj[8] ;
  wire \la_data_in_mprj[90] ;
  wire \la_data_in_mprj[91] ;
  wire \la_data_in_mprj[92] ;
  wire \la_data_in_mprj[93] ;
  wire \la_data_in_mprj[94] ;
  wire \la_data_in_mprj[95] ;
  wire \la_data_in_mprj[96] ;
  wire \la_data_in_mprj[97] ;
  wire \la_data_in_mprj[98] ;
  wire \la_data_in_mprj[99] ;
  wire \la_data_in_mprj[9] ;
  wire \la_data_in_user[0] ;
  wire \la_data_in_user[100] ;
  wire \la_data_in_user[101] ;
  wire \la_data_in_user[102] ;
  wire \la_data_in_user[103] ;
  wire \la_data_in_user[104] ;
  wire \la_data_in_user[105] ;
  wire \la_data_in_user[106] ;
  wire \la_data_in_user[107] ;
  wire \la_data_in_user[108] ;
  wire \la_data_in_user[109] ;
  wire \la_data_in_user[10] ;
  wire \la_data_in_user[110] ;
  wire \la_data_in_user[111] ;
  wire \la_data_in_user[112] ;
  wire \la_data_in_user[113] ;
  wire \la_data_in_user[114] ;
  wire \la_data_in_user[115] ;
  wire \la_data_in_user[116] ;
  wire \la_data_in_user[117] ;
  wire \la_data_in_user[118] ;
  wire \la_data_in_user[119] ;
  wire \la_data_in_user[11] ;
  wire \la_data_in_user[120] ;
  wire \la_data_in_user[121] ;
  wire \la_data_in_user[122] ;
  wire \la_data_in_user[123] ;
  wire \la_data_in_user[124] ;
  wire \la_data_in_user[125] ;
  wire \la_data_in_user[126] ;
  wire \la_data_in_user[127] ;
  wire \la_data_in_user[12] ;
  wire \la_data_in_user[13] ;
  wire \la_data_in_user[14] ;
  wire \la_data_in_user[15] ;
  wire \la_data_in_user[16] ;
  wire \la_data_in_user[17] ;
  wire \la_data_in_user[18] ;
  wire \la_data_in_user[19] ;
  wire \la_data_in_user[1] ;
  wire \la_data_in_user[20] ;
  wire \la_data_in_user[21] ;
  wire \la_data_in_user[22] ;
  wire \la_data_in_user[23] ;
  wire \la_data_in_user[24] ;
  wire \la_data_in_user[25] ;
  wire \la_data_in_user[26] ;
  wire \la_data_in_user[27] ;
  wire \la_data_in_user[28] ;
  wire \la_data_in_user[29] ;
  wire \la_data_in_user[2] ;
  wire \la_data_in_user[30] ;
  wire \la_data_in_user[31] ;
  wire \la_data_in_user[32] ;
  wire \la_data_in_user[33] ;
  wire \la_data_in_user[34] ;
  wire \la_data_in_user[35] ;
  wire \la_data_in_user[36] ;
  wire \la_data_in_user[37] ;
  wire \la_data_in_user[38] ;
  wire \la_data_in_user[39] ;
  wire \la_data_in_user[3] ;
  wire \la_data_in_user[40] ;
  wire \la_data_in_user[41] ;
  wire \la_data_in_user[42] ;
  wire \la_data_in_user[43] ;
  wire \la_data_in_user[44] ;
  wire \la_data_in_user[45] ;
  wire \la_data_in_user[46] ;
  wire \la_data_in_user[47] ;
  wire \la_data_in_user[48] ;
  wire \la_data_in_user[49] ;
  wire \la_data_in_user[4] ;
  wire \la_data_in_user[50] ;
  wire \la_data_in_user[51] ;
  wire \la_data_in_user[52] ;
  wire \la_data_in_user[53] ;
  wire \la_data_in_user[54] ;
  wire \la_data_in_user[55] ;
  wire \la_data_in_user[56] ;
  wire \la_data_in_user[57] ;
  wire \la_data_in_user[58] ;
  wire \la_data_in_user[59] ;
  wire \la_data_in_user[5] ;
  wire \la_data_in_user[60] ;
  wire \la_data_in_user[61] ;
  wire \la_data_in_user[62] ;
  wire \la_data_in_user[63] ;
  wire \la_data_in_user[64] ;
  wire \la_data_in_user[65] ;
  wire \la_data_in_user[66] ;
  wire \la_data_in_user[67] ;
  wire \la_data_in_user[68] ;
  wire \la_data_in_user[69] ;
  wire \la_data_in_user[6] ;
  wire \la_data_in_user[70] ;
  wire \la_data_in_user[71] ;
  wire \la_data_in_user[72] ;
  wire \la_data_in_user[73] ;
  wire \la_data_in_user[74] ;
  wire \la_data_in_user[75] ;
  wire \la_data_in_user[76] ;
  wire \la_data_in_user[77] ;
  wire \la_data_in_user[78] ;
  wire \la_data_in_user[79] ;
  wire \la_data_in_user[7] ;
  wire \la_data_in_user[80] ;
  wire \la_data_in_user[81] ;
  wire \la_data_in_user[82] ;
  wire \la_data_in_user[83] ;
  wire \la_data_in_user[84] ;
  wire \la_data_in_user[85] ;
  wire \la_data_in_user[86] ;
  wire \la_data_in_user[87] ;
  wire \la_data_in_user[88] ;
  wire \la_data_in_user[89] ;
  wire \la_data_in_user[8] ;
  wire \la_data_in_user[90] ;
  wire \la_data_in_user[91] ;
  wire \la_data_in_user[92] ;
  wire \la_data_in_user[93] ;
  wire \la_data_in_user[94] ;
  wire \la_data_in_user[95] ;
  wire \la_data_in_user[96] ;
  wire \la_data_in_user[97] ;
  wire \la_data_in_user[98] ;
  wire \la_data_in_user[99] ;
  wire \la_data_in_user[9] ;
  wire \la_data_out_mprj[0] ;
  wire \la_data_out_mprj[100] ;
  wire \la_data_out_mprj[101] ;
  wire \la_data_out_mprj[102] ;
  wire \la_data_out_mprj[103] ;
  wire \la_data_out_mprj[104] ;
  wire \la_data_out_mprj[105] ;
  wire \la_data_out_mprj[106] ;
  wire \la_data_out_mprj[107] ;
  wire \la_data_out_mprj[108] ;
  wire \la_data_out_mprj[109] ;
  wire \la_data_out_mprj[10] ;
  wire \la_data_out_mprj[110] ;
  wire \la_data_out_mprj[111] ;
  wire \la_data_out_mprj[112] ;
  wire \la_data_out_mprj[113] ;
  wire \la_data_out_mprj[114] ;
  wire \la_data_out_mprj[115] ;
  wire \la_data_out_mprj[116] ;
  wire \la_data_out_mprj[117] ;
  wire \la_data_out_mprj[118] ;
  wire \la_data_out_mprj[119] ;
  wire \la_data_out_mprj[11] ;
  wire \la_data_out_mprj[120] ;
  wire \la_data_out_mprj[121] ;
  wire \la_data_out_mprj[122] ;
  wire \la_data_out_mprj[123] ;
  wire \la_data_out_mprj[124] ;
  wire \la_data_out_mprj[125] ;
  wire \la_data_out_mprj[126] ;
  wire \la_data_out_mprj[127] ;
  wire \la_data_out_mprj[12] ;
  wire \la_data_out_mprj[13] ;
  wire \la_data_out_mprj[14] ;
  wire \la_data_out_mprj[15] ;
  wire \la_data_out_mprj[16] ;
  wire \la_data_out_mprj[17] ;
  wire \la_data_out_mprj[18] ;
  wire \la_data_out_mprj[19] ;
  wire \la_data_out_mprj[1] ;
  wire \la_data_out_mprj[20] ;
  wire \la_data_out_mprj[21] ;
  wire \la_data_out_mprj[22] ;
  wire \la_data_out_mprj[23] ;
  wire \la_data_out_mprj[24] ;
  wire \la_data_out_mprj[25] ;
  wire \la_data_out_mprj[26] ;
  wire \la_data_out_mprj[27] ;
  wire \la_data_out_mprj[28] ;
  wire \la_data_out_mprj[29] ;
  wire \la_data_out_mprj[2] ;
  wire \la_data_out_mprj[30] ;
  wire \la_data_out_mprj[31] ;
  wire \la_data_out_mprj[32] ;
  wire \la_data_out_mprj[33] ;
  wire \la_data_out_mprj[34] ;
  wire \la_data_out_mprj[35] ;
  wire \la_data_out_mprj[36] ;
  wire \la_data_out_mprj[37] ;
  wire \la_data_out_mprj[38] ;
  wire \la_data_out_mprj[39] ;
  wire \la_data_out_mprj[3] ;
  wire \la_data_out_mprj[40] ;
  wire \la_data_out_mprj[41] ;
  wire \la_data_out_mprj[42] ;
  wire \la_data_out_mprj[43] ;
  wire \la_data_out_mprj[44] ;
  wire \la_data_out_mprj[45] ;
  wire \la_data_out_mprj[46] ;
  wire \la_data_out_mprj[47] ;
  wire \la_data_out_mprj[48] ;
  wire \la_data_out_mprj[49] ;
  wire \la_data_out_mprj[4] ;
  wire \la_data_out_mprj[50] ;
  wire \la_data_out_mprj[51] ;
  wire \la_data_out_mprj[52] ;
  wire \la_data_out_mprj[53] ;
  wire \la_data_out_mprj[54] ;
  wire \la_data_out_mprj[55] ;
  wire \la_data_out_mprj[56] ;
  wire \la_data_out_mprj[57] ;
  wire \la_data_out_mprj[58] ;
  wire \la_data_out_mprj[59] ;
  wire \la_data_out_mprj[5] ;
  wire \la_data_out_mprj[60] ;
  wire \la_data_out_mprj[61] ;
  wire \la_data_out_mprj[62] ;
  wire \la_data_out_mprj[63] ;
  wire \la_data_out_mprj[64] ;
  wire \la_data_out_mprj[65] ;
  wire \la_data_out_mprj[66] ;
  wire \la_data_out_mprj[67] ;
  wire \la_data_out_mprj[68] ;
  wire \la_data_out_mprj[69] ;
  wire \la_data_out_mprj[6] ;
  wire \la_data_out_mprj[70] ;
  wire \la_data_out_mprj[71] ;
  wire \la_data_out_mprj[72] ;
  wire \la_data_out_mprj[73] ;
  wire \la_data_out_mprj[74] ;
  wire \la_data_out_mprj[75] ;
  wire \la_data_out_mprj[76] ;
  wire \la_data_out_mprj[77] ;
  wire \la_data_out_mprj[78] ;
  wire \la_data_out_mprj[79] ;
  wire \la_data_out_mprj[7] ;
  wire \la_data_out_mprj[80] ;
  wire \la_data_out_mprj[81] ;
  wire \la_data_out_mprj[82] ;
  wire \la_data_out_mprj[83] ;
  wire \la_data_out_mprj[84] ;
  wire \la_data_out_mprj[85] ;
  wire \la_data_out_mprj[86] ;
  wire \la_data_out_mprj[87] ;
  wire \la_data_out_mprj[88] ;
  wire \la_data_out_mprj[89] ;
  wire \la_data_out_mprj[8] ;
  wire \la_data_out_mprj[90] ;
  wire \la_data_out_mprj[91] ;
  wire \la_data_out_mprj[92] ;
  wire \la_data_out_mprj[93] ;
  wire \la_data_out_mprj[94] ;
  wire \la_data_out_mprj[95] ;
  wire \la_data_out_mprj[96] ;
  wire \la_data_out_mprj[97] ;
  wire \la_data_out_mprj[98] ;
  wire \la_data_out_mprj[99] ;
  wire \la_data_out_mprj[9] ;
  wire \la_data_out_user[0] ;
  wire \la_data_out_user[100] ;
  wire \la_data_out_user[101] ;
  wire \la_data_out_user[102] ;
  wire \la_data_out_user[103] ;
  wire \la_data_out_user[104] ;
  wire \la_data_out_user[105] ;
  wire \la_data_out_user[106] ;
  wire \la_data_out_user[107] ;
  wire \la_data_out_user[108] ;
  wire \la_data_out_user[109] ;
  wire \la_data_out_user[10] ;
  wire \la_data_out_user[110] ;
  wire \la_data_out_user[111] ;
  wire \la_data_out_user[112] ;
  wire \la_data_out_user[113] ;
  wire \la_data_out_user[114] ;
  wire \la_data_out_user[115] ;
  wire \la_data_out_user[116] ;
  wire \la_data_out_user[117] ;
  wire \la_data_out_user[118] ;
  wire \la_data_out_user[119] ;
  wire \la_data_out_user[11] ;
  wire \la_data_out_user[120] ;
  wire \la_data_out_user[121] ;
  wire \la_data_out_user[122] ;
  wire \la_data_out_user[123] ;
  wire \la_data_out_user[124] ;
  wire \la_data_out_user[125] ;
  wire \la_data_out_user[126] ;
  wire \la_data_out_user[127] ;
  wire \la_data_out_user[12] ;
  wire \la_data_out_user[13] ;
  wire \la_data_out_user[14] ;
  wire \la_data_out_user[15] ;
  wire \la_data_out_user[16] ;
  wire \la_data_out_user[17] ;
  wire \la_data_out_user[18] ;
  wire \la_data_out_user[19] ;
  wire \la_data_out_user[1] ;
  wire \la_data_out_user[20] ;
  wire \la_data_out_user[21] ;
  wire \la_data_out_user[22] ;
  wire \la_data_out_user[23] ;
  wire \la_data_out_user[24] ;
  wire \la_data_out_user[25] ;
  wire \la_data_out_user[26] ;
  wire \la_data_out_user[27] ;
  wire \la_data_out_user[28] ;
  wire \la_data_out_user[29] ;
  wire \la_data_out_user[2] ;
  wire \la_data_out_user[30] ;
  wire \la_data_out_user[31] ;
  wire \la_data_out_user[32] ;
  wire \la_data_out_user[33] ;
  wire \la_data_out_user[34] ;
  wire \la_data_out_user[35] ;
  wire \la_data_out_user[36] ;
  wire \la_data_out_user[37] ;
  wire \la_data_out_user[38] ;
  wire \la_data_out_user[39] ;
  wire \la_data_out_user[3] ;
  wire \la_data_out_user[40] ;
  wire \la_data_out_user[41] ;
  wire \la_data_out_user[42] ;
  wire \la_data_out_user[43] ;
  wire \la_data_out_user[44] ;
  wire \la_data_out_user[45] ;
  wire \la_data_out_user[46] ;
  wire \la_data_out_user[47] ;
  wire \la_data_out_user[48] ;
  wire \la_data_out_user[49] ;
  wire \la_data_out_user[4] ;
  wire \la_data_out_user[50] ;
  wire \la_data_out_user[51] ;
  wire \la_data_out_user[52] ;
  wire \la_data_out_user[53] ;
  wire \la_data_out_user[54] ;
  wire \la_data_out_user[55] ;
  wire \la_data_out_user[56] ;
  wire \la_data_out_user[57] ;
  wire \la_data_out_user[58] ;
  wire \la_data_out_user[59] ;
  wire \la_data_out_user[5] ;
  wire \la_data_out_user[60] ;
  wire \la_data_out_user[61] ;
  wire \la_data_out_user[62] ;
  wire \la_data_out_user[63] ;
  wire \la_data_out_user[64] ;
  wire \la_data_out_user[65] ;
  wire \la_data_out_user[66] ;
  wire \la_data_out_user[67] ;
  wire \la_data_out_user[68] ;
  wire \la_data_out_user[69] ;
  wire \la_data_out_user[6] ;
  wire \la_data_out_user[70] ;
  wire \la_data_out_user[71] ;
  wire \la_data_out_user[72] ;
  wire \la_data_out_user[73] ;
  wire \la_data_out_user[74] ;
  wire \la_data_out_user[75] ;
  wire \la_data_out_user[76] ;
  wire \la_data_out_user[77] ;
  wire \la_data_out_user[78] ;
  wire \la_data_out_user[79] ;
  wire \la_data_out_user[7] ;
  wire \la_data_out_user[80] ;
  wire \la_data_out_user[81] ;
  wire \la_data_out_user[82] ;
  wire \la_data_out_user[83] ;
  wire \la_data_out_user[84] ;
  wire \la_data_out_user[85] ;
  wire \la_data_out_user[86] ;
  wire \la_data_out_user[87] ;
  wire \la_data_out_user[88] ;
  wire \la_data_out_user[89] ;
  wire \la_data_out_user[8] ;
  wire \la_data_out_user[90] ;
  wire \la_data_out_user[91] ;
  wire \la_data_out_user[92] ;
  wire \la_data_out_user[93] ;
  wire \la_data_out_user[94] ;
  wire \la_data_out_user[95] ;
  wire \la_data_out_user[96] ;
  wire \la_data_out_user[97] ;
  wire \la_data_out_user[98] ;
  wire \la_data_out_user[99] ;
  wire \la_data_out_user[9] ;
  wire \la_oen_mprj[0] ;
  wire \la_oen_mprj[100] ;
  wire \la_oen_mprj[101] ;
  wire \la_oen_mprj[102] ;
  wire \la_oen_mprj[103] ;
  wire \la_oen_mprj[104] ;
  wire \la_oen_mprj[105] ;
  wire \la_oen_mprj[106] ;
  wire \la_oen_mprj[107] ;
  wire \la_oen_mprj[108] ;
  wire \la_oen_mprj[109] ;
  wire \la_oen_mprj[10] ;
  wire \la_oen_mprj[110] ;
  wire \la_oen_mprj[111] ;
  wire \la_oen_mprj[112] ;
  wire \la_oen_mprj[113] ;
  wire \la_oen_mprj[114] ;
  wire \la_oen_mprj[115] ;
  wire \la_oen_mprj[116] ;
  wire \la_oen_mprj[117] ;
  wire \la_oen_mprj[118] ;
  wire \la_oen_mprj[119] ;
  wire \la_oen_mprj[11] ;
  wire \la_oen_mprj[120] ;
  wire \la_oen_mprj[121] ;
  wire \la_oen_mprj[122] ;
  wire \la_oen_mprj[123] ;
  wire \la_oen_mprj[124] ;
  wire \la_oen_mprj[125] ;
  wire \la_oen_mprj[126] ;
  wire \la_oen_mprj[127] ;
  wire \la_oen_mprj[12] ;
  wire \la_oen_mprj[13] ;
  wire \la_oen_mprj[14] ;
  wire \la_oen_mprj[15] ;
  wire \la_oen_mprj[16] ;
  wire \la_oen_mprj[17] ;
  wire \la_oen_mprj[18] ;
  wire \la_oen_mprj[19] ;
  wire \la_oen_mprj[1] ;
  wire \la_oen_mprj[20] ;
  wire \la_oen_mprj[21] ;
  wire \la_oen_mprj[22] ;
  wire \la_oen_mprj[23] ;
  wire \la_oen_mprj[24] ;
  wire \la_oen_mprj[25] ;
  wire \la_oen_mprj[26] ;
  wire \la_oen_mprj[27] ;
  wire \la_oen_mprj[28] ;
  wire \la_oen_mprj[29] ;
  wire \la_oen_mprj[2] ;
  wire \la_oen_mprj[30] ;
  wire \la_oen_mprj[31] ;
  wire \la_oen_mprj[32] ;
  wire \la_oen_mprj[33] ;
  wire \la_oen_mprj[34] ;
  wire \la_oen_mprj[35] ;
  wire \la_oen_mprj[36] ;
  wire \la_oen_mprj[37] ;
  wire \la_oen_mprj[38] ;
  wire \la_oen_mprj[39] ;
  wire \la_oen_mprj[3] ;
  wire \la_oen_mprj[40] ;
  wire \la_oen_mprj[41] ;
  wire \la_oen_mprj[42] ;
  wire \la_oen_mprj[43] ;
  wire \la_oen_mprj[44] ;
  wire \la_oen_mprj[45] ;
  wire \la_oen_mprj[46] ;
  wire \la_oen_mprj[47] ;
  wire \la_oen_mprj[48] ;
  wire \la_oen_mprj[49] ;
  wire \la_oen_mprj[4] ;
  wire \la_oen_mprj[50] ;
  wire \la_oen_mprj[51] ;
  wire \la_oen_mprj[52] ;
  wire \la_oen_mprj[53] ;
  wire \la_oen_mprj[54] ;
  wire \la_oen_mprj[55] ;
  wire \la_oen_mprj[56] ;
  wire \la_oen_mprj[57] ;
  wire \la_oen_mprj[58] ;
  wire \la_oen_mprj[59] ;
  wire \la_oen_mprj[5] ;
  wire \la_oen_mprj[60] ;
  wire \la_oen_mprj[61] ;
  wire \la_oen_mprj[62] ;
  wire \la_oen_mprj[63] ;
  wire \la_oen_mprj[64] ;
  wire \la_oen_mprj[65] ;
  wire \la_oen_mprj[66] ;
  wire \la_oen_mprj[67] ;
  wire \la_oen_mprj[68] ;
  wire \la_oen_mprj[69] ;
  wire \la_oen_mprj[6] ;
  wire \la_oen_mprj[70] ;
  wire \la_oen_mprj[71] ;
  wire \la_oen_mprj[72] ;
  wire \la_oen_mprj[73] ;
  wire \la_oen_mprj[74] ;
  wire \la_oen_mprj[75] ;
  wire \la_oen_mprj[76] ;
  wire \la_oen_mprj[77] ;
  wire \la_oen_mprj[78] ;
  wire \la_oen_mprj[79] ;
  wire \la_oen_mprj[7] ;
  wire \la_oen_mprj[80] ;
  wire \la_oen_mprj[81] ;
  wire \la_oen_mprj[82] ;
  wire \la_oen_mprj[83] ;
  wire \la_oen_mprj[84] ;
  wire \la_oen_mprj[85] ;
  wire \la_oen_mprj[86] ;
  wire \la_oen_mprj[87] ;
  wire \la_oen_mprj[88] ;
  wire \la_oen_mprj[89] ;
  wire \la_oen_mprj[8] ;
  wire \la_oen_mprj[90] ;
  wire \la_oen_mprj[91] ;
  wire \la_oen_mprj[92] ;
  wire \la_oen_mprj[93] ;
  wire \la_oen_mprj[94] ;
  wire \la_oen_mprj[95] ;
  wire \la_oen_mprj[96] ;
  wire \la_oen_mprj[97] ;
  wire \la_oen_mprj[98] ;
  wire \la_oen_mprj[99] ;
  wire \la_oen_mprj[9] ;
  wire \la_oen_user[0] ;
  wire \la_oen_user[100] ;
  wire \la_oen_user[101] ;
  wire \la_oen_user[102] ;
  wire \la_oen_user[103] ;
  wire \la_oen_user[104] ;
  wire \la_oen_user[105] ;
  wire \la_oen_user[106] ;
  wire \la_oen_user[107] ;
  wire \la_oen_user[108] ;
  wire \la_oen_user[109] ;
  wire \la_oen_user[10] ;
  wire \la_oen_user[110] ;
  wire \la_oen_user[111] ;
  wire \la_oen_user[112] ;
  wire \la_oen_user[113] ;
  wire \la_oen_user[114] ;
  wire \la_oen_user[115] ;
  wire \la_oen_user[116] ;
  wire \la_oen_user[117] ;
  wire \la_oen_user[118] ;
  wire \la_oen_user[119] ;
  wire \la_oen_user[11] ;
  wire \la_oen_user[120] ;
  wire \la_oen_user[121] ;
  wire \la_oen_user[122] ;
  wire \la_oen_user[123] ;
  wire \la_oen_user[124] ;
  wire \la_oen_user[125] ;
  wire \la_oen_user[126] ;
  wire \la_oen_user[127] ;
  wire \la_oen_user[12] ;
  wire \la_oen_user[13] ;
  wire \la_oen_user[14] ;
  wire \la_oen_user[15] ;
  wire \la_oen_user[16] ;
  wire \la_oen_user[17] ;
  wire \la_oen_user[18] ;
  wire \la_oen_user[19] ;
  wire \la_oen_user[1] ;
  wire \la_oen_user[20] ;
  wire \la_oen_user[21] ;
  wire \la_oen_user[22] ;
  wire \la_oen_user[23] ;
  wire \la_oen_user[24] ;
  wire \la_oen_user[25] ;
  wire \la_oen_user[26] ;
  wire \la_oen_user[27] ;
  wire \la_oen_user[28] ;
  wire \la_oen_user[29] ;
  wire \la_oen_user[2] ;
  wire \la_oen_user[30] ;
  wire \la_oen_user[31] ;
  wire \la_oen_user[32] ;
  wire \la_oen_user[33] ;
  wire \la_oen_user[34] ;
  wire \la_oen_user[35] ;
  wire \la_oen_user[36] ;
  wire \la_oen_user[37] ;
  wire \la_oen_user[38] ;
  wire \la_oen_user[39] ;
  wire \la_oen_user[3] ;
  wire \la_oen_user[40] ;
  wire \la_oen_user[41] ;
  wire \la_oen_user[42] ;
  wire \la_oen_user[43] ;
  wire \la_oen_user[44] ;
  wire \la_oen_user[45] ;
  wire \la_oen_user[46] ;
  wire \la_oen_user[47] ;
  wire \la_oen_user[48] ;
  wire \la_oen_user[49] ;
  wire \la_oen_user[4] ;
  wire \la_oen_user[50] ;
  wire \la_oen_user[51] ;
  wire \la_oen_user[52] ;
  wire \la_oen_user[53] ;
  wire \la_oen_user[54] ;
  wire \la_oen_user[55] ;
  wire \la_oen_user[56] ;
  wire \la_oen_user[57] ;
  wire \la_oen_user[58] ;
  wire \la_oen_user[59] ;
  wire \la_oen_user[5] ;
  wire \la_oen_user[60] ;
  wire \la_oen_user[61] ;
  wire \la_oen_user[62] ;
  wire \la_oen_user[63] ;
  wire \la_oen_user[64] ;
  wire \la_oen_user[65] ;
  wire \la_oen_user[66] ;
  wire \la_oen_user[67] ;
  wire \la_oen_user[68] ;
  wire \la_oen_user[69] ;
  wire \la_oen_user[6] ;
  wire \la_oen_user[70] ;
  wire \la_oen_user[71] ;
  wire \la_oen_user[72] ;
  wire \la_oen_user[73] ;
  wire \la_oen_user[74] ;
  wire \la_oen_user[75] ;
  wire \la_oen_user[76] ;
  wire \la_oen_user[77] ;
  wire \la_oen_user[78] ;
  wire \la_oen_user[79] ;
  wire \la_oen_user[7] ;
  wire \la_oen_user[80] ;
  wire \la_oen_user[81] ;
  wire \la_oen_user[82] ;
  wire \la_oen_user[83] ;
  wire \la_oen_user[84] ;
  wire \la_oen_user[85] ;
  wire \la_oen_user[86] ;
  wire \la_oen_user[87] ;
  wire \la_oen_user[88] ;
  wire \la_oen_user[89] ;
  wire \la_oen_user[8] ;
  wire \la_oen_user[90] ;
  wire \la_oen_user[91] ;
  wire \la_oen_user[92] ;
  wire \la_oen_user[93] ;
  wire \la_oen_user[94] ;
  wire \la_oen_user[95] ;
  wire \la_oen_user[96] ;
  wire \la_oen_user[97] ;
  wire \la_oen_user[98] ;
  wire \la_oen_user[99] ;
  wire \la_oen_user[9] ;
  wire \mask_rev[0] ;
  wire \mask_rev[10] ;
  wire \mask_rev[11] ;
  wire \mask_rev[12] ;
  wire \mask_rev[13] ;
  wire \mask_rev[14] ;
  wire \mask_rev[15] ;
  wire \mask_rev[16] ;
  wire \mask_rev[17] ;
  wire \mask_rev[18] ;
  wire \mask_rev[19] ;
  wire \mask_rev[1] ;
  wire \mask_rev[20] ;
  wire \mask_rev[21] ;
  wire \mask_rev[22] ;
  wire \mask_rev[23] ;
  wire \mask_rev[24] ;
  wire \mask_rev[25] ;
  wire \mask_rev[26] ;
  wire \mask_rev[27] ;
  wire \mask_rev[28] ;
  wire \mask_rev[29] ;
  wire \mask_rev[2] ;
  wire \mask_rev[30] ;
  wire \mask_rev[31] ;
  wire \mask_rev[3] ;
  wire \mask_rev[4] ;
  wire \mask_rev[5] ;
  wire \mask_rev[6] ;
  wire \mask_rev[7] ;
  wire \mask_rev[8] ;
  wire \mask_rev[9] ;
  wire \mgmt_addr[0] ;
  wire \mgmt_addr[1] ;
  wire \mgmt_addr[2] ;
  wire \mgmt_addr[3] ;
  wire \mgmt_addr[4] ;
  wire \mgmt_addr[5] ;
  wire \mgmt_addr[6] ;
  wire \mgmt_addr[7] ;
  wire \mgmt_addr_ro[0] ;
  wire \mgmt_addr_ro[1] ;
  wire \mgmt_addr_ro[2] ;
  wire \mgmt_addr_ro[3] ;
  wire \mgmt_addr_ro[4] ;
  wire \mgmt_addr_ro[5] ;
  wire \mgmt_addr_ro[6] ;
  wire \mgmt_addr_ro[7] ;
  wire \mgmt_ena[0] ;
  wire \mgmt_ena[1] ;
  wire mgmt_ena_ro;
  wire \mgmt_io_in[0] ;
  wire \mgmt_io_in[10] ;
  wire \mgmt_io_in[11] ;
  wire \mgmt_io_in[12] ;
  wire \mgmt_io_in[13] ;
  wire \mgmt_io_in[14] ;
  wire \mgmt_io_in[15] ;
  wire \mgmt_io_in[16] ;
  wire \mgmt_io_in[17] ;
  wire \mgmt_io_in[18] ;
  wire \mgmt_io_in[19] ;
  wire \mgmt_io_in[1] ;
  wire \mgmt_io_in[20] ;
  wire \mgmt_io_in[21] ;
  wire \mgmt_io_in[22] ;
  wire \mgmt_io_in[23] ;
  wire \mgmt_io_in[24] ;
  wire \mgmt_io_in[25] ;
  wire \mgmt_io_in[26] ;
  wire \mgmt_io_in[27] ;
  wire \mgmt_io_in[28] ;
  wire \mgmt_io_in[29] ;
  wire \mgmt_io_in[2] ;
  wire \mgmt_io_in[30] ;
  wire \mgmt_io_in[31] ;
  wire \mgmt_io_in[32] ;
  wire \mgmt_io_in[33] ;
  wire \mgmt_io_in[34] ;
  wire \mgmt_io_in[35] ;
  wire \mgmt_io_in[36] ;
  wire \mgmt_io_in[37] ;
  wire \mgmt_io_in[3] ;
  wire \mgmt_io_in[4] ;
  wire \mgmt_io_in[5] ;
  wire \mgmt_io_in[6] ;
  wire \mgmt_io_in[7] ;
  wire \mgmt_io_in[8] ;
  wire \mgmt_io_in[9] ;
  wire \mgmt_io_nc1[0] ;
  wire \mgmt_io_nc1[10] ;
  wire \mgmt_io_nc1[11] ;
  wire \mgmt_io_nc1[12] ;
  wire \mgmt_io_nc1[13] ;
  wire \mgmt_io_nc1[14] ;
  wire \mgmt_io_nc1[15] ;
  wire \mgmt_io_nc1[16] ;
  wire \mgmt_io_nc1[17] ;
  wire \mgmt_io_nc1[18] ;
  wire \mgmt_io_nc1[19] ;
  wire \mgmt_io_nc1[1] ;
  wire \mgmt_io_nc1[20] ;
  wire \mgmt_io_nc1[21] ;
  wire \mgmt_io_nc1[22] ;
  wire \mgmt_io_nc1[23] ;
  wire \mgmt_io_nc1[24] ;
  wire \mgmt_io_nc1[25] ;
  wire \mgmt_io_nc1[26] ;
  wire \mgmt_io_nc1[27] ;
  wire \mgmt_io_nc1[28] ;
  wire \mgmt_io_nc1[29] ;
  wire \mgmt_io_nc1[2] ;
  wire \mgmt_io_nc1[30] ;
  wire \mgmt_io_nc1[31] ;
  wire \mgmt_io_nc1[32] ;
  wire \mgmt_io_nc1[33] ;
  wire \mgmt_io_nc1[34] ;
  wire \mgmt_io_nc1[35] ;
  wire \mgmt_io_nc1[3] ;
  wire \mgmt_io_nc1[4] ;
  wire \mgmt_io_nc1[5] ;
  wire \mgmt_io_nc1[6] ;
  wire \mgmt_io_nc1[7] ;
  wire \mgmt_io_nc1[8] ;
  wire \mgmt_io_nc1[9] ;
  wire \mgmt_io_nc2[0] ;
  wire \mgmt_io_nc2[1] ;
  wire \mgmt_io_nc3[0] ;
  wire \mgmt_io_nc3[10] ;
  wire \mgmt_io_nc3[11] ;
  wire \mgmt_io_nc3[12] ;
  wire \mgmt_io_nc3[13] ;
  wire \mgmt_io_nc3[14] ;
  wire \mgmt_io_nc3[15] ;
  wire \mgmt_io_nc3[16] ;
  wire \mgmt_io_nc3[17] ;
  wire \mgmt_io_nc3[18] ;
  wire \mgmt_io_nc3[19] ;
  wire \mgmt_io_nc3[1] ;
  wire \mgmt_io_nc3[20] ;
  wire \mgmt_io_nc3[21] ;
  wire \mgmt_io_nc3[22] ;
  wire \mgmt_io_nc3[23] ;
  wire \mgmt_io_nc3[24] ;
  wire \mgmt_io_nc3[25] ;
  wire \mgmt_io_nc3[26] ;
  wire \mgmt_io_nc3[27] ;
  wire \mgmt_io_nc3[28] ;
  wire \mgmt_io_nc3[29] ;
  wire \mgmt_io_nc3[2] ;
  wire \mgmt_io_nc3[30] ;
  wire \mgmt_io_nc3[31] ;
  wire \mgmt_io_nc3[32] ;
  wire \mgmt_io_nc3[33] ;
  wire \mgmt_io_nc3[34] ;
  wire \mgmt_io_nc3[35] ;
  wire \mgmt_io_nc3[3] ;
  wire \mgmt_io_nc3[4] ;
  wire \mgmt_io_nc3[5] ;
  wire \mgmt_io_nc3[6] ;
  wire \mgmt_io_nc3[7] ;
  wire \mgmt_io_nc3[8] ;
  wire \mgmt_io_nc3[9] ;
  wire \mgmt_rdata[0] ;
  wire \mgmt_rdata[10] ;
  wire \mgmt_rdata[11] ;
  wire \mgmt_rdata[12] ;
  wire \mgmt_rdata[13] ;
  wire \mgmt_rdata[14] ;
  wire \mgmt_rdata[15] ;
  wire \mgmt_rdata[16] ;
  wire \mgmt_rdata[17] ;
  wire \mgmt_rdata[18] ;
  wire \mgmt_rdata[19] ;
  wire \mgmt_rdata[1] ;
  wire \mgmt_rdata[20] ;
  wire \mgmt_rdata[21] ;
  wire \mgmt_rdata[22] ;
  wire \mgmt_rdata[23] ;
  wire \mgmt_rdata[24] ;
  wire \mgmt_rdata[25] ;
  wire \mgmt_rdata[26] ;
  wire \mgmt_rdata[27] ;
  wire \mgmt_rdata[28] ;
  wire \mgmt_rdata[29] ;
  wire \mgmt_rdata[2] ;
  wire \mgmt_rdata[30] ;
  wire \mgmt_rdata[31] ;
  wire \mgmt_rdata[32] ;
  wire \mgmt_rdata[33] ;
  wire \mgmt_rdata[34] ;
  wire \mgmt_rdata[35] ;
  wire \mgmt_rdata[36] ;
  wire \mgmt_rdata[37] ;
  wire \mgmt_rdata[38] ;
  wire \mgmt_rdata[39] ;
  wire \mgmt_rdata[3] ;
  wire \mgmt_rdata[40] ;
  wire \mgmt_rdata[41] ;
  wire \mgmt_rdata[42] ;
  wire \mgmt_rdata[43] ;
  wire \mgmt_rdata[44] ;
  wire \mgmt_rdata[45] ;
  wire \mgmt_rdata[46] ;
  wire \mgmt_rdata[47] ;
  wire \mgmt_rdata[48] ;
  wire \mgmt_rdata[49] ;
  wire \mgmt_rdata[4] ;
  wire \mgmt_rdata[50] ;
  wire \mgmt_rdata[51] ;
  wire \mgmt_rdata[52] ;
  wire \mgmt_rdata[53] ;
  wire \mgmt_rdata[54] ;
  wire \mgmt_rdata[55] ;
  wire \mgmt_rdata[56] ;
  wire \mgmt_rdata[57] ;
  wire \mgmt_rdata[58] ;
  wire \mgmt_rdata[59] ;
  wire \mgmt_rdata[5] ;
  wire \mgmt_rdata[60] ;
  wire \mgmt_rdata[61] ;
  wire \mgmt_rdata[62] ;
  wire \mgmt_rdata[63] ;
  wire \mgmt_rdata[6] ;
  wire \mgmt_rdata[7] ;
  wire \mgmt_rdata[8] ;
  wire \mgmt_rdata[9] ;
  wire \mgmt_rdata_ro[0] ;
  wire \mgmt_rdata_ro[10] ;
  wire \mgmt_rdata_ro[11] ;
  wire \mgmt_rdata_ro[12] ;
  wire \mgmt_rdata_ro[13] ;
  wire \mgmt_rdata_ro[14] ;
  wire \mgmt_rdata_ro[15] ;
  wire \mgmt_rdata_ro[16] ;
  wire \mgmt_rdata_ro[17] ;
  wire \mgmt_rdata_ro[18] ;
  wire \mgmt_rdata_ro[19] ;
  wire \mgmt_rdata_ro[1] ;
  wire \mgmt_rdata_ro[20] ;
  wire \mgmt_rdata_ro[21] ;
  wire \mgmt_rdata_ro[22] ;
  wire \mgmt_rdata_ro[23] ;
  wire \mgmt_rdata_ro[24] ;
  wire \mgmt_rdata_ro[25] ;
  wire \mgmt_rdata_ro[26] ;
  wire \mgmt_rdata_ro[27] ;
  wire \mgmt_rdata_ro[28] ;
  wire \mgmt_rdata_ro[29] ;
  wire \mgmt_rdata_ro[2] ;
  wire \mgmt_rdata_ro[30] ;
  wire \mgmt_rdata_ro[31] ;
  wire \mgmt_rdata_ro[3] ;
  wire \mgmt_rdata_ro[4] ;
  wire \mgmt_rdata_ro[5] ;
  wire \mgmt_rdata_ro[6] ;
  wire \mgmt_rdata_ro[7] ;
  wire \mgmt_rdata_ro[8] ;
  wire \mgmt_rdata_ro[9] ;
  wire mgmt_serial_clock;
  wire mgmt_serial_resetn;
  wire \mgmt_wdata[0] ;
  wire \mgmt_wdata[10] ;
  wire \mgmt_wdata[11] ;
  wire \mgmt_wdata[12] ;
  wire \mgmt_wdata[13] ;
  wire \mgmt_wdata[14] ;
  wire \mgmt_wdata[15] ;
  wire \mgmt_wdata[16] ;
  wire \mgmt_wdata[17] ;
  wire \mgmt_wdata[18] ;
  wire \mgmt_wdata[19] ;
  wire \mgmt_wdata[1] ;
  wire \mgmt_wdata[20] ;
  wire \mgmt_wdata[21] ;
  wire \mgmt_wdata[22] ;
  wire \mgmt_wdata[23] ;
  wire \mgmt_wdata[24] ;
  wire \mgmt_wdata[25] ;
  wire \mgmt_wdata[26] ;
  wire \mgmt_wdata[27] ;
  wire \mgmt_wdata[28] ;
  wire \mgmt_wdata[29] ;
  wire \mgmt_wdata[2] ;
  wire \mgmt_wdata[30] ;
  wire \mgmt_wdata[31] ;
  wire \mgmt_wdata[3] ;
  wire \mgmt_wdata[4] ;
  wire \mgmt_wdata[5] ;
  wire \mgmt_wdata[6] ;
  wire \mgmt_wdata[7] ;
  wire \mgmt_wdata[8] ;
  wire \mgmt_wdata[9] ;
  wire \mgmt_wen[0] ;
  wire \mgmt_wen[1] ;
  wire \mgmt_wen_mask[0] ;
  wire \mgmt_wen_mask[1] ;
  wire \mgmt_wen_mask[2] ;
  wire \mgmt_wen_mask[3] ;
  wire \mgmt_wen_mask[4] ;
  wire \mgmt_wen_mask[5] ;
  wire \mgmt_wen_mask[6] ;
  wire \mgmt_wen_mask[7] ;
  wire mprj2_vcc_pwrgood;
  wire mprj2_vdd_pwrgood;
  wire mprj_ack_i_core;
  wire \mprj_adr_o_core[0] ;
  wire \mprj_adr_o_core[10] ;
  wire \mprj_adr_o_core[11] ;
  wire \mprj_adr_o_core[12] ;
  wire \mprj_adr_o_core[13] ;
  wire \mprj_adr_o_core[14] ;
  wire \mprj_adr_o_core[15] ;
  wire \mprj_adr_o_core[16] ;
  wire \mprj_adr_o_core[17] ;
  wire \mprj_adr_o_core[18] ;
  wire \mprj_adr_o_core[19] ;
  wire \mprj_adr_o_core[1] ;
  wire \mprj_adr_o_core[20] ;
  wire \mprj_adr_o_core[21] ;
  wire \mprj_adr_o_core[22] ;
  wire \mprj_adr_o_core[23] ;
  wire \mprj_adr_o_core[24] ;
  wire \mprj_adr_o_core[25] ;
  wire \mprj_adr_o_core[26] ;
  wire \mprj_adr_o_core[27] ;
  wire \mprj_adr_o_core[28] ;
  wire \mprj_adr_o_core[29] ;
  wire \mprj_adr_o_core[2] ;
  wire \mprj_adr_o_core[30] ;
  wire \mprj_adr_o_core[31] ;
  wire \mprj_adr_o_core[3] ;
  wire \mprj_adr_o_core[4] ;
  wire \mprj_adr_o_core[5] ;
  wire \mprj_adr_o_core[6] ;
  wire \mprj_adr_o_core[7] ;
  wire \mprj_adr_o_core[8] ;
  wire \mprj_adr_o_core[9] ;
  wire \mprj_adr_o_user[0] ;
  wire \mprj_adr_o_user[10] ;
  wire \mprj_adr_o_user[11] ;
  wire \mprj_adr_o_user[12] ;
  wire \mprj_adr_o_user[13] ;
  wire \mprj_adr_o_user[14] ;
  wire \mprj_adr_o_user[15] ;
  wire \mprj_adr_o_user[16] ;
  wire \mprj_adr_o_user[17] ;
  wire \mprj_adr_o_user[18] ;
  wire \mprj_adr_o_user[19] ;
  wire \mprj_adr_o_user[1] ;
  wire \mprj_adr_o_user[20] ;
  wire \mprj_adr_o_user[21] ;
  wire \mprj_adr_o_user[22] ;
  wire \mprj_adr_o_user[23] ;
  wire \mprj_adr_o_user[24] ;
  wire \mprj_adr_o_user[25] ;
  wire \mprj_adr_o_user[26] ;
  wire \mprj_adr_o_user[27] ;
  wire \mprj_adr_o_user[28] ;
  wire \mprj_adr_o_user[29] ;
  wire \mprj_adr_o_user[2] ;
  wire \mprj_adr_o_user[30] ;
  wire \mprj_adr_o_user[31] ;
  wire \mprj_adr_o_user[3] ;
  wire \mprj_adr_o_user[4] ;
  wire \mprj_adr_o_user[5] ;
  wire \mprj_adr_o_user[6] ;
  wire \mprj_adr_o_user[7] ;
  wire \mprj_adr_o_user[8] ;
  wire \mprj_adr_o_user[9] ;
  wire mprj_clock;
  wire mprj_clock2;
  wire mprj_cyc_o_core;
  wire mprj_cyc_o_user;
  wire \mprj_dat_i_core[0] ;
  wire \mprj_dat_i_core[10] ;
  wire \mprj_dat_i_core[11] ;
  wire \mprj_dat_i_core[12] ;
  wire \mprj_dat_i_core[13] ;
  wire \mprj_dat_i_core[14] ;
  wire \mprj_dat_i_core[15] ;
  wire \mprj_dat_i_core[16] ;
  wire \mprj_dat_i_core[17] ;
  wire \mprj_dat_i_core[18] ;
  wire \mprj_dat_i_core[19] ;
  wire \mprj_dat_i_core[1] ;
  wire \mprj_dat_i_core[20] ;
  wire \mprj_dat_i_core[21] ;
  wire \mprj_dat_i_core[22] ;
  wire \mprj_dat_i_core[23] ;
  wire \mprj_dat_i_core[24] ;
  wire \mprj_dat_i_core[25] ;
  wire \mprj_dat_i_core[26] ;
  wire \mprj_dat_i_core[27] ;
  wire \mprj_dat_i_core[28] ;
  wire \mprj_dat_i_core[29] ;
  wire \mprj_dat_i_core[2] ;
  wire \mprj_dat_i_core[30] ;
  wire \mprj_dat_i_core[31] ;
  wire \mprj_dat_i_core[3] ;
  wire \mprj_dat_i_core[4] ;
  wire \mprj_dat_i_core[5] ;
  wire \mprj_dat_i_core[6] ;
  wire \mprj_dat_i_core[7] ;
  wire \mprj_dat_i_core[8] ;
  wire \mprj_dat_i_core[9] ;
  wire \mprj_dat_o_core[0] ;
  wire \mprj_dat_o_core[10] ;
  wire \mprj_dat_o_core[11] ;
  wire \mprj_dat_o_core[12] ;
  wire \mprj_dat_o_core[13] ;
  wire \mprj_dat_o_core[14] ;
  wire \mprj_dat_o_core[15] ;
  wire \mprj_dat_o_core[16] ;
  wire \mprj_dat_o_core[17] ;
  wire \mprj_dat_o_core[18] ;
  wire \mprj_dat_o_core[19] ;
  wire \mprj_dat_o_core[1] ;
  wire \mprj_dat_o_core[20] ;
  wire \mprj_dat_o_core[21] ;
  wire \mprj_dat_o_core[22] ;
  wire \mprj_dat_o_core[23] ;
  wire \mprj_dat_o_core[24] ;
  wire \mprj_dat_o_core[25] ;
  wire \mprj_dat_o_core[26] ;
  wire \mprj_dat_o_core[27] ;
  wire \mprj_dat_o_core[28] ;
  wire \mprj_dat_o_core[29] ;
  wire \mprj_dat_o_core[2] ;
  wire \mprj_dat_o_core[30] ;
  wire \mprj_dat_o_core[31] ;
  wire \mprj_dat_o_core[3] ;
  wire \mprj_dat_o_core[4] ;
  wire \mprj_dat_o_core[5] ;
  wire \mprj_dat_o_core[6] ;
  wire \mprj_dat_o_core[7] ;
  wire \mprj_dat_o_core[8] ;
  wire \mprj_dat_o_core[9] ;
  wire \mprj_dat_o_user[0] ;
  wire \mprj_dat_o_user[10] ;
  wire \mprj_dat_o_user[11] ;
  wire \mprj_dat_o_user[12] ;
  wire \mprj_dat_o_user[13] ;
  wire \mprj_dat_o_user[14] ;
  wire \mprj_dat_o_user[15] ;
  wire \mprj_dat_o_user[16] ;
  wire \mprj_dat_o_user[17] ;
  wire \mprj_dat_o_user[18] ;
  wire \mprj_dat_o_user[19] ;
  wire \mprj_dat_o_user[1] ;
  wire \mprj_dat_o_user[20] ;
  wire \mprj_dat_o_user[21] ;
  wire \mprj_dat_o_user[22] ;
  wire \mprj_dat_o_user[23] ;
  wire \mprj_dat_o_user[24] ;
  wire \mprj_dat_o_user[25] ;
  wire \mprj_dat_o_user[26] ;
  wire \mprj_dat_o_user[27] ;
  wire \mprj_dat_o_user[28] ;
  wire \mprj_dat_o_user[29] ;
  wire \mprj_dat_o_user[2] ;
  wire \mprj_dat_o_user[30] ;
  wire \mprj_dat_o_user[31] ;
  wire \mprj_dat_o_user[3] ;
  wire \mprj_dat_o_user[4] ;
  wire \mprj_dat_o_user[5] ;
  wire \mprj_dat_o_user[6] ;
  wire \mprj_dat_o_user[7] ;
  wire \mprj_dat_o_user[8] ;
  wire \mprj_dat_o_user[9] ;
  inout [37:0] mprj_io;
  wire \mprj_io_analog_en[0] ;
  wire \mprj_io_analog_en[10] ;
  wire \mprj_io_analog_en[11] ;
  wire \mprj_io_analog_en[12] ;
  wire \mprj_io_analog_en[13] ;
  wire \mprj_io_analog_en[14] ;
  wire \mprj_io_analog_en[15] ;
  wire \mprj_io_analog_en[16] ;
  wire \mprj_io_analog_en[17] ;
  wire \mprj_io_analog_en[18] ;
  wire \mprj_io_analog_en[19] ;
  wire \mprj_io_analog_en[1] ;
  wire \mprj_io_analog_en[20] ;
  wire \mprj_io_analog_en[21] ;
  wire \mprj_io_analog_en[22] ;
  wire \mprj_io_analog_en[23] ;
  wire \mprj_io_analog_en[24] ;
  wire \mprj_io_analog_en[25] ;
  wire \mprj_io_analog_en[26] ;
  wire \mprj_io_analog_en[27] ;
  wire \mprj_io_analog_en[28] ;
  wire \mprj_io_analog_en[29] ;
  wire \mprj_io_analog_en[2] ;
  wire \mprj_io_analog_en[30] ;
  wire \mprj_io_analog_en[31] ;
  wire \mprj_io_analog_en[32] ;
  wire \mprj_io_analog_en[33] ;
  wire \mprj_io_analog_en[34] ;
  wire \mprj_io_analog_en[35] ;
  wire \mprj_io_analog_en[36] ;
  wire \mprj_io_analog_en[37] ;
  wire \mprj_io_analog_en[3] ;
  wire \mprj_io_analog_en[4] ;
  wire \mprj_io_analog_en[5] ;
  wire \mprj_io_analog_en[6] ;
  wire \mprj_io_analog_en[7] ;
  wire \mprj_io_analog_en[8] ;
  wire \mprj_io_analog_en[9] ;
  wire \mprj_io_analog_pol[0] ;
  wire \mprj_io_analog_pol[10] ;
  wire \mprj_io_analog_pol[11] ;
  wire \mprj_io_analog_pol[12] ;
  wire \mprj_io_analog_pol[13] ;
  wire \mprj_io_analog_pol[14] ;
  wire \mprj_io_analog_pol[15] ;
  wire \mprj_io_analog_pol[16] ;
  wire \mprj_io_analog_pol[17] ;
  wire \mprj_io_analog_pol[18] ;
  wire \mprj_io_analog_pol[19] ;
  wire \mprj_io_analog_pol[1] ;
  wire \mprj_io_analog_pol[20] ;
  wire \mprj_io_analog_pol[21] ;
  wire \mprj_io_analog_pol[22] ;
  wire \mprj_io_analog_pol[23] ;
  wire \mprj_io_analog_pol[24] ;
  wire \mprj_io_analog_pol[25] ;
  wire \mprj_io_analog_pol[26] ;
  wire \mprj_io_analog_pol[27] ;
  wire \mprj_io_analog_pol[28] ;
  wire \mprj_io_analog_pol[29] ;
  wire \mprj_io_analog_pol[2] ;
  wire \mprj_io_analog_pol[30] ;
  wire \mprj_io_analog_pol[31] ;
  wire \mprj_io_analog_pol[32] ;
  wire \mprj_io_analog_pol[33] ;
  wire \mprj_io_analog_pol[34] ;
  wire \mprj_io_analog_pol[35] ;
  wire \mprj_io_analog_pol[36] ;
  wire \mprj_io_analog_pol[37] ;
  wire \mprj_io_analog_pol[3] ;
  wire \mprj_io_analog_pol[4] ;
  wire \mprj_io_analog_pol[5] ;
  wire \mprj_io_analog_pol[6] ;
  wire \mprj_io_analog_pol[7] ;
  wire \mprj_io_analog_pol[8] ;
  wire \mprj_io_analog_pol[9] ;
  wire \mprj_io_analog_sel[0] ;
  wire \mprj_io_analog_sel[10] ;
  wire \mprj_io_analog_sel[11] ;
  wire \mprj_io_analog_sel[12] ;
  wire \mprj_io_analog_sel[13] ;
  wire \mprj_io_analog_sel[14] ;
  wire \mprj_io_analog_sel[15] ;
  wire \mprj_io_analog_sel[16] ;
  wire \mprj_io_analog_sel[17] ;
  wire \mprj_io_analog_sel[18] ;
  wire \mprj_io_analog_sel[19] ;
  wire \mprj_io_analog_sel[1] ;
  wire \mprj_io_analog_sel[20] ;
  wire \mprj_io_analog_sel[21] ;
  wire \mprj_io_analog_sel[22] ;
  wire \mprj_io_analog_sel[23] ;
  wire \mprj_io_analog_sel[24] ;
  wire \mprj_io_analog_sel[25] ;
  wire \mprj_io_analog_sel[26] ;
  wire \mprj_io_analog_sel[27] ;
  wire \mprj_io_analog_sel[28] ;
  wire \mprj_io_analog_sel[29] ;
  wire \mprj_io_analog_sel[2] ;
  wire \mprj_io_analog_sel[30] ;
  wire \mprj_io_analog_sel[31] ;
  wire \mprj_io_analog_sel[32] ;
  wire \mprj_io_analog_sel[33] ;
  wire \mprj_io_analog_sel[34] ;
  wire \mprj_io_analog_sel[35] ;
  wire \mprj_io_analog_sel[36] ;
  wire \mprj_io_analog_sel[37] ;
  wire \mprj_io_analog_sel[3] ;
  wire \mprj_io_analog_sel[4] ;
  wire \mprj_io_analog_sel[5] ;
  wire \mprj_io_analog_sel[6] ;
  wire \mprj_io_analog_sel[7] ;
  wire \mprj_io_analog_sel[8] ;
  wire \mprj_io_analog_sel[9] ;
  wire \mprj_io_dm[0] ;
  wire \mprj_io_dm[100] ;
  wire \mprj_io_dm[101] ;
  wire \mprj_io_dm[102] ;
  wire \mprj_io_dm[103] ;
  wire \mprj_io_dm[104] ;
  wire \mprj_io_dm[105] ;
  wire \mprj_io_dm[106] ;
  wire \mprj_io_dm[107] ;
  wire \mprj_io_dm[108] ;
  wire \mprj_io_dm[109] ;
  wire \mprj_io_dm[10] ;
  wire \mprj_io_dm[110] ;
  wire \mprj_io_dm[111] ;
  wire \mprj_io_dm[112] ;
  wire \mprj_io_dm[113] ;
  wire \mprj_io_dm[11] ;
  wire \mprj_io_dm[12] ;
  wire \mprj_io_dm[13] ;
  wire \mprj_io_dm[14] ;
  wire \mprj_io_dm[15] ;
  wire \mprj_io_dm[16] ;
  wire \mprj_io_dm[17] ;
  wire \mprj_io_dm[18] ;
  wire \mprj_io_dm[19] ;
  wire \mprj_io_dm[1] ;
  wire \mprj_io_dm[20] ;
  wire \mprj_io_dm[21] ;
  wire \mprj_io_dm[22] ;
  wire \mprj_io_dm[23] ;
  wire \mprj_io_dm[24] ;
  wire \mprj_io_dm[25] ;
  wire \mprj_io_dm[26] ;
  wire \mprj_io_dm[27] ;
  wire \mprj_io_dm[28] ;
  wire \mprj_io_dm[29] ;
  wire \mprj_io_dm[2] ;
  wire \mprj_io_dm[30] ;
  wire \mprj_io_dm[31] ;
  wire \mprj_io_dm[32] ;
  wire \mprj_io_dm[33] ;
  wire \mprj_io_dm[34] ;
  wire \mprj_io_dm[35] ;
  wire \mprj_io_dm[36] ;
  wire \mprj_io_dm[37] ;
  wire \mprj_io_dm[38] ;
  wire \mprj_io_dm[39] ;
  wire \mprj_io_dm[3] ;
  wire \mprj_io_dm[40] ;
  wire \mprj_io_dm[41] ;
  wire \mprj_io_dm[42] ;
  wire \mprj_io_dm[43] ;
  wire \mprj_io_dm[44] ;
  wire \mprj_io_dm[45] ;
  wire \mprj_io_dm[46] ;
  wire \mprj_io_dm[47] ;
  wire \mprj_io_dm[48] ;
  wire \mprj_io_dm[49] ;
  wire \mprj_io_dm[4] ;
  wire \mprj_io_dm[50] ;
  wire \mprj_io_dm[51] ;
  wire \mprj_io_dm[52] ;
  wire \mprj_io_dm[53] ;
  wire \mprj_io_dm[54] ;
  wire \mprj_io_dm[55] ;
  wire \mprj_io_dm[56] ;
  wire \mprj_io_dm[57] ;
  wire \mprj_io_dm[58] ;
  wire \mprj_io_dm[59] ;
  wire \mprj_io_dm[5] ;
  wire \mprj_io_dm[60] ;
  wire \mprj_io_dm[61] ;
  wire \mprj_io_dm[62] ;
  wire \mprj_io_dm[63] ;
  wire \mprj_io_dm[64] ;
  wire \mprj_io_dm[65] ;
  wire \mprj_io_dm[66] ;
  wire \mprj_io_dm[67] ;
  wire \mprj_io_dm[68] ;
  wire \mprj_io_dm[69] ;
  wire \mprj_io_dm[6] ;
  wire \mprj_io_dm[70] ;
  wire \mprj_io_dm[71] ;
  wire \mprj_io_dm[72] ;
  wire \mprj_io_dm[73] ;
  wire \mprj_io_dm[74] ;
  wire \mprj_io_dm[75] ;
  wire \mprj_io_dm[76] ;
  wire \mprj_io_dm[77] ;
  wire \mprj_io_dm[78] ;
  wire \mprj_io_dm[79] ;
  wire \mprj_io_dm[7] ;
  wire \mprj_io_dm[80] ;
  wire \mprj_io_dm[81] ;
  wire \mprj_io_dm[82] ;
  wire \mprj_io_dm[83] ;
  wire \mprj_io_dm[84] ;
  wire \mprj_io_dm[85] ;
  wire \mprj_io_dm[86] ;
  wire \mprj_io_dm[87] ;
  wire \mprj_io_dm[88] ;
  wire \mprj_io_dm[89] ;
  wire \mprj_io_dm[8] ;
  wire \mprj_io_dm[90] ;
  wire \mprj_io_dm[91] ;
  wire \mprj_io_dm[92] ;
  wire \mprj_io_dm[93] ;
  wire \mprj_io_dm[94] ;
  wire \mprj_io_dm[95] ;
  wire \mprj_io_dm[96] ;
  wire \mprj_io_dm[97] ;
  wire \mprj_io_dm[98] ;
  wire \mprj_io_dm[99] ;
  wire \mprj_io_dm[9] ;
  wire \mprj_io_enh[0] ;
  wire \mprj_io_enh[10] ;
  wire \mprj_io_enh[11] ;
  wire \mprj_io_enh[12] ;
  wire \mprj_io_enh[13] ;
  wire \mprj_io_enh[14] ;
  wire \mprj_io_enh[15] ;
  wire \mprj_io_enh[16] ;
  wire \mprj_io_enh[17] ;
  wire \mprj_io_enh[18] ;
  wire \mprj_io_enh[19] ;
  wire \mprj_io_enh[1] ;
  wire \mprj_io_enh[20] ;
  wire \mprj_io_enh[21] ;
  wire \mprj_io_enh[22] ;
  wire \mprj_io_enh[23] ;
  wire \mprj_io_enh[24] ;
  wire \mprj_io_enh[25] ;
  wire \mprj_io_enh[26] ;
  wire \mprj_io_enh[27] ;
  wire \mprj_io_enh[28] ;
  wire \mprj_io_enh[29] ;
  wire \mprj_io_enh[2] ;
  wire \mprj_io_enh[30] ;
  wire \mprj_io_enh[31] ;
  wire \mprj_io_enh[32] ;
  wire \mprj_io_enh[33] ;
  wire \mprj_io_enh[34] ;
  wire \mprj_io_enh[35] ;
  wire \mprj_io_enh[36] ;
  wire \mprj_io_enh[37] ;
  wire \mprj_io_enh[3] ;
  wire \mprj_io_enh[4] ;
  wire \mprj_io_enh[5] ;
  wire \mprj_io_enh[6] ;
  wire \mprj_io_enh[7] ;
  wire \mprj_io_enh[8] ;
  wire \mprj_io_enh[9] ;
  wire \mprj_io_hldh_n[0] ;
  wire \mprj_io_hldh_n[10] ;
  wire \mprj_io_hldh_n[11] ;
  wire \mprj_io_hldh_n[12] ;
  wire \mprj_io_hldh_n[13] ;
  wire \mprj_io_hldh_n[14] ;
  wire \mprj_io_hldh_n[15] ;
  wire \mprj_io_hldh_n[16] ;
  wire \mprj_io_hldh_n[17] ;
  wire \mprj_io_hldh_n[18] ;
  wire \mprj_io_hldh_n[19] ;
  wire \mprj_io_hldh_n[1] ;
  wire \mprj_io_hldh_n[20] ;
  wire \mprj_io_hldh_n[21] ;
  wire \mprj_io_hldh_n[22] ;
  wire \mprj_io_hldh_n[23] ;
  wire \mprj_io_hldh_n[24] ;
  wire \mprj_io_hldh_n[25] ;
  wire \mprj_io_hldh_n[26] ;
  wire \mprj_io_hldh_n[27] ;
  wire \mprj_io_hldh_n[28] ;
  wire \mprj_io_hldh_n[29] ;
  wire \mprj_io_hldh_n[2] ;
  wire \mprj_io_hldh_n[30] ;
  wire \mprj_io_hldh_n[31] ;
  wire \mprj_io_hldh_n[32] ;
  wire \mprj_io_hldh_n[33] ;
  wire \mprj_io_hldh_n[34] ;
  wire \mprj_io_hldh_n[35] ;
  wire \mprj_io_hldh_n[36] ;
  wire \mprj_io_hldh_n[37] ;
  wire \mprj_io_hldh_n[3] ;
  wire \mprj_io_hldh_n[4] ;
  wire \mprj_io_hldh_n[5] ;
  wire \mprj_io_hldh_n[6] ;
  wire \mprj_io_hldh_n[7] ;
  wire \mprj_io_hldh_n[8] ;
  wire \mprj_io_hldh_n[9] ;
  wire \mprj_io_holdover[0] ;
  wire \mprj_io_holdover[10] ;
  wire \mprj_io_holdover[11] ;
  wire \mprj_io_holdover[12] ;
  wire \mprj_io_holdover[13] ;
  wire \mprj_io_holdover[14] ;
  wire \mprj_io_holdover[15] ;
  wire \mprj_io_holdover[16] ;
  wire \mprj_io_holdover[17] ;
  wire \mprj_io_holdover[18] ;
  wire \mprj_io_holdover[19] ;
  wire \mprj_io_holdover[1] ;
  wire \mprj_io_holdover[20] ;
  wire \mprj_io_holdover[21] ;
  wire \mprj_io_holdover[22] ;
  wire \mprj_io_holdover[23] ;
  wire \mprj_io_holdover[24] ;
  wire \mprj_io_holdover[25] ;
  wire \mprj_io_holdover[26] ;
  wire \mprj_io_holdover[27] ;
  wire \mprj_io_holdover[28] ;
  wire \mprj_io_holdover[29] ;
  wire \mprj_io_holdover[2] ;
  wire \mprj_io_holdover[30] ;
  wire \mprj_io_holdover[31] ;
  wire \mprj_io_holdover[32] ;
  wire \mprj_io_holdover[33] ;
  wire \mprj_io_holdover[34] ;
  wire \mprj_io_holdover[35] ;
  wire \mprj_io_holdover[36] ;
  wire \mprj_io_holdover[37] ;
  wire \mprj_io_holdover[3] ;
  wire \mprj_io_holdover[4] ;
  wire \mprj_io_holdover[5] ;
  wire \mprj_io_holdover[6] ;
  wire \mprj_io_holdover[7] ;
  wire \mprj_io_holdover[8] ;
  wire \mprj_io_holdover[9] ;
  wire \mprj_io_ib_mode_sel[0] ;
  wire \mprj_io_ib_mode_sel[10] ;
  wire \mprj_io_ib_mode_sel[11] ;
  wire \mprj_io_ib_mode_sel[12] ;
  wire \mprj_io_ib_mode_sel[13] ;
  wire \mprj_io_ib_mode_sel[14] ;
  wire \mprj_io_ib_mode_sel[15] ;
  wire \mprj_io_ib_mode_sel[16] ;
  wire \mprj_io_ib_mode_sel[17] ;
  wire \mprj_io_ib_mode_sel[18] ;
  wire \mprj_io_ib_mode_sel[19] ;
  wire \mprj_io_ib_mode_sel[1] ;
  wire \mprj_io_ib_mode_sel[20] ;
  wire \mprj_io_ib_mode_sel[21] ;
  wire \mprj_io_ib_mode_sel[22] ;
  wire \mprj_io_ib_mode_sel[23] ;
  wire \mprj_io_ib_mode_sel[24] ;
  wire \mprj_io_ib_mode_sel[25] ;
  wire \mprj_io_ib_mode_sel[26] ;
  wire \mprj_io_ib_mode_sel[27] ;
  wire \mprj_io_ib_mode_sel[28] ;
  wire \mprj_io_ib_mode_sel[29] ;
  wire \mprj_io_ib_mode_sel[2] ;
  wire \mprj_io_ib_mode_sel[30] ;
  wire \mprj_io_ib_mode_sel[31] ;
  wire \mprj_io_ib_mode_sel[32] ;
  wire \mprj_io_ib_mode_sel[33] ;
  wire \mprj_io_ib_mode_sel[34] ;
  wire \mprj_io_ib_mode_sel[35] ;
  wire \mprj_io_ib_mode_sel[36] ;
  wire \mprj_io_ib_mode_sel[37] ;
  wire \mprj_io_ib_mode_sel[3] ;
  wire \mprj_io_ib_mode_sel[4] ;
  wire \mprj_io_ib_mode_sel[5] ;
  wire \mprj_io_ib_mode_sel[6] ;
  wire \mprj_io_ib_mode_sel[7] ;
  wire \mprj_io_ib_mode_sel[8] ;
  wire \mprj_io_ib_mode_sel[9] ;
  wire \mprj_io_in[0] ;
  wire \mprj_io_in[10] ;
  wire \mprj_io_in[11] ;
  wire \mprj_io_in[12] ;
  wire \mprj_io_in[13] ;
  wire \mprj_io_in[14] ;
  wire \mprj_io_in[15] ;
  wire \mprj_io_in[16] ;
  wire \mprj_io_in[17] ;
  wire \mprj_io_in[18] ;
  wire \mprj_io_in[19] ;
  wire \mprj_io_in[1] ;
  wire \mprj_io_in[20] ;
  wire \mprj_io_in[21] ;
  wire \mprj_io_in[22] ;
  wire \mprj_io_in[23] ;
  wire \mprj_io_in[24] ;
  wire \mprj_io_in[25] ;
  wire \mprj_io_in[26] ;
  wire \mprj_io_in[27] ;
  wire \mprj_io_in[28] ;
  wire \mprj_io_in[29] ;
  wire \mprj_io_in[2] ;
  wire \mprj_io_in[30] ;
  wire \mprj_io_in[31] ;
  wire \mprj_io_in[32] ;
  wire \mprj_io_in[33] ;
  wire \mprj_io_in[34] ;
  wire \mprj_io_in[35] ;
  wire \mprj_io_in[36] ;
  wire \mprj_io_in[37] ;
  wire \mprj_io_in[3] ;
  wire \mprj_io_in[4] ;
  wire \mprj_io_in[5] ;
  wire \mprj_io_in[6] ;
  wire \mprj_io_in[7] ;
  wire \mprj_io_in[8] ;
  wire \mprj_io_in[9] ;
  wire \mprj_io_inp_dis[0] ;
  wire \mprj_io_inp_dis[10] ;
  wire \mprj_io_inp_dis[11] ;
  wire \mprj_io_inp_dis[12] ;
  wire \mprj_io_inp_dis[13] ;
  wire \mprj_io_inp_dis[14] ;
  wire \mprj_io_inp_dis[15] ;
  wire \mprj_io_inp_dis[16] ;
  wire \mprj_io_inp_dis[17] ;
  wire \mprj_io_inp_dis[18] ;
  wire \mprj_io_inp_dis[19] ;
  wire \mprj_io_inp_dis[1] ;
  wire \mprj_io_inp_dis[20] ;
  wire \mprj_io_inp_dis[21] ;
  wire \mprj_io_inp_dis[22] ;
  wire \mprj_io_inp_dis[23] ;
  wire \mprj_io_inp_dis[24] ;
  wire \mprj_io_inp_dis[25] ;
  wire \mprj_io_inp_dis[26] ;
  wire \mprj_io_inp_dis[27] ;
  wire \mprj_io_inp_dis[28] ;
  wire \mprj_io_inp_dis[29] ;
  wire \mprj_io_inp_dis[2] ;
  wire \mprj_io_inp_dis[30] ;
  wire \mprj_io_inp_dis[31] ;
  wire \mprj_io_inp_dis[32] ;
  wire \mprj_io_inp_dis[33] ;
  wire \mprj_io_inp_dis[34] ;
  wire \mprj_io_inp_dis[35] ;
  wire \mprj_io_inp_dis[36] ;
  wire \mprj_io_inp_dis[37] ;
  wire \mprj_io_inp_dis[3] ;
  wire \mprj_io_inp_dis[4] ;
  wire \mprj_io_inp_dis[5] ;
  wire \mprj_io_inp_dis[6] ;
  wire \mprj_io_inp_dis[7] ;
  wire \mprj_io_inp_dis[8] ;
  wire \mprj_io_inp_dis[9] ;
  wire mprj_io_loader_clock;
  wire mprj_io_loader_data;
  wire mprj_io_loader_resetn;
  wire \mprj_io_oeb[0] ;
  wire \mprj_io_oeb[10] ;
  wire \mprj_io_oeb[11] ;
  wire \mprj_io_oeb[12] ;
  wire \mprj_io_oeb[13] ;
  wire \mprj_io_oeb[14] ;
  wire \mprj_io_oeb[15] ;
  wire \mprj_io_oeb[16] ;
  wire \mprj_io_oeb[17] ;
  wire \mprj_io_oeb[18] ;
  wire \mprj_io_oeb[19] ;
  wire \mprj_io_oeb[1] ;
  wire \mprj_io_oeb[20] ;
  wire \mprj_io_oeb[21] ;
  wire \mprj_io_oeb[22] ;
  wire \mprj_io_oeb[23] ;
  wire \mprj_io_oeb[24] ;
  wire \mprj_io_oeb[25] ;
  wire \mprj_io_oeb[26] ;
  wire \mprj_io_oeb[27] ;
  wire \mprj_io_oeb[28] ;
  wire \mprj_io_oeb[29] ;
  wire \mprj_io_oeb[2] ;
  wire \mprj_io_oeb[30] ;
  wire \mprj_io_oeb[31] ;
  wire \mprj_io_oeb[32] ;
  wire \mprj_io_oeb[33] ;
  wire \mprj_io_oeb[34] ;
  wire \mprj_io_oeb[35] ;
  wire \mprj_io_oeb[36] ;
  wire \mprj_io_oeb[37] ;
  wire \mprj_io_oeb[3] ;
  wire \mprj_io_oeb[4] ;
  wire \mprj_io_oeb[5] ;
  wire \mprj_io_oeb[6] ;
  wire \mprj_io_oeb[7] ;
  wire \mprj_io_oeb[8] ;
  wire \mprj_io_oeb[9] ;
  wire \mprj_io_out[0] ;
  wire \mprj_io_out[10] ;
  wire \mprj_io_out[11] ;
  wire \mprj_io_out[12] ;
  wire \mprj_io_out[13] ;
  wire \mprj_io_out[14] ;
  wire \mprj_io_out[15] ;
  wire \mprj_io_out[16] ;
  wire \mprj_io_out[17] ;
  wire \mprj_io_out[18] ;
  wire \mprj_io_out[19] ;
  wire \mprj_io_out[1] ;
  wire \mprj_io_out[20] ;
  wire \mprj_io_out[21] ;
  wire \mprj_io_out[22] ;
  wire \mprj_io_out[23] ;
  wire \mprj_io_out[24] ;
  wire \mprj_io_out[25] ;
  wire \mprj_io_out[26] ;
  wire \mprj_io_out[27] ;
  wire \mprj_io_out[28] ;
  wire \mprj_io_out[29] ;
  wire \mprj_io_out[2] ;
  wire \mprj_io_out[30] ;
  wire \mprj_io_out[31] ;
  wire \mprj_io_out[32] ;
  wire \mprj_io_out[33] ;
  wire \mprj_io_out[34] ;
  wire \mprj_io_out[35] ;
  wire \mprj_io_out[36] ;
  wire \mprj_io_out[37] ;
  wire \mprj_io_out[3] ;
  wire \mprj_io_out[4] ;
  wire \mprj_io_out[5] ;
  wire \mprj_io_out[6] ;
  wire \mprj_io_out[7] ;
  wire \mprj_io_out[8] ;
  wire \mprj_io_out[9] ;
  wire \mprj_io_slow_sel[0] ;
  wire \mprj_io_slow_sel[10] ;
  wire \mprj_io_slow_sel[11] ;
  wire \mprj_io_slow_sel[12] ;
  wire \mprj_io_slow_sel[13] ;
  wire \mprj_io_slow_sel[14] ;
  wire \mprj_io_slow_sel[15] ;
  wire \mprj_io_slow_sel[16] ;
  wire \mprj_io_slow_sel[17] ;
  wire \mprj_io_slow_sel[18] ;
  wire \mprj_io_slow_sel[19] ;
  wire \mprj_io_slow_sel[1] ;
  wire \mprj_io_slow_sel[20] ;
  wire \mprj_io_slow_sel[21] ;
  wire \mprj_io_slow_sel[22] ;
  wire \mprj_io_slow_sel[23] ;
  wire \mprj_io_slow_sel[24] ;
  wire \mprj_io_slow_sel[25] ;
  wire \mprj_io_slow_sel[26] ;
  wire \mprj_io_slow_sel[27] ;
  wire \mprj_io_slow_sel[28] ;
  wire \mprj_io_slow_sel[29] ;
  wire \mprj_io_slow_sel[2] ;
  wire \mprj_io_slow_sel[30] ;
  wire \mprj_io_slow_sel[31] ;
  wire \mprj_io_slow_sel[32] ;
  wire \mprj_io_slow_sel[33] ;
  wire \mprj_io_slow_sel[34] ;
  wire \mprj_io_slow_sel[35] ;
  wire \mprj_io_slow_sel[36] ;
  wire \mprj_io_slow_sel[37] ;
  wire \mprj_io_slow_sel[3] ;
  wire \mprj_io_slow_sel[4] ;
  wire \mprj_io_slow_sel[5] ;
  wire \mprj_io_slow_sel[6] ;
  wire \mprj_io_slow_sel[7] ;
  wire \mprj_io_slow_sel[8] ;
  wire \mprj_io_slow_sel[9] ;
  wire \mprj_io_vtrip_sel[0] ;
  wire \mprj_io_vtrip_sel[10] ;
  wire \mprj_io_vtrip_sel[11] ;
  wire \mprj_io_vtrip_sel[12] ;
  wire \mprj_io_vtrip_sel[13] ;
  wire \mprj_io_vtrip_sel[14] ;
  wire \mprj_io_vtrip_sel[15] ;
  wire \mprj_io_vtrip_sel[16] ;
  wire \mprj_io_vtrip_sel[17] ;
  wire \mprj_io_vtrip_sel[18] ;
  wire \mprj_io_vtrip_sel[19] ;
  wire \mprj_io_vtrip_sel[1] ;
  wire \mprj_io_vtrip_sel[20] ;
  wire \mprj_io_vtrip_sel[21] ;
  wire \mprj_io_vtrip_sel[22] ;
  wire \mprj_io_vtrip_sel[23] ;
  wire \mprj_io_vtrip_sel[24] ;
  wire \mprj_io_vtrip_sel[25] ;
  wire \mprj_io_vtrip_sel[26] ;
  wire \mprj_io_vtrip_sel[27] ;
  wire \mprj_io_vtrip_sel[28] ;
  wire \mprj_io_vtrip_sel[29] ;
  wire \mprj_io_vtrip_sel[2] ;
  wire \mprj_io_vtrip_sel[30] ;
  wire \mprj_io_vtrip_sel[31] ;
  wire \mprj_io_vtrip_sel[32] ;
  wire \mprj_io_vtrip_sel[33] ;
  wire \mprj_io_vtrip_sel[34] ;
  wire \mprj_io_vtrip_sel[35] ;
  wire \mprj_io_vtrip_sel[36] ;
  wire \mprj_io_vtrip_sel[37] ;
  wire \mprj_io_vtrip_sel[3] ;
  wire \mprj_io_vtrip_sel[4] ;
  wire \mprj_io_vtrip_sel[5] ;
  wire \mprj_io_vtrip_sel[6] ;
  wire \mprj_io_vtrip_sel[7] ;
  wire \mprj_io_vtrip_sel[8] ;
  wire \mprj_io_vtrip_sel[9] ;
  wire mprj_reset;
  wire mprj_resetn;
  wire \mprj_sel_o_core[0] ;
  wire \mprj_sel_o_core[1] ;
  wire \mprj_sel_o_core[2] ;
  wire \mprj_sel_o_core[3] ;
  wire \mprj_sel_o_user[0] ;
  wire \mprj_sel_o_user[1] ;
  wire \mprj_sel_o_user[2] ;
  wire \mprj_sel_o_user[3] ;
  wire mprj_stb_o_core;
  wire mprj_stb_o_user;
  wire mprj_vcc_pwrgood;
  wire mprj_vdd_pwrgood;
  wire mprj_we_o_core;
  wire mprj_we_o_user;
  wire por_l;
  wire porb_h;
  wire porb_l;
  output [3:0] pwr_ctrl_out;
  input resetb;
  wire rstb_h;
  wire rstb_l;
  wire sdo_out;
  wire sdo_outenb;
  wire \spi_ro_config_core[0] ;
  wire \spi_ro_config_core[1] ;
  wire \spi_ro_config_core[2] ;
  wire \spi_ro_config_core[3] ;
  wire \spi_ro_config_core[4] ;
  wire \spi_ro_config_core[5] ;
  wire \spi_ro_config_core[6] ;
  wire \spi_ro_config_core[7] ;
  wire \user_analog_io[0] ;
  wire \user_analog_io[10] ;
  wire \user_analog_io[11] ;
  wire \user_analog_io[12] ;
  wire \user_analog_io[13] ;
  wire \user_analog_io[14] ;
  wire \user_analog_io[15] ;
  wire \user_analog_io[16] ;
  wire \user_analog_io[17] ;
  wire \user_analog_io[18] ;
  wire \user_analog_io[19] ;
  wire \user_analog_io[1] ;
  wire \user_analog_io[20] ;
  wire \user_analog_io[21] ;
  wire \user_analog_io[22] ;
  wire \user_analog_io[23] ;
  wire \user_analog_io[24] ;
  wire \user_analog_io[25] ;
  wire \user_analog_io[26] ;
  wire \user_analog_io[27] ;
  wire \user_analog_io[28] ;
  wire \user_analog_io[29] ;
  wire \user_analog_io[2] ;
  wire \user_analog_io[30] ;
  wire \user_analog_io[3] ;
  wire \user_analog_io[4] ;
  wire \user_analog_io[5] ;
  wire \user_analog_io[6] ;
  wire \user_analog_io[7] ;
  wire \user_analog_io[8] ;
  wire \user_analog_io[9] ;
  wire \user_io_in[0] ;
  wire \user_io_in[10] ;
  wire \user_io_in[11] ;
  wire \user_io_in[12] ;
  wire \user_io_in[13] ;
  wire \user_io_in[14] ;
  wire \user_io_in[15] ;
  wire \user_io_in[16] ;
  wire \user_io_in[17] ;
  wire \user_io_in[18] ;
  wire \user_io_in[19] ;
  wire \user_io_in[1] ;
  wire \user_io_in[20] ;
  wire \user_io_in[21] ;
  wire \user_io_in[22] ;
  wire \user_io_in[23] ;
  wire \user_io_in[24] ;
  wire \user_io_in[25] ;
  wire \user_io_in[26] ;
  wire \user_io_in[27] ;
  wire \user_io_in[28] ;
  wire \user_io_in[29] ;
  wire \user_io_in[2] ;
  wire \user_io_in[30] ;
  wire \user_io_in[31] ;
  wire \user_io_in[32] ;
  wire \user_io_in[33] ;
  wire \user_io_in[34] ;
  wire \user_io_in[35] ;
  wire \user_io_in[36] ;
  wire \user_io_in[37] ;
  wire \user_io_in[3] ;
  wire \user_io_in[4] ;
  wire \user_io_in[5] ;
  wire \user_io_in[6] ;
  wire \user_io_in[7] ;
  wire \user_io_in[8] ;
  wire \user_io_in[9] ;
  wire \user_io_oeb[0] ;
  wire \user_io_oeb[10] ;
  wire \user_io_oeb[11] ;
  wire \user_io_oeb[12] ;
  wire \user_io_oeb[13] ;
  wire \user_io_oeb[14] ;
  wire \user_io_oeb[15] ;
  wire \user_io_oeb[16] ;
  wire \user_io_oeb[17] ;
  wire \user_io_oeb[18] ;
  wire \user_io_oeb[19] ;
  wire \user_io_oeb[1] ;
  wire \user_io_oeb[20] ;
  wire \user_io_oeb[21] ;
  wire \user_io_oeb[22] ;
  wire \user_io_oeb[23] ;
  wire \user_io_oeb[24] ;
  wire \user_io_oeb[25] ;
  wire \user_io_oeb[26] ;
  wire \user_io_oeb[27] ;
  wire \user_io_oeb[28] ;
  wire \user_io_oeb[29] ;
  wire \user_io_oeb[2] ;
  wire \user_io_oeb[30] ;
  wire \user_io_oeb[31] ;
  wire \user_io_oeb[32] ;
  wire \user_io_oeb[33] ;
  wire \user_io_oeb[34] ;
  wire \user_io_oeb[35] ;
  wire \user_io_oeb[36] ;
  wire \user_io_oeb[37] ;
  wire \user_io_oeb[3] ;
  wire \user_io_oeb[4] ;
  wire \user_io_oeb[5] ;
  wire \user_io_oeb[6] ;
  wire \user_io_oeb[7] ;
  wire \user_io_oeb[8] ;
  wire \user_io_oeb[9] ;
  wire \user_io_out[0] ;
  wire \user_io_out[10] ;
  wire \user_io_out[11] ;
  wire \user_io_out[12] ;
  wire \user_io_out[13] ;
  wire \user_io_out[14] ;
  wire \user_io_out[15] ;
  wire \user_io_out[16] ;
  wire \user_io_out[17] ;
  wire \user_io_out[18] ;
  wire \user_io_out[19] ;
  wire \user_io_out[1] ;
  wire \user_io_out[20] ;
  wire \user_io_out[21] ;
  wire \user_io_out[22] ;
  wire \user_io_out[23] ;
  wire \user_io_out[24] ;
  wire \user_io_out[25] ;
  wire \user_io_out[26] ;
  wire \user_io_out[27] ;
  wire \user_io_out[28] ;
  wire \user_io_out[29] ;
  wire \user_io_out[2] ;
  wire \user_io_out[30] ;
  wire \user_io_out[31] ;
  wire \user_io_out[32] ;
  wire \user_io_out[33] ;
  wire \user_io_out[34] ;
  wire \user_io_out[35] ;
  wire \user_io_out[36] ;
  wire \user_io_out[37] ;
  wire \user_io_out[3] ;
  wire \user_io_out[4] ;
  wire \user_io_out[5] ;
  wire \user_io_out[6] ;
  wire \user_io_out[7] ;
  wire \user_io_out[8] ;
  wire \user_io_out[9] ;
  inout vccd;
  inout vccd1;
  inout vccd2;
  inout vdda;
  inout vdda1;
  inout vdda2;
  inout vddio;
  inout vssa;
  inout vssa1;
  inout vssa2;
  inout vssd;
  inout vssd1;
  inout vssd2;
  inout vssio;
  wire xbar_ack_i_core;
  wire \xbar_adr_o_core[0] ;
  wire \xbar_adr_o_core[10] ;
  wire \xbar_adr_o_core[11] ;
  wire \xbar_adr_o_core[12] ;
  wire \xbar_adr_o_core[13] ;
  wire \xbar_adr_o_core[14] ;
  wire \xbar_adr_o_core[15] ;
  wire \xbar_adr_o_core[16] ;
  wire \xbar_adr_o_core[17] ;
  wire \xbar_adr_o_core[18] ;
  wire \xbar_adr_o_core[19] ;
  wire \xbar_adr_o_core[1] ;
  wire \xbar_adr_o_core[20] ;
  wire \xbar_adr_o_core[21] ;
  wire \xbar_adr_o_core[22] ;
  wire \xbar_adr_o_core[23] ;
  wire \xbar_adr_o_core[24] ;
  wire \xbar_adr_o_core[25] ;
  wire \xbar_adr_o_core[26] ;
  wire \xbar_adr_o_core[27] ;
  wire \xbar_adr_o_core[28] ;
  wire \xbar_adr_o_core[29] ;
  wire \xbar_adr_o_core[2] ;
  wire \xbar_adr_o_core[30] ;
  wire \xbar_adr_o_core[31] ;
  wire \xbar_adr_o_core[3] ;
  wire \xbar_adr_o_core[4] ;
  wire \xbar_adr_o_core[5] ;
  wire \xbar_adr_o_core[6] ;
  wire \xbar_adr_o_core[7] ;
  wire \xbar_adr_o_core[8] ;
  wire \xbar_adr_o_core[9] ;
  wire xbar_cyc_o_core;
  wire \xbar_dat_i_core[0] ;
  wire \xbar_dat_i_core[10] ;
  wire \xbar_dat_i_core[11] ;
  wire \xbar_dat_i_core[12] ;
  wire \xbar_dat_i_core[13] ;
  wire \xbar_dat_i_core[14] ;
  wire \xbar_dat_i_core[15] ;
  wire \xbar_dat_i_core[16] ;
  wire \xbar_dat_i_core[17] ;
  wire \xbar_dat_i_core[18] ;
  wire \xbar_dat_i_core[19] ;
  wire \xbar_dat_i_core[1] ;
  wire \xbar_dat_i_core[20] ;
  wire \xbar_dat_i_core[21] ;
  wire \xbar_dat_i_core[22] ;
  wire \xbar_dat_i_core[23] ;
  wire \xbar_dat_i_core[24] ;
  wire \xbar_dat_i_core[25] ;
  wire \xbar_dat_i_core[26] ;
  wire \xbar_dat_i_core[27] ;
  wire \xbar_dat_i_core[28] ;
  wire \xbar_dat_i_core[29] ;
  wire \xbar_dat_i_core[2] ;
  wire \xbar_dat_i_core[30] ;
  wire \xbar_dat_i_core[31] ;
  wire \xbar_dat_i_core[3] ;
  wire \xbar_dat_i_core[4] ;
  wire \xbar_dat_i_core[5] ;
  wire \xbar_dat_i_core[6] ;
  wire \xbar_dat_i_core[7] ;
  wire \xbar_dat_i_core[8] ;
  wire \xbar_dat_i_core[9] ;
  wire \xbar_dat_o_core[0] ;
  wire \xbar_dat_o_core[10] ;
  wire \xbar_dat_o_core[11] ;
  wire \xbar_dat_o_core[12] ;
  wire \xbar_dat_o_core[13] ;
  wire \xbar_dat_o_core[14] ;
  wire \xbar_dat_o_core[15] ;
  wire \xbar_dat_o_core[16] ;
  wire \xbar_dat_o_core[17] ;
  wire \xbar_dat_o_core[18] ;
  wire \xbar_dat_o_core[19] ;
  wire \xbar_dat_o_core[1] ;
  wire \xbar_dat_o_core[20] ;
  wire \xbar_dat_o_core[21] ;
  wire \xbar_dat_o_core[22] ;
  wire \xbar_dat_o_core[23] ;
  wire \xbar_dat_o_core[24] ;
  wire \xbar_dat_o_core[25] ;
  wire \xbar_dat_o_core[26] ;
  wire \xbar_dat_o_core[27] ;
  wire \xbar_dat_o_core[28] ;
  wire \xbar_dat_o_core[29] ;
  wire \xbar_dat_o_core[2] ;
  wire \xbar_dat_o_core[30] ;
  wire \xbar_dat_o_core[31] ;
  wire \xbar_dat_o_core[3] ;
  wire \xbar_dat_o_core[4] ;
  wire \xbar_dat_o_core[5] ;
  wire \xbar_dat_o_core[6] ;
  wire \xbar_dat_o_core[7] ;
  wire \xbar_dat_o_core[8] ;
  wire \xbar_dat_o_core[9] ;
  wire \xbar_sel_o_core[0] ;
  wire \xbar_sel_o_core[1] ;
  wire \xbar_sel_o_core[2] ;
  wire \xbar_sel_o_core[3] ;
  wire xbar_stb_o_core;
  wire xbar_we_o_core;
  gpio_control_block \gpio_control_bidir[0]  (
    .mgmt_gpio_in(\mgmt_io_in[0] ),
    .mgmt_gpio_oeb(jtag_outenb),
    .mgmt_gpio_out(jtag_out),
    .pad_gpio_ana_en(\mprj_io_analog_en[0] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[0] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[0] ),
    .pad_gpio_dm({ \mprj_io_dm[2] , \mprj_io_dm[1] , \mprj_io_dm[0]  }),
    .pad_gpio_holdover(\mprj_io_holdover[0] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[0] ),
    .pad_gpio_in(\mprj_io_in[0] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[0] ),
    .pad_gpio_out(\mprj_io_out[0] ),
    .pad_gpio_outenb(\mprj_io_oeb[0] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[0] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[0] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link_shifted[0] ),
    .serial_data_out(\gpio_serial_link[0] ),
    .user_gpio_in(\user_io_in[0] ),
    .user_gpio_oeb(\user_io_oeb[0] ),
    .user_gpio_out(\user_io_out[0] )
  );
  gpio_control_block \gpio_control_bidir[1]  (
    .mgmt_gpio_in(\mgmt_io_in[1] ),
    .mgmt_gpio_oeb(sdo_outenb),
    .mgmt_gpio_out(sdo_out),
    .pad_gpio_ana_en(\mprj_io_analog_en[1] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[1] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[1] ),
    .pad_gpio_dm({ \mprj_io_dm[5] , \mprj_io_dm[4] , \mprj_io_dm[3]  }),
    .pad_gpio_holdover(\mprj_io_holdover[1] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[1] ),
    .pad_gpio_in(\mprj_io_in[1] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[1] ),
    .pad_gpio_out(\mprj_io_out[1] ),
    .pad_gpio_outenb(\mprj_io_oeb[1] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[1] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[1] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[0] ),
    .serial_data_out(\gpio_serial_link[1] ),
    .user_gpio_in(\user_io_in[1] ),
    .user_gpio_oeb(\user_io_oeb[1] ),
    .user_gpio_out(\user_io_out[1] )
  );
  gpio_control_block \gpio_control_in[10]  (
    .mgmt_gpio_in(\mgmt_io_in[10] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[10] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[10] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[10] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[10] ),
    .pad_gpio_dm({ \mprj_io_dm[32] , \mprj_io_dm[31] , \mprj_io_dm[30]  }),
    .pad_gpio_holdover(\mprj_io_holdover[10] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[10] ),
    .pad_gpio_in(\mprj_io_in[10] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[10] ),
    .pad_gpio_out(\mprj_io_out[10] ),
    .pad_gpio_outenb(\mprj_io_oeb[10] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[10] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[10] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[9] ),
    .serial_data_out(\gpio_serial_link[10] ),
    .user_gpio_in(\user_io_in[10] ),
    .user_gpio_oeb(\user_io_oeb[10] ),
    .user_gpio_out(\user_io_out[10] )
  );
  gpio_control_block \gpio_control_in[11]  (
    .mgmt_gpio_in(\mgmt_io_in[11] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[11] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[11] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[11] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[11] ),
    .pad_gpio_dm({ \mprj_io_dm[35] , \mprj_io_dm[34] , \mprj_io_dm[33]  }),
    .pad_gpio_holdover(\mprj_io_holdover[11] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[11] ),
    .pad_gpio_in(\mprj_io_in[11] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[11] ),
    .pad_gpio_out(\mprj_io_out[11] ),
    .pad_gpio_outenb(\mprj_io_oeb[11] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[11] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[11] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[10] ),
    .serial_data_out(\gpio_serial_link[11] ),
    .user_gpio_in(\user_io_in[11] ),
    .user_gpio_oeb(\user_io_oeb[11] ),
    .user_gpio_out(\user_io_out[11] )
  );
  gpio_control_block \gpio_control_in[12]  (
    .mgmt_gpio_in(\mgmt_io_in[12] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[12] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[12] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[12] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[12] ),
    .pad_gpio_dm({ \mprj_io_dm[38] , \mprj_io_dm[37] , \mprj_io_dm[36]  }),
    .pad_gpio_holdover(\mprj_io_holdover[12] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[12] ),
    .pad_gpio_in(\mprj_io_in[12] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[12] ),
    .pad_gpio_out(\mprj_io_out[12] ),
    .pad_gpio_outenb(\mprj_io_oeb[12] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[12] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[12] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[11] ),
    .serial_data_out(\gpio_serial_link[12] ),
    .user_gpio_in(\user_io_in[12] ),
    .user_gpio_oeb(\user_io_oeb[12] ),
    .user_gpio_out(\user_io_out[12] )
  );
  gpio_control_block \gpio_control_in[13]  (
    .mgmt_gpio_in(\mgmt_io_in[13] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[13] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[13] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[13] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[13] ),
    .pad_gpio_dm({ \mprj_io_dm[41] , \mprj_io_dm[40] , \mprj_io_dm[39]  }),
    .pad_gpio_holdover(\mprj_io_holdover[13] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[13] ),
    .pad_gpio_in(\mprj_io_in[13] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[13] ),
    .pad_gpio_out(\mprj_io_out[13] ),
    .pad_gpio_outenb(\mprj_io_oeb[13] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[13] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[13] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[12] ),
    .serial_data_out(\gpio_serial_link[13] ),
    .user_gpio_in(\user_io_in[13] ),
    .user_gpio_oeb(\user_io_oeb[13] ),
    .user_gpio_out(\user_io_out[13] )
  );
  gpio_control_block \gpio_control_in[14]  (
    .mgmt_gpio_in(\mgmt_io_in[14] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[14] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[14] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[14] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[14] ),
    .pad_gpio_dm({ \mprj_io_dm[44] , \mprj_io_dm[43] , \mprj_io_dm[42]  }),
    .pad_gpio_holdover(\mprj_io_holdover[14] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[14] ),
    .pad_gpio_in(\mprj_io_in[14] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[14] ),
    .pad_gpio_out(\mprj_io_out[14] ),
    .pad_gpio_outenb(\mprj_io_oeb[14] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[14] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[14] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[13] ),
    .serial_data_out(\gpio_serial_link[14] ),
    .user_gpio_in(\user_io_in[14] ),
    .user_gpio_oeb(\user_io_oeb[14] ),
    .user_gpio_out(\user_io_out[14] )
  );
  gpio_control_block \gpio_control_in[15]  (
    .mgmt_gpio_in(\mgmt_io_in[15] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[15] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[15] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[15] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[15] ),
    .pad_gpio_dm({ \mprj_io_dm[47] , \mprj_io_dm[46] , \mprj_io_dm[45]  }),
    .pad_gpio_holdover(\mprj_io_holdover[15] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[15] ),
    .pad_gpio_in(\mprj_io_in[15] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[15] ),
    .pad_gpio_out(\mprj_io_out[15] ),
    .pad_gpio_outenb(\mprj_io_oeb[15] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[15] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[15] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[14] ),
    .serial_data_out(\gpio_serial_link[15] ),
    .user_gpio_in(\user_io_in[15] ),
    .user_gpio_oeb(\user_io_oeb[15] ),
    .user_gpio_out(\user_io_out[15] )
  );
  gpio_control_block \gpio_control_in[16]  (
    .mgmt_gpio_in(\mgmt_io_in[16] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[16] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[16] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[16] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[16] ),
    .pad_gpio_dm({ \mprj_io_dm[50] , \mprj_io_dm[49] , \mprj_io_dm[48]  }),
    .pad_gpio_holdover(\mprj_io_holdover[16] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[16] ),
    .pad_gpio_in(\mprj_io_in[16] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[16] ),
    .pad_gpio_out(\mprj_io_out[16] ),
    .pad_gpio_outenb(\mprj_io_oeb[16] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[16] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[16] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[15] ),
    .serial_data_out(\gpio_serial_link[16] ),
    .user_gpio_in(\user_io_in[16] ),
    .user_gpio_oeb(\user_io_oeb[16] ),
    .user_gpio_out(\user_io_out[16] )
  );
  gpio_control_block \gpio_control_in[17]  (
    .mgmt_gpio_in(\mgmt_io_in[17] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[17] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[17] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[17] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[17] ),
    .pad_gpio_dm({ \mprj_io_dm[53] , \mprj_io_dm[52] , \mprj_io_dm[51]  }),
    .pad_gpio_holdover(\mprj_io_holdover[17] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[17] ),
    .pad_gpio_in(\mprj_io_in[17] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[17] ),
    .pad_gpio_out(\mprj_io_out[17] ),
    .pad_gpio_outenb(\mprj_io_oeb[17] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[17] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[17] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[16] ),
    .serial_data_out(\gpio_serial_link[17] ),
    .user_gpio_in(\user_io_in[17] ),
    .user_gpio_oeb(\user_io_oeb[17] ),
    .user_gpio_out(\user_io_out[17] )
  );
  gpio_control_block \gpio_control_in[18]  (
    .mgmt_gpio_in(\mgmt_io_in[18] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[18] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[18] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[18] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[18] ),
    .pad_gpio_dm({ \mprj_io_dm[56] , \mprj_io_dm[55] , \mprj_io_dm[54]  }),
    .pad_gpio_holdover(\mprj_io_holdover[18] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[18] ),
    .pad_gpio_in(\mprj_io_in[18] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[18] ),
    .pad_gpio_out(\mprj_io_out[18] ),
    .pad_gpio_outenb(\mprj_io_oeb[18] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[18] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[18] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[17] ),
    .serial_data_out(\gpio_serial_link[18] ),
    .user_gpio_in(\user_io_in[18] ),
    .user_gpio_oeb(\user_io_oeb[18] ),
    .user_gpio_out(\user_io_out[18] )
  );
  gpio_control_block \gpio_control_in[19]  (
    .mgmt_gpio_in(\mgmt_io_in[19] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[19] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[19] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[19] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[19] ),
    .pad_gpio_dm({ \mprj_io_dm[59] , \mprj_io_dm[58] , \mprj_io_dm[57]  }),
    .pad_gpio_holdover(\mprj_io_holdover[19] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[19] ),
    .pad_gpio_in(\mprj_io_in[19] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[19] ),
    .pad_gpio_out(\mprj_io_out[19] ),
    .pad_gpio_outenb(\mprj_io_oeb[19] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[19] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[19] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[18] ),
    .serial_data_out(\gpio_serial_link[19] ),
    .user_gpio_in(\user_io_in[19] ),
    .user_gpio_oeb(\user_io_oeb[19] ),
    .user_gpio_out(\user_io_out[19] )
  );
  gpio_control_block \gpio_control_in[20]  (
    .mgmt_gpio_in(\mgmt_io_in[20] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[20] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[20] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[20] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[20] ),
    .pad_gpio_dm({ \mprj_io_dm[62] , \mprj_io_dm[61] , \mprj_io_dm[60]  }),
    .pad_gpio_holdover(\mprj_io_holdover[20] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[20] ),
    .pad_gpio_in(\mprj_io_in[20] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[20] ),
    .pad_gpio_out(\mprj_io_out[20] ),
    .pad_gpio_outenb(\mprj_io_oeb[20] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[20] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[20] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[19] ),
    .serial_data_out(\gpio_serial_link[20] ),
    .user_gpio_in(\user_io_in[20] ),
    .user_gpio_oeb(\user_io_oeb[20] ),
    .user_gpio_out(\user_io_out[20] )
  );
  gpio_control_block \gpio_control_in[21]  (
    .mgmt_gpio_in(\mgmt_io_in[21] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[21] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[21] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[21] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[21] ),
    .pad_gpio_dm({ \mprj_io_dm[65] , \mprj_io_dm[64] , \mprj_io_dm[63]  }),
    .pad_gpio_holdover(\mprj_io_holdover[21] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[21] ),
    .pad_gpio_in(\mprj_io_in[21] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[21] ),
    .pad_gpio_out(\mprj_io_out[21] ),
    .pad_gpio_outenb(\mprj_io_oeb[21] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[21] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[21] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[20] ),
    .serial_data_out(\gpio_serial_link[21] ),
    .user_gpio_in(\user_io_in[21] ),
    .user_gpio_oeb(\user_io_oeb[21] ),
    .user_gpio_out(\user_io_out[21] )
  );
  gpio_control_block \gpio_control_in[22]  (
    .mgmt_gpio_in(\mgmt_io_in[22] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[22] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[22] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[22] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[22] ),
    .pad_gpio_dm({ \mprj_io_dm[68] , \mprj_io_dm[67] , \mprj_io_dm[66]  }),
    .pad_gpio_holdover(\mprj_io_holdover[22] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[22] ),
    .pad_gpio_in(\mprj_io_in[22] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[22] ),
    .pad_gpio_out(\mprj_io_out[22] ),
    .pad_gpio_outenb(\mprj_io_oeb[22] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[22] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[22] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[21] ),
    .serial_data_out(\gpio_serial_link[22] ),
    .user_gpio_in(\user_io_in[22] ),
    .user_gpio_oeb(\user_io_oeb[22] ),
    .user_gpio_out(\user_io_out[22] )
  );
  gpio_control_block \gpio_control_in[23]  (
    .mgmt_gpio_in(\mgmt_io_in[23] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[23] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[23] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[23] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[23] ),
    .pad_gpio_dm({ \mprj_io_dm[71] , \mprj_io_dm[70] , \mprj_io_dm[69]  }),
    .pad_gpio_holdover(\mprj_io_holdover[23] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[23] ),
    .pad_gpio_in(\mprj_io_in[23] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[23] ),
    .pad_gpio_out(\mprj_io_out[23] ),
    .pad_gpio_outenb(\mprj_io_oeb[23] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[23] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[23] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[22] ),
    .serial_data_out(\gpio_serial_link[23] ),
    .user_gpio_in(\user_io_in[23] ),
    .user_gpio_oeb(\user_io_oeb[23] ),
    .user_gpio_out(\user_io_out[23] )
  );
  gpio_control_block \gpio_control_in[24]  (
    .mgmt_gpio_in(\mgmt_io_in[24] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[24] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[24] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[24] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[24] ),
    .pad_gpio_dm({ \mprj_io_dm[74] , \mprj_io_dm[73] , \mprj_io_dm[72]  }),
    .pad_gpio_holdover(\mprj_io_holdover[24] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[24] ),
    .pad_gpio_in(\mprj_io_in[24] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[24] ),
    .pad_gpio_out(\mprj_io_out[24] ),
    .pad_gpio_outenb(\mprj_io_oeb[24] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[24] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[24] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[23] ),
    .serial_data_out(\gpio_serial_link[24] ),
    .user_gpio_in(\user_io_in[24] ),
    .user_gpio_oeb(\user_io_oeb[24] ),
    .user_gpio_out(\user_io_out[24] )
  );
  gpio_control_block \gpio_control_in[25]  (
    .mgmt_gpio_in(\mgmt_io_in[25] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[25] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[25] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[25] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[25] ),
    .pad_gpio_dm({ \mprj_io_dm[77] , \mprj_io_dm[76] , \mprj_io_dm[75]  }),
    .pad_gpio_holdover(\mprj_io_holdover[25] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[25] ),
    .pad_gpio_in(\mprj_io_in[25] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[25] ),
    .pad_gpio_out(\mprj_io_out[25] ),
    .pad_gpio_outenb(\mprj_io_oeb[25] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[25] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[25] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[24] ),
    .serial_data_out(\gpio_serial_link[25] ),
    .user_gpio_in(\user_io_in[25] ),
    .user_gpio_oeb(\user_io_oeb[25] ),
    .user_gpio_out(\user_io_out[25] )
  );
  gpio_control_block \gpio_control_in[26]  (
    .mgmt_gpio_in(\mgmt_io_in[26] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[26] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[26] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[26] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[26] ),
    .pad_gpio_dm({ \mprj_io_dm[80] , \mprj_io_dm[79] , \mprj_io_dm[78]  }),
    .pad_gpio_holdover(\mprj_io_holdover[26] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[26] ),
    .pad_gpio_in(\mprj_io_in[26] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[26] ),
    .pad_gpio_out(\mprj_io_out[26] ),
    .pad_gpio_outenb(\mprj_io_oeb[26] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[26] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[26] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[25] ),
    .serial_data_out(\gpio_serial_link[26] ),
    .user_gpio_in(\user_io_in[26] ),
    .user_gpio_oeb(\user_io_oeb[26] ),
    .user_gpio_out(\user_io_out[26] )
  );
  gpio_control_block \gpio_control_in[27]  (
    .mgmt_gpio_in(\mgmt_io_in[27] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[27] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[27] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[27] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[27] ),
    .pad_gpio_dm({ \mprj_io_dm[83] , \mprj_io_dm[82] , \mprj_io_dm[81]  }),
    .pad_gpio_holdover(\mprj_io_holdover[27] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[27] ),
    .pad_gpio_in(\mprj_io_in[27] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[27] ),
    .pad_gpio_out(\mprj_io_out[27] ),
    .pad_gpio_outenb(\mprj_io_oeb[27] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[27] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[27] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[26] ),
    .serial_data_out(\gpio_serial_link[27] ),
    .user_gpio_in(\user_io_in[27] ),
    .user_gpio_oeb(\user_io_oeb[27] ),
    .user_gpio_out(\user_io_out[27] )
  );
  gpio_control_block \gpio_control_in[28]  (
    .mgmt_gpio_in(\mgmt_io_in[28] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[28] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[28] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[28] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[28] ),
    .pad_gpio_dm({ \mprj_io_dm[86] , \mprj_io_dm[85] , \mprj_io_dm[84]  }),
    .pad_gpio_holdover(\mprj_io_holdover[28] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[28] ),
    .pad_gpio_in(\mprj_io_in[28] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[28] ),
    .pad_gpio_out(\mprj_io_out[28] ),
    .pad_gpio_outenb(\mprj_io_oeb[28] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[28] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[28] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[27] ),
    .serial_data_out(\gpio_serial_link[28] ),
    .user_gpio_in(\user_io_in[28] ),
    .user_gpio_oeb(\user_io_oeb[28] ),
    .user_gpio_out(\user_io_out[28] )
  );
  gpio_control_block \gpio_control_in[29]  (
    .mgmt_gpio_in(\mgmt_io_in[29] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[29] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[29] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[29] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[29] ),
    .pad_gpio_dm({ \mprj_io_dm[89] , \mprj_io_dm[88] , \mprj_io_dm[87]  }),
    .pad_gpio_holdover(\mprj_io_holdover[29] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[29] ),
    .pad_gpio_in(\mprj_io_in[29] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[29] ),
    .pad_gpio_out(\mprj_io_out[29] ),
    .pad_gpio_outenb(\mprj_io_oeb[29] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[29] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[29] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[28] ),
    .serial_data_out(\gpio_serial_link[29] ),
    .user_gpio_in(\user_io_in[29] ),
    .user_gpio_oeb(\user_io_oeb[29] ),
    .user_gpio_out(\user_io_out[29] )
  );
  gpio_control_block \gpio_control_in[2]  (
    .mgmt_gpio_in(\mgmt_io_in[2] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[2] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[2] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[2] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[2] ),
    .pad_gpio_dm({ \mprj_io_dm[8] , \mprj_io_dm[7] , \mprj_io_dm[6]  }),
    .pad_gpio_holdover(\mprj_io_holdover[2] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[2] ),
    .pad_gpio_in(\mprj_io_in[2] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[2] ),
    .pad_gpio_out(\mprj_io_out[2] ),
    .pad_gpio_outenb(\mprj_io_oeb[2] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[2] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[2] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[1] ),
    .serial_data_out(\gpio_serial_link[2] ),
    .user_gpio_in(\user_io_in[2] ),
    .user_gpio_oeb(\user_io_oeb[2] ),
    .user_gpio_out(\user_io_out[2] )
  );
  gpio_control_block \gpio_control_in[30]  (
    .mgmt_gpio_in(\mgmt_io_in[30] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[30] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[30] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[30] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[30] ),
    .pad_gpio_dm({ \mprj_io_dm[92] , \mprj_io_dm[91] , \mprj_io_dm[90]  }),
    .pad_gpio_holdover(\mprj_io_holdover[30] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[30] ),
    .pad_gpio_in(\mprj_io_in[30] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[30] ),
    .pad_gpio_out(\mprj_io_out[30] ),
    .pad_gpio_outenb(\mprj_io_oeb[30] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[30] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[30] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[29] ),
    .serial_data_out(\gpio_serial_link[30] ),
    .user_gpio_in(\user_io_in[30] ),
    .user_gpio_oeb(\user_io_oeb[30] ),
    .user_gpio_out(\user_io_out[30] )
  );
  gpio_control_block \gpio_control_in[31]  (
    .mgmt_gpio_in(\mgmt_io_in[31] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[31] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[31] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[31] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[31] ),
    .pad_gpio_dm({ \mprj_io_dm[95] , \mprj_io_dm[94] , \mprj_io_dm[93]  }),
    .pad_gpio_holdover(\mprj_io_holdover[31] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[31] ),
    .pad_gpio_in(\mprj_io_in[31] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[31] ),
    .pad_gpio_out(\mprj_io_out[31] ),
    .pad_gpio_outenb(\mprj_io_oeb[31] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[31] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[31] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[30] ),
    .serial_data_out(\gpio_serial_link[31] ),
    .user_gpio_in(\user_io_in[31] ),
    .user_gpio_oeb(\user_io_oeb[31] ),
    .user_gpio_out(\user_io_out[31] )
  );
  gpio_control_block \gpio_control_in[32]  (
    .mgmt_gpio_in(\mgmt_io_in[32] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[32] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[32] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[32] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[32] ),
    .pad_gpio_dm({ \mprj_io_dm[98] , \mprj_io_dm[97] , \mprj_io_dm[96]  }),
    .pad_gpio_holdover(\mprj_io_holdover[32] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[32] ),
    .pad_gpio_in(\mprj_io_in[32] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[32] ),
    .pad_gpio_out(\mprj_io_out[32] ),
    .pad_gpio_outenb(\mprj_io_oeb[32] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[32] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[32] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[31] ),
    .serial_data_out(\gpio_serial_link[32] ),
    .user_gpio_in(\user_io_in[32] ),
    .user_gpio_oeb(\user_io_oeb[32] ),
    .user_gpio_out(\user_io_out[32] )
  );
  gpio_control_block \gpio_control_in[33]  (
    .mgmt_gpio_in(\mgmt_io_in[33] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[33] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[33] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[33] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[33] ),
    .pad_gpio_dm({ \mprj_io_dm[101] , \mprj_io_dm[100] , \mprj_io_dm[99]  }),
    .pad_gpio_holdover(\mprj_io_holdover[33] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[33] ),
    .pad_gpio_in(\mprj_io_in[33] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[33] ),
    .pad_gpio_out(\mprj_io_out[33] ),
    .pad_gpio_outenb(\mprj_io_oeb[33] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[33] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[33] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[32] ),
    .serial_data_out(\gpio_serial_link[33] ),
    .user_gpio_in(\user_io_in[33] ),
    .user_gpio_oeb(\user_io_oeb[33] ),
    .user_gpio_out(\user_io_out[33] )
  );
  gpio_control_block \gpio_control_in[34]  (
    .mgmt_gpio_in(\mgmt_io_in[34] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[34] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[34] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[34] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[34] ),
    .pad_gpio_dm({ \mprj_io_dm[104] , \mprj_io_dm[103] , \mprj_io_dm[102]  }),
    .pad_gpio_holdover(\mprj_io_holdover[34] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[34] ),
    .pad_gpio_in(\mprj_io_in[34] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[34] ),
    .pad_gpio_out(\mprj_io_out[34] ),
    .pad_gpio_outenb(\mprj_io_oeb[34] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[34] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[34] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[33] ),
    .serial_data_out(\gpio_serial_link[34] ),
    .user_gpio_in(\user_io_in[34] ),
    .user_gpio_oeb(\user_io_oeb[34] ),
    .user_gpio_out(\user_io_out[34] )
  );
  gpio_control_block \gpio_control_in[35]  (
    .mgmt_gpio_in(\mgmt_io_in[35] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[35] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[35] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[35] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[35] ),
    .pad_gpio_dm({ \mprj_io_dm[107] , \mprj_io_dm[106] , \mprj_io_dm[105]  }),
    .pad_gpio_holdover(\mprj_io_holdover[35] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[35] ),
    .pad_gpio_in(\mprj_io_in[35] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[35] ),
    .pad_gpio_out(\mprj_io_out[35] ),
    .pad_gpio_outenb(\mprj_io_oeb[35] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[35] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[35] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[34] ),
    .serial_data_out(\gpio_serial_link[35] ),
    .user_gpio_in(\user_io_in[35] ),
    .user_gpio_oeb(\user_io_oeb[35] ),
    .user_gpio_out(\user_io_out[35] )
  );
  gpio_control_block \gpio_control_in[36]  (
    .mgmt_gpio_in(\mgmt_io_in[36] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[36] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[36] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[36] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[36] ),
    .pad_gpio_dm({ \mprj_io_dm[110] , \mprj_io_dm[109] , \mprj_io_dm[108]  }),
    .pad_gpio_holdover(\mprj_io_holdover[36] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[36] ),
    .pad_gpio_in(\mprj_io_in[36] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[36] ),
    .pad_gpio_out(\mprj_io_out[36] ),
    .pad_gpio_outenb(\mprj_io_oeb[36] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[36] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[36] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[35] ),
    .serial_data_out(\gpio_serial_link[36] ),
    .user_gpio_in(\user_io_in[36] ),
    .user_gpio_oeb(\user_io_oeb[36] ),
    .user_gpio_out(\user_io_out[36] )
  );
  gpio_control_block \gpio_control_in[37]  (
    .mgmt_gpio_in(\mgmt_io_in[37] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[37] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[37] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[37] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[37] ),
    .pad_gpio_dm({ \mprj_io_dm[113] , \mprj_io_dm[112] , \mprj_io_dm[111]  }),
    .pad_gpio_holdover(\mprj_io_holdover[37] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[37] ),
    .pad_gpio_in(\mprj_io_in[37] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[37] ),
    .pad_gpio_out(\mprj_io_out[37] ),
    .pad_gpio_outenb(\mprj_io_oeb[37] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[37] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[37] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[36] ),
    .serial_data_out(\gpio_serial_link[37] ),
    .user_gpio_in(\user_io_in[37] ),
    .user_gpio_oeb(\user_io_oeb[37] ),
    .user_gpio_out(\user_io_out[37] )
  );
  gpio_control_block \gpio_control_in[3]  (
    .mgmt_gpio_in(\mgmt_io_in[3] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[3] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[3] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[3] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[3] ),
    .pad_gpio_dm({ \mprj_io_dm[11] , \mprj_io_dm[10] , \mprj_io_dm[9]  }),
    .pad_gpio_holdover(\mprj_io_holdover[3] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[3] ),
    .pad_gpio_in(\mprj_io_in[3] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[3] ),
    .pad_gpio_out(\mprj_io_out[3] ),
    .pad_gpio_outenb(\mprj_io_oeb[3] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[3] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[3] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[2] ),
    .serial_data_out(\gpio_serial_link[3] ),
    .user_gpio_in(\user_io_in[3] ),
    .user_gpio_oeb(\user_io_oeb[3] ),
    .user_gpio_out(\user_io_out[3] )
  );
  gpio_control_block \gpio_control_in[4]  (
    .mgmt_gpio_in(\mgmt_io_in[4] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[4] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[4] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[4] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[4] ),
    .pad_gpio_dm({ \mprj_io_dm[14] , \mprj_io_dm[13] , \mprj_io_dm[12]  }),
    .pad_gpio_holdover(\mprj_io_holdover[4] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[4] ),
    .pad_gpio_in(\mprj_io_in[4] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[4] ),
    .pad_gpio_out(\mprj_io_out[4] ),
    .pad_gpio_outenb(\mprj_io_oeb[4] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[4] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[4] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[3] ),
    .serial_data_out(\gpio_serial_link[4] ),
    .user_gpio_in(\user_io_in[4] ),
    .user_gpio_oeb(\user_io_oeb[4] ),
    .user_gpio_out(\user_io_out[4] )
  );
  gpio_control_block \gpio_control_in[5]  (
    .mgmt_gpio_in(\mgmt_io_in[5] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[5] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[5] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[5] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[5] ),
    .pad_gpio_dm({ \mprj_io_dm[17] , \mprj_io_dm[16] , \mprj_io_dm[15]  }),
    .pad_gpio_holdover(\mprj_io_holdover[5] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[5] ),
    .pad_gpio_in(\mprj_io_in[5] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[5] ),
    .pad_gpio_out(\mprj_io_out[5] ),
    .pad_gpio_outenb(\mprj_io_oeb[5] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[5] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[5] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[4] ),
    .serial_data_out(\gpio_serial_link[5] ),
    .user_gpio_in(\user_io_in[5] ),
    .user_gpio_oeb(\user_io_oeb[5] ),
    .user_gpio_out(\user_io_out[5] )
  );
  gpio_control_block \gpio_control_in[6]  (
    .mgmt_gpio_in(\mgmt_io_in[6] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[6] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[6] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[6] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[6] ),
    .pad_gpio_dm({ \mprj_io_dm[20] , \mprj_io_dm[19] , \mprj_io_dm[18]  }),
    .pad_gpio_holdover(\mprj_io_holdover[6] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[6] ),
    .pad_gpio_in(\mprj_io_in[6] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[6] ),
    .pad_gpio_out(\mprj_io_out[6] ),
    .pad_gpio_outenb(\mprj_io_oeb[6] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[6] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[6] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[5] ),
    .serial_data_out(\gpio_serial_link[6] ),
    .user_gpio_in(\user_io_in[6] ),
    .user_gpio_oeb(\user_io_oeb[6] ),
    .user_gpio_out(\user_io_out[6] )
  );
  gpio_control_block \gpio_control_in[7]  (
    .mgmt_gpio_in(\mgmt_io_in[7] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[7] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[7] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[7] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[7] ),
    .pad_gpio_dm({ \mprj_io_dm[23] , \mprj_io_dm[22] , \mprj_io_dm[21]  }),
    .pad_gpio_holdover(\mprj_io_holdover[7] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[7] ),
    .pad_gpio_in(\mprj_io_in[7] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[7] ),
    .pad_gpio_out(\mprj_io_out[7] ),
    .pad_gpio_outenb(\mprj_io_oeb[7] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[7] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[7] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[6] ),
    .serial_data_out(\gpio_serial_link[7] ),
    .user_gpio_in(\user_io_in[7] ),
    .user_gpio_oeb(\user_io_oeb[7] ),
    .user_gpio_out(\user_io_out[7] )
  );
  gpio_control_block \gpio_control_in[8]  (
    .mgmt_gpio_in(\mgmt_io_in[8] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[8] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[8] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[8] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[8] ),
    .pad_gpio_dm({ \mprj_io_dm[26] , \mprj_io_dm[25] , \mprj_io_dm[24]  }),
    .pad_gpio_holdover(\mprj_io_holdover[8] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[8] ),
    .pad_gpio_in(\mprj_io_in[8] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[8] ),
    .pad_gpio_out(\mprj_io_out[8] ),
    .pad_gpio_outenb(\mprj_io_oeb[8] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[8] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[8] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[7] ),
    .serial_data_out(\gpio_serial_link[8] ),
    .user_gpio_in(\user_io_in[8] ),
    .user_gpio_oeb(\user_io_oeb[8] ),
    .user_gpio_out(\user_io_out[8] )
  );
  gpio_control_block \gpio_control_in[9]  (
    .mgmt_gpio_in(\mgmt_io_in[9] ),
    .mgmt_gpio_oeb(1'b1),
    .mgmt_gpio_out(\mgmt_io_in[9] ),
    .pad_gpio_ana_en(\mprj_io_analog_en[9] ),
    .pad_gpio_ana_pol(\mprj_io_analog_pol[9] ),
    .pad_gpio_ana_sel(\mprj_io_analog_sel[9] ),
    .pad_gpio_dm({ \mprj_io_dm[29] , \mprj_io_dm[28] , \mprj_io_dm[27]  }),
    .pad_gpio_holdover(\mprj_io_holdover[9] ),
    .pad_gpio_ib_mode_sel(\mprj_io_ib_mode_sel[9] ),
    .pad_gpio_in(\mprj_io_in[9] ),
    .pad_gpio_inenb(\mprj_io_inp_dis[9] ),
    .pad_gpio_out(\mprj_io_out[9] ),
    .pad_gpio_outenb(\mprj_io_oeb[9] ),
    .pad_gpio_slow_sel(\mprj_io_slow_sel[9] ),
    .pad_gpio_vtrip_sel(\mprj_io_vtrip_sel[9] ),
    .resetn(mprj_io_loader_resetn),
    .serial_clock(mprj_io_loader_clock),
    .serial_data_in(\gpio_serial_link[8] ),
    .serial_data_out(\gpio_serial_link[9] ),
    .user_gpio_in(\user_io_in[9] ),
    .user_gpio_oeb(\user_io_oeb[9] ),
    .user_gpio_out(\user_io_out[9] )
  );
  mgmt_protect mgmt_buffers (
    .caravel_clk(caravel_clk),
    .caravel_clk2(caravel_clk2),
    .caravel_rstn(caravel_rstn),
    .la_data_in_core({ \la_data_in_user[127] , \la_data_in_user[126] , \la_data_in_user[125] , \la_data_in_user[124] , \la_data_in_user[123] , \la_data_in_user[122] , \la_data_in_user[121] , \la_data_in_user[120] , \la_data_in_user[119] , \la_data_in_user[118] , \la_data_in_user[117] , \la_data_in_user[116] , \la_data_in_user[115] , \la_data_in_user[114] , \la_data_in_user[113] , \la_data_in_user[112] , \la_data_in_user[111] , \la_data_in_user[110] , \la_data_in_user[109] , \la_data_in_user[108] , \la_data_in_user[107] , \la_data_in_user[106] , \la_data_in_user[105] , \la_data_in_user[104] , \la_data_in_user[103] , \la_data_in_user[102] , \la_data_in_user[101] , \la_data_in_user[100] , \la_data_in_user[99] , \la_data_in_user[98] , \la_data_in_user[97] , \la_data_in_user[96] , \la_data_in_user[95] , \la_data_in_user[94] , \la_data_in_user[93] , \la_data_in_user[92] , \la_data_in_user[91] , \la_data_in_user[90] , \la_data_in_user[89] , \la_data_in_user[88] , \la_data_in_user[87] , \la_data_in_user[86] , \la_data_in_user[85] , \la_data_in_user[84] , \la_data_in_user[83] , \la_data_in_user[82] , \la_data_in_user[81] , \la_data_in_user[80] , \la_data_in_user[79] , \la_data_in_user[78] , \la_data_in_user[77] , \la_data_in_user[76] , \la_data_in_user[75] , \la_data_in_user[74] , \la_data_in_user[73] , \la_data_in_user[72] , \la_data_in_user[71] , \la_data_in_user[70] , \la_data_in_user[69] , \la_data_in_user[68] , \la_data_in_user[67] , \la_data_in_user[66] , \la_data_in_user[65] , \la_data_in_user[64] , \la_data_in_user[63] , \la_data_in_user[62] , \la_data_in_user[61] , \la_data_in_user[60] , \la_data_in_user[59] , \la_data_in_user[58] , \la_data_in_user[57] , \la_data_in_user[56] , \la_data_in_user[55] , \la_data_in_user[54] , \la_data_in_user[53] , \la_data_in_user[52] , \la_data_in_user[51] , \la_data_in_user[50] , \la_data_in_user[49] , \la_data_in_user[48] , \la_data_in_user[47] , \la_data_in_user[46] , \la_data_in_user[45] , \la_data_in_user[44] , \la_data_in_user[43] , \la_data_in_user[42] , \la_data_in_user[41] , \la_data_in_user[40] , \la_data_in_user[39] , \la_data_in_user[38] , \la_data_in_user[37] , \la_data_in_user[36] , \la_data_in_user[35] , \la_data_in_user[34] , \la_data_in_user[33] , \la_data_in_user[32] , \la_data_in_user[31] , \la_data_in_user[30] , \la_data_in_user[29] , \la_data_in_user[28] , \la_data_in_user[27] , \la_data_in_user[26] , \la_data_in_user[25] , \la_data_in_user[24] , \la_data_in_user[23] , \la_data_in_user[22] , \la_data_in_user[21] , \la_data_in_user[20] , \la_data_in_user[19] , \la_data_in_user[18] , \la_data_in_user[17] , \la_data_in_user[16] , \la_data_in_user[15] , \la_data_in_user[14] , \la_data_in_user[13] , \la_data_in_user[12] , \la_data_in_user[11] , \la_data_in_user[10] , \la_data_in_user[9] , \la_data_in_user[8] , \la_data_in_user[7] , \la_data_in_user[6] , \la_data_in_user[5] , \la_data_in_user[4] , \la_data_in_user[3] , \la_data_in_user[2] , \la_data_in_user[1] , \la_data_in_user[0]  }),
    .la_data_in_mprj({ \la_data_in_mprj[127] , \la_data_in_mprj[126] , \la_data_in_mprj[125] , \la_data_in_mprj[124] , \la_data_in_mprj[123] , \la_data_in_mprj[122] , \la_data_in_mprj[121] , \la_data_in_mprj[120] , \la_data_in_mprj[119] , \la_data_in_mprj[118] , \la_data_in_mprj[117] , \la_data_in_mprj[116] , \la_data_in_mprj[115] , \la_data_in_mprj[114] , \la_data_in_mprj[113] , \la_data_in_mprj[112] , \la_data_in_mprj[111] , \la_data_in_mprj[110] , \la_data_in_mprj[109] , \la_data_in_mprj[108] , \la_data_in_mprj[107] , \la_data_in_mprj[106] , \la_data_in_mprj[105] , \la_data_in_mprj[104] , \la_data_in_mprj[103] , \la_data_in_mprj[102] , \la_data_in_mprj[101] , \la_data_in_mprj[100] , \la_data_in_mprj[99] , \la_data_in_mprj[98] , \la_data_in_mprj[97] , \la_data_in_mprj[96] , \la_data_in_mprj[95] , \la_data_in_mprj[94] , \la_data_in_mprj[93] , \la_data_in_mprj[92] , \la_data_in_mprj[91] , \la_data_in_mprj[90] , \la_data_in_mprj[89] , \la_data_in_mprj[88] , \la_data_in_mprj[87] , \la_data_in_mprj[86] , \la_data_in_mprj[85] , \la_data_in_mprj[84] , \la_data_in_mprj[83] , \la_data_in_mprj[82] , \la_data_in_mprj[81] , \la_data_in_mprj[80] , \la_data_in_mprj[79] , \la_data_in_mprj[78] , \la_data_in_mprj[77] , \la_data_in_mprj[76] , \la_data_in_mprj[75] , \la_data_in_mprj[74] , \la_data_in_mprj[73] , \la_data_in_mprj[72] , \la_data_in_mprj[71] , \la_data_in_mprj[70] , \la_data_in_mprj[69] , \la_data_in_mprj[68] , \la_data_in_mprj[67] , \la_data_in_mprj[66] , \la_data_in_mprj[65] , \la_data_in_mprj[64] , \la_data_in_mprj[63] , \la_data_in_mprj[62] , \la_data_in_mprj[61] , \la_data_in_mprj[60] , \la_data_in_mprj[59] , \la_data_in_mprj[58] , \la_data_in_mprj[57] , \la_data_in_mprj[56] , \la_data_in_mprj[55] , \la_data_in_mprj[54] , \la_data_in_mprj[53] , \la_data_in_mprj[52] , \la_data_in_mprj[51] , \la_data_in_mprj[50] , \la_data_in_mprj[49] , \la_data_in_mprj[48] , \la_data_in_mprj[47] , \la_data_in_mprj[46] , \la_data_in_mprj[45] , \la_data_in_mprj[44] , \la_data_in_mprj[43] , \la_data_in_mprj[42] , \la_data_in_mprj[41] , \la_data_in_mprj[40] , \la_data_in_mprj[39] , \la_data_in_mprj[38] , \la_data_in_mprj[37] , \la_data_in_mprj[36] , \la_data_in_mprj[35] , \la_data_in_mprj[34] , \la_data_in_mprj[33] , \la_data_in_mprj[32] , \la_data_in_mprj[31] , \la_data_in_mprj[30] , \la_data_in_mprj[29] , \la_data_in_mprj[28] , \la_data_in_mprj[27] , \la_data_in_mprj[26] , \la_data_in_mprj[25] , \la_data_in_mprj[24] , \la_data_in_mprj[23] , \la_data_in_mprj[22] , \la_data_in_mprj[21] , \la_data_in_mprj[20] , \la_data_in_mprj[19] , \la_data_in_mprj[18] , \la_data_in_mprj[17] , \la_data_in_mprj[16] , \la_data_in_mprj[15] , \la_data_in_mprj[14] , \la_data_in_mprj[13] , \la_data_in_mprj[12] , \la_data_in_mprj[11] , \la_data_in_mprj[10] , \la_data_in_mprj[9] , \la_data_in_mprj[8] , \la_data_in_mprj[7] , \la_data_in_mprj[6] , \la_data_in_mprj[5] , \la_data_in_mprj[4] , \la_data_in_mprj[3] , \la_data_in_mprj[2] , \la_data_in_mprj[1] , \la_data_in_mprj[0]  }),
    .la_data_out_core({ \la_data_out_user[127] , \la_data_out_user[126] , \la_data_out_user[125] , \la_data_out_user[124] , \la_data_out_user[123] , \la_data_out_user[122] , \la_data_out_user[121] , \la_data_out_user[120] , \la_data_out_user[119] , \la_data_out_user[118] , \la_data_out_user[117] , \la_data_out_user[116] , \la_data_out_user[115] , \la_data_out_user[114] , \la_data_out_user[113] , \la_data_out_user[112] , \la_data_out_user[111] , \la_data_out_user[110] , \la_data_out_user[109] , \la_data_out_user[108] , \la_data_out_user[107] , \la_data_out_user[106] , \la_data_out_user[105] , \la_data_out_user[104] , \la_data_out_user[103] , \la_data_out_user[102] , \la_data_out_user[101] , \la_data_out_user[100] , \la_data_out_user[99] , \la_data_out_user[98] , \la_data_out_user[97] , \la_data_out_user[96] , \la_data_out_user[95] , \la_data_out_user[94] , \la_data_out_user[93] , \la_data_out_user[92] , \la_data_out_user[91] , \la_data_out_user[90] , \la_data_out_user[89] , \la_data_out_user[88] , \la_data_out_user[87] , \la_data_out_user[86] , \la_data_out_user[85] , \la_data_out_user[84] , \la_data_out_user[83] , \la_data_out_user[82] , \la_data_out_user[81] , \la_data_out_user[80] , \la_data_out_user[79] , \la_data_out_user[78] , \la_data_out_user[77] , \la_data_out_user[76] , \la_data_out_user[75] , \la_data_out_user[74] , \la_data_out_user[73] , \la_data_out_user[72] , \la_data_out_user[71] , \la_data_out_user[70] , \la_data_out_user[69] , \la_data_out_user[68] , \la_data_out_user[67] , \la_data_out_user[66] , \la_data_out_user[65] , \la_data_out_user[64] , \la_data_out_user[63] , \la_data_out_user[62] , \la_data_out_user[61] , \la_data_out_user[60] , \la_data_out_user[59] , \la_data_out_user[58] , \la_data_out_user[57] , \la_data_out_user[56] , \la_data_out_user[55] , \la_data_out_user[54] , \la_data_out_user[53] , \la_data_out_user[52] , \la_data_out_user[51] , \la_data_out_user[50] , \la_data_out_user[49] , \la_data_out_user[48] , \la_data_out_user[47] , \la_data_out_user[46] , \la_data_out_user[45] , \la_data_out_user[44] , \la_data_out_user[43] , \la_data_out_user[42] , \la_data_out_user[41] , \la_data_out_user[40] , \la_data_out_user[39] , \la_data_out_user[38] , \la_data_out_user[37] , \la_data_out_user[36] , \la_data_out_user[35] , \la_data_out_user[34] , \la_data_out_user[33] , \la_data_out_user[32] , \la_data_out_user[31] , \la_data_out_user[30] , \la_data_out_user[29] , \la_data_out_user[28] , \la_data_out_user[27] , \la_data_out_user[26] , \la_data_out_user[25] , \la_data_out_user[24] , \la_data_out_user[23] , \la_data_out_user[22] , \la_data_out_user[21] , \la_data_out_user[20] , \la_data_out_user[19] , \la_data_out_user[18] , \la_data_out_user[17] , \la_data_out_user[16] , \la_data_out_user[15] , \la_data_out_user[14] , \la_data_out_user[13] , \la_data_out_user[12] , \la_data_out_user[11] , \la_data_out_user[10] , \la_data_out_user[9] , \la_data_out_user[8] , \la_data_out_user[7] , \la_data_out_user[6] , \la_data_out_user[5] , \la_data_out_user[4] , \la_data_out_user[3] , \la_data_out_user[2] , \la_data_out_user[1] , \la_data_out_user[0]  }),
    .la_data_out_mprj({ \la_data_out_mprj[127] , \la_data_out_mprj[126] , \la_data_out_mprj[125] , \la_data_out_mprj[124] , \la_data_out_mprj[123] , \la_data_out_mprj[122] , \la_data_out_mprj[121] , \la_data_out_mprj[120] , \la_data_out_mprj[119] , \la_data_out_mprj[118] , \la_data_out_mprj[117] , \la_data_out_mprj[116] , \la_data_out_mprj[115] , \la_data_out_mprj[114] , \la_data_out_mprj[113] , \la_data_out_mprj[112] , \la_data_out_mprj[111] , \la_data_out_mprj[110] , \la_data_out_mprj[109] , \la_data_out_mprj[108] , \la_data_out_mprj[107] , \la_data_out_mprj[106] , \la_data_out_mprj[105] , \la_data_out_mprj[104] , \la_data_out_mprj[103] , \la_data_out_mprj[102] , \la_data_out_mprj[101] , \la_data_out_mprj[100] , \la_data_out_mprj[99] , \la_data_out_mprj[98] , \la_data_out_mprj[97] , \la_data_out_mprj[96] , \la_data_out_mprj[95] , \la_data_out_mprj[94] , \la_data_out_mprj[93] , \la_data_out_mprj[92] , \la_data_out_mprj[91] , \la_data_out_mprj[90] , \la_data_out_mprj[89] , \la_data_out_mprj[88] , \la_data_out_mprj[87] , \la_data_out_mprj[86] , \la_data_out_mprj[85] , \la_data_out_mprj[84] , \la_data_out_mprj[83] , \la_data_out_mprj[82] , \la_data_out_mprj[81] , \la_data_out_mprj[80] , \la_data_out_mprj[79] , \la_data_out_mprj[78] , \la_data_out_mprj[77] , \la_data_out_mprj[76] , \la_data_out_mprj[75] , \la_data_out_mprj[74] , \la_data_out_mprj[73] , \la_data_out_mprj[72] , \la_data_out_mprj[71] , \la_data_out_mprj[70] , \la_data_out_mprj[69] , \la_data_out_mprj[68] , \la_data_out_mprj[67] , \la_data_out_mprj[66] , \la_data_out_mprj[65] , \la_data_out_mprj[64] , \la_data_out_mprj[63] , \la_data_out_mprj[62] , \la_data_out_mprj[61] , \la_data_out_mprj[60] , \la_data_out_mprj[59] , \la_data_out_mprj[58] , \la_data_out_mprj[57] , \la_data_out_mprj[56] , \la_data_out_mprj[55] , \la_data_out_mprj[54] , \la_data_out_mprj[53] , \la_data_out_mprj[52] , \la_data_out_mprj[51] , \la_data_out_mprj[50] , \la_data_out_mprj[49] , \la_data_out_mprj[48] , \la_data_out_mprj[47] , \la_data_out_mprj[46] , \la_data_out_mprj[45] , \la_data_out_mprj[44] , \la_data_out_mprj[43] , \la_data_out_mprj[42] , \la_data_out_mprj[41] , \la_data_out_mprj[40] , \la_data_out_mprj[39] , \la_data_out_mprj[38] , \la_data_out_mprj[37] , \la_data_out_mprj[36] , \la_data_out_mprj[35] , \la_data_out_mprj[34] , \la_data_out_mprj[33] , \la_data_out_mprj[32] , \la_data_out_mprj[31] , \la_data_out_mprj[30] , \la_data_out_mprj[29] , \la_data_out_mprj[28] , \la_data_out_mprj[27] , \la_data_out_mprj[26] , \la_data_out_mprj[25] , \la_data_out_mprj[24] , \la_data_out_mprj[23] , \la_data_out_mprj[22] , \la_data_out_mprj[21] , \la_data_out_mprj[20] , \la_data_out_mprj[19] , \la_data_out_mprj[18] , \la_data_out_mprj[17] , \la_data_out_mprj[16] , \la_data_out_mprj[15] , \la_data_out_mprj[14] , \la_data_out_mprj[13] , \la_data_out_mprj[12] , \la_data_out_mprj[11] , \la_data_out_mprj[10] , \la_data_out_mprj[9] , \la_data_out_mprj[8] , \la_data_out_mprj[7] , \la_data_out_mprj[6] , \la_data_out_mprj[5] , \la_data_out_mprj[4] , \la_data_out_mprj[3] , \la_data_out_mprj[2] , \la_data_out_mprj[1] , \la_data_out_mprj[0]  }),
    .la_oen_core({ \la_oen_user[127] , \la_oen_user[126] , \la_oen_user[125] , \la_oen_user[124] , \la_oen_user[123] , \la_oen_user[122] , \la_oen_user[121] , \la_oen_user[120] , \la_oen_user[119] , \la_oen_user[118] , \la_oen_user[117] , \la_oen_user[116] , \la_oen_user[115] , \la_oen_user[114] , \la_oen_user[113] , \la_oen_user[112] , \la_oen_user[111] , \la_oen_user[110] , \la_oen_user[109] , \la_oen_user[108] , \la_oen_user[107] , \la_oen_user[106] , \la_oen_user[105] , \la_oen_user[104] , \la_oen_user[103] , \la_oen_user[102] , \la_oen_user[101] , \la_oen_user[100] , \la_oen_user[99] , \la_oen_user[98] , \la_oen_user[97] , \la_oen_user[96] , \la_oen_user[95] , \la_oen_user[94] , \la_oen_user[93] , \la_oen_user[92] , \la_oen_user[91] , \la_oen_user[90] , \la_oen_user[89] , \la_oen_user[88] , \la_oen_user[87] , \la_oen_user[86] , \la_oen_user[85] , \la_oen_user[84] , \la_oen_user[83] , \la_oen_user[82] , \la_oen_user[81] , \la_oen_user[80] , \la_oen_user[79] , \la_oen_user[78] , \la_oen_user[77] , \la_oen_user[76] , \la_oen_user[75] , \la_oen_user[74] , \la_oen_user[73] , \la_oen_user[72] , \la_oen_user[71] , \la_oen_user[70] , \la_oen_user[69] , \la_oen_user[68] , \la_oen_user[67] , \la_oen_user[66] , \la_oen_user[65] , \la_oen_user[64] , \la_oen_user[63] , \la_oen_user[62] , \la_oen_user[61] , \la_oen_user[60] , \la_oen_user[59] , \la_oen_user[58] , \la_oen_user[57] , \la_oen_user[56] , \la_oen_user[55] , \la_oen_user[54] , \la_oen_user[53] , \la_oen_user[52] , \la_oen_user[51] , \la_oen_user[50] , \la_oen_user[49] , \la_oen_user[48] , \la_oen_user[47] , \la_oen_user[46] , \la_oen_user[45] , \la_oen_user[44] , \la_oen_user[43] , \la_oen_user[42] , \la_oen_user[41] , \la_oen_user[40] , \la_oen_user[39] , \la_oen_user[38] , \la_oen_user[37] , \la_oen_user[36] , \la_oen_user[35] , \la_oen_user[34] , \la_oen_user[33] , \la_oen_user[32] , \la_oen_user[31] , \la_oen_user[30] , \la_oen_user[29] , \la_oen_user[28] , \la_oen_user[27] , \la_oen_user[26] , \la_oen_user[25] , \la_oen_user[24] , \la_oen_user[23] , \la_oen_user[22] , \la_oen_user[21] , \la_oen_user[20] , \la_oen_user[19] , \la_oen_user[18] , \la_oen_user[17] , \la_oen_user[16] , \la_oen_user[15] , \la_oen_user[14] , \la_oen_user[13] , \la_oen_user[12] , \la_oen_user[11] , \la_oen_user[10] , \la_oen_user[9] , \la_oen_user[8] , \la_oen_user[7] , \la_oen_user[6] , \la_oen_user[5] , \la_oen_user[4] , \la_oen_user[3] , \la_oen_user[2] , \la_oen_user[1] , \la_oen_user[0]  }),
    .la_oen_mprj({ \la_oen_mprj[127] , \la_oen_mprj[126] , \la_oen_mprj[125] , \la_oen_mprj[124] , \la_oen_mprj[123] , \la_oen_mprj[122] , \la_oen_mprj[121] , \la_oen_mprj[120] , \la_oen_mprj[119] , \la_oen_mprj[118] , \la_oen_mprj[117] , \la_oen_mprj[116] , \la_oen_mprj[115] , \la_oen_mprj[114] , \la_oen_mprj[113] , \la_oen_mprj[112] , \la_oen_mprj[111] , \la_oen_mprj[110] , \la_oen_mprj[109] , \la_oen_mprj[108] , \la_oen_mprj[107] , \la_oen_mprj[106] , \la_oen_mprj[105] , \la_oen_mprj[104] , \la_oen_mprj[103] , \la_oen_mprj[102] , \la_oen_mprj[101] , \la_oen_mprj[100] , \la_oen_mprj[99] , \la_oen_mprj[98] , \la_oen_mprj[97] , \la_oen_mprj[96] , \la_oen_mprj[95] , \la_oen_mprj[94] , \la_oen_mprj[93] , \la_oen_mprj[92] , \la_oen_mprj[91] , \la_oen_mprj[90] , \la_oen_mprj[89] , \la_oen_mprj[88] , \la_oen_mprj[87] , \la_oen_mprj[86] , \la_oen_mprj[85] , \la_oen_mprj[84] , \la_oen_mprj[83] , \la_oen_mprj[82] , \la_oen_mprj[81] , \la_oen_mprj[80] , \la_oen_mprj[79] , \la_oen_mprj[78] , \la_oen_mprj[77] , \la_oen_mprj[76] , \la_oen_mprj[75] , \la_oen_mprj[74] , \la_oen_mprj[73] , \la_oen_mprj[72] , \la_oen_mprj[71] , \la_oen_mprj[70] , \la_oen_mprj[69] , \la_oen_mprj[68] , \la_oen_mprj[67] , \la_oen_mprj[66] , \la_oen_mprj[65] , \la_oen_mprj[64] , \la_oen_mprj[63] , \la_oen_mprj[62] , \la_oen_mprj[61] , \la_oen_mprj[60] , \la_oen_mprj[59] , \la_oen_mprj[58] , \la_oen_mprj[57] , \la_oen_mprj[56] , \la_oen_mprj[55] , \la_oen_mprj[54] , \la_oen_mprj[53] , \la_oen_mprj[52] , \la_oen_mprj[51] , \la_oen_mprj[50] , \la_oen_mprj[49] , \la_oen_mprj[48] , \la_oen_mprj[47] , \la_oen_mprj[46] , \la_oen_mprj[45] , \la_oen_mprj[44] , \la_oen_mprj[43] , \la_oen_mprj[42] , \la_oen_mprj[41] , \la_oen_mprj[40] , \la_oen_mprj[39] , \la_oen_mprj[38] , \la_oen_mprj[37] , \la_oen_mprj[36] , \la_oen_mprj[35] , \la_oen_mprj[34] , \la_oen_mprj[33] , \la_oen_mprj[32] , \la_oen_mprj[31] , \la_oen_mprj[30] , \la_oen_mprj[29] , \la_oen_mprj[28] , \la_oen_mprj[27] , \la_oen_mprj[26] , \la_oen_mprj[25] , \la_oen_mprj[24] , \la_oen_mprj[23] , \la_oen_mprj[22] , \la_oen_mprj[21] , \la_oen_mprj[20] , \la_oen_mprj[19] , \la_oen_mprj[18] , \la_oen_mprj[17] , \la_oen_mprj[16] , \la_oen_mprj[15] , \la_oen_mprj[14] , \la_oen_mprj[13] , \la_oen_mprj[12] , \la_oen_mprj[11] , \la_oen_mprj[10] , \la_oen_mprj[9] , \la_oen_mprj[8] , \la_oen_mprj[7] , \la_oen_mprj[6] , \la_oen_mprj[5] , \la_oen_mprj[4] , \la_oen_mprj[3] , \la_oen_mprj[2] , \la_oen_mprj[1] , \la_oen_mprj[0]  }),
    .mprj_adr_o_core({ \mprj_adr_o_core[31] , \mprj_adr_o_core[30] , \mprj_adr_o_core[29] , \mprj_adr_o_core[28] , \mprj_adr_o_core[27] , \mprj_adr_o_core[26] , \mprj_adr_o_core[25] , \mprj_adr_o_core[24] , \mprj_adr_o_core[23] , \mprj_adr_o_core[22] , \mprj_adr_o_core[21] , \mprj_adr_o_core[20] , \mprj_adr_o_core[19] , \mprj_adr_o_core[18] , \mprj_adr_o_core[17] , \mprj_adr_o_core[16] , \mprj_adr_o_core[15] , \mprj_adr_o_core[14] , \mprj_adr_o_core[13] , \mprj_adr_o_core[12] , \mprj_adr_o_core[11] , \mprj_adr_o_core[10] , \mprj_adr_o_core[9] , \mprj_adr_o_core[8] , \mprj_adr_o_core[7] , \mprj_adr_o_core[6] , \mprj_adr_o_core[5] , \mprj_adr_o_core[4] , \mprj_adr_o_core[3] , \mprj_adr_o_core[2] , \mprj_adr_o_core[1] , \mprj_adr_o_core[0]  }),
    .mprj_adr_o_user({ \mprj_adr_o_user[31] , \mprj_adr_o_user[30] , \mprj_adr_o_user[29] , \mprj_adr_o_user[28] , \mprj_adr_o_user[27] , \mprj_adr_o_user[26] , \mprj_adr_o_user[25] , \mprj_adr_o_user[24] , \mprj_adr_o_user[23] , \mprj_adr_o_user[22] , \mprj_adr_o_user[21] , \mprj_adr_o_user[20] , \mprj_adr_o_user[19] , \mprj_adr_o_user[18] , \mprj_adr_o_user[17] , \mprj_adr_o_user[16] , \mprj_adr_o_user[15] , \mprj_adr_o_user[14] , \mprj_adr_o_user[13] , \mprj_adr_o_user[12] , \mprj_adr_o_user[11] , \mprj_adr_o_user[10] , \mprj_adr_o_user[9] , \mprj_adr_o_user[8] , \mprj_adr_o_user[7] , \mprj_adr_o_user[6] , \mprj_adr_o_user[5] , \mprj_adr_o_user[4] , \mprj_adr_o_user[3] , \mprj_adr_o_user[2] , \mprj_adr_o_user[1] , \mprj_adr_o_user[0]  }),
    .mprj_cyc_o_core(mprj_cyc_o_core),
    .mprj_cyc_o_user(mprj_cyc_o_user),
    .mprj_dat_o_core({ \mprj_dat_o_core[31] , \mprj_dat_o_core[30] , \mprj_dat_o_core[29] , \mprj_dat_o_core[28] , \mprj_dat_o_core[27] , \mprj_dat_o_core[26] , \mprj_dat_o_core[25] , \mprj_dat_o_core[24] , \mprj_dat_o_core[23] , \mprj_dat_o_core[22] , \mprj_dat_o_core[21] , \mprj_dat_o_core[20] , \mprj_dat_o_core[19] , \mprj_dat_o_core[18] , \mprj_dat_o_core[17] , \mprj_dat_o_core[16] , \mprj_dat_o_core[15] , \mprj_dat_o_core[14] , \mprj_dat_o_core[13] , \mprj_dat_o_core[12] , \mprj_dat_o_core[11] , \mprj_dat_o_core[10] , \mprj_dat_o_core[9] , \mprj_dat_o_core[8] , \mprj_dat_o_core[7] , \mprj_dat_o_core[6] , \mprj_dat_o_core[5] , \mprj_dat_o_core[4] , \mprj_dat_o_core[3] , \mprj_dat_o_core[2] , \mprj_dat_o_core[1] , \mprj_dat_o_core[0]  }),
    .mprj_dat_o_user({ \mprj_dat_o_user[31] , \mprj_dat_o_user[30] , \mprj_dat_o_user[29] , \mprj_dat_o_user[28] , \mprj_dat_o_user[27] , \mprj_dat_o_user[26] , \mprj_dat_o_user[25] , \mprj_dat_o_user[24] , \mprj_dat_o_user[23] , \mprj_dat_o_user[22] , \mprj_dat_o_user[21] , \mprj_dat_o_user[20] , \mprj_dat_o_user[19] , \mprj_dat_o_user[18] , \mprj_dat_o_user[17] , \mprj_dat_o_user[16] , \mprj_dat_o_user[15] , \mprj_dat_o_user[14] , \mprj_dat_o_user[13] , \mprj_dat_o_user[12] , \mprj_dat_o_user[11] , \mprj_dat_o_user[10] , \mprj_dat_o_user[9] , \mprj_dat_o_user[8] , \mprj_dat_o_user[7] , \mprj_dat_o_user[6] , \mprj_dat_o_user[5] , \mprj_dat_o_user[4] , \mprj_dat_o_user[3] , \mprj_dat_o_user[2] , \mprj_dat_o_user[1] , \mprj_dat_o_user[0]  }),
    .mprj_sel_o_core({ \mprj_sel_o_core[3] , \mprj_sel_o_core[2] , \mprj_sel_o_core[1] , \mprj_sel_o_core[0]  }),
    .mprj_sel_o_user({ \mprj_sel_o_user[3] , \mprj_sel_o_user[2] , \mprj_sel_o_user[1] , \mprj_sel_o_user[0]  }),
    .mprj_stb_o_core(mprj_stb_o_core),
    .mprj_stb_o_user(mprj_stb_o_user),
    .mprj_we_o_core(mprj_we_o_core),
    .mprj_we_o_user(mprj_we_o_user),
    .user1_vcc_powergood(mprj_vcc_pwrgood),
    .user1_vdd_powergood(mprj_vdd_pwrgood),
    .user2_vcc_powergood(mprj2_vcc_pwrgood),
    .user2_vdd_powergood(mprj2_vdd_pwrgood),
    .user_clock(mprj_clock),
    .user_clock2(mprj_clock2),
    .user_reset(mprj_reset),
    .user_resetn(mprj_resetn)
  );
  user_project_wrapper mprj (
    .analog_io({ \user_analog_io[30] , \user_analog_io[29] , \user_analog_io[28] , \user_analog_io[27] , \user_analog_io[26] , \user_analog_io[25] , \user_analog_io[24] , \user_analog_io[23] , \user_analog_io[22] , \user_analog_io[21] , \user_analog_io[20] , \user_analog_io[19] , \user_analog_io[18] , \user_analog_io[17] , \user_analog_io[16] , \user_analog_io[15] , \user_analog_io[14] , \user_analog_io[13] , \user_analog_io[12] , \user_analog_io[11] , \user_analog_io[10] , \user_analog_io[9] , \user_analog_io[8] , \user_analog_io[7] , \user_analog_io[6] , \user_analog_io[5] , \user_analog_io[4] , \user_analog_io[3] , \user_analog_io[2] , \user_analog_io[1] , \user_analog_io[0]  }),
    .io_in({ \user_io_in[37] , \user_io_in[36] , \user_io_in[35] , \user_io_in[34] , \user_io_in[33] , \user_io_in[32] , \user_io_in[31] , \user_io_in[30] , \user_io_in[29] , \user_io_in[28] , \user_io_in[27] , \user_io_in[26] , \user_io_in[25] , \user_io_in[24] , \user_io_in[23] , \user_io_in[22] , \user_io_in[21] , \user_io_in[20] , \user_io_in[19] , \user_io_in[18] , \user_io_in[17] , \user_io_in[16] , \user_io_in[15] , \user_io_in[14] , \user_io_in[13] , \user_io_in[12] , \user_io_in[11] , \user_io_in[10] , \user_io_in[9] , \user_io_in[8] , \user_io_in[7] , \user_io_in[6] , \user_io_in[5] , \user_io_in[4] , \user_io_in[3] , \user_io_in[2] , \user_io_in[1] , \user_io_in[0]  }),
    .io_oeb({ \user_io_oeb[37] , \user_io_oeb[36] , \user_io_oeb[35] , \user_io_oeb[34] , \user_io_oeb[33] , \user_io_oeb[32] , \user_io_oeb[31] , \user_io_oeb[30] , \user_io_oeb[29] , \user_io_oeb[28] , \user_io_oeb[27] , \user_io_oeb[26] , \user_io_oeb[25] , \user_io_oeb[24] , \user_io_oeb[23] , \user_io_oeb[22] , \user_io_oeb[21] , \user_io_oeb[20] , \user_io_oeb[19] , \user_io_oeb[18] , \user_io_oeb[17] , \user_io_oeb[16] , \user_io_oeb[15] , \user_io_oeb[14] , \user_io_oeb[13] , \user_io_oeb[12] , \user_io_oeb[11] , \user_io_oeb[10] , \user_io_oeb[9] , \user_io_oeb[8] , \user_io_oeb[7] , \user_io_oeb[6] , \user_io_oeb[5] , \user_io_oeb[4] , \user_io_oeb[3] , \user_io_oeb[2] , \user_io_oeb[1] , \user_io_oeb[0]  }),
    .io_out({ \user_io_out[37] , \user_io_out[36] , \user_io_out[35] , \user_io_out[34] , \user_io_out[33] , \user_io_out[32] , \user_io_out[31] , \user_io_out[30] , \user_io_out[29] , \user_io_out[28] , \user_io_out[27] , \user_io_out[26] , \user_io_out[25] , \user_io_out[24] , \user_io_out[23] , \user_io_out[22] , \user_io_out[21] , \user_io_out[20] , \user_io_out[19] , \user_io_out[18] , \user_io_out[17] , \user_io_out[16] , \user_io_out[15] , \user_io_out[14] , \user_io_out[13] , \user_io_out[12] , \user_io_out[11] , \user_io_out[10] , \user_io_out[9] , \user_io_out[8] , \user_io_out[7] , \user_io_out[6] , \user_io_out[5] , \user_io_out[4] , \user_io_out[3] , \user_io_out[2] , \user_io_out[1] , \user_io_out[0]  }),
    .la_data_in({ \la_data_in_user[127] , \la_data_in_user[126] , \la_data_in_user[125] , \la_data_in_user[124] , \la_data_in_user[123] , \la_data_in_user[122] , \la_data_in_user[121] , \la_data_in_user[120] , \la_data_in_user[119] , \la_data_in_user[118] , \la_data_in_user[117] , \la_data_in_user[116] , \la_data_in_user[115] , \la_data_in_user[114] , \la_data_in_user[113] , \la_data_in_user[112] , \la_data_in_user[111] , \la_data_in_user[110] , \la_data_in_user[109] , \la_data_in_user[108] , \la_data_in_user[107] , \la_data_in_user[106] , \la_data_in_user[105] , \la_data_in_user[104] , \la_data_in_user[103] , \la_data_in_user[102] , \la_data_in_user[101] , \la_data_in_user[100] , \la_data_in_user[99] , \la_data_in_user[98] , \la_data_in_user[97] , \la_data_in_user[96] , \la_data_in_user[95] , \la_data_in_user[94] , \la_data_in_user[93] , \la_data_in_user[92] , \la_data_in_user[91] , \la_data_in_user[90] , \la_data_in_user[89] , \la_data_in_user[88] , \la_data_in_user[87] , \la_data_in_user[86] , \la_data_in_user[85] , \la_data_in_user[84] , \la_data_in_user[83] , \la_data_in_user[82] , \la_data_in_user[81] , \la_data_in_user[80] , \la_data_in_user[79] , \la_data_in_user[78] , \la_data_in_user[77] , \la_data_in_user[76] , \la_data_in_user[75] , \la_data_in_user[74] , \la_data_in_user[73] , \la_data_in_user[72] , \la_data_in_user[71] , \la_data_in_user[70] , \la_data_in_user[69] , \la_data_in_user[68] , \la_data_in_user[67] , \la_data_in_user[66] , \la_data_in_user[65] , \la_data_in_user[64] , \la_data_in_user[63] , \la_data_in_user[62] , \la_data_in_user[61] , \la_data_in_user[60] , \la_data_in_user[59] , \la_data_in_user[58] , \la_data_in_user[57] , \la_data_in_user[56] , \la_data_in_user[55] , \la_data_in_user[54] , \la_data_in_user[53] , \la_data_in_user[52] , \la_data_in_user[51] , \la_data_in_user[50] , \la_data_in_user[49] , \la_data_in_user[48] , \la_data_in_user[47] , \la_data_in_user[46] , \la_data_in_user[45] , \la_data_in_user[44] , \la_data_in_user[43] , \la_data_in_user[42] , \la_data_in_user[41] , \la_data_in_user[40] , \la_data_in_user[39] , \la_data_in_user[38] , \la_data_in_user[37] , \la_data_in_user[36] , \la_data_in_user[35] , \la_data_in_user[34] , \la_data_in_user[33] , \la_data_in_user[32] , \la_data_in_user[31] , \la_data_in_user[30] , \la_data_in_user[29] , \la_data_in_user[28] , \la_data_in_user[27] , \la_data_in_user[26] , \la_data_in_user[25] , \la_data_in_user[24] , \la_data_in_user[23] , \la_data_in_user[22] , \la_data_in_user[21] , \la_data_in_user[20] , \la_data_in_user[19] , \la_data_in_user[18] , \la_data_in_user[17] , \la_data_in_user[16] , \la_data_in_user[15] , \la_data_in_user[14] , \la_data_in_user[13] , \la_data_in_user[12] , \la_data_in_user[11] , \la_data_in_user[10] , \la_data_in_user[9] , \la_data_in_user[8] , \la_data_in_user[7] , \la_data_in_user[6] , \la_data_in_user[5] , \la_data_in_user[4] , \la_data_in_user[3] , \la_data_in_user[2] , \la_data_in_user[1] , \la_data_in_user[0]  }),
    .la_data_out({ \la_data_out_user[127] , \la_data_out_user[126] , \la_data_out_user[125] , \la_data_out_user[124] , \la_data_out_user[123] , \la_data_out_user[122] , \la_data_out_user[121] , \la_data_out_user[120] , \la_data_out_user[119] , \la_data_out_user[118] , \la_data_out_user[117] , \la_data_out_user[116] , \la_data_out_user[115] , \la_data_out_user[114] , \la_data_out_user[113] , \la_data_out_user[112] , \la_data_out_user[111] , \la_data_out_user[110] , \la_data_out_user[109] , \la_data_out_user[108] , \la_data_out_user[107] , \la_data_out_user[106] , \la_data_out_user[105] , \la_data_out_user[104] , \la_data_out_user[103] , \la_data_out_user[102] , \la_data_out_user[101] , \la_data_out_user[100] , \la_data_out_user[99] , \la_data_out_user[98] , \la_data_out_user[97] , \la_data_out_user[96] , \la_data_out_user[95] , \la_data_out_user[94] , \la_data_out_user[93] , \la_data_out_user[92] , \la_data_out_user[91] , \la_data_out_user[90] , \la_data_out_user[89] , \la_data_out_user[88] , \la_data_out_user[87] , \la_data_out_user[86] , \la_data_out_user[85] , \la_data_out_user[84] , \la_data_out_user[83] , \la_data_out_user[82] , \la_data_out_user[81] , \la_data_out_user[80] , \la_data_out_user[79] , \la_data_out_user[78] , \la_data_out_user[77] , \la_data_out_user[76] , \la_data_out_user[75] , \la_data_out_user[74] , \la_data_out_user[73] , \la_data_out_user[72] , \la_data_out_user[71] , \la_data_out_user[70] , \la_data_out_user[69] , \la_data_out_user[68] , \la_data_out_user[67] , \la_data_out_user[66] , \la_data_out_user[65] , \la_data_out_user[64] , \la_data_out_user[63] , \la_data_out_user[62] , \la_data_out_user[61] , \la_data_out_user[60] , \la_data_out_user[59] , \la_data_out_user[58] , \la_data_out_user[57] , \la_data_out_user[56] , \la_data_out_user[55] , \la_data_out_user[54] , \la_data_out_user[53] , \la_data_out_user[52] , \la_data_out_user[51] , \la_data_out_user[50] , \la_data_out_user[49] , \la_data_out_user[48] , \la_data_out_user[47] , \la_data_out_user[46] , \la_data_out_user[45] , \la_data_out_user[44] , \la_data_out_user[43] , \la_data_out_user[42] , \la_data_out_user[41] , \la_data_out_user[40] , \la_data_out_user[39] , \la_data_out_user[38] , \la_data_out_user[37] , \la_data_out_user[36] , \la_data_out_user[35] , \la_data_out_user[34] , \la_data_out_user[33] , \la_data_out_user[32] , \la_data_out_user[31] , \la_data_out_user[30] , \la_data_out_user[29] , \la_data_out_user[28] , \la_data_out_user[27] , \la_data_out_user[26] , \la_data_out_user[25] , \la_data_out_user[24] , \la_data_out_user[23] , \la_data_out_user[22] , \la_data_out_user[21] , \la_data_out_user[20] , \la_data_out_user[19] , \la_data_out_user[18] , \la_data_out_user[17] , \la_data_out_user[16] , \la_data_out_user[15] , \la_data_out_user[14] , \la_data_out_user[13] , \la_data_out_user[12] , \la_data_out_user[11] , \la_data_out_user[10] , \la_data_out_user[9] , \la_data_out_user[8] , \la_data_out_user[7] , \la_data_out_user[6] , \la_data_out_user[5] , \la_data_out_user[4] , \la_data_out_user[3] , \la_data_out_user[2] , \la_data_out_user[1] , \la_data_out_user[0]  }),
    .la_oen({ \la_oen_user[127] , \la_oen_user[126] , \la_oen_user[125] , \la_oen_user[124] , \la_oen_user[123] , \la_oen_user[122] , \la_oen_user[121] , \la_oen_user[120] , \la_oen_user[119] , \la_oen_user[118] , \la_oen_user[117] , \la_oen_user[116] , \la_oen_user[115] , \la_oen_user[114] , \la_oen_user[113] , \la_oen_user[112] , \la_oen_user[111] , \la_oen_user[110] , \la_oen_user[109] , \la_oen_user[108] , \la_oen_user[107] , \la_oen_user[106] , \la_oen_user[105] , \la_oen_user[104] , \la_oen_user[103] , \la_oen_user[102] , \la_oen_user[101] , \la_oen_user[100] , \la_oen_user[99] , \la_oen_user[98] , \la_oen_user[97] , \la_oen_user[96] , \la_oen_user[95] , \la_oen_user[94] , \la_oen_user[93] , \la_oen_user[92] , \la_oen_user[91] , \la_oen_user[90] , \la_oen_user[89] , \la_oen_user[88] , \la_oen_user[87] , \la_oen_user[86] , \la_oen_user[85] , \la_oen_user[84] , \la_oen_user[83] , \la_oen_user[82] , \la_oen_user[81] , \la_oen_user[80] , \la_oen_user[79] , \la_oen_user[78] , \la_oen_user[77] , \la_oen_user[76] , \la_oen_user[75] , \la_oen_user[74] , \la_oen_user[73] , \la_oen_user[72] , \la_oen_user[71] , \la_oen_user[70] , \la_oen_user[69] , \la_oen_user[68] , \la_oen_user[67] , \la_oen_user[66] , \la_oen_user[65] , \la_oen_user[64] , \la_oen_user[63] , \la_oen_user[62] , \la_oen_user[61] , \la_oen_user[60] , \la_oen_user[59] , \la_oen_user[58] , \la_oen_user[57] , \la_oen_user[56] , \la_oen_user[55] , \la_oen_user[54] , \la_oen_user[53] , \la_oen_user[52] , \la_oen_user[51] , \la_oen_user[50] , \la_oen_user[49] , \la_oen_user[48] , \la_oen_user[47] , \la_oen_user[46] , \la_oen_user[45] , \la_oen_user[44] , \la_oen_user[43] , \la_oen_user[42] , \la_oen_user[41] , \la_oen_user[40] , \la_oen_user[39] , \la_oen_user[38] , \la_oen_user[37] , \la_oen_user[36] , \la_oen_user[35] , \la_oen_user[34] , \la_oen_user[33] , \la_oen_user[32] , \la_oen_user[31] , \la_oen_user[30] , \la_oen_user[29] , \la_oen_user[28] , \la_oen_user[27] , \la_oen_user[26] , \la_oen_user[25] , \la_oen_user[24] , \la_oen_user[23] , \la_oen_user[22] , \la_oen_user[21] , \la_oen_user[20] , \la_oen_user[19] , \la_oen_user[18] , \la_oen_user[17] , \la_oen_user[16] , \la_oen_user[15] , \la_oen_user[14] , \la_oen_user[13] , \la_oen_user[12] , \la_oen_user[11] , \la_oen_user[10] , \la_oen_user[9] , \la_oen_user[8] , \la_oen_user[7] , \la_oen_user[6] , \la_oen_user[5] , \la_oen_user[4] , \la_oen_user[3] , \la_oen_user[2] , \la_oen_user[1] , \la_oen_user[0]  }),
    .user_clock2(mprj_clock2),
    .wb_clk_i(mprj_clock),
    .wb_rst_i(mprj_reset),
    .wbs_ack_o(mprj_ack_i_core),
    .wbs_adr_i({ \mprj_adr_o_user[31] , \mprj_adr_o_user[30] , \mprj_adr_o_user[29] , \mprj_adr_o_user[28] , \mprj_adr_o_user[27] , \mprj_adr_o_user[26] , \mprj_adr_o_user[25] , \mprj_adr_o_user[24] , \mprj_adr_o_user[23] , \mprj_adr_o_user[22] , \mprj_adr_o_user[21] , \mprj_adr_o_user[20] , \mprj_adr_o_user[19] , \mprj_adr_o_user[18] , \mprj_adr_o_user[17] , \mprj_adr_o_user[16] , \mprj_adr_o_user[15] , \mprj_adr_o_user[14] , \mprj_adr_o_user[13] , \mprj_adr_o_user[12] , \mprj_adr_o_user[11] , \mprj_adr_o_user[10] , \mprj_adr_o_user[9] , \mprj_adr_o_user[8] , \mprj_adr_o_user[7] , \mprj_adr_o_user[6] , \mprj_adr_o_user[5] , \mprj_adr_o_user[4] , \mprj_adr_o_user[3] , \mprj_adr_o_user[2] , \mprj_adr_o_user[1] , \mprj_adr_o_user[0]  }),
    .wbs_cyc_i(mprj_cyc_o_user),
    .wbs_dat_i({ \mprj_dat_o_user[31] , \mprj_dat_o_user[30] , \mprj_dat_o_user[29] , \mprj_dat_o_user[28] , \mprj_dat_o_user[27] , \mprj_dat_o_user[26] , \mprj_dat_o_user[25] , \mprj_dat_o_user[24] , \mprj_dat_o_user[23] , \mprj_dat_o_user[22] , \mprj_dat_o_user[21] , \mprj_dat_o_user[20] , \mprj_dat_o_user[19] , \mprj_dat_o_user[18] , \mprj_dat_o_user[17] , \mprj_dat_o_user[16] , \mprj_dat_o_user[15] , \mprj_dat_o_user[14] , \mprj_dat_o_user[13] , \mprj_dat_o_user[12] , \mprj_dat_o_user[11] , \mprj_dat_o_user[10] , \mprj_dat_o_user[9] , \mprj_dat_o_user[8] , \mprj_dat_o_user[7] , \mprj_dat_o_user[6] , \mprj_dat_o_user[5] , \mprj_dat_o_user[4] , \mprj_dat_o_user[3] , \mprj_dat_o_user[2] , \mprj_dat_o_user[1] , \mprj_dat_o_user[0]  }),
    .wbs_dat_o({ \mprj_dat_i_core[31] , \mprj_dat_i_core[30] , \mprj_dat_i_core[29] , \mprj_dat_i_core[28] , \mprj_dat_i_core[27] , \mprj_dat_i_core[26] , \mprj_dat_i_core[25] , \mprj_dat_i_core[24] , \mprj_dat_i_core[23] , \mprj_dat_i_core[22] , \mprj_dat_i_core[21] , \mprj_dat_i_core[20] , \mprj_dat_i_core[19] , \mprj_dat_i_core[18] , \mprj_dat_i_core[17] , \mprj_dat_i_core[16] , \mprj_dat_i_core[15] , \mprj_dat_i_core[14] , \mprj_dat_i_core[13] , \mprj_dat_i_core[12] , \mprj_dat_i_core[11] , \mprj_dat_i_core[10] , \mprj_dat_i_core[9] , \mprj_dat_i_core[8] , \mprj_dat_i_core[7] , \mprj_dat_i_core[6] , \mprj_dat_i_core[5] , \mprj_dat_i_core[4] , \mprj_dat_i_core[3] , \mprj_dat_i_core[2] , \mprj_dat_i_core[1] , \mprj_dat_i_core[0]  }),
    .wbs_sel_i({ \mprj_sel_o_user[3] , \mprj_sel_o_user[2] , \mprj_sel_o_user[1] , \mprj_sel_o_user[0]  }),
    .wbs_stb_i(mprj_stb_o_user),
    .wbs_we_i(mprj_we_o_user)
  );
  chip_io padframe (
    .clock(clock),
    .clock_core(clock_core),
    .flash_clk(flash_clk),
    .flash_clk_core(flash_clk_core),
    .flash_clk_ieb_core(flash_clk_ieb_core),
    .flash_clk_oeb_core(flash_clk_oeb_core),
    .flash_csb(flash_csb),
    .flash_csb_core(flash_csb_core),
    .flash_csb_ieb_core(flash_csb_ieb_core),
    .flash_csb_oeb_core(flash_csb_oeb_core),
    .flash_io0(flash_io0),
    .flash_io0_di_core(flash_io0_di_core),
    .flash_io0_do_core(flash_io0_do_core),
    .flash_io0_ieb_core(flash_io0_ieb_core),
    .flash_io0_oeb_core(flash_io0_oeb_core),
    .flash_io1(flash_io1),
    .flash_io1_di_core(flash_io1_di_core),
    .flash_io1_do_core(flash_io1_do_core),
    .flash_io1_ieb_core(flash_io1_ieb_core),
    .flash_io1_oeb_core(flash_io1_oeb_core),
    .gpio(gpio),
    .gpio_in_core(gpio_in_core),
    .gpio_inenb_core(gpio_inenb_core),
    .gpio_mode0_core(gpio_mode0_core),
    .gpio_mode1_core(gpio_mode1_core),
    .gpio_out_core(gpio_out_core),
    .gpio_outenb_core(gpio_outenb_core),
    .mprj_analog_io({ \user_analog_io[30] , \user_analog_io[29] , \user_analog_io[28] , \user_analog_io[27] , \user_analog_io[26] , \user_analog_io[25] , \user_analog_io[24] , \user_analog_io[23] , \user_analog_io[22] , \user_analog_io[21] , \user_analog_io[20] , \user_analog_io[19] , \user_analog_io[18] , \user_analog_io[17] , \user_analog_io[16] , \user_analog_io[15] , \user_analog_io[14] , \user_analog_io[13] , \user_analog_io[12] , \user_analog_io[11] , \user_analog_io[10] , \user_analog_io[9] , \user_analog_io[8] , \user_analog_io[7] , \user_analog_io[6] , \user_analog_io[5] , \user_analog_io[4] , \user_analog_io[3] , \user_analog_io[2] , \user_analog_io[1] , \user_analog_io[0]  }),
    .mprj_io(mprj_io),
    .mprj_io_analog_en({ \mprj_io_analog_en[37] , \mprj_io_analog_en[36] , \mprj_io_analog_en[35] , \mprj_io_analog_en[34] , \mprj_io_analog_en[33] , \mprj_io_analog_en[32] , \mprj_io_analog_en[31] , \mprj_io_analog_en[30] , \mprj_io_analog_en[29] , \mprj_io_analog_en[28] , \mprj_io_analog_en[27] , \mprj_io_analog_en[26] , \mprj_io_analog_en[25] , \mprj_io_analog_en[24] , \mprj_io_analog_en[23] , \mprj_io_analog_en[22] , \mprj_io_analog_en[21] , \mprj_io_analog_en[20] , \mprj_io_analog_en[19] , \mprj_io_analog_en[18] , \mprj_io_analog_en[17] , \mprj_io_analog_en[16] , \mprj_io_analog_en[15] , \mprj_io_analog_en[14] , \mprj_io_analog_en[13] , \mprj_io_analog_en[12] , \mprj_io_analog_en[11] , \mprj_io_analog_en[10] , \mprj_io_analog_en[9] , \mprj_io_analog_en[8] , \mprj_io_analog_en[7] , \mprj_io_analog_en[6] , \mprj_io_analog_en[5] , \mprj_io_analog_en[4] , \mprj_io_analog_en[3] , \mprj_io_analog_en[2] , \mprj_io_analog_en[1] , \mprj_io_analog_en[0]  }),
    .mprj_io_analog_pol({ \mprj_io_analog_pol[37] , \mprj_io_analog_pol[36] , \mprj_io_analog_pol[35] , \mprj_io_analog_pol[34] , \mprj_io_analog_pol[33] , \mprj_io_analog_pol[32] , \mprj_io_analog_pol[31] , \mprj_io_analog_pol[30] , \mprj_io_analog_pol[29] , \mprj_io_analog_pol[28] , \mprj_io_analog_pol[27] , \mprj_io_analog_pol[26] , \mprj_io_analog_pol[25] , \mprj_io_analog_pol[24] , \mprj_io_analog_pol[23] , \mprj_io_analog_pol[22] , \mprj_io_analog_pol[21] , \mprj_io_analog_pol[20] , \mprj_io_analog_pol[19] , \mprj_io_analog_pol[18] , \mprj_io_analog_pol[17] , \mprj_io_analog_pol[16] , \mprj_io_analog_pol[15] , \mprj_io_analog_pol[14] , \mprj_io_analog_pol[13] , \mprj_io_analog_pol[12] , \mprj_io_analog_pol[11] , \mprj_io_analog_pol[10] , \mprj_io_analog_pol[9] , \mprj_io_analog_pol[8] , \mprj_io_analog_pol[7] , \mprj_io_analog_pol[6] , \mprj_io_analog_pol[5] , \mprj_io_analog_pol[4] , \mprj_io_analog_pol[3] , \mprj_io_analog_pol[2] , \mprj_io_analog_pol[1] , \mprj_io_analog_pol[0]  }),
    .mprj_io_analog_sel({ \mprj_io_analog_sel[37] , \mprj_io_analog_sel[36] , \mprj_io_analog_sel[35] , \mprj_io_analog_sel[34] , \mprj_io_analog_sel[33] , \mprj_io_analog_sel[32] , \mprj_io_analog_sel[31] , \mprj_io_analog_sel[30] , \mprj_io_analog_sel[29] , \mprj_io_analog_sel[28] , \mprj_io_analog_sel[27] , \mprj_io_analog_sel[26] , \mprj_io_analog_sel[25] , \mprj_io_analog_sel[24] , \mprj_io_analog_sel[23] , \mprj_io_analog_sel[22] , \mprj_io_analog_sel[21] , \mprj_io_analog_sel[20] , \mprj_io_analog_sel[19] , \mprj_io_analog_sel[18] , \mprj_io_analog_sel[17] , \mprj_io_analog_sel[16] , \mprj_io_analog_sel[15] , \mprj_io_analog_sel[14] , \mprj_io_analog_sel[13] , \mprj_io_analog_sel[12] , \mprj_io_analog_sel[11] , \mprj_io_analog_sel[10] , \mprj_io_analog_sel[9] , \mprj_io_analog_sel[8] , \mprj_io_analog_sel[7] , \mprj_io_analog_sel[6] , \mprj_io_analog_sel[5] , \mprj_io_analog_sel[4] , \mprj_io_analog_sel[3] , \mprj_io_analog_sel[2] , \mprj_io_analog_sel[1] , \mprj_io_analog_sel[0]  }),
    .mprj_io_dm({ \mprj_io_dm[113] , \mprj_io_dm[112] , \mprj_io_dm[111] , \mprj_io_dm[110] , \mprj_io_dm[109] , \mprj_io_dm[108] , \mprj_io_dm[107] , \mprj_io_dm[106] , \mprj_io_dm[105] , \mprj_io_dm[104] , \mprj_io_dm[103] , \mprj_io_dm[102] , \mprj_io_dm[101] , \mprj_io_dm[100] , \mprj_io_dm[99] , \mprj_io_dm[98] , \mprj_io_dm[97] , \mprj_io_dm[96] , \mprj_io_dm[95] , \mprj_io_dm[94] , \mprj_io_dm[93] , \mprj_io_dm[92] , \mprj_io_dm[91] , \mprj_io_dm[90] , \mprj_io_dm[89] , \mprj_io_dm[88] , \mprj_io_dm[87] , \mprj_io_dm[86] , \mprj_io_dm[85] , \mprj_io_dm[84] , \mprj_io_dm[83] , \mprj_io_dm[82] , \mprj_io_dm[81] , \mprj_io_dm[80] , \mprj_io_dm[79] , \mprj_io_dm[78] , \mprj_io_dm[77] , \mprj_io_dm[76] , \mprj_io_dm[75] , \mprj_io_dm[74] , \mprj_io_dm[73] , \mprj_io_dm[72] , \mprj_io_dm[71] , \mprj_io_dm[70] , \mprj_io_dm[69] , \mprj_io_dm[68] , \mprj_io_dm[67] , \mprj_io_dm[66] , \mprj_io_dm[65] , \mprj_io_dm[64] , \mprj_io_dm[63] , \mprj_io_dm[62] , \mprj_io_dm[61] , \mprj_io_dm[60] , \mprj_io_dm[59] , \mprj_io_dm[58] , \mprj_io_dm[57] , \mprj_io_dm[56] , \mprj_io_dm[55] , \mprj_io_dm[54] , \mprj_io_dm[53] , \mprj_io_dm[52] , \mprj_io_dm[51] , \mprj_io_dm[50] , \mprj_io_dm[49] , \mprj_io_dm[48] , \mprj_io_dm[47] , \mprj_io_dm[46] , \mprj_io_dm[45] , \mprj_io_dm[44] , \mprj_io_dm[43] , \mprj_io_dm[42] , \mprj_io_dm[41] , \mprj_io_dm[40] , \mprj_io_dm[39] , \mprj_io_dm[38] , \mprj_io_dm[37] , \mprj_io_dm[36] , \mprj_io_dm[35] , \mprj_io_dm[34] , \mprj_io_dm[33] , \mprj_io_dm[32] , \mprj_io_dm[31] , \mprj_io_dm[30] , \mprj_io_dm[29] , \mprj_io_dm[28] , \mprj_io_dm[27] , \mprj_io_dm[26] , \mprj_io_dm[25] , \mprj_io_dm[24] , \mprj_io_dm[23] , \mprj_io_dm[22] , \mprj_io_dm[21] , \mprj_io_dm[20] , \mprj_io_dm[19] , \mprj_io_dm[18] , \mprj_io_dm[17] , \mprj_io_dm[16] , \mprj_io_dm[15] , \mprj_io_dm[14] , \mprj_io_dm[13] , \mprj_io_dm[12] , \mprj_io_dm[11] , \mprj_io_dm[10] , \mprj_io_dm[9] , \mprj_io_dm[8] , \mprj_io_dm[7] , \mprj_io_dm[6] , \mprj_io_dm[5] , \mprj_io_dm[4] , \mprj_io_dm[3] , \mprj_io_dm[2] , \mprj_io_dm[1] , \mprj_io_dm[0]  }),
    .mprj_io_enh({ \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0] , \mprj_io_enh[0]  }),
    .mprj_io_hldh_n({ vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio, vddio }),
    .mprj_io_holdover({ \mprj_io_holdover[37] , \mprj_io_holdover[36] , \mprj_io_holdover[35] , \mprj_io_holdover[34] , \mprj_io_holdover[33] , \mprj_io_holdover[32] , \mprj_io_holdover[31] , \mprj_io_holdover[30] , \mprj_io_holdover[29] , \mprj_io_holdover[28] , \mprj_io_holdover[27] , \mprj_io_holdover[26] , \mprj_io_holdover[25] , \mprj_io_holdover[24] , \mprj_io_holdover[23] , \mprj_io_holdover[22] , \mprj_io_holdover[21] , \mprj_io_holdover[20] , \mprj_io_holdover[19] , \mprj_io_holdover[18] , \mprj_io_holdover[17] , \mprj_io_holdover[16] , \mprj_io_holdover[15] , \mprj_io_holdover[14] , \mprj_io_holdover[13] , \mprj_io_holdover[12] , \mprj_io_holdover[11] , \mprj_io_holdover[10] , \mprj_io_holdover[9] , \mprj_io_holdover[8] , \mprj_io_holdover[7] , \mprj_io_holdover[6] , \mprj_io_holdover[5] , \mprj_io_holdover[4] , \mprj_io_holdover[3] , \mprj_io_holdover[2] , \mprj_io_holdover[1] , \mprj_io_holdover[0]  }),
    .mprj_io_ib_mode_sel({ \mprj_io_ib_mode_sel[37] , \mprj_io_ib_mode_sel[36] , \mprj_io_ib_mode_sel[35] , \mprj_io_ib_mode_sel[34] , \mprj_io_ib_mode_sel[33] , \mprj_io_ib_mode_sel[32] , \mprj_io_ib_mode_sel[31] , \mprj_io_ib_mode_sel[30] , \mprj_io_ib_mode_sel[29] , \mprj_io_ib_mode_sel[28] , \mprj_io_ib_mode_sel[27] , \mprj_io_ib_mode_sel[26] , \mprj_io_ib_mode_sel[25] , \mprj_io_ib_mode_sel[24] , \mprj_io_ib_mode_sel[23] , \mprj_io_ib_mode_sel[22] , \mprj_io_ib_mode_sel[21] , \mprj_io_ib_mode_sel[20] , \mprj_io_ib_mode_sel[19] , \mprj_io_ib_mode_sel[18] , \mprj_io_ib_mode_sel[17] , \mprj_io_ib_mode_sel[16] , \mprj_io_ib_mode_sel[15] , \mprj_io_ib_mode_sel[14] , \mprj_io_ib_mode_sel[13] , \mprj_io_ib_mode_sel[12] , \mprj_io_ib_mode_sel[11] , \mprj_io_ib_mode_sel[10] , \mprj_io_ib_mode_sel[9] , \mprj_io_ib_mode_sel[8] , \mprj_io_ib_mode_sel[7] , \mprj_io_ib_mode_sel[6] , \mprj_io_ib_mode_sel[5] , \mprj_io_ib_mode_sel[4] , \mprj_io_ib_mode_sel[3] , \mprj_io_ib_mode_sel[2] , \mprj_io_ib_mode_sel[1] , \mprj_io_ib_mode_sel[0]  }),
    .mprj_io_in({ \mprj_io_in[37] , \mprj_io_in[36] , \mprj_io_in[35] , \mprj_io_in[34] , \mprj_io_in[33] , \mprj_io_in[32] , \mprj_io_in[31] , \mprj_io_in[30] , \mprj_io_in[29] , \mprj_io_in[28] , \mprj_io_in[27] , \mprj_io_in[26] , \mprj_io_in[25] , \mprj_io_in[24] , \mprj_io_in[23] , \mprj_io_in[22] , \mprj_io_in[21] , \mprj_io_in[20] , \mprj_io_in[19] , \mprj_io_in[18] , \mprj_io_in[17] , \mprj_io_in[16] , \mprj_io_in[15] , \mprj_io_in[14] , \mprj_io_in[13] , \mprj_io_in[12] , \mprj_io_in[11] , \mprj_io_in[10] , \mprj_io_in[9] , \mprj_io_in[8] , \mprj_io_in[7] , \mprj_io_in[6] , \mprj_io_in[5] , \mprj_io_in[4] , \mprj_io_in[3] , \mprj_io_in[2] , \mprj_io_in[1] , \mprj_io_in[0]  }),
    .mprj_io_inp_dis({ \mprj_io_inp_dis[37] , \mprj_io_inp_dis[36] , \mprj_io_inp_dis[35] , \mprj_io_inp_dis[34] , \mprj_io_inp_dis[33] , \mprj_io_inp_dis[32] , \mprj_io_inp_dis[31] , \mprj_io_inp_dis[30] , \mprj_io_inp_dis[29] , \mprj_io_inp_dis[28] , \mprj_io_inp_dis[27] , \mprj_io_inp_dis[26] , \mprj_io_inp_dis[25] , \mprj_io_inp_dis[24] , \mprj_io_inp_dis[23] , \mprj_io_inp_dis[22] , \mprj_io_inp_dis[21] , \mprj_io_inp_dis[20] , \mprj_io_inp_dis[19] , \mprj_io_inp_dis[18] , \mprj_io_inp_dis[17] , \mprj_io_inp_dis[16] , \mprj_io_inp_dis[15] , \mprj_io_inp_dis[14] , \mprj_io_inp_dis[13] , \mprj_io_inp_dis[12] , \mprj_io_inp_dis[11] , \mprj_io_inp_dis[10] , \mprj_io_inp_dis[9] , \mprj_io_inp_dis[8] , \mprj_io_inp_dis[7] , \mprj_io_inp_dis[6] , \mprj_io_inp_dis[5] , \mprj_io_inp_dis[4] , \mprj_io_inp_dis[3] , \mprj_io_inp_dis[2] , \mprj_io_inp_dis[1] , \mprj_io_inp_dis[0]  }),
    .mprj_io_oeb({ \mprj_io_oeb[37] , \mprj_io_oeb[36] , \mprj_io_oeb[35] , \mprj_io_oeb[34] , \mprj_io_oeb[33] , \mprj_io_oeb[32] , \mprj_io_oeb[31] , \mprj_io_oeb[30] , \mprj_io_oeb[29] , \mprj_io_oeb[28] , \mprj_io_oeb[27] , \mprj_io_oeb[26] , \mprj_io_oeb[25] , \mprj_io_oeb[24] , \mprj_io_oeb[23] , \mprj_io_oeb[22] , \mprj_io_oeb[21] , \mprj_io_oeb[20] , \mprj_io_oeb[19] , \mprj_io_oeb[18] , \mprj_io_oeb[17] , \mprj_io_oeb[16] , \mprj_io_oeb[15] , \mprj_io_oeb[14] , \mprj_io_oeb[13] , \mprj_io_oeb[12] , \mprj_io_oeb[11] , \mprj_io_oeb[10] , \mprj_io_oeb[9] , \mprj_io_oeb[8] , \mprj_io_oeb[7] , \mprj_io_oeb[6] , \mprj_io_oeb[5] , \mprj_io_oeb[4] , \mprj_io_oeb[3] , \mprj_io_oeb[2] , \mprj_io_oeb[1] , \mprj_io_oeb[0]  }),
    .mprj_io_out({ \mprj_io_out[37] , \mprj_io_out[36] , \mprj_io_out[35] , \mprj_io_out[34] , \mprj_io_out[33] , \mprj_io_out[32] , \mprj_io_out[31] , \mprj_io_out[30] , \mprj_io_out[29] , \mprj_io_out[28] , \mprj_io_out[27] , \mprj_io_out[26] , \mprj_io_out[25] , \mprj_io_out[24] , \mprj_io_out[23] , \mprj_io_out[22] , \mprj_io_out[21] , \mprj_io_out[20] , \mprj_io_out[19] , \mprj_io_out[18] , \mprj_io_out[17] , \mprj_io_out[16] , \mprj_io_out[15] , \mprj_io_out[14] , \mprj_io_out[13] , \mprj_io_out[12] , \mprj_io_out[11] , \mprj_io_out[10] , \mprj_io_out[9] , \mprj_io_out[8] , \mprj_io_out[7] , \mprj_io_out[6] , \mprj_io_out[5] , \mprj_io_out[4] , \mprj_io_out[3] , \mprj_io_out[2] , \mprj_io_out[1] , \mprj_io_out[0]  }),
    .mprj_io_slow_sel({ \mprj_io_slow_sel[37] , \mprj_io_slow_sel[36] , \mprj_io_slow_sel[35] , \mprj_io_slow_sel[34] , \mprj_io_slow_sel[33] , \mprj_io_slow_sel[32] , \mprj_io_slow_sel[31] , \mprj_io_slow_sel[30] , \mprj_io_slow_sel[29] , \mprj_io_slow_sel[28] , \mprj_io_slow_sel[27] , \mprj_io_slow_sel[26] , \mprj_io_slow_sel[25] , \mprj_io_slow_sel[24] , \mprj_io_slow_sel[23] , \mprj_io_slow_sel[22] , \mprj_io_slow_sel[21] , \mprj_io_slow_sel[20] , \mprj_io_slow_sel[19] , \mprj_io_slow_sel[18] , \mprj_io_slow_sel[17] , \mprj_io_slow_sel[16] , \mprj_io_slow_sel[15] , \mprj_io_slow_sel[14] , \mprj_io_slow_sel[13] , \mprj_io_slow_sel[12] , \mprj_io_slow_sel[11] , \mprj_io_slow_sel[10] , \mprj_io_slow_sel[9] , \mprj_io_slow_sel[8] , \mprj_io_slow_sel[7] , \mprj_io_slow_sel[6] , \mprj_io_slow_sel[5] , \mprj_io_slow_sel[4] , \mprj_io_slow_sel[3] , \mprj_io_slow_sel[2] , \mprj_io_slow_sel[1] , \mprj_io_slow_sel[0]  }),
    .mprj_io_vtrip_sel({ \mprj_io_vtrip_sel[37] , \mprj_io_vtrip_sel[36] , \mprj_io_vtrip_sel[35] , \mprj_io_vtrip_sel[34] , \mprj_io_vtrip_sel[33] , \mprj_io_vtrip_sel[32] , \mprj_io_vtrip_sel[31] , \mprj_io_vtrip_sel[30] , \mprj_io_vtrip_sel[29] , \mprj_io_vtrip_sel[28] , \mprj_io_vtrip_sel[27] , \mprj_io_vtrip_sel[26] , \mprj_io_vtrip_sel[25] , \mprj_io_vtrip_sel[24] , \mprj_io_vtrip_sel[23] , \mprj_io_vtrip_sel[22] , \mprj_io_vtrip_sel[21] , \mprj_io_vtrip_sel[20] , \mprj_io_vtrip_sel[19] , \mprj_io_vtrip_sel[18] , \mprj_io_vtrip_sel[17] , \mprj_io_vtrip_sel[16] , \mprj_io_vtrip_sel[15] , \mprj_io_vtrip_sel[14] , \mprj_io_vtrip_sel[13] , \mprj_io_vtrip_sel[12] , \mprj_io_vtrip_sel[11] , \mprj_io_vtrip_sel[10] , \mprj_io_vtrip_sel[9] , \mprj_io_vtrip_sel[8] , \mprj_io_vtrip_sel[7] , \mprj_io_vtrip_sel[6] , \mprj_io_vtrip_sel[5] , \mprj_io_vtrip_sel[4] , \mprj_io_vtrip_sel[3] , \mprj_io_vtrip_sel[2] , \mprj_io_vtrip_sel[1] , \mprj_io_vtrip_sel[0]  }),
    .por(por_l),
    .porb_h(\mprj_io_enh[0] ),
    .resetb(resetb),
    .resetb_core_h(rstb_h),
    .vccd(vccd),
    .vccd1(vccd1),
    .vccd2(vccd2),
    .vdda(vdda),
    .vdda1(vdda1),
    .vdda2(vdda2),
    .vddio(vddio),
    .vssa(vssa),
    .vssa1(vssa1),
    .vssa2(vssa2),
    .vssd(vssd),
    .vssd1(vssd1),
    .vssd2(vssd2),
    .vssio(vssio)
  );
  simple_por por (
    .por_l(por_l),
    .porb_h(\mprj_io_enh[0] ),
    .porb_l(porb_l)
  );
  sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped rstb_level (
    .A(rstb_h),
    .X(rstb_l)
  );
  mgmt_core soc (
    .clock(clock_core),
    .core_clk(caravel_clk),
    .core_rstn(caravel_rstn),
    .flash_clk(flash_clk_core),
    .flash_clk_ieb(flash_clk_ieb_core),
    .flash_clk_oeb(flash_clk_oeb_core),
    .flash_csb(flash_csb_core),
    .flash_csb_ieb(flash_csb_ieb_core),
    .flash_csb_oeb(flash_csb_oeb_core),
    .flash_io0_di(flash_io0_di_core),
    .flash_io0_do(flash_io0_do_core),
    .flash_io0_ieb(flash_io0_ieb_core),
    .flash_io0_oeb(flash_io0_oeb_core),
    .flash_io1_di(flash_io1_di_core),
    .flash_io1_do(flash_io1_do_core),
    .flash_io1_ieb(flash_io1_ieb_core),
    .flash_io1_oeb(flash_io1_oeb_core),
    .gpio_in_pad(gpio_in_core),
    .gpio_inenb_pad(gpio_inenb_core),
    .gpio_mode0_pad(gpio_mode0_core),
    .gpio_mode1_pad(gpio_mode1_core),
    .gpio_out_pad(gpio_out_core),
    .gpio_outenb_pad(gpio_outenb_core),
    .jtag_out(jtag_out),
    .jtag_outenb(jtag_outenb),
    .la_input({ \la_data_in_mprj[127] , \la_data_in_mprj[126] , \la_data_in_mprj[125] , \la_data_in_mprj[124] , \la_data_in_mprj[123] , \la_data_in_mprj[122] , \la_data_in_mprj[121] , \la_data_in_mprj[120] , \la_data_in_mprj[119] , \la_data_in_mprj[118] , \la_data_in_mprj[117] , \la_data_in_mprj[116] , \la_data_in_mprj[115] , \la_data_in_mprj[114] , \la_data_in_mprj[113] , \la_data_in_mprj[112] , \la_data_in_mprj[111] , \la_data_in_mprj[110] , \la_data_in_mprj[109] , \la_data_in_mprj[108] , \la_data_in_mprj[107] , \la_data_in_mprj[106] , \la_data_in_mprj[105] , \la_data_in_mprj[104] , \la_data_in_mprj[103] , \la_data_in_mprj[102] , \la_data_in_mprj[101] , \la_data_in_mprj[100] , \la_data_in_mprj[99] , \la_data_in_mprj[98] , \la_data_in_mprj[97] , \la_data_in_mprj[96] , \la_data_in_mprj[95] , \la_data_in_mprj[94] , \la_data_in_mprj[93] , \la_data_in_mprj[92] , \la_data_in_mprj[91] , \la_data_in_mprj[90] , \la_data_in_mprj[89] , \la_data_in_mprj[88] , \la_data_in_mprj[87] , \la_data_in_mprj[86] , \la_data_in_mprj[85] , \la_data_in_mprj[84] , \la_data_in_mprj[83] , \la_data_in_mprj[82] , \la_data_in_mprj[81] , \la_data_in_mprj[80] , \la_data_in_mprj[79] , \la_data_in_mprj[78] , \la_data_in_mprj[77] , \la_data_in_mprj[76] , \la_data_in_mprj[75] , \la_data_in_mprj[74] , \la_data_in_mprj[73] , \la_data_in_mprj[72] , \la_data_in_mprj[71] , \la_data_in_mprj[70] , \la_data_in_mprj[69] , \la_data_in_mprj[68] , \la_data_in_mprj[67] , \la_data_in_mprj[66] , \la_data_in_mprj[65] , \la_data_in_mprj[64] , \la_data_in_mprj[63] , \la_data_in_mprj[62] , \la_data_in_mprj[61] , \la_data_in_mprj[60] , \la_data_in_mprj[59] , \la_data_in_mprj[58] , \la_data_in_mprj[57] , \la_data_in_mprj[56] , \la_data_in_mprj[55] , \la_data_in_mprj[54] , \la_data_in_mprj[53] , \la_data_in_mprj[52] , \la_data_in_mprj[51] , \la_data_in_mprj[50] , \la_data_in_mprj[49] , \la_data_in_mprj[48] , \la_data_in_mprj[47] , \la_data_in_mprj[46] , \la_data_in_mprj[45] , \la_data_in_mprj[44] , \la_data_in_mprj[43] , \la_data_in_mprj[42] , \la_data_in_mprj[41] , \la_data_in_mprj[40] , \la_data_in_mprj[39] , \la_data_in_mprj[38] , \la_data_in_mprj[37] , \la_data_in_mprj[36] , \la_data_in_mprj[35] , \la_data_in_mprj[34] , \la_data_in_mprj[33] , \la_data_in_mprj[32] , \la_data_in_mprj[31] , \la_data_in_mprj[30] , \la_data_in_mprj[29] , \la_data_in_mprj[28] , \la_data_in_mprj[27] , \la_data_in_mprj[26] , \la_data_in_mprj[25] , \la_data_in_mprj[24] , \la_data_in_mprj[23] , \la_data_in_mprj[22] , \la_data_in_mprj[21] , \la_data_in_mprj[20] , \la_data_in_mprj[19] , \la_data_in_mprj[18] , \la_data_in_mprj[17] , \la_data_in_mprj[16] , \la_data_in_mprj[15] , \la_data_in_mprj[14] , \la_data_in_mprj[13] , \la_data_in_mprj[12] , \la_data_in_mprj[11] , \la_data_in_mprj[10] , \la_data_in_mprj[9] , \la_data_in_mprj[8] , \la_data_in_mprj[7] , \la_data_in_mprj[6] , \la_data_in_mprj[5] , \la_data_in_mprj[4] , \la_data_in_mprj[3] , \la_data_in_mprj[2] , \la_data_in_mprj[1] , \la_data_in_mprj[0]  }),
    .la_oen({ \la_oen_mprj[127] , \la_oen_mprj[126] , \la_oen_mprj[125] , \la_oen_mprj[124] , \la_oen_mprj[123] , \la_oen_mprj[122] , \la_oen_mprj[121] , \la_oen_mprj[120] , \la_oen_mprj[119] , \la_oen_mprj[118] , \la_oen_mprj[117] , \la_oen_mprj[116] , \la_oen_mprj[115] , \la_oen_mprj[114] , \la_oen_mprj[113] , \la_oen_mprj[112] , \la_oen_mprj[111] , \la_oen_mprj[110] , \la_oen_mprj[109] , \la_oen_mprj[108] , \la_oen_mprj[107] , \la_oen_mprj[106] , \la_oen_mprj[105] , \la_oen_mprj[104] , \la_oen_mprj[103] , \la_oen_mprj[102] , \la_oen_mprj[101] , \la_oen_mprj[100] , \la_oen_mprj[99] , \la_oen_mprj[98] , \la_oen_mprj[97] , \la_oen_mprj[96] , \la_oen_mprj[95] , \la_oen_mprj[94] , \la_oen_mprj[93] , \la_oen_mprj[92] , \la_oen_mprj[91] , \la_oen_mprj[90] , \la_oen_mprj[89] , \la_oen_mprj[88] , \la_oen_mprj[87] , \la_oen_mprj[86] , \la_oen_mprj[85] , \la_oen_mprj[84] , \la_oen_mprj[83] , \la_oen_mprj[82] , \la_oen_mprj[81] , \la_oen_mprj[80] , \la_oen_mprj[79] , \la_oen_mprj[78] , \la_oen_mprj[77] , \la_oen_mprj[76] , \la_oen_mprj[75] , \la_oen_mprj[74] , \la_oen_mprj[73] , \la_oen_mprj[72] , \la_oen_mprj[71] , \la_oen_mprj[70] , \la_oen_mprj[69] , \la_oen_mprj[68] , \la_oen_mprj[67] , \la_oen_mprj[66] , \la_oen_mprj[65] , \la_oen_mprj[64] , \la_oen_mprj[63] , \la_oen_mprj[62] , \la_oen_mprj[61] , \la_oen_mprj[60] , \la_oen_mprj[59] , \la_oen_mprj[58] , \la_oen_mprj[57] , \la_oen_mprj[56] , \la_oen_mprj[55] , \la_oen_mprj[54] , \la_oen_mprj[53] , \la_oen_mprj[52] , \la_oen_mprj[51] , \la_oen_mprj[50] , \la_oen_mprj[49] , \la_oen_mprj[48] , \la_oen_mprj[47] , \la_oen_mprj[46] , \la_oen_mprj[45] , \la_oen_mprj[44] , \la_oen_mprj[43] , \la_oen_mprj[42] , \la_oen_mprj[41] , \la_oen_mprj[40] , \la_oen_mprj[39] , \la_oen_mprj[38] , \la_oen_mprj[37] , \la_oen_mprj[36] , \la_oen_mprj[35] , \la_oen_mprj[34] , \la_oen_mprj[33] , \la_oen_mprj[32] , \la_oen_mprj[31] , \la_oen_mprj[30] , \la_oen_mprj[29] , \la_oen_mprj[28] , \la_oen_mprj[27] , \la_oen_mprj[26] , \la_oen_mprj[25] , \la_oen_mprj[24] , \la_oen_mprj[23] , \la_oen_mprj[22] , \la_oen_mprj[21] , \la_oen_mprj[20] , \la_oen_mprj[19] , \la_oen_mprj[18] , \la_oen_mprj[17] , \la_oen_mprj[16] , \la_oen_mprj[15] , \la_oen_mprj[14] , \la_oen_mprj[13] , \la_oen_mprj[12] , \la_oen_mprj[11] , \la_oen_mprj[10] , \la_oen_mprj[9] , \la_oen_mprj[8] , \la_oen_mprj[7] , \la_oen_mprj[6] , \la_oen_mprj[5] , \la_oen_mprj[4] , \la_oen_mprj[3] , \la_oen_mprj[2] , \la_oen_mprj[1] , \la_oen_mprj[0]  }),
    .la_output({ \la_data_out_mprj[127] , \la_data_out_mprj[126] , \la_data_out_mprj[125] , \la_data_out_mprj[124] , \la_data_out_mprj[123] , \la_data_out_mprj[122] , \la_data_out_mprj[121] , \la_data_out_mprj[120] , \la_data_out_mprj[119] , \la_data_out_mprj[118] , \la_data_out_mprj[117] , \la_data_out_mprj[116] , \la_data_out_mprj[115] , \la_data_out_mprj[114] , \la_data_out_mprj[113] , \la_data_out_mprj[112] , \la_data_out_mprj[111] , \la_data_out_mprj[110] , \la_data_out_mprj[109] , \la_data_out_mprj[108] , \la_data_out_mprj[107] , \la_data_out_mprj[106] , \la_data_out_mprj[105] , \la_data_out_mprj[104] , \la_data_out_mprj[103] , \la_data_out_mprj[102] , \la_data_out_mprj[101] , \la_data_out_mprj[100] , \la_data_out_mprj[99] , \la_data_out_mprj[98] , \la_data_out_mprj[97] , \la_data_out_mprj[96] , \la_data_out_mprj[95] , \la_data_out_mprj[94] , \la_data_out_mprj[93] , \la_data_out_mprj[92] , \la_data_out_mprj[91] , \la_data_out_mprj[90] , \la_data_out_mprj[89] , \la_data_out_mprj[88] , \la_data_out_mprj[87] , \la_data_out_mprj[86] , \la_data_out_mprj[85] , \la_data_out_mprj[84] , \la_data_out_mprj[83] , \la_data_out_mprj[82] , \la_data_out_mprj[81] , \la_data_out_mprj[80] , \la_data_out_mprj[79] , \la_data_out_mprj[78] , \la_data_out_mprj[77] , \la_data_out_mprj[76] , \la_data_out_mprj[75] , \la_data_out_mprj[74] , \la_data_out_mprj[73] , \la_data_out_mprj[72] , \la_data_out_mprj[71] , \la_data_out_mprj[70] , \la_data_out_mprj[69] , \la_data_out_mprj[68] , \la_data_out_mprj[67] , \la_data_out_mprj[66] , \la_data_out_mprj[65] , \la_data_out_mprj[64] , \la_data_out_mprj[63] , \la_data_out_mprj[62] , \la_data_out_mprj[61] , \la_data_out_mprj[60] , \la_data_out_mprj[59] , \la_data_out_mprj[58] , \la_data_out_mprj[57] , \la_data_out_mprj[56] , \la_data_out_mprj[55] , \la_data_out_mprj[54] , \la_data_out_mprj[53] , \la_data_out_mprj[52] , \la_data_out_mprj[51] , \la_data_out_mprj[50] , \la_data_out_mprj[49] , \la_data_out_mprj[48] , \la_data_out_mprj[47] , \la_data_out_mprj[46] , \la_data_out_mprj[45] , \la_data_out_mprj[44] , \la_data_out_mprj[43] , \la_data_out_mprj[42] , \la_data_out_mprj[41] , \la_data_out_mprj[40] , \la_data_out_mprj[39] , \la_data_out_mprj[38] , \la_data_out_mprj[37] , \la_data_out_mprj[36] , \la_data_out_mprj[35] , \la_data_out_mprj[34] , \la_data_out_mprj[33] , \la_data_out_mprj[32] , \la_data_out_mprj[31] , \la_data_out_mprj[30] , \la_data_out_mprj[29] , \la_data_out_mprj[28] , \la_data_out_mprj[27] , \la_data_out_mprj[26] , \la_data_out_mprj[25] , \la_data_out_mprj[24] , \la_data_out_mprj[23] , \la_data_out_mprj[22] , \la_data_out_mprj[21] , \la_data_out_mprj[20] , \la_data_out_mprj[19] , \la_data_out_mprj[18] , \la_data_out_mprj[17] , \la_data_out_mprj[16] , \la_data_out_mprj[15] , \la_data_out_mprj[14] , \la_data_out_mprj[13] , \la_data_out_mprj[12] , \la_data_out_mprj[11] , \la_data_out_mprj[10] , \la_data_out_mprj[9] , \la_data_out_mprj[8] , \la_data_out_mprj[7] , \la_data_out_mprj[6] , \la_data_out_mprj[5] , \la_data_out_mprj[4] , \la_data_out_mprj[3] , \la_data_out_mprj[2] , \la_data_out_mprj[1] , \la_data_out_mprj[0]  }),
    .mask_rev({ \mask_rev[31] , \mask_rev[30] , \mask_rev[29] , \mask_rev[28] , \mask_rev[27] , \mask_rev[26] , \mask_rev[25] , \mask_rev[24] , \mask_rev[23] , \mask_rev[22] , \mask_rev[21] , \mask_rev[20] , \mask_rev[19] , \mask_rev[18] , \mask_rev[17] , \mask_rev[16] , \mask_rev[15] , \mask_rev[14] , \mask_rev[13] , \mask_rev[12] , \mask_rev[11] , \mask_rev[10] , \mask_rev[9] , \mask_rev[8] , \mask_rev[7] , \mask_rev[6] , \mask_rev[5] , \mask_rev[4] , \mask_rev[3] , \mask_rev[2] , \mask_rev[1] , \mask_rev[0]  }),
    .mgmt_addr({ \mgmt_addr[7] , \mgmt_addr[6] , \mgmt_addr[5] , \mgmt_addr[4] , \mgmt_addr[3] , \mgmt_addr[2] , \mgmt_addr[1] , \mgmt_addr[0]  }),
    .mgmt_addr_ro({ \mgmt_addr_ro[7] , \mgmt_addr_ro[6] , \mgmt_addr_ro[5] , \mgmt_addr_ro[4] , \mgmt_addr_ro[3] , \mgmt_addr_ro[2] , \mgmt_addr_ro[1] , \mgmt_addr_ro[0]  }),
    .mgmt_ena({ \mgmt_ena[1] , \mgmt_ena[0]  }),
    .mgmt_ena_ro(mgmt_ena_ro),
    .mgmt_in_data({ \mgmt_io_in[37] , \mgmt_io_in[36] , \mgmt_io_in[35] , \mgmt_io_in[34] , \mgmt_io_in[33] , \mgmt_io_in[32] , \mgmt_io_in[31] , \mgmt_io_in[30] , \mgmt_io_in[29] , \mgmt_io_in[28] , \mgmt_io_in[27] , \mgmt_io_in[26] , \mgmt_io_in[25] , \mgmt_io_in[24] , \mgmt_io_in[23] , \mgmt_io_in[22] , \mgmt_io_in[21] , \mgmt_io_in[20] , \mgmt_io_in[19] , \mgmt_io_in[18] , \mgmt_io_in[17] , \mgmt_io_in[16] , \mgmt_io_in[15] , \mgmt_io_in[14] , \mgmt_io_in[13] , \mgmt_io_in[12] , \mgmt_io_in[11] , \mgmt_io_in[10] , \mgmt_io_in[9] , \mgmt_io_in[8] , \mgmt_io_in[7] , \mgmt_io_in[6] , \mgmt_io_in[5] , \mgmt_io_in[4] , \mgmt_io_in[3] , \mgmt_io_in[2] , \mgmt_io_in[1] , \mgmt_io_in[0]  }),
    .mgmt_out_data({ \mgmt_io_in[37] , \mgmt_io_in[36] , \mgmt_io_in[35] , \mgmt_io_in[34] , \mgmt_io_in[33] , \mgmt_io_in[32] , \mgmt_io_in[31] , \mgmt_io_in[30] , \mgmt_io_in[29] , \mgmt_io_in[28] , \mgmt_io_in[27] , \mgmt_io_in[26] , \mgmt_io_in[25] , \mgmt_io_in[24] , \mgmt_io_in[23] , \mgmt_io_in[22] , \mgmt_io_in[21] , \mgmt_io_in[20] , \mgmt_io_in[19] , \mgmt_io_in[18] , \mgmt_io_in[17] , \mgmt_io_in[16] , \mgmt_io_in[15] , \mgmt_io_in[14] , \mgmt_io_in[13] , \mgmt_io_in[12] , \mgmt_io_in[11] , \mgmt_io_in[10] , \mgmt_io_in[9] , \mgmt_io_in[8] , \mgmt_io_in[7] , \mgmt_io_in[6] , \mgmt_io_in[5] , \mgmt_io_in[4] , \mgmt_io_in[3] , \mgmt_io_in[2] , \mgmt_io_nc2[1] , \mgmt_io_nc2[0]  }),
    .mgmt_rdata({ \mgmt_rdata[63] , \mgmt_rdata[62] , \mgmt_rdata[61] , \mgmt_rdata[60] , \mgmt_rdata[59] , \mgmt_rdata[58] , \mgmt_rdata[57] , \mgmt_rdata[56] , \mgmt_rdata[55] , \mgmt_rdata[54] , \mgmt_rdata[53] , \mgmt_rdata[52] , \mgmt_rdata[51] , \mgmt_rdata[50] , \mgmt_rdata[49] , \mgmt_rdata[48] , \mgmt_rdata[47] , \mgmt_rdata[46] , \mgmt_rdata[45] , \mgmt_rdata[44] , \mgmt_rdata[43] , \mgmt_rdata[42] , \mgmt_rdata[41] , \mgmt_rdata[40] , \mgmt_rdata[39] , \mgmt_rdata[38] , \mgmt_rdata[37] , \mgmt_rdata[36] , \mgmt_rdata[35] , \mgmt_rdata[34] , \mgmt_rdata[33] , \mgmt_rdata[32] , \mgmt_rdata[31] , \mgmt_rdata[30] , \mgmt_rdata[29] , \mgmt_rdata[28] , \mgmt_rdata[27] , \mgmt_rdata[26] , \mgmt_rdata[25] , \mgmt_rdata[24] , \mgmt_rdata[23] , \mgmt_rdata[22] , \mgmt_rdata[21] , \mgmt_rdata[20] , \mgmt_rdata[19] , \mgmt_rdata[18] , \mgmt_rdata[17] , \mgmt_rdata[16] , \mgmt_rdata[15] , \mgmt_rdata[14] , \mgmt_rdata[13] , \mgmt_rdata[12] , \mgmt_rdata[11] , \mgmt_rdata[10] , \mgmt_rdata[9] , \mgmt_rdata[8] , \mgmt_rdata[7] , \mgmt_rdata[6] , \mgmt_rdata[5] , \mgmt_rdata[4] , \mgmt_rdata[3] , \mgmt_rdata[2] , \mgmt_rdata[1] , \mgmt_rdata[0]  }),
    .mgmt_rdata_ro({ \mgmt_rdata_ro[31] , \mgmt_rdata_ro[30] , \mgmt_rdata_ro[29] , \mgmt_rdata_ro[28] , \mgmt_rdata_ro[27] , \mgmt_rdata_ro[26] , \mgmt_rdata_ro[25] , \mgmt_rdata_ro[24] , \mgmt_rdata_ro[23] , \mgmt_rdata_ro[22] , \mgmt_rdata_ro[21] , \mgmt_rdata_ro[20] , \mgmt_rdata_ro[19] , \mgmt_rdata_ro[18] , \mgmt_rdata_ro[17] , \mgmt_rdata_ro[16] , \mgmt_rdata_ro[15] , \mgmt_rdata_ro[14] , \mgmt_rdata_ro[13] , \mgmt_rdata_ro[12] , \mgmt_rdata_ro[11] , \mgmt_rdata_ro[10] , \mgmt_rdata_ro[9] , \mgmt_rdata_ro[8] , \mgmt_rdata_ro[7] , \mgmt_rdata_ro[6] , \mgmt_rdata_ro[5] , \mgmt_rdata_ro[4] , \mgmt_rdata_ro[3] , \mgmt_rdata_ro[2] , \mgmt_rdata_ro[1] , \mgmt_rdata_ro[0]  }),
    .mgmt_wdata({ \mgmt_wdata[31] , \mgmt_wdata[30] , \mgmt_wdata[29] , \mgmt_wdata[28] , \mgmt_wdata[27] , \mgmt_wdata[26] , \mgmt_wdata[25] , \mgmt_wdata[24] , \mgmt_wdata[23] , \mgmt_wdata[22] , \mgmt_wdata[21] , \mgmt_wdata[20] , \mgmt_wdata[19] , \mgmt_wdata[18] , \mgmt_wdata[17] , \mgmt_wdata[16] , \mgmt_wdata[15] , \mgmt_wdata[14] , \mgmt_wdata[13] , \mgmt_wdata[12] , \mgmt_wdata[11] , \mgmt_wdata[10] , \mgmt_wdata[9] , \mgmt_wdata[8] , \mgmt_wdata[7] , \mgmt_wdata[6] , \mgmt_wdata[5] , \mgmt_wdata[4] , \mgmt_wdata[3] , \mgmt_wdata[2] , \mgmt_wdata[1] , \mgmt_wdata[0]  }),
    .mgmt_wen({ \mgmt_wen[1] , \mgmt_wen[0]  }),
    .mgmt_wen_mask({ \mgmt_wen_mask[7] , \mgmt_wen_mask[6] , \mgmt_wen_mask[5] , \mgmt_wen_mask[4] , \mgmt_wen_mask[3] , \mgmt_wen_mask[2] , \mgmt_wen_mask[1] , \mgmt_wen_mask[0]  }),
    .mprj2_vcc_pwrgood(mprj2_vcc_pwrgood),
    .mprj2_vdd_pwrgood(mprj2_vdd_pwrgood),
    .mprj_ack_i(mprj_ack_i_core),
    .mprj_adr_o({ \mprj_adr_o_core[31] , \mprj_adr_o_core[30] , \mprj_adr_o_core[29] , \mprj_adr_o_core[28] , \mprj_adr_o_core[27] , \mprj_adr_o_core[26] , \mprj_adr_o_core[25] , \mprj_adr_o_core[24] , \mprj_adr_o_core[23] , \mprj_adr_o_core[22] , \mprj_adr_o_core[21] , \mprj_adr_o_core[20] , \mprj_adr_o_core[19] , \mprj_adr_o_core[18] , \mprj_adr_o_core[17] , \mprj_adr_o_core[16] , \mprj_adr_o_core[15] , \mprj_adr_o_core[14] , \mprj_adr_o_core[13] , \mprj_adr_o_core[12] , \mprj_adr_o_core[11] , \mprj_adr_o_core[10] , \mprj_adr_o_core[9] , \mprj_adr_o_core[8] , \mprj_adr_o_core[7] , \mprj_adr_o_core[6] , \mprj_adr_o_core[5] , \mprj_adr_o_core[4] , \mprj_adr_o_core[3] , \mprj_adr_o_core[2] , \mprj_adr_o_core[1] , \mprj_adr_o_core[0]  }),
    .mprj_cyc_o(mprj_cyc_o_core),
    .mprj_dat_i({ \mprj_dat_i_core[31] , \mprj_dat_i_core[30] , \mprj_dat_i_core[29] , \mprj_dat_i_core[28] , \mprj_dat_i_core[27] , \mprj_dat_i_core[26] , \mprj_dat_i_core[25] , \mprj_dat_i_core[24] , \mprj_dat_i_core[23] , \mprj_dat_i_core[22] , \mprj_dat_i_core[21] , \mprj_dat_i_core[20] , \mprj_dat_i_core[19] , \mprj_dat_i_core[18] , \mprj_dat_i_core[17] , \mprj_dat_i_core[16] , \mprj_dat_i_core[15] , \mprj_dat_i_core[14] , \mprj_dat_i_core[13] , \mprj_dat_i_core[12] , \mprj_dat_i_core[11] , \mprj_dat_i_core[10] , \mprj_dat_i_core[9] , \mprj_dat_i_core[8] , \mprj_dat_i_core[7] , \mprj_dat_i_core[6] , \mprj_dat_i_core[5] , \mprj_dat_i_core[4] , \mprj_dat_i_core[3] , \mprj_dat_i_core[2] , \mprj_dat_i_core[1] , \mprj_dat_i_core[0]  }),
    .mprj_dat_o({ \mprj_dat_o_core[31] , \mprj_dat_o_core[30] , \mprj_dat_o_core[29] , \mprj_dat_o_core[28] , \mprj_dat_o_core[27] , \mprj_dat_o_core[26] , \mprj_dat_o_core[25] , \mprj_dat_o_core[24] , \mprj_dat_o_core[23] , \mprj_dat_o_core[22] , \mprj_dat_o_core[21] , \mprj_dat_o_core[20] , \mprj_dat_o_core[19] , \mprj_dat_o_core[18] , \mprj_dat_o_core[17] , \mprj_dat_o_core[16] , \mprj_dat_o_core[15] , \mprj_dat_o_core[14] , \mprj_dat_o_core[13] , \mprj_dat_o_core[12] , \mprj_dat_o_core[11] , \mprj_dat_o_core[10] , \mprj_dat_o_core[9] , \mprj_dat_o_core[8] , \mprj_dat_o_core[7] , \mprj_dat_o_core[6] , \mprj_dat_o_core[5] , \mprj_dat_o_core[4] , \mprj_dat_o_core[3] , \mprj_dat_o_core[2] , \mprj_dat_o_core[1] , \mprj_dat_o_core[0]  }),
    .mprj_io_loader_clock(mprj_io_loader_clock),
    .mprj_io_loader_data(\gpio_serial_link_shifted[0] ),
    .mprj_io_loader_resetn(mprj_io_loader_resetn),
    .mprj_sel_o({ \mprj_sel_o_core[3] , \mprj_sel_o_core[2] , \mprj_sel_o_core[1] , \mprj_sel_o_core[0]  }),
    .mprj_stb_o(mprj_stb_o_core),
    .mprj_vcc_pwrgood(mprj_vcc_pwrgood),
    .mprj_vdd_pwrgood(mprj_vdd_pwrgood),
    .mprj_we_o(mprj_we_o_core),
    .porb(porb_l),
    .pwr_ctrl_out(pwr_ctrl_out),
    .resetb(rstb_l),
    .sdo_out(sdo_out),
    .sdo_outenb(sdo_outenb),
    .user_clk(caravel_clk2)
  );
  storage storage (
    .mgmt_addr({ \mgmt_addr[7] , \mgmt_addr[6] , \mgmt_addr[5] , \mgmt_addr[4] , \mgmt_addr[3] , \mgmt_addr[2] , \mgmt_addr[1] , \mgmt_addr[0]  }),
    .mgmt_addr_ro({ \mgmt_addr_ro[7] , \mgmt_addr_ro[6] , \mgmt_addr_ro[5] , \mgmt_addr_ro[4] , \mgmt_addr_ro[3] , \mgmt_addr_ro[2] , \mgmt_addr_ro[1] , \mgmt_addr_ro[0]  }),
    .mgmt_clk(caravel_clk),
    .mgmt_ena({ \mgmt_ena[1] , \mgmt_ena[0]  }),
    .mgmt_ena_ro(mgmt_ena_ro),
    .mgmt_rdata({ \mgmt_rdata[63] , \mgmt_rdata[62] , \mgmt_rdata[61] , \mgmt_rdata[60] , \mgmt_rdata[59] , \mgmt_rdata[58] , \mgmt_rdata[57] , \mgmt_rdata[56] , \mgmt_rdata[55] , \mgmt_rdata[54] , \mgmt_rdata[53] , \mgmt_rdata[52] , \mgmt_rdata[51] , \mgmt_rdata[50] , \mgmt_rdata[49] , \mgmt_rdata[48] , \mgmt_rdata[47] , \mgmt_rdata[46] , \mgmt_rdata[45] , \mgmt_rdata[44] , \mgmt_rdata[43] , \mgmt_rdata[42] , \mgmt_rdata[41] , \mgmt_rdata[40] , \mgmt_rdata[39] , \mgmt_rdata[38] , \mgmt_rdata[37] , \mgmt_rdata[36] , \mgmt_rdata[35] , \mgmt_rdata[34] , \mgmt_rdata[33] , \mgmt_rdata[32] , \mgmt_rdata[31] , \mgmt_rdata[30] , \mgmt_rdata[29] , \mgmt_rdata[28] , \mgmt_rdata[27] , \mgmt_rdata[26] , \mgmt_rdata[25] , \mgmt_rdata[24] , \mgmt_rdata[23] , \mgmt_rdata[22] , \mgmt_rdata[21] , \mgmt_rdata[20] , \mgmt_rdata[19] , \mgmt_rdata[18] , \mgmt_rdata[17] , \mgmt_rdata[16] , \mgmt_rdata[15] , \mgmt_rdata[14] , \mgmt_rdata[13] , \mgmt_rdata[12] , \mgmt_rdata[11] , \mgmt_rdata[10] , \mgmt_rdata[9] , \mgmt_rdata[8] , \mgmt_rdata[7] , \mgmt_rdata[6] , \mgmt_rdata[5] , \mgmt_rdata[4] , \mgmt_rdata[3] , \mgmt_rdata[2] , \mgmt_rdata[1] , \mgmt_rdata[0]  }),
    .mgmt_rdata_ro({ \mgmt_rdata_ro[31] , \mgmt_rdata_ro[30] , \mgmt_rdata_ro[29] , \mgmt_rdata_ro[28] , \mgmt_rdata_ro[27] , \mgmt_rdata_ro[26] , \mgmt_rdata_ro[25] , \mgmt_rdata_ro[24] , \mgmt_rdata_ro[23] , \mgmt_rdata_ro[22] , \mgmt_rdata_ro[21] , \mgmt_rdata_ro[20] , \mgmt_rdata_ro[19] , \mgmt_rdata_ro[18] , \mgmt_rdata_ro[17] , \mgmt_rdata_ro[16] , \mgmt_rdata_ro[15] , \mgmt_rdata_ro[14] , \mgmt_rdata_ro[13] , \mgmt_rdata_ro[12] , \mgmt_rdata_ro[11] , \mgmt_rdata_ro[10] , \mgmt_rdata_ro[9] , \mgmt_rdata_ro[8] , \mgmt_rdata_ro[7] , \mgmt_rdata_ro[6] , \mgmt_rdata_ro[5] , \mgmt_rdata_ro[4] , \mgmt_rdata_ro[3] , \mgmt_rdata_ro[2] , \mgmt_rdata_ro[1] , \mgmt_rdata_ro[0]  }),
    .mgmt_wdata({ \mgmt_wdata[31] , \mgmt_wdata[30] , \mgmt_wdata[29] , \mgmt_wdata[28] , \mgmt_wdata[27] , \mgmt_wdata[26] , \mgmt_wdata[25] , \mgmt_wdata[24] , \mgmt_wdata[23] , \mgmt_wdata[22] , \mgmt_wdata[21] , \mgmt_wdata[20] , \mgmt_wdata[19] , \mgmt_wdata[18] , \mgmt_wdata[17] , \mgmt_wdata[16] , \mgmt_wdata[15] , \mgmt_wdata[14] , \mgmt_wdata[13] , \mgmt_wdata[12] , \mgmt_wdata[11] , \mgmt_wdata[10] , \mgmt_wdata[9] , \mgmt_wdata[8] , \mgmt_wdata[7] , \mgmt_wdata[6] , \mgmt_wdata[5] , \mgmt_wdata[4] , \mgmt_wdata[3] , \mgmt_wdata[2] , \mgmt_wdata[1] , \mgmt_wdata[0]  }),
    .mgmt_wen({ \mgmt_wen[1] , \mgmt_wen[0]  }),
    .mgmt_wen_mask({ \mgmt_wen_mask[7] , \mgmt_wen_mask[6] , \mgmt_wen_mask[5] , \mgmt_wen_mask[4] , \mgmt_wen_mask[3] , \mgmt_wen_mask[2] , \mgmt_wen_mask[1] , \mgmt_wen_mask[0]  })
  );
  user_id_programming user_id_value (
    .mask_rev({ \mask_rev[31] , \mask_rev[30] , \mask_rev[29] , \mask_rev[28] , \mask_rev[27] , \mask_rev[26] , \mask_rev[25] , \mask_rev[24] , \mask_rev[23] , \mask_rev[22] , \mask_rev[21] , \mask_rev[20] , \mask_rev[19] , \mask_rev[18] , \mask_rev[17] , \mask_rev[16] , \mask_rev[15] , \mask_rev[14] , \mask_rev[13] , \mask_rev[12] , \mask_rev[11] , \mask_rev[10] , \mask_rev[9] , \mask_rev[8] , \mask_rev[7] , \mask_rev[6] , \mask_rev[5] , \mask_rev[4] , \mask_rev[3] , \mask_rev[2] , \mask_rev[1] , \mask_rev[0]  })
  );
  assign \gpio_serial_link_shifted[37]  = \gpio_serial_link[36] ;
  assign \gpio_serial_link_shifted[36]  = \gpio_serial_link[35] ;
  assign \gpio_serial_link_shifted[35]  = \gpio_serial_link[34] ;
  assign \gpio_serial_link_shifted[34]  = \gpio_serial_link[33] ;
  assign \gpio_serial_link_shifted[33]  = \gpio_serial_link[32] ;
  assign \gpio_serial_link_shifted[32]  = \gpio_serial_link[31] ;
  assign \gpio_serial_link_shifted[31]  = \gpio_serial_link[30] ;
  assign \gpio_serial_link_shifted[30]  = \gpio_serial_link[29] ;
  assign \gpio_serial_link_shifted[29]  = \gpio_serial_link[28] ;
  assign \gpio_serial_link_shifted[28]  = \gpio_serial_link[27] ;
  assign \gpio_serial_link_shifted[27]  = \gpio_serial_link[26] ;
  assign \gpio_serial_link_shifted[26]  = \gpio_serial_link[25] ;
  assign \gpio_serial_link_shifted[25]  = \gpio_serial_link[24] ;
  assign \gpio_serial_link_shifted[24]  = \gpio_serial_link[23] ;
  assign \gpio_serial_link_shifted[23]  = \gpio_serial_link[22] ;
  assign \gpio_serial_link_shifted[22]  = \gpio_serial_link[21] ;
  assign \gpio_serial_link_shifted[21]  = \gpio_serial_link[20] ;
  assign \gpio_serial_link_shifted[20]  = \gpio_serial_link[19] ;
  assign \gpio_serial_link_shifted[19]  = \gpio_serial_link[18] ;
  assign \gpio_serial_link_shifted[18]  = \gpio_serial_link[17] ;
  assign \gpio_serial_link_shifted[17]  = \gpio_serial_link[16] ;
  assign \gpio_serial_link_shifted[16]  = \gpio_serial_link[15] ;
  assign \gpio_serial_link_shifted[15]  = \gpio_serial_link[14] ;
  assign \gpio_serial_link_shifted[14]  = \gpio_serial_link[13] ;
  assign \gpio_serial_link_shifted[13]  = \gpio_serial_link[12] ;
  assign \gpio_serial_link_shifted[12]  = \gpio_serial_link[11] ;
  assign \gpio_serial_link_shifted[11]  = \gpio_serial_link[10] ;
  assign \gpio_serial_link_shifted[10]  = \gpio_serial_link[9] ;
  assign \gpio_serial_link_shifted[9]  = \gpio_serial_link[8] ;
  assign \gpio_serial_link_shifted[8]  = \gpio_serial_link[7] ;
  assign \gpio_serial_link_shifted[7]  = \gpio_serial_link[6] ;
  assign \gpio_serial_link_shifted[6]  = \gpio_serial_link[5] ;
  assign \gpio_serial_link_shifted[5]  = \gpio_serial_link[4] ;
  assign \gpio_serial_link_shifted[4]  = \gpio_serial_link[3] ;
  assign \gpio_serial_link_shifted[3]  = \gpio_serial_link[2] ;
  assign \gpio_serial_link_shifted[2]  = \gpio_serial_link[1] ;
  assign \gpio_serial_link_shifted[1]  = \gpio_serial_link[0] ;
  assign \mprj_io_hldh_n[37]  = vddio;
  assign \mprj_io_hldh_n[36]  = vddio;
  assign \mprj_io_hldh_n[35]  = vddio;
  assign \mprj_io_hldh_n[34]  = vddio;
  assign \mprj_io_hldh_n[33]  = vddio;
  assign \mprj_io_hldh_n[32]  = vddio;
  assign \mprj_io_hldh_n[31]  = vddio;
  assign \mprj_io_hldh_n[30]  = vddio;
  assign \mprj_io_hldh_n[29]  = vddio;
  assign \mprj_io_hldh_n[28]  = vddio;
  assign \mprj_io_hldh_n[27]  = vddio;
  assign \mprj_io_hldh_n[26]  = vddio;
  assign \mprj_io_hldh_n[25]  = vddio;
  assign \mprj_io_hldh_n[24]  = vddio;
  assign \mprj_io_hldh_n[23]  = vddio;
  assign \mprj_io_hldh_n[22]  = vddio;
  assign \mprj_io_hldh_n[21]  = vddio;
  assign \mprj_io_hldh_n[20]  = vddio;
  assign \mprj_io_hldh_n[19]  = vddio;
  assign \mprj_io_hldh_n[18]  = vddio;
  assign \mprj_io_hldh_n[17]  = vddio;
  assign \mprj_io_hldh_n[16]  = vddio;
  assign \mprj_io_hldh_n[15]  = vddio;
  assign \mprj_io_hldh_n[14]  = vddio;
  assign \mprj_io_hldh_n[13]  = vddio;
  assign \mprj_io_hldh_n[12]  = vddio;
  assign \mprj_io_hldh_n[11]  = vddio;
  assign \mprj_io_hldh_n[10]  = vddio;
  assign \mprj_io_hldh_n[9]  = vddio;
  assign \mprj_io_hldh_n[8]  = vddio;
  assign \mprj_io_hldh_n[7]  = vddio;
  assign \mprj_io_hldh_n[6]  = vddio;
  assign \mprj_io_hldh_n[5]  = vddio;
  assign \mprj_io_hldh_n[4]  = vddio;
  assign \mprj_io_hldh_n[3]  = vddio;
  assign \mprj_io_hldh_n[2]  = vddio;
  assign \mprj_io_hldh_n[1]  = vddio;
  assign \mprj_io_hldh_n[0]  = vddio;
  assign \mprj_io_enh[37]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[36]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[35]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[34]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[33]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[32]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[31]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[30]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[29]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[28]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[27]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[26]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[25]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[24]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[23]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[22]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[21]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[20]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[19]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[18]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[17]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[16]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[15]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[14]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[13]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[12]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[11]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[10]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[9]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[8]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[7]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[6]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[5]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[4]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[3]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[2]  = \mprj_io_enh[0] ;
  assign \mprj_io_enh[1]  = \mprj_io_enh[0] ;
  assign porb_h = \mprj_io_enh[0] ;
  assign mprj_io_loader_data = \gpio_serial_link_shifted[0] ;
endmodule
