magic
tech sky130A
magscale 1 2
timestamp 1623173305
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< metal1 >>
rect 434992 1008039 434998 1008091
rect 435050 1008079 435056 1008091
rect 470800 1008079 470806 1008091
rect 435050 1008051 470806 1008079
rect 435050 1008039 435056 1008051
rect 470800 1008039 470806 1008051
rect 470858 1008039 470864 1008091
rect 434704 1005523 434710 1005575
rect 434762 1005563 434768 1005575
rect 472144 1005563 472150 1005575
rect 434762 1005535 472150 1005563
rect 434762 1005523 434768 1005535
rect 472144 1005523 472150 1005535
rect 472202 1005523 472208 1005575
rect 367216 1005375 367222 1005427
rect 367274 1005415 367280 1005427
rect 383632 1005415 383638 1005427
rect 367274 1005387 383638 1005415
rect 367274 1005375 367280 1005387
rect 383632 1005375 383638 1005387
rect 383690 1005375 383696 1005427
rect 434896 1005375 434902 1005427
rect 434954 1005415 434960 1005427
rect 459280 1005415 459286 1005427
rect 434954 1005387 459286 1005415
rect 434954 1005375 434960 1005387
rect 459280 1005375 459286 1005387
rect 459338 1005375 459344 1005427
rect 436912 1005301 436918 1005353
rect 436970 1005341 436976 1005353
rect 471376 1005341 471382 1005353
rect 436970 1005313 471382 1005341
rect 436970 1005301 436976 1005313
rect 471376 1005301 471382 1005313
rect 471434 1005301 471440 1005353
rect 164272 1005227 164278 1005279
rect 164330 1005267 164336 1005279
rect 172816 1005267 172822 1005279
rect 164330 1005239 172822 1005267
rect 164330 1005227 164336 1005239
rect 172816 1005227 172822 1005239
rect 172874 1005227 172880 1005279
rect 316816 1005227 316822 1005279
rect 316874 1005267 316880 1005279
rect 331216 1005267 331222 1005279
rect 316874 1005239 331222 1005267
rect 316874 1005227 316880 1005239
rect 331216 1005227 331222 1005239
rect 331274 1005227 331280 1005279
rect 434608 1005227 434614 1005279
rect 434666 1005267 434672 1005279
rect 472240 1005267 472246 1005279
rect 434666 1005239 472246 1005267
rect 434666 1005227 434672 1005239
rect 472240 1005227 472246 1005239
rect 472298 1005227 472304 1005279
rect 218800 1005153 218806 1005205
rect 218858 1005193 218864 1005205
rect 222736 1005193 222742 1005205
rect 218858 1005165 222742 1005193
rect 218858 1005153 218864 1005165
rect 222736 1005153 222742 1005165
rect 222794 1005153 222800 1005205
rect 434800 1005153 434806 1005205
rect 434858 1005193 434864 1005205
rect 443728 1005193 443734 1005205
rect 434858 1005165 443734 1005193
rect 434858 1005153 434864 1005165
rect 443728 1005153 443734 1005165
rect 443786 1005153 443792 1005205
rect 443536 1003673 443542 1003725
rect 443594 1003713 443600 1003725
rect 463792 1003713 463798 1003725
rect 443594 1003685 463798 1003713
rect 443594 1003673 443600 1003685
rect 463792 1003673 463798 1003685
rect 463850 1003673 463856 1003725
rect 377680 1003269 377686 1003281
rect 359074 1003241 377686 1003269
rect 359074 1003207 359102 1003241
rect 377680 1003229 377686 1003241
rect 377738 1003229 377744 1003281
rect 467056 1003269 467062 1003281
rect 426082 1003241 467062 1003269
rect 426082 1003207 426110 1003241
rect 467056 1003229 467062 1003241
rect 467114 1003229 467120 1003281
rect 518608 1003269 518614 1003281
rect 502402 1003241 518614 1003269
rect 160432 1003155 160438 1003207
rect 160490 1003195 160496 1003207
rect 164272 1003195 164278 1003207
rect 160490 1003167 164278 1003195
rect 160490 1003155 160496 1003167
rect 164272 1003155 164278 1003167
rect 164330 1003155 164336 1003207
rect 211792 1003155 211798 1003207
rect 211850 1003195 211856 1003207
rect 213808 1003195 213814 1003207
rect 211850 1003167 213814 1003195
rect 211850 1003155 211856 1003167
rect 213808 1003155 213814 1003167
rect 213866 1003155 213872 1003207
rect 359056 1003155 359062 1003207
rect 359114 1003155 359120 1003207
rect 362512 1003155 362518 1003207
rect 362570 1003195 362576 1003207
rect 367216 1003195 367222 1003207
rect 362570 1003167 367222 1003195
rect 362570 1003155 362576 1003167
rect 367216 1003155 367222 1003167
rect 367274 1003155 367280 1003207
rect 426064 1003155 426070 1003207
rect 426122 1003155 426128 1003207
rect 429232 1003155 429238 1003207
rect 429290 1003195 429296 1003207
rect 434608 1003195 434614 1003207
rect 429290 1003167 434614 1003195
rect 429290 1003155 429296 1003167
rect 434608 1003155 434614 1003167
rect 434666 1003155 434672 1003207
rect 439216 1003155 439222 1003207
rect 439274 1003195 439280 1003207
rect 466576 1003195 466582 1003207
rect 439274 1003167 466582 1003195
rect 439274 1003155 439280 1003167
rect 466576 1003155 466582 1003167
rect 466634 1003155 466640 1003207
rect 502402 1003133 502430 1003241
rect 518608 1003229 518614 1003241
rect 518666 1003229 518672 1003281
rect 518800 1003195 518806 1003207
rect 502882 1003167 518806 1003195
rect 449200 1003081 449206 1003133
rect 449258 1003121 449264 1003133
rect 467824 1003121 467830 1003133
rect 449258 1003093 467830 1003121
rect 449258 1003081 449264 1003093
rect 467824 1003081 467830 1003093
rect 467882 1003081 467888 1003133
rect 502384 1003081 502390 1003133
rect 502442 1003081 502448 1003133
rect 425392 1003007 425398 1003059
rect 425450 1003047 425456 1003059
rect 430192 1003047 430198 1003059
rect 425450 1003019 430198 1003047
rect 425450 1003007 425456 1003019
rect 430192 1003007 430198 1003019
rect 430250 1003007 430256 1003059
rect 430288 1003007 430294 1003059
rect 430346 1003047 430352 1003059
rect 434896 1003047 434902 1003059
rect 430346 1003019 434902 1003047
rect 430346 1003007 430352 1003019
rect 434896 1003007 434902 1003019
rect 434954 1003007 434960 1003059
rect 439120 1003007 439126 1003059
rect 439178 1003047 439184 1003059
rect 463504 1003047 463510 1003059
rect 439178 1003019 463510 1003047
rect 439178 1003007 439184 1003019
rect 463504 1003007 463510 1003019
rect 463562 1003007 463568 1003059
rect 501328 1003007 501334 1003059
rect 501386 1003047 501392 1003059
rect 502882 1003047 502910 1003167
rect 518800 1003155 518806 1003167
rect 518858 1003155 518864 1003207
rect 502960 1003081 502966 1003133
rect 503018 1003121 503024 1003133
rect 518704 1003121 518710 1003133
rect 503018 1003093 518710 1003121
rect 503018 1003081 503024 1003093
rect 518704 1003081 518710 1003093
rect 518762 1003081 518768 1003133
rect 501386 1003019 502910 1003047
rect 501386 1003007 501392 1003019
rect 504016 1003007 504022 1003059
rect 504074 1003047 504080 1003059
rect 518416 1003047 518422 1003059
rect 504074 1003019 518422 1003047
rect 504074 1003007 504080 1003019
rect 518416 1003007 518422 1003019
rect 518474 1003007 518480 1003059
rect 424336 1002933 424342 1002985
rect 424394 1002973 424400 1002985
rect 463600 1002973 463606 1002985
rect 424394 1002945 463606 1002973
rect 424394 1002933 424400 1002945
rect 463600 1002933 463606 1002945
rect 463658 1002933 463664 1002985
rect 554896 1002933 554902 1002985
rect 554954 1002973 554960 1002985
rect 573040 1002973 573046 1002985
rect 554954 1002945 573046 1002973
rect 554954 1002933 554960 1002945
rect 573040 1002933 573046 1002945
rect 573098 1002933 573104 1002985
rect 299344 1002859 299350 1002911
rect 299402 1002899 299408 1002911
rect 308848 1002899 308854 1002911
rect 299402 1002871 308854 1002899
rect 299402 1002859 299408 1002871
rect 308848 1002859 308854 1002871
rect 308906 1002859 308912 1002911
rect 428752 1002859 428758 1002911
rect 428810 1002899 428816 1002911
rect 434704 1002899 434710 1002911
rect 428810 1002871 434710 1002899
rect 428810 1002859 428816 1002871
rect 434704 1002859 434710 1002871
rect 434762 1002859 434768 1002911
rect 161488 1002785 161494 1002837
rect 161546 1002825 161552 1002837
rect 169936 1002825 169942 1002837
rect 161546 1002797 169942 1002825
rect 161546 1002785 161552 1002797
rect 169936 1002785 169942 1002797
rect 169994 1002785 170000 1002837
rect 299440 1002785 299446 1002837
rect 299498 1002825 299504 1002837
rect 309328 1002825 309334 1002837
rect 299498 1002797 309334 1002825
rect 299498 1002785 299504 1002797
rect 309328 1002785 309334 1002797
rect 309386 1002785 309392 1002837
rect 428272 1002785 428278 1002837
rect 428330 1002825 428336 1002837
rect 434800 1002825 434806 1002837
rect 428330 1002797 434806 1002825
rect 428330 1002785 428336 1002797
rect 434800 1002785 434806 1002797
rect 434858 1002785 434864 1002837
rect 554320 1002785 554326 1002837
rect 554378 1002825 554384 1002837
rect 572848 1002825 572854 1002837
rect 554378 1002797 572854 1002825
rect 554378 1002785 554384 1002797
rect 572848 1002785 572854 1002797
rect 572906 1002785 572912 1002837
rect 299248 1002711 299254 1002763
rect 299306 1002751 299312 1002763
rect 308272 1002751 308278 1002763
rect 299306 1002723 308278 1002751
rect 299306 1002711 299312 1002723
rect 308272 1002711 308278 1002723
rect 308330 1002711 308336 1002763
rect 423760 1002711 423766 1002763
rect 423818 1002751 423824 1002763
rect 439120 1002751 439126 1002763
rect 423818 1002723 439126 1002751
rect 423818 1002711 423824 1002723
rect 439120 1002711 439126 1002723
rect 439178 1002711 439184 1002763
rect 424816 1002637 424822 1002689
rect 424874 1002677 424880 1002689
rect 439216 1002677 439222 1002689
rect 424874 1002649 439222 1002677
rect 424874 1002637 424880 1002649
rect 439216 1002637 439222 1002649
rect 439274 1002637 439280 1002689
rect 361264 1002563 361270 1002615
rect 361322 1002603 361328 1002615
rect 368848 1002603 368854 1002615
rect 361322 1002575 368854 1002603
rect 361322 1002563 361328 1002575
rect 368848 1002563 368854 1002575
rect 368906 1002563 368912 1002615
rect 427696 1002563 427702 1002615
rect 427754 1002603 427760 1002615
rect 435184 1002603 435190 1002615
rect 427754 1002575 435190 1002603
rect 427754 1002563 427760 1002575
rect 435184 1002563 435190 1002575
rect 435242 1002563 435248 1002615
rect 553744 1002563 553750 1002615
rect 553802 1002603 553808 1002615
rect 572944 1002603 572950 1002615
rect 553802 1002575 572950 1002603
rect 553802 1002563 553808 1002575
rect 572944 1002563 572950 1002575
rect 573002 1002563 573008 1002615
rect 361840 1002489 361846 1002541
rect 361898 1002529 361904 1002541
rect 368656 1002529 368662 1002541
rect 361898 1002501 368662 1002529
rect 361898 1002489 361904 1002501
rect 368656 1002489 368662 1002501
rect 368714 1002489 368720 1002541
rect 426640 1002489 426646 1002541
rect 426698 1002529 426704 1002541
rect 435088 1002529 435094 1002541
rect 426698 1002501 435094 1002529
rect 426698 1002489 426704 1002501
rect 435088 1002489 435094 1002501
rect 435146 1002489 435152 1002541
rect 151120 1002455 151126 1002467
rect 143842 1002427 151126 1002455
rect 143728 1002341 143734 1002393
rect 143786 1002381 143792 1002393
rect 143842 1002381 143870 1002427
rect 151120 1002415 151126 1002427
rect 151178 1002415 151184 1002467
rect 427120 1002415 427126 1002467
rect 427178 1002455 427184 1002467
rect 443632 1002455 443638 1002467
rect 427178 1002427 443638 1002455
rect 427178 1002415 427184 1002427
rect 443632 1002415 443638 1002427
rect 443690 1002415 443696 1002467
rect 143786 1002353 143870 1002381
rect 143786 1002341 143792 1002353
rect 146800 1002341 146806 1002393
rect 146858 1002381 146864 1002393
rect 152752 1002381 152758 1002393
rect 146858 1002353 152758 1002381
rect 146858 1002341 146864 1002353
rect 152752 1002341 152758 1002353
rect 152810 1002341 152816 1002393
rect 255472 1002381 255478 1002393
rect 246568 1002353 255478 1002381
rect 143920 1002267 143926 1002319
rect 143978 1002307 143984 1002319
rect 175696 1002307 175702 1002319
rect 143978 1002279 175702 1002307
rect 143978 1002267 143984 1002279
rect 175696 1002267 175702 1002279
rect 175754 1002267 175760 1002319
rect 246568 1002245 246596 1002353
rect 255472 1002341 255478 1002353
rect 255530 1002341 255536 1002393
rect 363472 1002341 363478 1002393
rect 363530 1002381 363536 1002393
rect 377104 1002381 377110 1002393
rect 363530 1002353 377110 1002381
rect 363530 1002341 363536 1002353
rect 377104 1002341 377110 1002353
rect 377162 1002341 377168 1002393
rect 431920 1002341 431926 1002393
rect 431978 1002381 431984 1002393
rect 434992 1002381 434998 1002393
rect 431978 1002353 434998 1002381
rect 431978 1002341 431984 1002353
rect 434992 1002341 434998 1002353
rect 435050 1002341 435056 1002393
rect 503440 1002341 503446 1002393
rect 503498 1002381 503504 1002393
rect 514000 1002381 514006 1002393
rect 503498 1002353 514006 1002381
rect 503498 1002341 503504 1002353
rect 514000 1002341 514006 1002353
rect 514058 1002341 514064 1002393
rect 553264 1002341 553270 1002393
rect 553322 1002381 553328 1002393
rect 567472 1002381 567478 1002393
rect 553322 1002353 567478 1002381
rect 553322 1002341 553328 1002353
rect 567472 1002341 567478 1002353
rect 567530 1002341 567536 1002393
rect 246640 1002267 246646 1002319
rect 246698 1002307 246704 1002319
rect 253840 1002307 253846 1002319
rect 246698 1002279 253846 1002307
rect 246698 1002267 246704 1002279
rect 253840 1002267 253846 1002279
rect 253898 1002267 253904 1002319
rect 362896 1002267 362902 1002319
rect 362954 1002307 362960 1002319
rect 368752 1002307 368758 1002319
rect 362954 1002279 368758 1002307
rect 362954 1002267 362960 1002279
rect 368752 1002267 368758 1002279
rect 368810 1002267 368816 1002319
rect 377680 1002267 377686 1002319
rect 377738 1002307 377744 1002319
rect 383440 1002307 383446 1002319
rect 377738 1002279 383446 1002307
rect 377738 1002267 377744 1002279
rect 383440 1002267 383446 1002279
rect 383498 1002267 383504 1002319
rect 430192 1002267 430198 1002319
rect 430250 1002307 430256 1002319
rect 449200 1002307 449206 1002319
rect 430250 1002279 449206 1002307
rect 430250 1002267 430256 1002279
rect 449200 1002267 449206 1002279
rect 449258 1002267 449264 1002319
rect 489520 1002267 489526 1002319
rect 489578 1002307 489584 1002319
rect 519856 1002307 519862 1002319
rect 489578 1002279 519862 1002307
rect 489578 1002267 489584 1002279
rect 519856 1002267 519862 1002279
rect 519914 1002267 519920 1002319
rect 555376 1002267 555382 1002319
rect 555434 1002307 555440 1002319
rect 567376 1002307 567382 1002319
rect 555434 1002279 567382 1002307
rect 555434 1002267 555440 1002279
rect 567376 1002267 567382 1002279
rect 567434 1002267 567440 1002319
rect 246544 1002233 246550 1002245
rect 246541 1002205 246550 1002233
rect 246544 1002193 246550 1002205
rect 246602 1002193 246608 1002245
rect 506224 1001453 506230 1001505
rect 506282 1001493 506288 1001505
rect 518512 1001493 518518 1001505
rect 506282 1001465 518518 1001493
rect 506282 1001453 506288 1001465
rect 518512 1001453 518518 1001465
rect 518570 1001453 518576 1001505
rect 557776 1001305 557782 1001357
rect 557834 1001345 557840 1001357
rect 571024 1001345 571030 1001357
rect 557834 1001317 571030 1001345
rect 557834 1001305 557840 1001317
rect 571024 1001305 571030 1001317
rect 571082 1001305 571088 1001357
rect 465712 1001009 465718 1001061
rect 465770 1001049 465776 1001061
rect 472624 1001049 472630 1001061
rect 465770 1001021 472630 1001049
rect 465770 1001009 465776 1001021
rect 472624 1001009 472630 1001021
rect 472682 1001009 472688 1001061
rect 443632 1000935 443638 1000987
rect 443690 1000975 443696 1000987
rect 472432 1000975 472438 1000987
rect 443690 1000947 472438 1000975
rect 443690 1000935 443696 1000947
rect 472432 1000935 472438 1000947
rect 472490 1000935 472496 1000987
rect 507856 1000935 507862 1000987
rect 507914 1000975 507920 1000987
rect 512656 1000975 512662 1000987
rect 507914 1000947 512662 1000975
rect 507914 1000935 507920 1000947
rect 512656 1000935 512662 1000947
rect 512714 1000935 512720 1000987
rect 356368 1000861 356374 1000913
rect 356426 1000901 356432 1000913
rect 377200 1000901 377206 1000913
rect 356426 1000873 377206 1000901
rect 356426 1000861 356432 1000873
rect 377200 1000861 377206 1000873
rect 377258 1000861 377264 1000913
rect 429904 1000861 429910 1000913
rect 429962 1000901 429968 1000913
rect 472624 1000901 472630 1000913
rect 429962 1000873 472630 1000901
rect 429962 1000861 429968 1000873
rect 472624 1000861 472630 1000873
rect 472682 1000861 472688 1000913
rect 552304 1000861 552310 1000913
rect 552362 1000901 552368 1000913
rect 573232 1000901 573238 1000913
rect 552362 1000873 573238 1000901
rect 552362 1000861 552368 1000873
rect 573232 1000861 573238 1000873
rect 573290 1000861 573296 1000913
rect 143824 1000787 143830 1000839
rect 143882 1000827 143888 1000839
rect 157648 1000827 157654 1000839
rect 143882 1000799 157654 1000827
rect 143882 1000787 143888 1000799
rect 157648 1000787 157654 1000799
rect 157706 1000787 157712 1000839
rect 195184 1000787 195190 1000839
rect 195242 1000827 195248 1000839
rect 209104 1000827 209110 1000839
rect 195242 1000799 209110 1000827
rect 195242 1000787 195248 1000799
rect 209104 1000787 209110 1000799
rect 209162 1000787 209168 1000839
rect 360208 1000787 360214 1000839
rect 360266 1000827 360272 1000839
rect 383632 1000827 383638 1000839
rect 360266 1000799 383638 1000827
rect 360266 1000787 360272 1000799
rect 383632 1000787 383638 1000799
rect 383690 1000787 383696 1000839
rect 430960 1000787 430966 1000839
rect 431018 1000827 431024 1000839
rect 472528 1000827 472534 1000839
rect 431018 1000799 472534 1000827
rect 431018 1000787 431024 1000799
rect 472528 1000787 472534 1000799
rect 472586 1000787 472592 1000839
rect 500752 1000787 500758 1000839
rect 500810 1000827 500816 1000839
rect 523312 1000827 523318 1000839
rect 500810 1000799 523318 1000827
rect 500810 1000787 500816 1000799
rect 523312 1000787 523318 1000799
rect 523370 1000787 523376 1000839
rect 552976 1000787 552982 1000839
rect 553034 1000827 553040 1000839
rect 575152 1000827 575158 1000839
rect 553034 1000799 575158 1000827
rect 553034 1000787 553040 1000799
rect 575152 1000787 575158 1000799
rect 575210 1000787 575216 1000839
rect 506896 1000639 506902 1000691
rect 506954 1000679 506960 1000691
rect 512080 1000679 512086 1000691
rect 506954 1000651 512086 1000679
rect 506954 1000639 506960 1000651
rect 512080 1000639 512086 1000651
rect 512138 1000639 512144 1000691
rect 610672 999751 610678 999803
rect 610730 999791 610736 999803
rect 625840 999791 625846 999803
rect 610730 999763 625846 999791
rect 610730 999751 610736 999763
rect 625840 999751 625846 999763
rect 625898 999751 625904 999803
rect 502000 999677 502006 999729
rect 502058 999717 502064 999729
rect 512080 999717 512086 999729
rect 502058 999689 512086 999717
rect 502058 999677 502064 999689
rect 512080 999677 512086 999689
rect 512138 999677 512144 999729
rect 609040 999677 609046 999729
rect 609098 999717 609104 999729
rect 625744 999717 625750 999729
rect 609098 999689 625750 999717
rect 609098 999677 609104 999689
rect 625744 999677 625750 999689
rect 625802 999677 625808 999729
rect 247024 999603 247030 999655
rect 247082 999643 247088 999655
rect 258832 999643 258838 999655
rect 247082 999615 258838 999643
rect 247082 999603 247088 999615
rect 258832 999603 258838 999615
rect 258890 999603 258896 999655
rect 610576 999603 610582 999655
rect 610634 999643 610640 999655
rect 625648 999643 625654 999655
rect 610634 999615 625654 999643
rect 610634 999603 610640 999615
rect 625648 999603 625654 999615
rect 625706 999603 625712 999655
rect 246736 999529 246742 999581
rect 246794 999569 246800 999581
rect 258352 999569 258358 999581
rect 246794 999541 258358 999569
rect 246794 999529 246800 999541
rect 258352 999529 258358 999541
rect 258410 999529 258416 999581
rect 298288 999529 298294 999581
rect 298346 999569 298352 999581
rect 312112 999569 312118 999581
rect 298346 999541 312118 999569
rect 298346 999529 298352 999541
rect 312112 999529 312118 999541
rect 312170 999529 312176 999581
rect 504688 999529 504694 999581
rect 504746 999569 504752 999581
rect 512080 999569 512086 999581
rect 504746 999541 512086 999569
rect 504746 999529 504752 999541
rect 512080 999529 512086 999541
rect 512138 999529 512144 999581
rect 596272 999529 596278 999581
rect 596330 999569 596336 999581
rect 625552 999569 625558 999581
rect 596330 999541 625558 999569
rect 596330 999529 596336 999541
rect 625552 999529 625558 999541
rect 625610 999529 625616 999581
rect 92560 999455 92566 999507
rect 92618 999495 92624 999507
rect 92618 999467 106430 999495
rect 92618 999455 92624 999467
rect 92368 999381 92374 999433
rect 92426 999421 92432 999433
rect 106288 999421 106294 999433
rect 92426 999393 106294 999421
rect 92426 999381 92432 999393
rect 106288 999381 106294 999393
rect 106346 999381 106352 999433
rect 106402 999421 106430 999467
rect 143728 999455 143734 999507
rect 143786 999495 143792 999507
rect 155536 999495 155542 999507
rect 143786 999467 155542 999495
rect 143786 999455 143792 999467
rect 155536 999455 155542 999467
rect 155594 999455 155600 999507
rect 246832 999455 246838 999507
rect 246890 999495 246896 999507
rect 260464 999495 260470 999507
rect 246890 999467 260470 999495
rect 246890 999455 246896 999467
rect 260464 999455 260470 999467
rect 260522 999455 260528 999507
rect 298384 999455 298390 999507
rect 298442 999495 298448 999507
rect 310480 999495 310486 999507
rect 298442 999467 310486 999495
rect 298442 999455 298448 999467
rect 310480 999455 310486 999467
rect 310538 999455 310544 999507
rect 593296 999455 593302 999507
rect 593354 999495 593360 999507
rect 625840 999495 625846 999507
rect 593354 999467 625846 999495
rect 593354 999455 593360 999467
rect 625840 999455 625846 999467
rect 625898 999455 625904 999507
rect 126640 999421 126646 999433
rect 106402 999393 126646 999421
rect 126640 999381 126646 999393
rect 126698 999381 126704 999433
rect 144016 999381 144022 999433
rect 144074 999421 144080 999433
rect 146800 999421 146806 999433
rect 144074 999393 146806 999421
rect 144074 999381 144080 999393
rect 146800 999381 146806 999393
rect 146858 999381 146864 999433
rect 195088 999381 195094 999433
rect 195146 999421 195152 999433
rect 206896 999421 206902 999433
rect 195146 999393 206902 999421
rect 195146 999381 195152 999393
rect 206896 999381 206902 999393
rect 206954 999381 206960 999433
rect 246928 999381 246934 999433
rect 246986 999421 246992 999433
rect 279280 999421 279286 999433
rect 246986 999393 279286 999421
rect 246986 999381 246992 999393
rect 279280 999381 279286 999393
rect 279338 999381 279344 999433
rect 298096 999381 298102 999433
rect 298154 999421 298160 999433
rect 309904 999421 309910 999433
rect 298154 999393 309910 999421
rect 298154 999381 298160 999393
rect 309904 999381 309910 999393
rect 309962 999381 309968 999433
rect 357136 999381 357142 999433
rect 357194 999421 357200 999433
rect 357194 999393 376382 999421
rect 357194 999381 357200 999393
rect 313744 999307 313750 999359
rect 313802 999347 313808 999359
rect 331120 999347 331126 999359
rect 313802 999319 331126 999347
rect 313802 999307 313808 999319
rect 331120 999307 331126 999319
rect 331178 999307 331184 999359
rect 376354 999347 376382 999393
rect 377104 999381 377110 999433
rect 377162 999421 377168 999433
rect 383536 999421 383542 999433
rect 377162 999393 383542 999421
rect 377162 999381 377168 999393
rect 383536 999381 383542 999393
rect 383594 999381 383600 999433
rect 459280 999381 459286 999433
rect 459338 999421 459344 999433
rect 459338 999393 462302 999421
rect 459338 999381 459344 999393
rect 383152 999347 383158 999359
rect 376354 999319 383158 999347
rect 383152 999307 383158 999319
rect 383210 999307 383216 999359
rect 462274 999347 462302 999393
rect 500176 999381 500182 999433
rect 500234 999421 500240 999433
rect 515824 999421 515830 999433
rect 500234 999393 515830 999421
rect 500234 999381 500240 999393
rect 515824 999381 515830 999393
rect 515882 999381 515888 999433
rect 596176 999381 596182 999433
rect 596234 999421 596240 999433
rect 625456 999421 625462 999433
rect 596234 999393 625462 999421
rect 596234 999381 596240 999393
rect 625456 999381 625462 999393
rect 625514 999381 625520 999433
rect 464752 999347 464758 999359
rect 462274 999319 464758 999347
rect 464752 999307 464758 999319
rect 464810 999307 464816 999359
rect 302992 999233 302998 999285
rect 303050 999273 303056 999285
rect 304336 999273 304342 999285
rect 303050 999245 304342 999273
rect 303050 999233 303056 999245
rect 304336 999233 304342 999245
rect 304394 999273 304400 999285
rect 304912 999273 304918 999285
rect 304394 999245 304918 999273
rect 304394 999233 304400 999245
rect 304912 999233 304918 999245
rect 304970 999233 304976 999285
rect 364528 999159 364534 999211
rect 364586 999199 364592 999211
rect 380176 999199 380182 999211
rect 364586 999171 380182 999199
rect 364586 999159 364592 999171
rect 380176 999159 380182 999171
rect 380234 999159 380240 999211
rect 557200 999085 557206 999137
rect 557258 999125 557264 999137
rect 573808 999125 573814 999137
rect 557258 999097 573814 999125
rect 557258 999085 557264 999097
rect 573808 999085 573814 999097
rect 573866 999085 573872 999137
rect 558832 998937 558838 998989
rect 558890 998977 558896 998989
rect 573520 998977 573526 998989
rect 558890 998949 573526 998977
rect 558890 998937 558896 998949
rect 573520 998937 573526 998949
rect 573578 998937 573584 998989
rect 368848 998641 368854 998693
rect 368906 998681 368912 998693
rect 374512 998681 374518 998693
rect 368906 998653 374518 998681
rect 368906 998641 368912 998653
rect 374512 998641 374518 998653
rect 374570 998641 374576 998693
rect 377200 997827 377206 997879
rect 377258 997867 377264 997879
rect 383056 997867 383062 997879
rect 377258 997839 383062 997867
rect 377258 997827 377264 997839
rect 383056 997827 383062 997839
rect 383114 997827 383120 997879
rect 314800 997679 314806 997731
rect 314858 997719 314864 997731
rect 365200 997719 365206 997731
rect 314858 997691 365206 997719
rect 314858 997679 314864 997691
rect 365200 997679 365206 997691
rect 365258 997679 365264 997731
rect 555952 997679 555958 997731
rect 556010 997719 556016 997731
rect 593296 997719 593302 997731
rect 556010 997691 593302 997719
rect 556010 997679 556016 997691
rect 593296 997679 593302 997691
rect 593354 997679 593360 997731
rect 331120 997605 331126 997657
rect 331178 997645 331184 997657
rect 364528 997645 364534 997657
rect 331178 997617 364534 997645
rect 331178 997605 331184 997617
rect 364528 997605 364534 997617
rect 364586 997605 364592 997657
rect 567472 997605 567478 997657
rect 567530 997645 567536 997657
rect 596176 997645 596182 997657
rect 567530 997617 596182 997645
rect 567530 997605 567536 997617
rect 596176 997605 596182 997617
rect 596234 997605 596240 997657
rect 567376 997531 567382 997583
rect 567434 997571 567440 997583
rect 596272 997571 596278 997583
rect 567434 997543 596278 997571
rect 567434 997531 567440 997543
rect 596272 997531 596278 997543
rect 596330 997531 596336 997583
rect 571024 997457 571030 997509
rect 571082 997497 571088 997509
rect 610576 997497 610582 997509
rect 571082 997469 610582 997497
rect 571082 997457 571088 997469
rect 610576 997457 610582 997469
rect 610634 997457 610640 997509
rect 558160 997383 558166 997435
rect 558218 997423 558224 997435
rect 609040 997423 609046 997435
rect 558218 997395 609046 997423
rect 558218 997383 558224 997395
rect 609040 997383 609046 997395
rect 609098 997383 609104 997435
rect 559408 997309 559414 997361
rect 559466 997349 559472 997361
rect 610672 997349 610678 997361
rect 559466 997321 610678 997349
rect 559466 997309 559472 997321
rect 610672 997309 610678 997321
rect 610730 997309 610736 997361
rect 463504 997161 463510 997213
rect 463562 997201 463568 997213
rect 465328 997201 465334 997213
rect 463562 997173 465334 997201
rect 463562 997161 463568 997173
rect 465328 997161 465334 997173
rect 465386 997161 465392 997213
rect 298096 997087 298102 997139
rect 298154 997127 298160 997139
rect 313744 997127 313750 997139
rect 298154 997099 313750 997127
rect 298154 997087 298160 997099
rect 313744 997087 313750 997099
rect 313802 997087 313808 997139
rect 368752 997087 368758 997139
rect 368810 997127 368816 997139
rect 377104 997127 377110 997139
rect 368810 997099 377110 997127
rect 368810 997087 368816 997099
rect 377104 997087 377110 997099
rect 377162 997087 377168 997139
rect 507280 996569 507286 996621
rect 507338 996609 507344 996621
rect 523408 996609 523414 996621
rect 507338 996581 523414 996609
rect 507338 996569 507344 996581
rect 523408 996569 523414 996581
rect 523466 996569 523472 996621
rect 144112 996495 144118 996547
rect 144170 996535 144176 996547
rect 156016 996535 156022 996547
rect 144170 996507 156022 996535
rect 144170 996495 144176 996507
rect 156016 996495 156022 996507
rect 156074 996495 156080 996547
rect 195760 996495 195766 996547
rect 195818 996535 195824 996547
rect 205264 996535 205270 996547
rect 195818 996507 205270 996535
rect 195818 996495 195824 996507
rect 205264 996495 205270 996507
rect 205322 996495 205328 996547
rect 247120 996495 247126 996547
rect 247178 996535 247184 996547
rect 259984 996535 259990 996547
rect 247178 996507 259990 996535
rect 247178 996495 247184 996507
rect 259984 996495 259990 996507
rect 260042 996495 260048 996547
rect 368656 996495 368662 996547
rect 368714 996535 368720 996547
rect 377200 996535 377206 996547
rect 368714 996507 377206 996535
rect 368714 996495 368720 996507
rect 377200 996495 377206 996507
rect 377258 996495 377264 996547
rect 505648 996495 505654 996547
rect 505706 996535 505712 996547
rect 521200 996535 521206 996547
rect 505706 996507 521206 996535
rect 505706 996495 505712 996507
rect 521200 996495 521206 996507
rect 521258 996495 521264 996547
rect 210160 996421 210166 996473
rect 210218 996461 210224 996473
rect 225424 996461 225430 996473
rect 210218 996433 225430 996461
rect 210218 996421 210224 996433
rect 225424 996421 225430 996433
rect 225482 996421 225488 996473
rect 313168 996421 313174 996473
rect 313226 996461 313232 996473
rect 363952 996461 363958 996473
rect 313226 996433 363958 996461
rect 313226 996421 313232 996433
rect 363952 996421 363958 996433
rect 364010 996421 364016 996473
rect 280240 996239 280246 996251
rect 262114 996211 280246 996239
rect 262114 996177 262142 996211
rect 280240 996199 280246 996211
rect 280298 996199 280304 996251
rect 432592 996239 432598 996251
rect 430978 996211 432598 996239
rect 107920 996125 107926 996177
rect 107978 996165 107984 996177
rect 159760 996165 159766 996177
rect 107978 996137 159766 996165
rect 107978 996125 107984 996137
rect 159760 996125 159766 996137
rect 159818 996165 159824 996177
rect 178480 996165 178486 996177
rect 159818 996137 178486 996165
rect 159818 996125 159824 996137
rect 178480 996125 178486 996137
rect 178538 996125 178544 996177
rect 198640 996125 198646 996177
rect 198698 996165 198704 996177
rect 204016 996165 204022 996177
rect 198698 996137 204022 996165
rect 198698 996125 198704 996137
rect 204016 996125 204022 996137
rect 204074 996125 204080 996177
rect 262096 996165 262102 996177
rect 210658 996137 262102 996165
rect 107536 996051 107542 996103
rect 107594 996091 107600 996103
rect 159184 996091 159190 996103
rect 107594 996063 159190 996091
rect 107594 996051 107600 996063
rect 159184 996051 159190 996063
rect 159242 996091 159248 996103
rect 210160 996091 210166 996103
rect 159242 996063 210166 996091
rect 159242 996051 159248 996063
rect 210160 996051 210166 996063
rect 210218 996051 210224 996103
rect 210658 996029 210686 996137
rect 262096 996125 262102 996137
rect 262154 996125 262160 996177
rect 263056 996125 263062 996177
rect 263114 996165 263120 996177
rect 314800 996165 314806 996177
rect 263114 996137 314806 996165
rect 263114 996125 263120 996137
rect 314800 996125 314806 996137
rect 314858 996125 314864 996177
rect 368656 996125 368662 996177
rect 368714 996165 368720 996177
rect 430978 996165 431006 996211
rect 432592 996199 432598 996211
rect 432650 996199 432656 996251
rect 508336 996199 508342 996251
rect 508394 996239 508400 996251
rect 508394 996211 509726 996239
rect 508394 996199 508400 996211
rect 368714 996137 431006 996165
rect 368714 996125 368720 996137
rect 432496 996125 432502 996177
rect 432554 996165 432560 996177
rect 509584 996165 509590 996177
rect 432554 996137 509590 996165
rect 432554 996125 432560 996137
rect 509584 996125 509590 996137
rect 509642 996125 509648 996177
rect 225424 996051 225430 996103
rect 225482 996091 225488 996103
rect 262000 996091 262006 996103
rect 225482 996063 262006 996091
rect 225482 996051 225488 996063
rect 262000 996051 262006 996063
rect 262058 996091 262064 996103
rect 313168 996091 313174 996103
rect 262058 996063 313174 996091
rect 262058 996051 262064 996063
rect 313168 996051 313174 996063
rect 313226 996051 313232 996103
rect 380176 996051 380182 996103
rect 380234 996091 380240 996103
rect 434992 996091 434998 996103
rect 380234 996063 434998 996091
rect 380234 996051 380240 996063
rect 434992 996051 434998 996063
rect 435050 996051 435056 996103
rect 470800 996051 470806 996103
rect 470858 996091 470864 996103
rect 508528 996091 508534 996103
rect 470858 996063 508534 996091
rect 470858 996051 470864 996063
rect 508528 996051 508534 996063
rect 508586 996051 508592 996103
rect 509698 996091 509726 996211
rect 518416 996125 518422 996177
rect 518474 996165 518480 996177
rect 561040 996165 561046 996177
rect 518474 996137 561046 996165
rect 518474 996125 518480 996137
rect 561040 996125 561046 996137
rect 561098 996125 561104 996177
rect 559792 996091 559798 996103
rect 509698 996063 559798 996091
rect 559792 996051 559798 996063
rect 559850 996051 559856 996103
rect 108976 995977 108982 996029
rect 109034 996017 109040 996029
rect 160432 996017 160438 996029
rect 109034 995989 160438 996017
rect 109034 995977 109040 995989
rect 160432 995977 160438 995989
rect 160490 995977 160496 996029
rect 178480 995977 178486 996029
rect 178538 996017 178544 996029
rect 210640 996017 210646 996029
rect 178538 995989 210646 996017
rect 178538 995977 178544 995989
rect 210640 995977 210646 995989
rect 210698 995977 210704 996029
rect 222736 995977 222742 996029
rect 222794 996017 222800 996029
rect 263248 996017 263254 996029
rect 222794 995989 263254 996017
rect 222794 995977 222800 995989
rect 263248 995977 263254 995989
rect 263306 995977 263312 996029
rect 299440 996017 299446 996029
rect 283810 995989 299446 996017
rect 94960 995903 94966 995955
rect 95018 995943 95024 995955
rect 102928 995943 102934 995955
rect 95018 995915 102934 995943
rect 95018 995903 95024 995915
rect 102928 995903 102934 995915
rect 102986 995903 102992 995955
rect 146800 995903 146806 995955
rect 146858 995943 146864 995955
rect 152080 995943 152086 995955
rect 146858 995915 152086 995943
rect 146858 995903 146864 995915
rect 152080 995903 152086 995915
rect 152138 995903 152144 995955
rect 172816 995903 172822 995955
rect 172874 995943 172880 995955
rect 211792 995943 211798 995955
rect 172874 995915 211798 995943
rect 172874 995903 172880 995915
rect 211792 995903 211798 995915
rect 211850 995903 211856 995955
rect 97840 995869 97846 995881
rect 82306 995841 97846 995869
rect 82306 995807 82334 995841
rect 97840 995829 97846 995841
rect 97898 995829 97904 995881
rect 144016 995869 144022 995881
rect 137410 995841 144022 995869
rect 137410 995807 137438 995841
rect 144016 995829 144022 995841
rect 144074 995829 144080 995881
rect 183778 995841 195806 995869
rect 183778 995807 183806 995841
rect 82288 995755 82294 995807
rect 82346 995755 82352 995807
rect 91504 995755 91510 995807
rect 91562 995795 91568 995807
rect 92272 995795 92278 995807
rect 91562 995767 92278 995795
rect 91562 995755 91568 995767
rect 92272 995755 92278 995767
rect 92330 995755 92336 995807
rect 93520 995755 93526 995807
rect 93578 995795 93584 995807
rect 97936 995795 97942 995807
rect 93578 995767 97942 995795
rect 93578 995755 93584 995767
rect 97936 995755 97942 995767
rect 97994 995755 98000 995807
rect 137392 995755 137398 995807
rect 137450 995755 137456 995807
rect 137968 995755 137974 995807
rect 138026 995795 138032 995807
rect 143632 995795 143638 995807
rect 138026 995767 143638 995795
rect 138026 995755 138032 995767
rect 143632 995755 143638 995767
rect 143690 995755 143696 995807
rect 149584 995755 149590 995807
rect 149642 995795 149648 995807
rect 154864 995795 154870 995807
rect 149642 995767 154870 995795
rect 149642 995755 149648 995767
rect 154864 995755 154870 995767
rect 154922 995755 154928 995807
rect 183760 995755 183766 995807
rect 183818 995755 183824 995807
rect 195778 995795 195806 995841
rect 198640 995829 198646 995881
rect 198698 995869 198704 995881
rect 202480 995869 202486 995881
rect 198698 995841 202486 995869
rect 198698 995829 198704 995841
rect 202480 995829 202486 995841
rect 202538 995829 202544 995881
rect 254512 995869 254518 995881
rect 239554 995841 254518 995869
rect 239554 995807 239582 995841
rect 254512 995829 254518 995841
rect 254570 995829 254576 995881
rect 283810 995807 283838 995989
rect 299440 995977 299446 995989
rect 299498 995977 299504 996029
rect 363952 995977 363958 996029
rect 364010 996017 364016 996029
rect 430960 996017 430966 996029
rect 364010 995989 430966 996017
rect 364010 995977 364016 995989
rect 430960 995977 430966 995989
rect 431018 996017 431024 996029
rect 436912 996017 436918 996029
rect 431018 995989 436918 996017
rect 431018 995977 431024 995989
rect 436912 995977 436918 995989
rect 436970 995977 436976 996029
rect 508546 996017 508574 996051
rect 560176 996017 560182 996029
rect 508546 995989 560182 996017
rect 560176 995977 560182 995989
rect 560234 995977 560240 996029
rect 471376 995903 471382 995955
rect 471434 995943 471440 995955
rect 508336 995943 508342 995955
rect 471434 995915 508342 995943
rect 471434 995903 471440 995915
rect 508336 995903 508342 995915
rect 508394 995903 508400 995955
rect 510544 995903 510550 995955
rect 510602 995943 510608 995955
rect 515728 995943 515734 995955
rect 510602 995915 515734 995943
rect 510602 995903 510608 995915
rect 515728 995903 515734 995915
rect 515786 995903 515792 995955
rect 523696 995903 523702 995955
rect 523754 995943 523760 995955
rect 523754 995915 529886 995943
rect 523754 995903 523760 995915
rect 299248 995869 299254 995881
rect 290722 995841 299254 995869
rect 290722 995807 290750 995841
rect 299248 995829 299254 995841
rect 299306 995829 299312 995881
rect 383440 995829 383446 995881
rect 383498 995869 383504 995881
rect 383498 995841 388862 995869
rect 383498 995829 383504 995841
rect 388834 995807 388862 995841
rect 472432 995829 472438 995881
rect 472490 995869 472496 995881
rect 472490 995841 476990 995869
rect 472490 995829 472496 995841
rect 476962 995807 476990 995841
rect 523888 995829 523894 995881
rect 523946 995869 523952 995881
rect 523946 995841 528446 995869
rect 523946 995829 523952 995841
rect 528418 995807 528446 995841
rect 529858 995807 529886 995915
rect 561904 995903 561910 995955
rect 561962 995943 561968 995955
rect 569776 995943 569782 995955
rect 561962 995915 569782 995943
rect 561962 995903 561968 995915
rect 569776 995903 569782 995915
rect 569834 995903 569840 995955
rect 625456 995903 625462 995955
rect 625514 995943 625520 995955
rect 625514 995915 631550 995943
rect 625514 995903 625520 995915
rect 625648 995829 625654 995881
rect 625706 995869 625712 995881
rect 625706 995841 629630 995869
rect 625706 995829 625712 995841
rect 629602 995807 629630 995841
rect 631522 995807 631550 995915
rect 205648 995795 205654 995807
rect 195778 995767 205654 995795
rect 205648 995755 205654 995767
rect 205706 995755 205712 995807
rect 239536 995755 239542 995807
rect 239594 995755 239600 995807
rect 240880 995755 240886 995807
rect 240938 995795 240944 995807
rect 246640 995795 246646 995807
rect 240938 995767 246646 995795
rect 240938 995755 240944 995767
rect 246640 995755 246646 995767
rect 246698 995755 246704 995807
rect 246928 995755 246934 995807
rect 246986 995795 246992 995807
rect 257680 995795 257686 995807
rect 246986 995767 257686 995795
rect 246986 995755 246992 995767
rect 257680 995755 257686 995767
rect 257738 995755 257744 995807
rect 283792 995755 283798 995807
rect 283850 995755 283856 995807
rect 290704 995755 290710 995807
rect 290762 995755 290768 995807
rect 291184 995755 291190 995807
rect 291242 995795 291248 995807
rect 306064 995795 306070 995807
rect 291242 995767 306070 995795
rect 291242 995755 291248 995767
rect 306064 995755 306070 995767
rect 306122 995755 306128 995807
rect 366736 995755 366742 995807
rect 366794 995795 366800 995807
rect 371632 995795 371638 995807
rect 366794 995767 371638 995795
rect 366794 995755 366800 995767
rect 371632 995755 371638 995767
rect 371690 995755 371696 995807
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384976 995795 384982 995807
rect 383690 995767 384982 995795
rect 383690 995755 383696 995767
rect 384976 995755 384982 995767
rect 385034 995755 385040 995807
rect 388816 995755 388822 995807
rect 388874 995755 388880 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 473296 995795 473302 995807
rect 472682 995767 473302 995795
rect 472682 995755 472688 995767
rect 473296 995755 473302 995767
rect 473354 995755 473360 995807
rect 476944 995755 476950 995807
rect 477002 995755 477008 995807
rect 511120 995755 511126 995807
rect 511178 995795 511184 995807
rect 515632 995795 515638 995807
rect 511178 995767 515638 995795
rect 511178 995755 511184 995767
rect 515632 995755 515638 995767
rect 515690 995755 515696 995807
rect 524176 995755 524182 995807
rect 524234 995795 524240 995807
rect 525328 995795 525334 995807
rect 524234 995767 525334 995795
rect 524234 995755 524240 995767
rect 525328 995755 525334 995767
rect 525386 995755 525392 995807
rect 528400 995755 528406 995807
rect 528458 995755 528464 995807
rect 529840 995755 529846 995807
rect 529898 995755 529904 995807
rect 559792 995755 559798 995807
rect 559850 995795 559856 995807
rect 564592 995795 564598 995807
rect 559850 995767 564598 995795
rect 559850 995755 559856 995767
rect 564592 995755 564598 995767
rect 564650 995755 564656 995807
rect 625840 995755 625846 995807
rect 625898 995795 625904 995807
rect 627088 995795 627094 995807
rect 625898 995767 627094 995795
rect 625898 995755 625904 995767
rect 627088 995755 627094 995767
rect 627146 995755 627152 995807
rect 629584 995755 629590 995807
rect 629642 995755 629648 995807
rect 631504 995755 631510 995807
rect 631562 995755 631568 995807
rect 89776 995681 89782 995733
rect 89834 995721 89840 995733
rect 92368 995721 92374 995733
rect 89834 995693 92374 995721
rect 89834 995681 89840 995693
rect 92368 995681 92374 995693
rect 92426 995681 92432 995733
rect 136720 995681 136726 995733
rect 136778 995721 136784 995733
rect 151696 995721 151702 995733
rect 136778 995693 151702 995721
rect 136778 995681 136784 995693
rect 151696 995681 151702 995693
rect 151754 995681 151760 995733
rect 175696 995681 175702 995733
rect 175754 995721 175760 995733
rect 185200 995721 185206 995733
rect 175754 995693 185206 995721
rect 175754 995681 175760 995693
rect 185200 995681 185206 995693
rect 185258 995681 185264 995733
rect 194416 995681 194422 995733
rect 194474 995721 194480 995733
rect 195088 995721 195094 995733
rect 194474 995693 195094 995721
rect 194474 995681 194480 995693
rect 195088 995681 195094 995693
rect 195146 995681 195152 995733
rect 198448 995681 198454 995733
rect 198506 995721 198512 995733
rect 202960 995721 202966 995733
rect 198506 995693 202966 995721
rect 198506 995681 198512 995693
rect 202960 995681 202966 995693
rect 203018 995681 203024 995733
rect 240304 995681 240310 995733
rect 240362 995721 240368 995733
rect 246544 995721 246550 995733
rect 240362 995693 246550 995721
rect 240362 995681 240368 995693
rect 246544 995681 246550 995693
rect 246602 995681 246608 995733
rect 247600 995681 247606 995733
rect 247658 995721 247664 995733
rect 256144 995721 256150 995733
rect 247658 995693 256150 995721
rect 247658 995681 247664 995693
rect 256144 995681 256150 995693
rect 256202 995681 256208 995733
rect 291760 995681 291766 995733
rect 291818 995721 291824 995733
rect 306448 995721 306454 995733
rect 291818 995693 306454 995721
rect 291818 995681 291824 995693
rect 306448 995681 306454 995693
rect 306506 995681 306512 995733
rect 366160 995681 366166 995733
rect 366218 995721 366224 995733
rect 371728 995721 371734 995733
rect 366218 995693 371734 995721
rect 366218 995681 366224 995693
rect 371728 995681 371734 995693
rect 371786 995681 371792 995733
rect 383536 995681 383542 995733
rect 383594 995721 383600 995733
rect 386032 995721 386038 995733
rect 383594 995693 386038 995721
rect 383594 995681 383600 995693
rect 386032 995681 386038 995693
rect 386090 995681 386096 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 474640 995721 474646 995733
rect 472586 995693 474646 995721
rect 472586 995681 472592 995693
rect 474640 995681 474646 995693
rect 474698 995681 474704 995733
rect 523984 995681 523990 995733
rect 524042 995721 524048 995733
rect 524752 995721 524758 995733
rect 524042 995693 524758 995721
rect 524042 995681 524048 995693
rect 524752 995681 524758 995693
rect 524810 995681 524816 995733
rect 625744 995681 625750 995733
rect 625802 995721 625808 995733
rect 626512 995721 626518 995733
rect 625802 995693 626518 995721
rect 625802 995681 625808 995693
rect 626512 995681 626518 995693
rect 626570 995681 626576 995733
rect 93808 995607 93814 995659
rect 93866 995647 93872 995659
rect 98992 995647 98998 995659
rect 93866 995619 98998 995647
rect 93866 995607 93872 995619
rect 98992 995607 98998 995619
rect 99050 995607 99056 995659
rect 142960 995607 142966 995659
rect 143018 995647 143024 995659
rect 143728 995647 143734 995659
rect 143018 995619 143734 995647
rect 143018 995607 143024 995619
rect 143728 995607 143734 995619
rect 143786 995607 143792 995659
rect 192496 995607 192502 995659
rect 192554 995647 192560 995659
rect 195184 995647 195190 995659
rect 192554 995619 195190 995647
rect 192554 995607 192560 995619
rect 195184 995607 195190 995619
rect 195242 995607 195248 995659
rect 297328 995607 297334 995659
rect 297386 995647 297392 995659
rect 298000 995647 298006 995659
rect 297386 995619 298006 995647
rect 297386 995607 297392 995619
rect 298000 995607 298006 995619
rect 298058 995607 298064 995659
rect 383728 995607 383734 995659
rect 383786 995647 383792 995659
rect 384400 995647 384406 995659
rect 383786 995619 384406 995647
rect 383786 995607 383792 995619
rect 384400 995607 384406 995619
rect 384458 995607 384464 995659
rect 472720 995607 472726 995659
rect 472778 995647 472784 995659
rect 474064 995647 474070 995659
rect 472778 995619 474070 995647
rect 472778 995607 472784 995619
rect 474064 995607 474070 995619
rect 474122 995607 474128 995659
rect 478384 995647 478390 995659
rect 474178 995619 478390 995647
rect 141040 995533 141046 995585
rect 141098 995573 141104 995585
rect 143824 995573 143830 995585
rect 141098 995545 143830 995573
rect 141098 995533 141104 995545
rect 143824 995533 143830 995545
rect 143882 995533 143888 995585
rect 185104 995533 185110 995585
rect 185162 995573 185168 995585
rect 198640 995573 198646 995585
rect 185162 995545 198646 995573
rect 185162 995533 185168 995545
rect 198640 995533 198646 995545
rect 198698 995533 198704 995585
rect 286768 995533 286774 995585
rect 286826 995573 286832 995585
rect 286826 995545 295358 995573
rect 286826 995533 286832 995545
rect 81616 995459 81622 995511
rect 81674 995499 81680 995511
rect 102448 995499 102454 995511
rect 81674 995471 102454 995499
rect 81674 995459 81680 995471
rect 102448 995459 102454 995471
rect 102506 995459 102512 995511
rect 184048 995459 184054 995511
rect 184106 995499 184112 995511
rect 195760 995499 195766 995511
rect 184106 995471 195766 995499
rect 184106 995459 184112 995471
rect 195760 995459 195766 995471
rect 195818 995459 195824 995511
rect 245680 995459 245686 995511
rect 245738 995499 245744 995511
rect 246736 995499 246742 995511
rect 245738 995471 246742 995499
rect 245738 995459 245744 995471
rect 246736 995459 246742 995471
rect 246794 995459 246800 995511
rect 287440 995459 287446 995511
rect 287498 995499 287504 995511
rect 290704 995499 290710 995511
rect 287498 995471 290710 995499
rect 287498 995459 287504 995471
rect 290704 995459 290710 995471
rect 290762 995459 290768 995511
rect 295330 995499 295358 995545
rect 295408 995533 295414 995585
rect 295466 995573 295472 995585
rect 298288 995573 298294 995585
rect 295466 995545 298294 995573
rect 295466 995533 295472 995545
rect 298288 995533 298294 995545
rect 298346 995533 298352 995585
rect 383152 995533 383158 995585
rect 383210 995573 383216 995585
rect 392368 995573 392374 995585
rect 383210 995545 392374 995573
rect 383210 995533 383216 995545
rect 392368 995533 392374 995545
rect 392426 995533 392432 995585
rect 466576 995533 466582 995585
rect 466634 995573 466640 995585
rect 474178 995573 474206 995619
rect 478384 995607 478390 995619
rect 478442 995607 478448 995659
rect 523792 995607 523798 995659
rect 523850 995647 523856 995659
rect 526096 995647 526102 995659
rect 523850 995619 526102 995647
rect 523850 995607 523856 995619
rect 526096 995607 526102 995619
rect 526154 995607 526160 995659
rect 560176 995607 560182 995659
rect 560234 995647 560240 995659
rect 564496 995647 564502 995659
rect 560234 995619 564502 995647
rect 560234 995607 560240 995619
rect 564496 995607 564502 995619
rect 564554 995607 564560 995659
rect 625552 995607 625558 995659
rect 625610 995647 625616 995659
rect 630160 995647 630166 995659
rect 625610 995619 630166 995647
rect 625610 995607 625616 995619
rect 630160 995607 630166 995619
rect 630218 995607 630224 995659
rect 466634 995545 474206 995573
rect 466634 995533 466640 995545
rect 523600 995533 523606 995585
rect 523658 995573 523664 995585
rect 527824 995573 527830 995585
rect 523658 995545 527830 995573
rect 523658 995533 523664 995545
rect 527824 995533 527830 995545
rect 527882 995533 527888 995585
rect 625936 995533 625942 995585
rect 625994 995573 626000 995585
rect 627856 995573 627862 995585
rect 625994 995545 627862 995573
rect 625994 995533 626000 995545
rect 627856 995533 627862 995545
rect 627914 995533 627920 995585
rect 299344 995499 299350 995511
rect 295330 995471 299350 995499
rect 299344 995459 299350 995471
rect 299402 995459 299408 995511
rect 518800 995459 518806 995511
rect 518858 995499 518864 995511
rect 532816 995499 532822 995511
rect 518858 995471 532822 995499
rect 518858 995459 518864 995471
rect 532816 995459 532822 995471
rect 532874 995459 532880 995511
rect 287920 995385 287926 995437
rect 287978 995425 287984 995437
rect 306544 995425 306550 995437
rect 287978 995397 306550 995425
rect 287978 995385 287984 995397
rect 306544 995385 306550 995397
rect 306602 995385 306608 995437
rect 383152 995385 383158 995437
rect 383210 995425 383216 995437
rect 390448 995425 390454 995437
rect 383210 995397 390454 995425
rect 383210 995385 383216 995397
rect 390448 995385 390454 995397
rect 390506 995425 390512 995437
rect 403120 995425 403126 995437
rect 390506 995397 403126 995425
rect 390506 995385 390512 995397
rect 403120 995385 403126 995397
rect 403178 995385 403184 995437
rect 518608 995385 518614 995437
rect 518666 995425 518672 995437
rect 533392 995425 533398 995437
rect 518666 995397 533398 995425
rect 518666 995385 518672 995397
rect 533392 995385 533398 995397
rect 533450 995385 533456 995437
rect 518704 995311 518710 995363
rect 518762 995351 518768 995363
rect 535552 995351 535558 995363
rect 518762 995323 535558 995351
rect 518762 995311 518768 995323
rect 535552 995311 535558 995323
rect 535610 995311 535616 995363
rect 523408 995237 523414 995289
rect 523466 995277 523472 995289
rect 537376 995277 537382 995289
rect 523466 995249 537382 995277
rect 523466 995237 523472 995249
rect 537376 995237 537382 995249
rect 537434 995237 537440 995289
rect 523312 995163 523318 995215
rect 523370 995203 523376 995215
rect 534352 995203 534358 995215
rect 523370 995175 534358 995203
rect 523370 995163 523376 995175
rect 534352 995163 534358 995175
rect 534410 995163 534416 995215
rect 66832 995089 66838 995141
rect 66890 995129 66896 995141
rect 349648 995129 349654 995141
rect 66890 995101 349654 995129
rect 66890 995089 66896 995101
rect 349648 995089 349654 995101
rect 349706 995089 349712 995141
rect 519856 995089 519862 995141
rect 519914 995129 519920 995141
rect 530704 995129 530710 995141
rect 519914 995101 530710 995129
rect 519914 995089 519920 995101
rect 530704 995089 530710 995101
rect 530762 995129 530768 995141
rect 532720 995129 532726 995141
rect 530762 995101 532726 995129
rect 530762 995089 530768 995101
rect 532720 995089 532726 995101
rect 532778 995089 532784 995141
rect 555376 995089 555382 995141
rect 555434 995129 555440 995141
rect 649360 995129 649366 995141
rect 555434 995101 649366 995129
rect 555434 995089 555440 995101
rect 649360 995089 649366 995101
rect 649418 995089 649424 995141
rect 233296 995015 233302 995067
rect 233354 995055 233360 995067
rect 247792 995055 247798 995067
rect 233354 995027 247798 995055
rect 233354 995015 233360 995027
rect 247792 995015 247798 995027
rect 247850 995015 247856 995067
rect 279280 995015 279286 995067
rect 279338 995055 279344 995067
rect 609040 995055 609046 995067
rect 279338 995027 609046 995055
rect 279338 995015 279344 995027
rect 609040 995015 609046 995027
rect 609098 995015 609104 995067
rect 524080 994645 524086 994697
rect 524138 994685 524144 994697
rect 531184 994685 531190 994697
rect 524138 994657 531190 994685
rect 524138 994645 524144 994657
rect 531184 994645 531190 994657
rect 531242 994645 531248 994697
rect 290896 994275 290902 994327
rect 290954 994315 290960 994327
rect 299152 994315 299158 994327
rect 290954 994287 299158 994315
rect 290954 994275 290960 994287
rect 299152 994275 299158 994287
rect 299210 994275 299216 994327
rect 463696 994127 463702 994179
rect 463754 994167 463760 994179
rect 479152 994167 479158 994179
rect 463754 994139 479158 994167
rect 463754 994127 463760 994139
rect 479152 994127 479158 994139
rect 479210 994127 479216 994179
rect 235792 993979 235798 994031
rect 235850 994019 235856 994031
rect 247600 994019 247606 994031
rect 235850 993991 247606 994019
rect 235850 993979 235856 993991
rect 247600 993979 247606 993991
rect 247658 993979 247664 994031
rect 180496 993905 180502 993957
rect 180554 993945 180560 993957
rect 198640 993945 198646 993957
rect 180554 993917 198646 993945
rect 180554 993905 180560 993917
rect 198640 993905 198646 993917
rect 198698 993905 198704 993957
rect 234928 993905 234934 993957
rect 234986 993945 234992 993957
rect 250480 993945 250486 993957
rect 234986 993917 250486 993945
rect 234986 993905 234992 993917
rect 250480 993905 250486 993917
rect 250538 993905 250544 993957
rect 77680 993831 77686 993883
rect 77738 993871 77744 993883
rect 97840 993871 97846 993883
rect 77738 993843 97846 993871
rect 77738 993831 77744 993843
rect 97840 993831 97846 993843
rect 97898 993831 97904 993883
rect 132112 993831 132118 993883
rect 132170 993871 132176 993883
rect 149680 993871 149686 993883
rect 132170 993843 149686 993871
rect 132170 993831 132176 993843
rect 149680 993831 149686 993843
rect 149738 993831 149744 993883
rect 182992 993831 182998 993883
rect 183050 993871 183056 993883
rect 208144 993871 208150 993883
rect 183050 993843 208150 993871
rect 183050 993831 183056 993843
rect 208144 993831 208150 993843
rect 208202 993831 208208 993883
rect 232144 993831 232150 993883
rect 232202 993871 232208 993883
rect 246928 993871 246934 993883
rect 232202 993843 246934 993871
rect 232202 993831 232208 993843
rect 246928 993831 246934 993843
rect 246986 993831 246992 993883
rect 561616 993831 561622 993883
rect 561674 993871 561680 993883
rect 641008 993871 641014 993883
rect 561674 993843 641014 993871
rect 561674 993831 561680 993843
rect 641008 993831 641014 993843
rect 641066 993831 641072 993883
rect 80176 993757 80182 993809
rect 80234 993797 80240 993809
rect 105328 993797 105334 993809
rect 80234 993769 105334 993797
rect 80234 993757 80240 993769
rect 105328 993757 105334 993769
rect 105386 993757 105392 993809
rect 129328 993757 129334 993809
rect 129386 993797 129392 993809
rect 149584 993797 149590 993809
rect 129386 993769 149590 993797
rect 129386 993757 129392 993769
rect 149584 993757 149590 993769
rect 149642 993757 149648 993809
rect 181360 993757 181366 993809
rect 181418 993797 181424 993809
rect 209776 993797 209782 993809
rect 181418 993769 209782 993797
rect 181418 993757 181424 993769
rect 209776 993757 209782 993769
rect 209834 993757 209840 993809
rect 231472 993757 231478 993809
rect 231530 993797 231536 993809
rect 247120 993797 247126 993809
rect 231530 993769 247126 993797
rect 231530 993757 231536 993769
rect 247120 993757 247126 993769
rect 247178 993757 247184 993809
rect 521296 993757 521302 993809
rect 521354 993797 521360 993809
rect 538960 993797 538966 993809
rect 521354 993769 538966 993797
rect 521354 993757 521360 993769
rect 538960 993757 538966 993769
rect 539018 993757 539024 993809
rect 78352 993683 78358 993735
rect 78410 993723 78416 993735
rect 106960 993723 106966 993735
rect 78410 993695 106966 993723
rect 78410 993683 78416 993695
rect 106960 993683 106966 993695
rect 107018 993683 107024 993735
rect 128464 993683 128470 993735
rect 128522 993723 128528 993735
rect 157264 993723 157270 993735
rect 128522 993695 157270 993723
rect 128522 993683 128528 993695
rect 157264 993683 157270 993695
rect 157322 993683 157328 993735
rect 179824 993683 179830 993735
rect 179882 993723 179888 993735
rect 208720 993723 208726 993735
rect 179882 993695 208726 993723
rect 179882 993683 179888 993695
rect 208720 993683 208726 993695
rect 208778 993683 208784 993735
rect 234352 993683 234358 993735
rect 234410 993723 234416 993735
rect 259408 993723 259414 993735
rect 234410 993695 259414 993723
rect 234410 993683 234416 993695
rect 259408 993683 259414 993695
rect 259466 993683 259472 993735
rect 282832 993683 282838 993735
rect 282890 993723 282896 993735
rect 311536 993723 311542 993735
rect 282890 993695 311542 993723
rect 282890 993683 282896 993695
rect 311536 993683 311542 993695
rect 311594 993683 311600 993735
rect 374512 993683 374518 993735
rect 374570 993723 374576 993735
rect 392080 993723 392086 993735
rect 374570 993695 392086 993723
rect 374570 993683 374576 993695
rect 392080 993683 392086 993695
rect 392138 993683 392144 993735
rect 532720 993683 532726 993735
rect 532778 993723 532784 993735
rect 632368 993723 632374 993735
rect 532778 993695 632374 993723
rect 532778 993683 532784 993695
rect 632368 993683 632374 993695
rect 632426 993683 632432 993735
rect 77296 993609 77302 993661
rect 77354 993649 77360 993661
rect 105904 993649 105910 993661
rect 77354 993621 105910 993649
rect 77354 993609 77360 993621
rect 105904 993609 105910 993621
rect 105962 993609 105968 993661
rect 129712 993609 129718 993661
rect 129770 993649 129776 993661
rect 158224 993649 158230 993661
rect 129770 993621 158230 993649
rect 129770 993609 129776 993621
rect 158224 993609 158230 993621
rect 158282 993609 158288 993661
rect 185392 993609 185398 993661
rect 185450 993649 185456 993661
rect 236752 993649 236758 993661
rect 185450 993621 236758 993649
rect 185450 993609 185456 993621
rect 236752 993609 236758 993621
rect 236810 993649 236816 993661
rect 236810 993621 282110 993649
rect 236810 993609 236816 993621
rect 61840 993535 61846 993587
rect 61898 993575 61904 993587
rect 82576 993575 82582 993587
rect 61898 993547 82582 993575
rect 61898 993535 61904 993547
rect 82576 993535 82582 993547
rect 82634 993575 82640 993587
rect 133936 993575 133942 993587
rect 82634 993547 133942 993575
rect 82634 993535 82640 993547
rect 133936 993535 133942 993547
rect 133994 993575 134000 993587
rect 143920 993575 143926 993587
rect 133994 993547 143926 993575
rect 133994 993535 134000 993547
rect 143920 993535 143926 993547
rect 143978 993535 143984 993587
rect 62032 993461 62038 993513
rect 62090 993501 62096 993513
rect 83440 993501 83446 993513
rect 62090 993473 83446 993501
rect 62090 993461 62096 993473
rect 83440 993461 83446 993473
rect 83498 993501 83504 993513
rect 92560 993501 92566 993513
rect 83498 993473 92566 993501
rect 83498 993461 83504 993473
rect 92560 993461 92566 993473
rect 92618 993461 92624 993513
rect 282082 993427 282110 993621
rect 284368 993609 284374 993661
rect 284426 993649 284432 993661
rect 312784 993649 312790 993661
rect 284426 993621 312790 993649
rect 284426 993609 284432 993621
rect 312784 993609 312790 993621
rect 312842 993609 312848 993661
rect 365776 993609 365782 993661
rect 365834 993649 365840 993661
rect 398800 993649 398806 993661
rect 365834 993621 398806 993649
rect 365834 993609 365840 993621
rect 398800 993609 398806 993621
rect 398858 993609 398864 993661
rect 443728 993609 443734 993661
rect 443786 993649 443792 993661
rect 487792 993649 487798 993661
rect 443786 993621 487798 993649
rect 443786 993609 443792 993621
rect 487792 993609 487798 993621
rect 487850 993609 487856 993661
rect 531184 993609 531190 993661
rect 531242 993649 531248 993661
rect 633040 993649 633046 993661
rect 531242 993621 633046 993649
rect 531242 993609 531248 993621
rect 633040 993609 633046 993621
rect 633098 993609 633104 993661
rect 328240 993575 328246 993587
rect 308290 993547 328246 993575
rect 308290 993501 308318 993547
rect 328240 993535 328246 993547
rect 328298 993535 328304 993587
rect 423376 993575 423382 993587
rect 412354 993547 423382 993575
rect 348400 993501 348406 993513
rect 308194 993473 308318 993501
rect 342754 993473 348406 993501
rect 288112 993427 288118 993439
rect 282082 993399 288118 993427
rect 288112 993387 288118 993399
rect 288170 993427 288176 993439
rect 308194 993427 308222 993473
rect 288170 993399 308222 993427
rect 288170 993387 288176 993399
rect 328432 993387 328438 993439
rect 328490 993427 328496 993439
rect 342754 993427 342782 993473
rect 348400 993461 348406 993473
rect 348458 993461 348464 993513
rect 362818 993473 362942 993501
rect 328490 993399 342782 993427
rect 328490 993387 328496 993399
rect 348496 993387 348502 993439
rect 348554 993427 348560 993439
rect 362818 993427 362846 993473
rect 348554 993399 362846 993427
rect 348554 993387 348560 993399
rect 362914 993365 362942 993473
rect 408976 993461 408982 993513
rect 409034 993501 409040 993513
rect 412354 993501 412382 993547
rect 423376 993535 423382 993547
rect 423434 993535 423440 993587
rect 409034 993473 412382 993501
rect 409034 993461 409040 993473
rect 443440 993461 443446 993513
rect 443498 993501 443504 993513
rect 449200 993501 449206 993513
rect 443498 993473 449206 993501
rect 443498 993461 443504 993473
rect 449200 993461 449206 993473
rect 449258 993461 449264 993513
rect 642256 993461 642262 993513
rect 642314 993501 642320 993513
rect 650320 993501 650326 993513
rect 642314 993473 650326 993501
rect 642314 993461 642320 993473
rect 650320 993461 650326 993473
rect 650378 993461 650384 993513
rect 403120 993387 403126 993439
rect 403178 993427 403184 993439
rect 408880 993427 408886 993439
rect 403178 993399 408886 993427
rect 403178 993387 403184 993399
rect 408880 993387 408886 993399
rect 408938 993387 408944 993439
rect 449392 993387 449398 993439
rect 449450 993427 449456 993439
rect 463696 993427 463702 993439
rect 449450 993399 463702 993427
rect 449450 993387 449456 993399
rect 463696 993387 463702 993399
rect 463754 993387 463760 993439
rect 479152 993387 479158 993439
rect 479210 993427 479216 993439
rect 489520 993427 489526 993439
rect 479210 993399 489526 993427
rect 479210 993387 479216 993399
rect 489520 993387 489526 993399
rect 489578 993387 489584 993439
rect 362896 993313 362902 993365
rect 362954 993313 362960 993365
rect 382960 993313 382966 993365
rect 383018 993353 383024 993365
rect 383018 993325 383102 993353
rect 383018 993313 383024 993325
rect 383074 993291 383102 993325
rect 383056 993239 383062 993291
rect 383114 993239 383120 993291
rect 422128 992721 422134 992773
rect 422186 992761 422192 992773
rect 426256 992761 426262 992773
rect 422186 992733 426262 992761
rect 422186 992721 422192 992733
rect 426256 992721 426262 992733
rect 426314 992721 426320 992773
rect 73456 992129 73462 992181
rect 73514 992169 73520 992181
rect 110224 992169 110230 992181
rect 73514 992141 110230 992169
rect 73514 992129 73520 992141
rect 110224 992129 110230 992141
rect 110282 992129 110288 992181
rect 604720 991907 604726 991959
rect 604778 991947 604784 991959
rect 605776 991947 605782 991959
rect 604778 991919 605782 991947
rect 604778 991907 604784 991919
rect 605776 991907 605782 991919
rect 605834 991907 605840 991959
rect 605776 991611 605782 991663
rect 605834 991651 605840 991663
rect 619792 991651 619798 991663
rect 605834 991623 619798 991651
rect 605834 991611 605840 991623
rect 619792 991611 619798 991623
rect 619850 991611 619856 991663
rect 105808 990427 105814 990479
rect 105866 990467 105872 990479
rect 109552 990467 109558 990479
rect 105866 990439 109558 990467
rect 105866 990427 105872 990439
rect 109552 990427 109558 990439
rect 109610 990427 109616 990479
rect 371632 989391 371638 989443
rect 371690 989431 371696 989443
rect 397840 989431 397846 989443
rect 371690 989403 397846 989431
rect 371690 989391 371696 989403
rect 397840 989391 397846 989403
rect 397898 989391 397904 989443
rect 437776 989391 437782 989443
rect 437834 989431 437840 989443
rect 462736 989431 462742 989443
rect 437834 989403 462742 989431
rect 437834 989391 437840 989403
rect 462736 989391 462742 989403
rect 462794 989391 462800 989443
rect 515632 989391 515638 989443
rect 515690 989431 515696 989443
rect 527632 989431 527638 989443
rect 515690 989403 527638 989431
rect 515690 989391 515696 989403
rect 527632 989391 527638 989403
rect 527690 989391 527696 989443
rect 569680 989391 569686 989443
rect 569738 989431 569744 989443
rect 592432 989431 592438 989443
rect 569738 989403 592438 989431
rect 569738 989391 569744 989403
rect 592432 989391 592438 989403
rect 592490 989391 592496 989443
rect 154480 989317 154486 989369
rect 154538 989357 154544 989369
rect 161680 989357 161686 989369
rect 154538 989329 161686 989357
rect 154538 989317 154544 989329
rect 161680 989317 161686 989329
rect 161738 989317 161744 989369
rect 203152 989317 203158 989369
rect 203210 989357 203216 989369
rect 213328 989357 213334 989369
rect 203210 989329 213334 989357
rect 203210 989317 203216 989329
rect 213328 989317 213334 989329
rect 213386 989317 213392 989369
rect 270736 989317 270742 989369
rect 270794 989357 270800 989369
rect 284272 989357 284278 989369
rect 270794 989329 284278 989357
rect 270794 989317 270800 989329
rect 284272 989317 284278 989329
rect 284330 989317 284336 989369
rect 319600 989317 319606 989369
rect 319658 989357 319664 989369
rect 349168 989357 349174 989369
rect 319658 989329 349174 989357
rect 319658 989317 319664 989329
rect 349168 989317 349174 989329
rect 349226 989317 349232 989369
rect 371536 989317 371542 989369
rect 371594 989357 371600 989369
rect 414064 989357 414070 989369
rect 371594 989329 414070 989357
rect 371594 989317 371600 989329
rect 414064 989317 414070 989329
rect 414122 989317 414128 989369
rect 437872 989317 437878 989369
rect 437930 989357 437936 989369
rect 478960 989357 478966 989369
rect 437930 989329 478966 989357
rect 437930 989317 437936 989329
rect 478960 989317 478966 989329
rect 479018 989317 479024 989369
rect 515536 989317 515542 989369
rect 515594 989357 515600 989369
rect 543760 989357 543766 989369
rect 515594 989329 543766 989357
rect 515594 989317 515600 989329
rect 543760 989317 543766 989329
rect 543818 989317 543824 989369
rect 569872 989317 569878 989369
rect 569930 989357 569936 989369
rect 608752 989357 608758 989369
rect 569930 989329 608758 989357
rect 569930 989317 569936 989329
rect 608752 989317 608758 989329
rect 608810 989317 608816 989369
rect 89584 989243 89590 989295
rect 89642 989283 89648 989295
rect 109360 989283 109366 989295
rect 89642 989255 109366 989283
rect 89642 989243 89648 989255
rect 109360 989243 109366 989255
rect 109418 989243 109424 989295
rect 138256 989243 138262 989295
rect 138314 989283 138320 989295
rect 161488 989283 161494 989295
rect 138314 989255 161494 989283
rect 138314 989243 138320 989255
rect 161488 989243 161494 989255
rect 161546 989243 161552 989295
rect 216016 989243 216022 989295
rect 216074 989283 216080 989295
rect 235600 989283 235606 989295
rect 216074 989255 235606 989283
rect 216074 989243 216080 989255
rect 235600 989243 235606 989255
rect 235658 989243 235664 989295
rect 267856 989243 267862 989295
rect 267914 989283 267920 989295
rect 300496 989283 300502 989295
rect 267914 989255 300502 989283
rect 267914 989243 267920 989255
rect 300496 989243 300502 989255
rect 300554 989243 300560 989295
rect 319696 989243 319702 989295
rect 319754 989283 319760 989295
rect 365392 989283 365398 989295
rect 319754 989255 365398 989283
rect 319754 989243 319760 989255
rect 365392 989243 365398 989255
rect 365450 989243 365456 989295
rect 371728 989243 371734 989295
rect 371786 989283 371792 989295
rect 430288 989283 430294 989295
rect 371786 989255 430294 989283
rect 371786 989243 371792 989255
rect 430288 989243 430294 989255
rect 430346 989243 430352 989295
rect 437968 989243 437974 989295
rect 438026 989283 438032 989295
rect 495184 989283 495190 989295
rect 438026 989255 495190 989283
rect 438026 989243 438032 989255
rect 495184 989243 495190 989255
rect 495242 989243 495248 989295
rect 515728 989243 515734 989295
rect 515786 989283 515792 989295
rect 560080 989283 560086 989295
rect 515786 989255 560086 989283
rect 515786 989243 515792 989255
rect 560080 989243 560086 989255
rect 560138 989243 560144 989295
rect 569776 989243 569782 989295
rect 569834 989283 569840 989295
rect 624976 989283 624982 989295
rect 569834 989255 624982 989283
rect 569834 989243 569840 989255
rect 624976 989243 624982 989255
rect 625034 989243 625040 989295
rect 634288 989243 634294 989295
rect 634346 989283 634352 989295
rect 649840 989283 649846 989295
rect 634346 989255 649846 989283
rect 634346 989243 634352 989255
rect 649840 989243 649846 989255
rect 649898 989243 649904 989295
rect 64816 988503 64822 988555
rect 64874 988543 64880 988555
rect 66832 988543 66838 988555
rect 64874 988515 66838 988543
rect 64874 988503 64880 988515
rect 66832 988503 66838 988515
rect 66890 988503 66896 988555
rect 50416 988281 50422 988333
rect 50474 988321 50480 988333
rect 122032 988321 122038 988333
rect 50474 988293 122038 988321
rect 50474 988281 50480 988293
rect 122032 988281 122038 988293
rect 122090 988281 122096 988333
rect 331216 988281 331222 988333
rect 331274 988321 331280 988333
rect 332560 988321 332566 988333
rect 331274 988293 332566 988321
rect 331274 988281 331280 988293
rect 332560 988281 332566 988293
rect 332618 988281 332624 988333
rect 47632 988207 47638 988259
rect 47690 988247 47696 988259
rect 186928 988247 186934 988259
rect 47690 988219 186934 988247
rect 47690 988207 47696 988219
rect 186928 988207 186934 988219
rect 186986 988207 186992 988259
rect 44752 988133 44758 988185
rect 44810 988173 44816 988185
rect 251824 988173 251830 988185
rect 44810 988145 251830 988173
rect 44810 988133 44816 988145
rect 251824 988133 251830 988145
rect 251882 988133 251888 988185
rect 44848 988059 44854 988111
rect 44906 988099 44912 988111
rect 316720 988099 316726 988111
rect 44906 988071 316726 988099
rect 44906 988059 44912 988071
rect 316720 988059 316726 988071
rect 316778 988059 316784 988111
rect 44944 987985 44950 988037
rect 45002 988025 45008 988037
rect 381616 988025 381622 988037
rect 45002 987997 381622 988025
rect 45002 987985 45008 987997
rect 381616 987985 381622 987997
rect 381674 987985 381680 988037
rect 45040 987911 45046 987963
rect 45098 987951 45104 987963
rect 446512 987951 446518 987963
rect 45098 987923 446518 987951
rect 45098 987911 45104 987923
rect 446512 987911 446518 987923
rect 446570 987911 446576 987963
rect 43120 987837 43126 987889
rect 43178 987877 43184 987889
rect 511408 987877 511414 987889
rect 43178 987849 511414 987877
rect 43178 987837 43184 987849
rect 511408 987837 511414 987849
rect 511466 987837 511472 987889
rect 65104 986727 65110 986779
rect 65162 986767 65168 986779
rect 93520 986767 93526 986779
rect 65162 986739 93526 986767
rect 65162 986727 65168 986739
rect 93520 986727 93526 986739
rect 93578 986727 93584 986779
rect 47536 986653 47542 986705
rect 47594 986693 47600 986705
rect 109168 986693 109174 986705
rect 47594 986665 109174 986693
rect 47594 986653 47600 986665
rect 109168 986653 109174 986665
rect 109226 986653 109232 986705
rect 619792 986653 619798 986705
rect 619850 986693 619856 986705
rect 650224 986693 650230 986705
rect 619850 986665 650230 986693
rect 619850 986653 619856 986665
rect 650224 986653 650230 986665
rect 650282 986653 650288 986705
rect 47440 986579 47446 986631
rect 47498 986619 47504 986631
rect 107536 986619 107542 986631
rect 47498 986591 107542 986619
rect 47498 986579 47504 986591
rect 107536 986579 107542 986591
rect 107594 986579 107600 986631
rect 609040 986579 609046 986631
rect 609098 986619 609104 986631
rect 650128 986619 650134 986631
rect 609098 986591 650134 986619
rect 609098 986579 609104 986591
rect 650128 986579 650134 986591
rect 650186 986579 650192 986631
rect 44560 986505 44566 986557
rect 44618 986545 44624 986557
rect 107920 986545 107926 986557
rect 44618 986517 107926 986545
rect 44618 986505 44624 986517
rect 107920 986505 107926 986517
rect 107978 986505 107984 986557
rect 564496 986505 564502 986557
rect 564554 986545 564560 986557
rect 658000 986545 658006 986557
rect 564554 986517 658006 986545
rect 564554 986505 564560 986517
rect 658000 986505 658006 986517
rect 658058 986505 658064 986557
rect 65200 986431 65206 986483
rect 65258 986471 65264 986483
rect 145360 986471 145366 986483
rect 65258 986443 145366 986471
rect 65258 986431 65264 986443
rect 145360 986431 145366 986443
rect 145418 986431 145424 986483
rect 565840 986431 565846 986483
rect 565898 986471 565904 986483
rect 658096 986471 658102 986483
rect 565898 986443 658102 986471
rect 565898 986431 565904 986443
rect 658096 986431 658102 986443
rect 658154 986431 658160 986483
rect 65008 986357 65014 986409
rect 65066 986397 65072 986409
rect 197200 986397 197206 986409
rect 65066 986369 197206 986397
rect 65066 986357 65072 986369
rect 197200 986357 197206 986369
rect 197258 986357 197264 986409
rect 267856 986357 267862 986409
rect 267914 986397 267920 986409
rect 290896 986397 290902 986409
rect 267914 986369 290902 986397
rect 267914 986357 267920 986369
rect 290896 986357 290902 986369
rect 290954 986357 290960 986409
rect 564592 986357 564598 986409
rect 564650 986397 564656 986409
rect 660880 986397 660886 986409
rect 564650 986369 660886 986397
rect 564650 986357 564656 986369
rect 660880 986357 660886 986369
rect 660938 986357 660944 986409
rect 225520 984951 225526 985003
rect 225578 984991 225584 985003
rect 233200 984991 233206 985003
rect 225578 984963 233206 984991
rect 225578 984951 225584 984963
rect 233200 984951 233206 984963
rect 233258 984951 233264 985003
rect 632368 983693 632374 983745
rect 632426 983733 632432 983745
rect 674512 983733 674518 983745
rect 632426 983705 674518 983733
rect 632426 983693 632432 983705
rect 674512 983693 674518 983705
rect 674570 983693 674576 983745
rect 633040 983619 633046 983671
rect 633098 983659 633104 983671
rect 674320 983659 674326 983671
rect 633098 983631 674326 983659
rect 633098 983619 633104 983631
rect 674320 983619 674326 983631
rect 674378 983619 674384 983671
rect 64720 983545 64726 983597
rect 64778 983585 64784 983597
rect 225520 983585 225526 983597
rect 64778 983557 225526 983585
rect 64778 983545 64784 983557
rect 225520 983545 225526 983557
rect 225578 983545 225584 983597
rect 515824 983545 515830 983597
rect 515882 983585 515888 983597
rect 649552 983585 649558 983597
rect 515882 983557 649558 983585
rect 515882 983545 515888 983557
rect 649552 983545 649558 983557
rect 649610 983545 649616 983597
rect 64912 983471 64918 983523
rect 64970 983511 64976 983523
rect 267856 983511 267862 983523
rect 64970 983483 267862 983511
rect 64970 983471 64976 983483
rect 267856 983471 267862 983483
rect 267914 983471 267920 983523
rect 426256 983471 426262 983523
rect 426314 983511 426320 983523
rect 649456 983511 649462 983523
rect 426314 983483 649462 983511
rect 426314 983471 426320 983483
rect 649456 983471 649462 983483
rect 649514 983471 649520 983523
rect 53680 973481 53686 973533
rect 53738 973521 53744 973533
rect 59440 973521 59446 973533
rect 53738 973493 59446 973521
rect 53738 973481 53744 973493
rect 59440 973481 59446 973493
rect 59498 973481 59504 973533
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 43120 967305 43126 967317
rect 42218 967277 43126 967305
rect 42218 967265 42224 967277
rect 43120 967265 43126 967277
rect 43178 967265 43184 967317
rect 42160 960901 42166 960953
rect 42218 960941 42224 960953
rect 42832 960941 42838 960953
rect 42218 960913 42838 960941
rect 42218 960901 42224 960913
rect 42832 960901 42838 960913
rect 42890 960901 42896 960953
rect 42736 959051 42742 959103
rect 42794 959091 42800 959103
rect 59536 959091 59542 959103
rect 42794 959063 59542 959091
rect 42794 959051 42800 959063
rect 59536 959051 59542 959063
rect 59594 959051 59600 959103
rect 675088 958385 675094 958437
rect 675146 958425 675152 958437
rect 675376 958425 675382 958437
rect 675146 958397 675382 958425
rect 675146 958385 675152 958397
rect 675376 958385 675382 958397
rect 675434 958385 675440 958437
rect 675184 956979 675190 957031
rect 675242 957019 675248 957031
rect 675472 957019 675478 957031
rect 675242 956991 675478 957019
rect 675242 956979 675248 956991
rect 675472 956979 675478 956991
rect 675530 956979 675536 957031
rect 669520 954685 669526 954737
rect 669578 954725 669584 954737
rect 675376 954725 675382 954737
rect 669578 954697 675382 954725
rect 669578 954685 669584 954697
rect 675376 954685 675382 954697
rect 675434 954685 675440 954737
rect 674128 953871 674134 953923
rect 674186 953911 674192 953923
rect 675472 953911 675478 953923
rect 674186 953883 675478 953911
rect 674186 953871 674192 953883
rect 675472 953871 675478 953883
rect 675530 953871 675536 953923
rect 42160 953205 42166 953257
rect 42218 953245 42224 953257
rect 42448 953245 42454 953257
rect 42218 953217 42454 953245
rect 42218 953205 42224 953217
rect 42448 953205 42454 953217
rect 42506 953205 42512 953257
rect 674032 952021 674038 952073
rect 674090 952061 674096 952073
rect 675472 952061 675478 952073
rect 674090 952033 675478 952061
rect 674090 952021 674096 952033
rect 675472 952021 675478 952033
rect 675530 952021 675536 952073
rect 42640 944621 42646 944673
rect 42698 944661 42704 944673
rect 59536 944661 59542 944673
rect 42698 944633 59542 944661
rect 42698 944621 42704 944633
rect 59536 944621 59542 944633
rect 59594 944621 59600 944673
rect 42640 944251 42646 944303
rect 42698 944291 42704 944303
rect 48880 944291 48886 944303
rect 42698 944263 48886 944291
rect 42698 944251 42704 944263
rect 48880 944251 48886 944263
rect 48938 944251 48944 944303
rect 42640 942697 42646 942749
rect 42698 942737 42704 942749
rect 47536 942737 47542 942749
rect 42698 942709 47542 942737
rect 42698 942697 42704 942709
rect 47536 942697 47542 942709
rect 47594 942697 47600 942749
rect 39952 942179 39958 942231
rect 40010 942219 40016 942231
rect 42640 942219 42646 942231
rect 40010 942191 42646 942219
rect 40010 942179 40016 942191
rect 42640 942179 42646 942191
rect 42698 942219 42704 942231
rect 44560 942219 44566 942231
rect 42698 942191 44566 942219
rect 42698 942179 42704 942191
rect 44560 942179 44566 942191
rect 44618 942179 44624 942231
rect 658096 939515 658102 939567
rect 658154 939555 658160 939567
rect 674416 939555 674422 939567
rect 658154 939527 674422 939555
rect 658154 939515 658160 939527
rect 674416 939515 674422 939527
rect 674474 939515 674480 939567
rect 655312 939367 655318 939419
rect 655370 939407 655376 939419
rect 674608 939407 674614 939419
rect 655370 939379 674614 939407
rect 655370 939367 655376 939379
rect 674608 939367 674614 939379
rect 674666 939367 674672 939419
rect 655216 939219 655222 939271
rect 655274 939259 655280 939271
rect 676816 939259 676822 939271
rect 655274 939231 676822 939259
rect 655274 939219 655280 939231
rect 676816 939219 676822 939231
rect 676874 939219 676880 939271
rect 655120 939071 655126 939123
rect 655178 939111 655184 939123
rect 676912 939111 676918 939123
rect 655178 939083 676918 939111
rect 655178 939071 655184 939083
rect 676912 939071 676918 939083
rect 676970 939071 676976 939123
rect 660880 937961 660886 938013
rect 660938 938001 660944 938013
rect 674416 938001 674422 938013
rect 660938 937973 674422 938001
rect 660938 937961 660944 937973
rect 674416 937961 674422 937973
rect 674474 937961 674480 938013
rect 658000 936111 658006 936163
rect 658058 936151 658064 936163
rect 676816 936151 676822 936163
rect 658058 936123 676822 936151
rect 658058 936111 658064 936123
rect 676816 936111 676822 936123
rect 676874 936111 676880 936163
rect 39952 933077 39958 933129
rect 40010 933117 40016 933129
rect 40144 933117 40150 933129
rect 40010 933089 40150 933117
rect 40010 933077 40016 933089
rect 40144 933077 40150 933089
rect 40202 933077 40208 933129
rect 42640 932115 42646 932167
rect 42698 932155 42704 932167
rect 53200 932155 53206 932167
rect 42698 932127 53206 932155
rect 42698 932115 42704 932127
rect 53200 932115 53206 932127
rect 53258 932115 53264 932167
rect 48880 930487 48886 930539
rect 48938 930527 48944 930539
rect 59536 930527 59542 930539
rect 48938 930499 59542 930527
rect 48938 930487 48944 930499
rect 59536 930487 59542 930499
rect 59594 930487 59600 930539
rect 654448 927453 654454 927505
rect 654506 927493 654512 927505
rect 666736 927493 666742 927505
rect 654506 927465 666742 927493
rect 654506 927453 654512 927465
rect 666736 927453 666742 927465
rect 666794 927453 666800 927505
rect 649648 927379 649654 927431
rect 649706 927419 649712 927431
rect 677008 927419 677014 927431
rect 649706 927391 677014 927419
rect 649706 927379 649712 927391
rect 677008 927379 677014 927391
rect 677066 927379 677072 927431
rect 47440 915835 47446 915887
rect 47498 915875 47504 915887
rect 59536 915875 59542 915887
rect 47498 915847 59542 915875
rect 47498 915835 47504 915847
rect 59536 915835 59542 915847
rect 59594 915835 59600 915887
rect 653968 915835 653974 915887
rect 654026 915875 654032 915887
rect 660976 915875 660982 915887
rect 654026 915847 660982 915875
rect 654026 915835 654032 915847
rect 660976 915835 660982 915847
rect 661034 915835 661040 915887
rect 39856 907177 39862 907229
rect 39914 907217 39920 907229
rect 40240 907217 40246 907229
rect 39914 907189 40246 907217
rect 39914 907177 39920 907189
rect 40240 907177 40246 907189
rect 40298 907177 40304 907229
rect 654448 904365 654454 904417
rect 654506 904405 654512 904417
rect 663952 904405 663958 904417
rect 654506 904377 663958 904405
rect 654506 904365 654512 904377
rect 663952 904365 663958 904377
rect 664010 904365 664016 904417
rect 53296 901479 53302 901531
rect 53354 901519 53360 901531
rect 59536 901519 59542 901531
rect 53354 901491 59542 901519
rect 53354 901479 53360 901491
rect 59536 901479 59542 901491
rect 59594 901479 59600 901531
rect 40240 892861 40246 892873
rect 40066 892833 40246 892861
rect 40066 892799 40094 892833
rect 40240 892821 40246 892833
rect 40298 892821 40304 892873
rect 40048 892747 40054 892799
rect 40106 892747 40112 892799
rect 50512 887123 50518 887175
rect 50570 887163 50576 887175
rect 59536 887163 59542 887175
rect 50570 887135 59542 887163
rect 50570 887123 50576 887135
rect 59536 887123 59542 887135
rect 59594 887123 59600 887175
rect 40048 886975 40054 887027
rect 40106 887015 40112 887027
rect 40144 887015 40150 887027
rect 40106 886987 40150 887015
rect 40106 886975 40112 886987
rect 40144 886975 40150 886987
rect 40202 886975 40208 887027
rect 653968 881277 653974 881329
rect 654026 881317 654032 881329
rect 660880 881317 660886 881329
rect 654026 881289 660886 881317
rect 654026 881277 654032 881289
rect 660880 881277 660886 881289
rect 660938 881277 660944 881329
rect 40144 872693 40150 872745
rect 40202 872693 40208 872745
rect 40162 872523 40190 872693
rect 41680 872619 41686 872671
rect 41738 872659 41744 872671
rect 59536 872659 59542 872671
rect 41738 872631 59542 872659
rect 41738 872619 41744 872631
rect 59536 872619 59542 872631
rect 59594 872619 59600 872671
rect 40144 872471 40150 872523
rect 40202 872471 40208 872523
rect 674608 872101 674614 872153
rect 674666 872141 674672 872153
rect 675472 872141 675478 872153
rect 674666 872113 675478 872141
rect 674666 872101 674672 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 675088 871435 675094 871487
rect 675146 871475 675152 871487
rect 675376 871475 675382 871487
rect 675146 871447 675382 871475
rect 675146 871435 675152 871447
rect 675376 871435 675382 871447
rect 675434 871435 675440 871487
rect 654448 869807 654454 869859
rect 654506 869847 654512 869859
rect 663760 869847 663766 869859
rect 654506 869819 663766 869847
rect 654506 869807 654512 869819
rect 663760 869807 663766 869819
rect 663818 869807 663824 869859
rect 674416 868993 674422 869045
rect 674474 869033 674480 869045
rect 675184 869033 675190 869045
rect 674474 869005 675190 869033
rect 674474 868993 674480 869005
rect 675184 868993 675190 869005
rect 675242 868993 675248 869045
rect 673360 866921 673366 866973
rect 673418 866961 673424 866973
rect 675184 866961 675190 866973
rect 673418 866933 675190 866961
rect 673418 866921 673424 866933
rect 675184 866921 675190 866933
rect 675242 866921 675248 866973
rect 674512 866477 674518 866529
rect 674570 866517 674576 866529
rect 675376 866517 675382 866529
rect 674570 866489 675382 866517
rect 674570 866477 674576 866489
rect 675376 866477 675382 866489
rect 675434 866477 675440 866529
rect 674320 864997 674326 865049
rect 674378 865037 674384 865049
rect 675088 865037 675094 865049
rect 674378 865009 675094 865037
rect 674378 864997 674384 865009
rect 675088 864997 675094 865009
rect 675146 864997 675152 865049
rect 666640 864035 666646 864087
rect 666698 864075 666704 864087
rect 675184 864075 675190 864087
rect 666698 864047 675190 864075
rect 666698 864035 666704 864047
rect 675184 864035 675190 864047
rect 675242 864035 675248 864087
rect 39856 863961 39862 864013
rect 39914 864001 39920 864013
rect 40144 864001 40150 864013
rect 39914 863973 40150 864001
rect 39914 863961 39920 863973
rect 40144 863961 40150 863973
rect 40202 863961 40208 864013
rect 674416 862037 674422 862089
rect 674474 862077 674480 862089
rect 674896 862077 674902 862089
rect 674474 862049 674902 862077
rect 674474 862037 674480 862049
rect 674896 862037 674902 862049
rect 674954 862037 674960 862089
rect 674992 861075 674998 861127
rect 675050 861115 675056 861127
rect 675184 861115 675190 861127
rect 675050 861087 675190 861115
rect 675050 861075 675056 861087
rect 675184 861075 675190 861087
rect 675242 861075 675248 861127
rect 50320 858263 50326 858315
rect 50378 858303 50384 858315
rect 58576 858303 58582 858315
rect 50378 858275 58582 858303
rect 50378 858263 50384 858275
rect 58576 858263 58582 858275
rect 58634 858263 58640 858315
rect 654160 858263 654166 858315
rect 654218 858303 654224 858315
rect 661072 858303 661078 858315
rect 654218 858275 661078 858303
rect 654218 858263 654224 858275
rect 661072 858263 661078 858275
rect 661130 858263 661136 858315
rect 39856 843833 39862 843885
rect 39914 843873 39920 843885
rect 40048 843873 40054 843885
rect 39914 843845 40054 843873
rect 39914 843833 39920 843845
rect 40048 843833 40054 843845
rect 40106 843833 40112 843885
rect 53392 843833 53398 843885
rect 53450 843873 53456 843885
rect 59536 843873 59542 843885
rect 53450 843845 59542 843873
rect 53450 843833 53456 843845
rect 59536 843833 59542 843845
rect 59594 843833 59600 843885
rect 653968 835175 653974 835227
rect 654026 835215 654032 835227
rect 666832 835215 666838 835227
rect 654026 835187 666838 835215
rect 654026 835175 654032 835187
rect 666832 835175 666838 835187
rect 666890 835175 666896 835227
rect 40048 832511 40054 832563
rect 40106 832551 40112 832563
rect 40106 832523 40286 832551
rect 40106 832511 40112 832523
rect 40258 832267 40286 832523
rect 40240 832215 40246 832267
rect 40298 832215 40304 832267
rect 50608 829477 50614 829529
rect 50666 829517 50672 829529
rect 59536 829517 59542 829529
rect 50666 829489 59542 829517
rect 50666 829477 50672 829489
rect 59536 829477 59542 829489
rect 59594 829477 59600 829529
rect 653968 823705 653974 823757
rect 654026 823745 654032 823757
rect 669808 823745 669814 823757
rect 654026 823717 669814 823745
rect 654026 823705 654032 823717
rect 669808 823705 669814 823717
rect 669866 823705 669872 823757
rect 42640 819117 42646 819169
rect 42698 819157 42704 819169
rect 50512 819157 50518 819169
rect 42698 819129 50518 819157
rect 42698 819117 42704 819129
rect 50512 819117 50518 819129
rect 50570 819117 50576 819169
rect 42640 818081 42646 818133
rect 42698 818121 42704 818133
rect 53296 818121 53302 818133
rect 42698 818093 53302 818121
rect 42698 818081 42704 818093
rect 53296 818081 53302 818093
rect 53354 818081 53360 818133
rect 47536 815047 47542 815099
rect 47594 815087 47600 815099
rect 59536 815087 59542 815099
rect 47594 815059 59542 815087
rect 47594 815047 47600 815059
rect 59536 815047 59542 815059
rect 59594 815047 59600 815099
rect 37360 814973 37366 815025
rect 37418 815013 37424 815025
rect 40240 815013 40246 815025
rect 37418 814985 40246 815013
rect 37418 814973 37424 814985
rect 40240 814973 40246 814985
rect 40298 814973 40304 815025
rect 654448 812161 654454 812213
rect 654506 812201 654512 812213
rect 664048 812201 664054 812213
rect 654506 812173 664054 812201
rect 654506 812161 654512 812173
rect 664048 812161 664054 812173
rect 664106 812161 664112 812213
rect 41968 802393 41974 802445
rect 42026 802433 42032 802445
rect 42928 802433 42934 802445
rect 42026 802405 42934 802433
rect 42026 802393 42032 802405
rect 42928 802393 42934 802405
rect 42986 802393 42992 802445
rect 41776 802171 41782 802223
rect 41834 802211 41840 802223
rect 41968 802211 41974 802223
rect 41834 802183 41974 802211
rect 41834 802171 41840 802183
rect 41968 802171 41974 802183
rect 42026 802171 42032 802223
rect 42736 800839 42742 800891
rect 42794 800879 42800 800891
rect 43408 800879 43414 800891
rect 42794 800851 43414 800879
rect 42794 800839 42800 800851
rect 43408 800839 43414 800851
rect 43466 800839 43472 800891
rect 44656 800617 44662 800669
rect 44714 800657 44720 800669
rect 59536 800657 59542 800669
rect 44714 800629 59542 800657
rect 44714 800617 44720 800629
rect 59536 800617 59542 800629
rect 59594 800617 59600 800669
rect 674992 800617 674998 800669
rect 675050 800657 675056 800669
rect 675184 800657 675190 800669
rect 675050 800629 675190 800657
rect 675050 800617 675056 800629
rect 675184 800617 675190 800629
rect 675242 800617 675248 800669
rect 41872 800287 41878 800299
rect 41698 800259 41878 800287
rect 41698 799991 41726 800259
rect 41872 800247 41878 800259
rect 41930 800247 41936 800299
rect 42160 800247 42166 800299
rect 42218 800287 42224 800299
rect 43504 800287 43510 800299
rect 42218 800259 43510 800287
rect 42218 800247 42224 800259
rect 43504 800247 43510 800259
rect 43562 800247 43568 800299
rect 41776 800173 41782 800225
rect 41834 800213 41840 800225
rect 43312 800213 43318 800225
rect 41834 800185 43318 800213
rect 41834 800173 41840 800185
rect 43312 800173 43318 800185
rect 43370 800173 43376 800225
rect 41872 799991 41878 800003
rect 41698 799963 41878 799991
rect 41872 799951 41878 799963
rect 41930 799951 41936 800003
rect 42160 798101 42166 798153
rect 42218 798141 42224 798153
rect 42640 798141 42646 798153
rect 42218 798113 42646 798141
rect 42218 798101 42224 798113
rect 42640 798101 42646 798113
rect 42698 798101 42704 798153
rect 42544 797583 42550 797635
rect 42602 797623 42608 797635
rect 43408 797623 43414 797635
rect 42602 797595 43414 797623
rect 42602 797583 42608 797595
rect 43408 797583 43414 797595
rect 43466 797583 43472 797635
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 45040 797327 45046 797339
rect 42122 797299 45046 797327
rect 42122 797287 42128 797299
rect 45040 797287 45046 797299
rect 45098 797287 45104 797339
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 43024 796291 43030 796303
rect 42218 796263 43030 796291
rect 42218 796251 42224 796263
rect 43024 796251 43030 796263
rect 43082 796251 43088 796303
rect 43024 796103 43030 796155
rect 43082 796143 43088 796155
rect 43312 796143 43318 796155
rect 43082 796115 43318 796143
rect 43082 796103 43088 796115
rect 43312 796103 43318 796115
rect 43370 796103 43376 796155
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 42832 795033 42838 795045
rect 42218 795005 42838 795033
rect 42218 794993 42224 795005
rect 42832 794993 42838 795005
rect 42890 794993 42896 795045
rect 42064 794253 42070 794305
rect 42122 794293 42128 794305
rect 42448 794293 42454 794305
rect 42122 794265 42454 794293
rect 42122 794253 42128 794265
rect 42448 794253 42454 794265
rect 42506 794253 42512 794305
rect 42160 793809 42166 793861
rect 42218 793849 42224 793861
rect 43120 793849 43126 793861
rect 42218 793821 43126 793849
rect 42218 793809 42224 793821
rect 43120 793809 43126 793821
rect 43178 793809 43184 793861
rect 43120 793661 43126 793713
rect 43178 793701 43184 793713
rect 43504 793701 43510 793713
rect 43178 793673 43510 793701
rect 43178 793661 43184 793673
rect 43504 793661 43510 793673
rect 43562 793661 43568 793713
rect 42160 793143 42166 793195
rect 42218 793183 42224 793195
rect 42928 793183 42934 793195
rect 42218 793155 42934 793183
rect 42218 793143 42224 793155
rect 42928 793143 42934 793155
rect 42986 793143 42992 793195
rect 42544 792921 42550 792973
rect 42602 792961 42608 792973
rect 43024 792961 43030 792973
rect 42602 792933 43030 792961
rect 42602 792921 42608 792933
rect 43024 792921 43030 792933
rect 43082 792921 43088 792973
rect 42160 790479 42166 790531
rect 42218 790519 42224 790531
rect 42544 790519 42550 790531
rect 42218 790491 42550 790519
rect 42218 790479 42224 790491
rect 42544 790479 42550 790491
rect 42602 790479 42608 790531
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 43120 789927 43126 789939
rect 42218 789899 43126 789927
rect 42218 789887 42224 789899
rect 43120 789887 43126 789899
rect 43178 789887 43184 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42544 789483 42550 789495
rect 42218 789455 42550 789483
rect 42218 789443 42224 789455
rect 42544 789443 42550 789455
rect 42602 789443 42608 789495
rect 42160 788703 42166 788755
rect 42218 788743 42224 788755
rect 42832 788743 42838 788755
rect 42218 788715 42838 788743
rect 42218 788703 42224 788715
rect 42832 788703 42838 788715
rect 42890 788703 42896 788755
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 43024 787041 43030 787053
rect 42218 787013 43030 787041
rect 42218 787001 42224 787013
rect 43024 787001 43030 787013
rect 43082 787001 43088 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42352 786449 42358 786461
rect 42218 786421 42358 786449
rect 42218 786409 42224 786421
rect 42352 786409 42358 786421
rect 42410 786409 42416 786461
rect 45040 786261 45046 786313
rect 45098 786301 45104 786313
rect 59536 786301 59542 786313
rect 45098 786273 59542 786301
rect 45098 786261 45104 786273
rect 59536 786261 59542 786273
rect 59594 786261 59600 786313
rect 654064 786261 654070 786313
rect 654122 786301 654128 786313
rect 669712 786301 669718 786313
rect 654122 786273 669718 786301
rect 654122 786261 654128 786273
rect 669712 786261 669718 786273
rect 669770 786261 669776 786313
rect 42064 785595 42070 785647
rect 42122 785635 42128 785647
rect 42448 785635 42454 785647
rect 42122 785607 42454 785635
rect 42122 785595 42128 785607
rect 42448 785595 42454 785607
rect 42506 785595 42512 785647
rect 672496 783449 672502 783501
rect 672554 783489 672560 783501
rect 675376 783489 675382 783501
rect 672554 783461 675382 783489
rect 672554 783449 672560 783461
rect 675376 783449 675382 783461
rect 675434 783449 675440 783501
rect 672976 783079 672982 783131
rect 673034 783119 673040 783131
rect 675088 783119 675094 783131
rect 673034 783091 675094 783119
rect 673034 783079 673040 783091
rect 675088 783079 675094 783091
rect 675146 783119 675152 783131
rect 675472 783119 675478 783131
rect 675146 783091 675478 783119
rect 675146 783079 675152 783091
rect 675472 783079 675478 783091
rect 675530 783079 675536 783131
rect 673264 782931 673270 782983
rect 673322 782971 673328 782983
rect 675376 782971 675382 782983
rect 673322 782943 675382 782971
rect 673322 782931 673328 782943
rect 675376 782931 675382 782943
rect 675434 782931 675440 782983
rect 674992 782487 674998 782539
rect 675050 782527 675056 782539
rect 675472 782527 675478 782539
rect 675050 782499 675478 782527
rect 675050 782487 675056 782499
rect 675472 782487 675478 782499
rect 675530 782487 675536 782539
rect 663856 780489 663862 780541
rect 663914 780529 663920 780541
rect 675088 780529 675094 780541
rect 663914 780501 675094 780529
rect 663914 780489 663920 780501
rect 675088 780489 675094 780501
rect 675146 780489 675152 780541
rect 673072 779749 673078 779801
rect 673130 779789 673136 779801
rect 675376 779789 675382 779801
rect 673130 779761 675382 779789
rect 673130 779749 673136 779761
rect 675376 779749 675382 779761
rect 675434 779749 675440 779801
rect 672880 779305 672886 779357
rect 672938 779345 672944 779357
rect 675472 779345 675478 779357
rect 672938 779317 675478 779345
rect 672938 779305 672944 779317
rect 675472 779305 675478 779317
rect 675530 779305 675536 779357
rect 673168 778565 673174 778617
rect 673226 778605 673232 778617
rect 675376 778605 675382 778617
rect 673226 778577 675382 778605
rect 673226 778565 673232 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 672592 777603 672598 777655
rect 672650 777643 672656 777655
rect 675472 777643 675478 777655
rect 672650 777615 675478 777643
rect 672650 777603 672656 777615
rect 675472 777603 675478 777615
rect 675530 777603 675536 777655
rect 675088 777011 675094 777063
rect 675146 777051 675152 777063
rect 675376 777051 675382 777063
rect 675146 777023 675382 777051
rect 675146 777011 675152 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 42448 776049 42454 776101
rect 42506 776089 42512 776101
rect 50608 776089 50614 776101
rect 42506 776061 50614 776089
rect 42506 776049 42512 776061
rect 50608 776049 50614 776061
rect 50666 776049 50672 776101
rect 674416 775457 674422 775509
rect 674474 775497 674480 775509
rect 675376 775497 675382 775509
rect 674474 775469 675382 775497
rect 674474 775457 674480 775469
rect 675376 775457 675382 775469
rect 675434 775457 675440 775509
rect 42832 775309 42838 775361
rect 42890 775349 42896 775361
rect 47536 775349 47542 775361
rect 42890 775321 47542 775349
rect 42890 775309 42896 775321
rect 47536 775309 47542 775321
rect 47594 775309 47600 775361
rect 42832 774791 42838 774843
rect 42890 774831 42896 774843
rect 53392 774831 53398 774843
rect 42890 774803 53398 774831
rect 42890 774791 42896 774803
rect 53392 774791 53398 774803
rect 53450 774791 53456 774843
rect 654064 774717 654070 774769
rect 654122 774757 654128 774769
rect 672400 774757 672406 774769
rect 654122 774729 672406 774757
rect 654122 774717 654128 774729
rect 672400 774717 672406 774729
rect 672458 774717 672464 774769
rect 674128 773607 674134 773659
rect 674186 773647 674192 773659
rect 675472 773647 675478 773659
rect 674186 773619 675478 773647
rect 674186 773607 674192 773619
rect 675472 773607 675478 773619
rect 675530 773607 675536 773659
rect 53392 771831 53398 771883
rect 53450 771871 53456 771883
rect 59536 771871 59542 771883
rect 53450 771843 59542 771871
rect 53450 771831 53456 771843
rect 59536 771831 59542 771843
rect 59594 771831 59600 771883
rect 653968 763247 653974 763299
rect 654026 763287 654032 763299
rect 661168 763287 661174 763299
rect 654026 763259 661174 763287
rect 654026 763247 654032 763259
rect 661168 763247 661174 763259
rect 661226 763247 661232 763299
rect 660976 762877 660982 762929
rect 661034 762917 661040 762929
rect 674320 762917 674326 762929
rect 661034 762889 674326 762917
rect 661034 762877 661040 762889
rect 674320 762877 674326 762889
rect 674378 762877 674384 762929
rect 666736 762285 666742 762337
rect 666794 762325 666800 762337
rect 674320 762325 674326 762337
rect 666794 762297 674326 762325
rect 666794 762285 666800 762297
rect 674320 762285 674326 762297
rect 674378 762285 674384 762337
rect 663952 761989 663958 762041
rect 664010 762029 664016 762041
rect 674608 762029 674614 762041
rect 664010 762001 674614 762029
rect 664010 761989 664016 762001
rect 674608 761989 674614 762001
rect 674666 761989 674672 762041
rect 672304 760435 672310 760487
rect 672362 760475 672368 760487
rect 673840 760475 673846 760487
rect 672362 760447 673846 760475
rect 672362 760435 672368 760447
rect 673840 760435 673846 760447
rect 673898 760435 673904 760487
rect 42928 757549 42934 757601
rect 42986 757589 42992 757601
rect 43600 757589 43606 757601
rect 42986 757561 43606 757589
rect 42986 757549 42992 757561
rect 43600 757549 43606 757561
rect 43658 757549 43664 757601
rect 44944 757515 44950 757527
rect 42946 757487 44950 757515
rect 42946 757453 42974 757487
rect 44944 757475 44950 757487
rect 45002 757475 45008 757527
rect 53584 757475 53590 757527
rect 53642 757515 53648 757527
rect 59536 757515 59542 757527
rect 53642 757487 59542 757515
rect 53642 757475 53648 757487
rect 59536 757475 59542 757487
rect 59594 757475 59600 757527
rect 42928 757401 42934 757453
rect 42986 757401 42992 757453
rect 41680 757253 41686 757305
rect 41738 757293 41744 757305
rect 43504 757293 43510 757305
rect 41738 757265 43510 757293
rect 41738 757253 41744 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 41776 757031 41782 757083
rect 41834 757071 41840 757083
rect 43312 757071 43318 757083
rect 41834 757043 43318 757071
rect 41834 757031 41840 757043
rect 43312 757031 43318 757043
rect 43370 757031 43376 757083
rect 42160 756735 42166 756787
rect 42218 756775 42224 756787
rect 42352 756775 42358 756787
rect 42218 756747 42358 756775
rect 42218 756735 42224 756747
rect 42352 756735 42358 756747
rect 42410 756735 42416 756787
rect 42928 754219 42934 754271
rect 42986 754219 42992 754271
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 42946 754111 42974 754219
rect 42218 754083 42974 754111
rect 42218 754071 42224 754083
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 43120 753075 43126 753087
rect 42122 753047 43126 753075
rect 42122 753035 42128 753047
rect 43120 753035 43126 753047
rect 43178 753035 43184 753087
rect 42832 751629 42838 751681
rect 42890 751669 42896 751681
rect 43504 751669 43510 751681
rect 42890 751641 43510 751669
rect 42890 751629 42896 751641
rect 43504 751629 43510 751641
rect 43562 751629 43568 751681
rect 42064 749779 42070 749831
rect 42122 749819 42128 749831
rect 42832 749819 42838 749831
rect 42122 749791 42838 749819
rect 42122 749779 42128 749791
rect 42832 749779 42838 749791
rect 42890 749779 42896 749831
rect 649744 748817 649750 748869
rect 649802 748857 649808 748869
rect 677008 748857 677014 748869
rect 649802 748829 677014 748857
rect 649802 748817 649808 748829
rect 677008 748817 677014 748829
rect 677066 748817 677072 748869
rect 42160 747263 42166 747315
rect 42218 747303 42224 747315
rect 43120 747303 43126 747315
rect 42218 747275 43126 747303
rect 42218 747263 42224 747275
rect 43120 747263 43126 747275
rect 43178 747263 43184 747315
rect 42160 746893 42166 746945
rect 42218 746933 42224 746945
rect 43600 746933 43606 746945
rect 42218 746905 43606 746933
rect 42218 746893 42224 746905
rect 43600 746893 43606 746905
rect 43658 746893 43664 746945
rect 42064 746227 42070 746279
rect 42122 746267 42128 746279
rect 42736 746267 42742 746279
rect 42122 746239 42742 746267
rect 42122 746227 42128 746239
rect 42736 746227 42742 746239
rect 42794 746227 42800 746279
rect 672976 745931 672982 745983
rect 673034 745971 673040 745983
rect 675088 745971 675094 745983
rect 673034 745943 675094 745971
rect 673034 745931 673040 745943
rect 675088 745931 675094 745943
rect 675146 745931 675152 745983
rect 42160 745487 42166 745539
rect 42218 745527 42224 745539
rect 43024 745527 43030 745539
rect 42218 745499 43030 745527
rect 42218 745487 42224 745499
rect 43024 745487 43030 745499
rect 43082 745487 43088 745539
rect 674128 745413 674134 745465
rect 674186 745453 674192 745465
rect 674512 745453 674518 745465
rect 674186 745425 674518 745453
rect 674186 745413 674192 745425
rect 674512 745413 674518 745425
rect 674570 745413 674576 745465
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 42832 743825 42838 743837
rect 42218 743797 42838 743825
rect 42218 743785 42224 743797
rect 42832 743785 42838 743797
rect 42890 743785 42896 743837
rect 42064 743193 42070 743245
rect 42122 743233 42128 743245
rect 42736 743233 42742 743245
rect 42122 743205 42742 743233
rect 42122 743193 42128 743205
rect 42736 743193 42742 743205
rect 42794 743193 42800 743245
rect 53488 743045 53494 743097
rect 53546 743085 53552 743097
rect 59536 743085 59542 743097
rect 53546 743057 59542 743085
rect 53546 743045 53552 743057
rect 59536 743045 59542 743057
rect 59594 743045 59600 743097
rect 42160 742379 42166 742431
rect 42218 742419 42224 742431
rect 43120 742419 43126 742431
rect 42218 742391 43126 742419
rect 42218 742379 42224 742391
rect 43120 742379 43126 742391
rect 43178 742379 43184 742431
rect 653968 740159 653974 740211
rect 654026 740199 654032 740211
rect 663952 740199 663958 740211
rect 654026 740171 663958 740199
rect 654026 740159 654032 740171
rect 663952 740159 663958 740171
rect 664010 740159 664016 740211
rect 672784 738087 672790 738139
rect 672842 738127 672848 738139
rect 675088 738127 675094 738139
rect 672842 738099 675094 738127
rect 672842 738087 672848 738099
rect 675088 738087 675094 738099
rect 675146 738127 675152 738139
rect 675472 738127 675478 738139
rect 675146 738099 675478 738127
rect 675146 738087 675152 738099
rect 675472 738087 675478 738099
rect 675530 738087 675536 738139
rect 672688 737865 672694 737917
rect 672746 737905 672752 737917
rect 675376 737905 675382 737917
rect 672746 737877 675382 737905
rect 672746 737865 672752 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 675184 737643 675190 737695
rect 675242 737683 675248 737695
rect 675376 737683 675382 737695
rect 675242 737655 675382 737683
rect 675242 737643 675248 737655
rect 675376 737643 675382 737655
rect 675434 737643 675440 737695
rect 660976 737273 660982 737325
rect 661034 737313 661040 737325
rect 675088 737313 675094 737325
rect 661034 737285 675094 737313
rect 661034 737273 661040 737285
rect 675088 737273 675094 737285
rect 675146 737273 675152 737325
rect 674224 735423 674230 735475
rect 674282 735463 674288 735475
rect 675472 735463 675478 735475
rect 674282 735435 675478 735463
rect 674282 735423 674288 735435
rect 675472 735423 675478 735435
rect 675530 735423 675536 735475
rect 673360 734905 673366 734957
rect 673418 734945 673424 734957
rect 675376 734945 675382 734957
rect 673418 734917 675382 734945
rect 673418 734905 673424 734917
rect 675376 734905 675382 734917
rect 675434 734905 675440 734957
rect 672976 733573 672982 733625
rect 673034 733613 673040 733625
rect 675472 733613 675478 733625
rect 673034 733585 675478 733613
rect 673034 733573 673040 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 42736 732685 42742 732737
rect 42794 732725 42800 732737
rect 53392 732725 53398 732737
rect 42794 732697 53398 732725
rect 42794 732685 42800 732697
rect 53392 732685 53398 732697
rect 53450 732685 53456 732737
rect 674896 732315 674902 732367
rect 674954 732355 674960 732367
rect 675472 732355 675478 732367
rect 674954 732327 675478 732355
rect 674954 732315 674960 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 42736 732093 42742 732145
rect 42794 732133 42800 732145
rect 53584 732133 53590 732145
rect 42794 732105 53590 732133
rect 42794 732093 42800 732105
rect 53584 732093 53590 732105
rect 53642 732093 53648 732145
rect 675088 732019 675094 732071
rect 675146 732059 675152 732071
rect 675376 732059 675382 732071
rect 675146 732031 675382 732059
rect 675146 732019 675152 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 42352 731797 42358 731849
rect 42410 731837 42416 731849
rect 45040 731837 45046 731849
rect 42410 731809 45046 731837
rect 42410 731797 42416 731809
rect 45040 731797 45046 731809
rect 45098 731797 45104 731849
rect 674608 730465 674614 730517
rect 674666 730505 674672 730517
rect 675472 730505 675478 730517
rect 674666 730477 675478 730505
rect 674666 730465 674672 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 674224 728911 674230 728963
rect 674282 728911 674288 728963
rect 674242 728741 674270 728911
rect 674224 728689 674230 728741
rect 674282 728689 674288 728741
rect 47536 728615 47542 728667
rect 47594 728655 47600 728667
rect 59536 728655 59542 728667
rect 47594 728627 59542 728655
rect 47594 728615 47600 728627
rect 59536 728615 59542 728627
rect 59594 728615 59600 728667
rect 674320 728615 674326 728667
rect 674378 728655 674384 728667
rect 675472 728655 675478 728667
rect 674378 728627 675478 728655
rect 674378 728615 674384 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 674992 725729 674998 725781
rect 675050 725769 675056 725781
rect 675376 725769 675382 725781
rect 675050 725741 675382 725769
rect 675050 725729 675056 725741
rect 675376 725729 675382 725741
rect 675434 725729 675440 725781
rect 42736 720623 42742 720675
rect 42794 720623 42800 720675
rect 42754 720453 42782 720623
rect 42736 720401 42742 720453
rect 42794 720401 42800 720453
rect 663760 717885 663766 717937
rect 663818 717925 663824 717937
rect 674416 717925 674422 717937
rect 663818 717897 674422 717925
rect 663818 717885 663824 717897
rect 674416 717885 674422 717897
rect 674474 717885 674480 717937
rect 660880 717293 660886 717345
rect 660938 717333 660944 717345
rect 674416 717333 674422 717345
rect 660938 717305 674422 717333
rect 660938 717293 660944 717305
rect 674416 717293 674422 717305
rect 674474 717293 674480 717345
rect 654256 717145 654262 717197
rect 654314 717185 654320 717197
rect 666928 717185 666934 717197
rect 654314 717157 666934 717185
rect 654314 717145 654320 717157
rect 666928 717145 666934 717157
rect 666986 717145 666992 717197
rect 43120 717071 43126 717123
rect 43178 717111 43184 717123
rect 44848 717111 44854 717123
rect 43178 717083 44854 717111
rect 43178 717071 43184 717083
rect 44848 717071 44854 717083
rect 44906 717071 44912 717123
rect 661072 716849 661078 716901
rect 661130 716889 661136 716901
rect 674416 716889 674422 716901
rect 661130 716861 674422 716889
rect 661130 716849 661136 716861
rect 674416 716849 674422 716861
rect 674474 716849 674480 716901
rect 672304 716257 672310 716309
rect 672362 716297 672368 716309
rect 674416 716297 674422 716309
rect 672362 716269 674422 716297
rect 672362 716257 672368 716269
rect 674416 716257 674422 716269
rect 674474 716257 674480 716309
rect 41680 714290 41732 714296
rect 44944 714259 44950 714311
rect 45002 714299 45008 714311
rect 59536 714299 59542 714311
rect 45002 714271 59542 714299
rect 45002 714259 45008 714271
rect 59536 714259 59542 714271
rect 59594 714259 59600 714311
rect 41680 714232 41732 714238
rect 41692 714077 41720 714232
rect 43504 714077 43510 714089
rect 41692 714049 43510 714077
rect 43504 714037 43510 714049
rect 43562 714037 43568 714089
rect 41776 713963 41782 714015
rect 41834 714003 41840 714015
rect 43408 714003 43414 714015
rect 41834 713975 43414 714003
rect 41834 713963 41840 713975
rect 43408 713963 43414 713975
rect 43466 713963 43472 714015
rect 42064 713519 42070 713571
rect 42122 713559 42128 713571
rect 42352 713559 42358 713571
rect 42122 713531 42358 713559
rect 42122 713519 42128 713531
rect 42352 713519 42358 713531
rect 42410 713519 42416 713571
rect 43408 711709 43414 711721
rect 43042 711681 43414 711709
rect 43042 711573 43070 711681
rect 43408 711669 43414 711681
rect 43466 711669 43472 711721
rect 43024 711521 43030 711573
rect 43082 711521 43088 711573
rect 43024 711003 43030 711055
rect 43082 711043 43088 711055
rect 43216 711043 43222 711055
rect 43082 711015 43222 711043
rect 43082 711003 43088 711015
rect 43216 711003 43222 711015
rect 43274 711003 43280 711055
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 43408 710895 43414 710907
rect 42218 710867 43414 710895
rect 42218 710855 42224 710867
rect 43408 710855 43414 710867
rect 43466 710855 43472 710907
rect 672496 709745 672502 709797
rect 672554 709785 672560 709797
rect 674416 709785 674422 709797
rect 672554 709757 674422 709785
rect 672554 709745 672560 709757
rect 674416 709745 674422 709757
rect 674474 709745 674480 709797
rect 672592 709153 672598 709205
rect 672650 709193 672656 709205
rect 674416 709193 674422 709205
rect 672650 709165 674422 709193
rect 672650 709153 672656 709165
rect 674416 709153 674422 709165
rect 674474 709153 674480 709205
rect 672880 708635 672886 708687
rect 672938 708675 672944 708687
rect 674416 708675 674422 708687
rect 672938 708647 674422 708675
rect 672938 708635 672944 708647
rect 674416 708635 674422 708647
rect 674474 708635 674480 708687
rect 42064 708561 42070 708613
rect 42122 708601 42128 708613
rect 43120 708601 43126 708613
rect 42122 708573 43126 708601
rect 42122 708561 42128 708573
rect 43120 708561 43126 708573
rect 43178 708561 43184 708613
rect 42160 708043 42166 708095
rect 42218 708083 42224 708095
rect 42448 708083 42454 708095
rect 42218 708055 42454 708083
rect 42218 708043 42224 708055
rect 42448 708043 42454 708055
rect 42506 708043 42512 708095
rect 42160 706563 42166 706615
rect 42218 706603 42224 706615
rect 43120 706603 43126 706615
rect 42218 706575 43126 706603
rect 42218 706563 42224 706575
rect 43120 706563 43126 706575
rect 43178 706563 43184 706615
rect 675184 705601 675190 705653
rect 675242 705641 675248 705653
rect 675376 705641 675382 705653
rect 675242 705613 675382 705641
rect 675242 705601 675248 705613
rect 675376 705601 675382 705613
rect 675434 705601 675440 705653
rect 43024 704269 43030 704321
rect 43082 704269 43088 704321
rect 43042 704235 43070 704269
rect 42274 704207 43070 704235
rect 42160 704047 42166 704099
rect 42218 704087 42224 704099
rect 42274 704087 42302 704207
rect 43024 704121 43030 704173
rect 43082 704161 43088 704173
rect 43504 704161 43510 704173
rect 43082 704133 43510 704161
rect 43082 704121 43088 704133
rect 43504 704121 43510 704133
rect 43562 704121 43568 704173
rect 42218 704059 42302 704087
rect 42218 704047 42224 704059
rect 42064 703529 42070 703581
rect 42122 703569 42128 703581
rect 42448 703569 42454 703581
rect 42122 703541 42454 703569
rect 42122 703529 42128 703541
rect 42448 703529 42454 703541
rect 42506 703529 42512 703581
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 43120 702903 43126 702915
rect 42218 702875 43126 702903
rect 42218 702863 42224 702875
rect 43120 702863 43126 702875
rect 43178 702863 43184 702915
rect 649840 702715 649846 702767
rect 649898 702755 649904 702767
rect 677008 702755 677014 702767
rect 649898 702727 677014 702755
rect 649898 702715 649904 702727
rect 677008 702715 677014 702727
rect 677066 702715 677072 702767
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 43024 702311 43030 702323
rect 42218 702283 43030 702311
rect 42218 702271 42224 702283
rect 43024 702271 43030 702283
rect 43082 702271 43088 702323
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42448 700091 42454 700103
rect 42218 700063 42454 700091
rect 42218 700051 42224 700063
rect 42448 700051 42454 700063
rect 42506 700051 42512 700103
rect 43120 699829 43126 699881
rect 43178 699869 43184 699881
rect 59536 699869 59542 699881
rect 43178 699841 59542 699869
rect 43178 699829 43184 699841
rect 59536 699829 59542 699841
rect 59594 699829 59600 699881
rect 672784 699829 672790 699881
rect 672842 699869 672848 699881
rect 673168 699869 673174 699881
rect 672842 699841 673174 699869
rect 672842 699829 672848 699841
rect 673168 699829 673174 699841
rect 673226 699829 673232 699881
rect 42160 699385 42166 699437
rect 42218 699425 42224 699437
rect 42352 699425 42358 699437
rect 42218 699397 42358 699425
rect 42218 699385 42224 699397
rect 42352 699385 42358 699397
rect 42410 699385 42416 699437
rect 654448 694057 654454 694109
rect 654506 694097 654512 694109
rect 672496 694097 672502 694109
rect 654506 694069 672502 694097
rect 654506 694057 654512 694069
rect 672496 694057 672502 694069
rect 672554 694057 672560 694109
rect 675088 693465 675094 693517
rect 675146 693505 675152 693517
rect 675472 693505 675478 693517
rect 675146 693477 675478 693505
rect 675146 693465 675152 693477
rect 675472 693465 675478 693477
rect 675530 693465 675536 693517
rect 673168 692947 673174 692999
rect 673226 692987 673232 692999
rect 675472 692987 675478 692999
rect 673226 692959 675478 692987
rect 673226 692947 673232 692959
rect 675472 692947 675478 692959
rect 675530 692947 675536 692999
rect 672784 692873 672790 692925
rect 672842 692913 672848 692925
rect 675376 692913 675382 692925
rect 672842 692885 675382 692913
rect 672842 692873 672848 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 675184 692651 675190 692703
rect 675242 692691 675248 692703
rect 675376 692691 675382 692703
rect 675242 692663 675382 692691
rect 675242 692651 675248 692663
rect 675376 692651 675382 692663
rect 675434 692651 675440 692703
rect 674992 690653 674998 690705
rect 675050 690693 675056 690705
rect 675472 690693 675478 690705
rect 675050 690665 675478 690693
rect 675050 690653 675056 690665
rect 675472 690653 675478 690665
rect 675530 690653 675536 690705
rect 673264 689765 673270 689817
rect 673322 689805 673328 689817
rect 675376 689805 675382 689817
rect 673322 689777 675382 689805
rect 673322 689765 673328 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 43216 689469 43222 689521
rect 43274 689509 43280 689521
rect 44944 689509 44950 689521
rect 43274 689481 44950 689509
rect 43274 689469 43280 689481
rect 44944 689469 44950 689481
rect 45002 689469 45008 689521
rect 673072 688581 673078 688633
rect 673130 688621 673136 688633
rect 675472 688621 675478 688633
rect 673130 688593 675478 688621
rect 673130 688581 673136 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 42832 688433 42838 688485
rect 42890 688473 42896 688485
rect 47536 688473 47542 688485
rect 42890 688445 47542 688473
rect 42890 688433 42896 688445
rect 47536 688433 47542 688445
rect 47594 688433 47600 688485
rect 675088 687323 675094 687375
rect 675146 687363 675152 687375
rect 675472 687363 675478 687375
rect 675146 687335 675478 687363
rect 675146 687323 675152 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 669616 686213 669622 686265
rect 669674 686253 669680 686265
rect 675376 686253 675382 686265
rect 669674 686225 675382 686253
rect 669674 686213 669680 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 47536 685473 47542 685525
rect 47594 685513 47600 685525
rect 59536 685513 59542 685525
rect 47594 685485 59542 685513
rect 47594 685473 47600 685485
rect 59536 685473 59542 685485
rect 59594 685473 59600 685525
rect 674320 685473 674326 685525
rect 674378 685513 674384 685525
rect 675472 685513 675478 685525
rect 674378 685485 675478 685513
rect 674378 685473 674384 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 674896 684067 674902 684119
rect 674954 684067 674960 684119
rect 674992 684067 674998 684119
rect 675050 684067 675056 684119
rect 674914 683823 674942 684067
rect 675010 683897 675038 684067
rect 674992 683845 674998 683897
rect 675050 683845 675056 683897
rect 674896 683771 674902 683823
rect 674954 683771 674960 683823
rect 675088 683623 675094 683675
rect 675146 683663 675152 683675
rect 675472 683663 675478 683675
rect 675146 683635 675478 683663
rect 675146 683623 675152 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 674992 680959 674998 681011
rect 675050 680999 675056 681011
rect 675184 680999 675190 681011
rect 675050 680971 675190 680999
rect 675050 680959 675056 680971
rect 675184 680959 675190 680971
rect 675242 680959 675248 681011
rect 42160 674003 42166 674055
rect 42218 674043 42224 674055
rect 43024 674043 43030 674055
rect 42218 674015 43030 674043
rect 42218 674003 42224 674015
rect 43024 674003 43030 674015
rect 43082 674003 43088 674055
rect 43408 673855 43414 673907
rect 43466 673895 43472 673907
rect 44752 673895 44758 673907
rect 43466 673867 44758 673895
rect 43466 673855 43472 673867
rect 44752 673855 44758 673867
rect 44810 673855 44816 673907
rect 669808 672671 669814 672723
rect 669866 672711 669872 672723
rect 674416 672711 674422 672723
rect 669866 672683 674422 672711
rect 669866 672671 669872 672683
rect 674416 672671 674422 672683
rect 674474 672671 674480 672723
rect 666832 672153 666838 672205
rect 666890 672193 666896 672205
rect 674416 672193 674422 672205
rect 666890 672165 674422 672193
rect 666890 672153 666896 672165
rect 674416 672153 674422 672165
rect 674474 672153 674480 672205
rect 41872 672079 41878 672131
rect 41930 672119 41936 672131
rect 42640 672119 42646 672131
rect 41930 672091 42646 672119
rect 41930 672079 41936 672091
rect 42640 672079 42646 672091
rect 42698 672079 42704 672131
rect 664048 671561 664054 671613
rect 664106 671601 664112 671613
rect 674416 671601 674422 671613
rect 664106 671573 674422 671601
rect 664106 671561 664112 671573
rect 674416 671561 674422 671573
rect 674474 671561 674480 671613
rect 44848 671043 44854 671095
rect 44906 671083 44912 671095
rect 59536 671083 59542 671095
rect 44906 671055 59542 671083
rect 44906 671043 44912 671055
rect 59536 671043 59542 671055
rect 59594 671043 59600 671095
rect 654448 671043 654454 671095
rect 654506 671083 654512 671095
rect 661072 671083 661078 671095
rect 654506 671055 661078 671083
rect 654506 671043 654512 671055
rect 661072 671043 661078 671055
rect 661130 671043 661136 671095
rect 43216 670895 43222 670947
rect 43274 670935 43280 670947
rect 43274 670907 43454 670935
rect 43274 670895 43280 670907
rect 43426 670873 43454 670907
rect 43408 670821 43414 670873
rect 43466 670821 43472 670873
rect 42640 670747 42646 670799
rect 42698 670787 42704 670799
rect 42928 670787 42934 670799
rect 42698 670759 42934 670787
rect 42698 670747 42704 670759
rect 42928 670747 42934 670759
rect 42986 670747 42992 670799
rect 41968 670673 41974 670725
rect 42026 670713 42032 670725
rect 43120 670713 43126 670725
rect 42026 670685 43126 670713
rect 42026 670673 42032 670685
rect 43120 670673 43126 670685
rect 43178 670673 43184 670725
rect 41776 670599 41782 670651
rect 41834 670639 41840 670651
rect 42640 670639 42646 670651
rect 41834 670611 42646 670639
rect 41834 670599 41840 670611
rect 42640 670599 42646 670611
rect 42698 670599 42704 670651
rect 42160 670303 42166 670355
rect 42218 670343 42224 670355
rect 42352 670343 42358 670355
rect 42218 670315 42358 670343
rect 42218 670303 42224 670315
rect 42352 670303 42358 670315
rect 42410 670303 42416 670355
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 42928 668567 42934 668579
rect 42218 668539 42934 668567
rect 42218 668527 42224 668539
rect 42928 668527 42934 668539
rect 42986 668527 42992 668579
rect 42928 668379 42934 668431
rect 42986 668419 42992 668431
rect 43216 668419 43222 668431
rect 42986 668391 43222 668419
rect 42986 668379 42992 668391
rect 43216 668379 43222 668391
rect 43274 668379 43280 668431
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43504 667901 43510 667913
rect 42218 667873 43510 667901
rect 42218 667861 42224 667873
rect 43504 667861 43510 667873
rect 43562 667861 43568 667913
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 42928 666717 42934 666729
rect 42218 666689 42934 666717
rect 42218 666677 42224 666689
rect 42928 666677 42934 666689
rect 42986 666677 42992 666729
rect 42928 665197 42934 665249
rect 42986 665237 42992 665249
rect 43408 665237 43414 665249
rect 42986 665209 43414 665237
rect 42986 665197 42992 665209
rect 43408 665197 43414 665209
rect 43466 665197 43472 665249
rect 672688 665197 672694 665249
rect 672746 665237 672752 665249
rect 673840 665237 673846 665249
rect 672746 665209 673846 665237
rect 672746 665197 672752 665209
rect 673840 665197 673846 665209
rect 673898 665197 673904 665249
rect 42064 664161 42070 664213
rect 42122 664201 42128 664213
rect 42640 664201 42646 664213
rect 42122 664173 42646 664201
rect 42122 664161 42128 664173
rect 42640 664161 42646 664173
rect 42698 664161 42704 664213
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 43024 663387 43030 663399
rect 42218 663359 43030 663387
rect 42218 663347 42224 663359
rect 43024 663347 43030 663359
rect 43082 663347 43088 663399
rect 672976 662311 672982 662363
rect 673034 662351 673040 662363
rect 673840 662351 673846 662363
rect 673034 662323 673846 662351
rect 673034 662311 673040 662323
rect 673840 662311 673846 662323
rect 673898 662311 673904 662363
rect 42064 661053 42070 661105
rect 42122 661093 42128 661105
rect 43120 661093 43126 661105
rect 42122 661065 43126 661093
rect 42122 661053 42128 661065
rect 43120 661053 43126 661065
rect 43178 661053 43184 661105
rect 674416 660979 674422 661031
rect 674474 661019 674480 661031
rect 675088 661019 675094 661031
rect 674474 660991 675094 661019
rect 674474 660979 674480 660991
rect 675088 660979 675094 660991
rect 675146 660979 675152 661031
rect 42064 660387 42070 660439
rect 42122 660427 42128 660439
rect 42928 660427 42934 660439
rect 42122 660399 42934 660427
rect 42122 660387 42128 660399
rect 42928 660387 42934 660399
rect 42986 660387 42992 660439
rect 42160 659647 42166 659699
rect 42218 659687 42224 659699
rect 42640 659687 42646 659699
rect 42218 659659 42646 659687
rect 42218 659647 42224 659659
rect 42640 659647 42646 659659
rect 42698 659647 42704 659699
rect 42640 659499 42646 659551
rect 42698 659539 42704 659551
rect 43696 659539 43702 659551
rect 42698 659511 43702 659539
rect 42698 659499 42704 659511
rect 43696 659499 43702 659511
rect 43754 659499 43760 659551
rect 649936 659499 649942 659551
rect 649994 659539 650000 659551
rect 674896 659539 674902 659551
rect 649994 659511 674902 659539
rect 649994 659499 650000 659511
rect 674896 659499 674902 659511
rect 674954 659499 674960 659551
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 42640 659095 42646 659107
rect 42122 659067 42646 659095
rect 42122 659055 42128 659067
rect 42640 659055 42646 659067
rect 42698 659055 42704 659107
rect 42064 657353 42070 657405
rect 42122 657393 42128 657405
rect 42352 657393 42358 657405
rect 42122 657365 42358 657393
rect 42122 657353 42128 657365
rect 42352 657353 42358 657365
rect 42410 657353 42416 657405
rect 42928 656687 42934 656739
rect 42986 656727 42992 656739
rect 59536 656727 59542 656739
rect 42986 656699 59542 656727
rect 42986 656687 42992 656699
rect 59536 656687 59542 656699
rect 59594 656687 59600 656739
rect 42160 656613 42166 656665
rect 42218 656653 42224 656665
rect 43024 656653 43030 656665
rect 42218 656625 43030 656653
rect 42218 656613 42224 656625
rect 43024 656613 43030 656625
rect 43082 656613 43088 656665
rect 42160 656169 42166 656221
rect 42218 656209 42224 656221
rect 43120 656209 43126 656221
rect 42218 656181 43126 656209
rect 42218 656169 42224 656181
rect 43120 656169 43126 656181
rect 43178 656169 43184 656221
rect 674608 655207 674614 655259
rect 674666 655247 674672 655259
rect 675184 655247 675190 655259
rect 674666 655219 675190 655247
rect 674666 655207 674672 655219
rect 675184 655207 675190 655219
rect 675242 655207 675248 655259
rect 673168 653727 673174 653779
rect 673226 653767 673232 653779
rect 675184 653767 675190 653779
rect 673226 653739 675190 653767
rect 673226 653727 673232 653739
rect 675184 653727 675190 653739
rect 675242 653727 675248 653779
rect 671728 648251 671734 648303
rect 671786 648291 671792 648303
rect 675376 648291 675382 648303
rect 671786 648263 675382 648291
rect 671786 648251 671792 648263
rect 675376 648251 675382 648263
rect 675434 648251 675440 648303
rect 654256 648029 654262 648081
rect 654314 648069 654320 648081
rect 664048 648069 664054 648081
rect 654314 648041 664054 648069
rect 654314 648029 654320 648041
rect 664048 648029 664054 648041
rect 664106 648029 664112 648081
rect 672304 648029 672310 648081
rect 672362 648069 672368 648081
rect 675376 648069 675382 648081
rect 672362 648041 675382 648069
rect 672362 648029 672368 648041
rect 675376 648029 675382 648041
rect 675434 648029 675440 648081
rect 43216 647733 43222 647785
rect 43274 647773 43280 647785
rect 44848 647773 44854 647785
rect 43274 647745 44854 647773
rect 43274 647733 43280 647745
rect 44848 647733 44854 647745
rect 44906 647733 44912 647785
rect 674512 647067 674518 647119
rect 674570 647107 674576 647119
rect 675184 647107 675190 647119
rect 674570 647079 675190 647107
rect 674570 647067 674576 647079
rect 675184 647067 675190 647079
rect 675242 647107 675248 647119
rect 675376 647107 675382 647119
rect 675242 647079 675382 647107
rect 675242 647067 675248 647079
rect 675376 647067 675382 647079
rect 675434 647067 675440 647119
rect 674224 646401 674230 646453
rect 674282 646441 674288 646453
rect 675088 646441 675094 646453
rect 674282 646413 675094 646441
rect 674282 646401 674288 646413
rect 675088 646401 675094 646413
rect 675146 646441 675152 646453
rect 675376 646441 675382 646453
rect 675146 646413 675382 646441
rect 675146 646401 675152 646413
rect 675376 646401 675382 646413
rect 675434 646401 675440 646453
rect 674608 645217 674614 645269
rect 674666 645257 674672 645269
rect 674896 645257 674902 645269
rect 674666 645229 674902 645257
rect 674666 645217 674672 645229
rect 674896 645217 674902 645229
rect 674954 645217 674960 645269
rect 666736 645143 666742 645195
rect 666794 645183 666800 645195
rect 675088 645183 675094 645195
rect 666794 645155 675094 645183
rect 666794 645143 666800 645155
rect 675088 645143 675094 645155
rect 675146 645143 675152 645195
rect 42352 645069 42358 645121
rect 42410 645109 42416 645121
rect 59536 645109 59542 645121
rect 42410 645081 59542 645109
rect 42410 645069 42416 645081
rect 59536 645069 59542 645081
rect 59594 645069 59600 645121
rect 672208 644551 672214 644603
rect 672266 644591 672272 644603
rect 675472 644591 675478 644603
rect 672266 644563 675478 644591
rect 672266 644551 672272 644563
rect 675472 644551 675478 644563
rect 675530 644551 675536 644603
rect 672592 644033 672598 644085
rect 672650 644073 672656 644085
rect 675472 644073 675478 644085
rect 672650 644045 675478 644073
rect 672650 644033 672656 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 672880 643367 672886 643419
rect 672938 643407 672944 643419
rect 675376 643407 675382 643419
rect 672938 643379 675382 643407
rect 672938 643367 672944 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 673360 642257 673366 642309
rect 673418 642297 673424 642309
rect 675472 642297 675478 642309
rect 673418 642269 675478 642297
rect 673418 642257 673424 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 675088 641813 675094 641865
rect 675146 641853 675152 641865
rect 675376 641853 675382 641865
rect 675146 641825 675382 641853
rect 675146 641813 675152 641825
rect 675376 641813 675382 641825
rect 675434 641813 675440 641865
rect 41776 631749 41782 631801
rect 41834 631789 41840 631801
rect 42640 631789 42646 631801
rect 41834 631761 42646 631789
rect 41834 631749 41840 631761
rect 42640 631749 42646 631761
rect 42698 631749 42704 631801
rect 42640 628271 42646 628323
rect 42698 628271 42704 628323
rect 42658 628027 42686 628271
rect 42640 627975 42646 628027
rect 42698 627975 42704 628027
rect 42448 627901 42454 627953
rect 42506 627941 42512 627953
rect 47632 627941 47638 627953
rect 42506 627913 47638 627941
rect 42506 627901 42512 627913
rect 47632 627901 47638 627913
rect 47690 627901 47696 627953
rect 44752 627827 44758 627879
rect 44810 627867 44816 627879
rect 59536 627867 59542 627879
rect 44810 627839 59542 627867
rect 44810 627827 44816 627839
rect 59536 627827 59542 627839
rect 59594 627827 59600 627879
rect 41008 627753 41014 627805
rect 41066 627793 41072 627805
rect 43408 627793 43414 627805
rect 41066 627765 43414 627793
rect 41066 627753 41072 627765
rect 43408 627753 43414 627765
rect 43466 627753 43472 627805
rect 672400 627753 672406 627805
rect 672458 627793 672464 627805
rect 673840 627793 673846 627805
rect 672458 627765 673846 627793
rect 672458 627753 672464 627765
rect 673840 627753 673846 627765
rect 673898 627753 673904 627805
rect 41584 627679 41590 627731
rect 41642 627719 41648 627731
rect 43120 627719 43126 627731
rect 41642 627691 43126 627719
rect 41642 627679 41648 627691
rect 43120 627679 43126 627691
rect 43178 627679 43184 627731
rect 41872 627383 41878 627435
rect 41930 627383 41936 627435
rect 41890 627213 41918 627383
rect 669712 627309 669718 627361
rect 669770 627349 669776 627361
rect 674608 627349 674614 627361
rect 669770 627321 674614 627349
rect 669770 627309 669776 627321
rect 674608 627309 674614 627321
rect 674666 627309 674672 627361
rect 41872 627161 41878 627213
rect 41930 627161 41936 627213
rect 661168 626865 661174 626917
rect 661226 626905 661232 626917
rect 674608 626905 674614 626917
rect 661226 626877 674614 626905
rect 661226 626865 661232 626877
rect 674608 626865 674614 626877
rect 674666 626865 674672 626917
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 42640 625351 42646 625363
rect 42218 625323 42646 625351
rect 42218 625311 42224 625323
rect 42640 625311 42646 625323
rect 42698 625311 42704 625363
rect 670960 625163 670966 625215
rect 671018 625203 671024 625215
rect 674608 625203 674614 625215
rect 671018 625175 674614 625203
rect 671018 625163 671024 625175
rect 674608 625163 674614 625175
rect 674666 625163 674672 625215
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 42448 624685 42454 624697
rect 42218 624657 42454 624685
rect 42218 624645 42224 624657
rect 42448 624645 42454 624657
rect 42506 624645 42512 624697
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 43216 623501 43222 623513
rect 42218 623473 43222 623501
rect 42218 623461 42224 623473
rect 43216 623461 43222 623473
rect 43274 623461 43280 623513
rect 42160 622203 42166 622255
rect 42218 622243 42224 622255
rect 42448 622243 42454 622255
rect 42218 622215 42454 622243
rect 42218 622203 42224 622215
rect 42448 622203 42454 622215
rect 42506 622203 42512 622255
rect 671920 622203 671926 622255
rect 671978 622243 671984 622255
rect 677200 622243 677206 622255
rect 671978 622215 677206 622243
rect 671978 622203 671984 622215
rect 677200 622203 677206 622215
rect 677258 622203 677264 622255
rect 654064 622129 654070 622181
rect 654122 622169 654128 622181
rect 672688 622169 672694 622181
rect 654122 622141 672694 622169
rect 654122 622129 654128 622141
rect 672688 622129 672694 622141
rect 672746 622129 672752 622181
rect 673744 622055 673750 622107
rect 673802 622095 673808 622107
rect 676816 622095 676822 622107
rect 673802 622067 676822 622095
rect 673802 622055 673808 622067
rect 676816 622055 676822 622067
rect 676874 622055 676880 622107
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 42640 621651 42646 621663
rect 42218 621623 42646 621651
rect 42218 621611 42224 621623
rect 42640 621611 42646 621623
rect 42698 621611 42704 621663
rect 42064 620871 42070 620923
rect 42122 620911 42128 620923
rect 43312 620911 43318 620923
rect 42122 620883 43318 620911
rect 42122 620871 42128 620883
rect 43312 620871 43318 620883
rect 43370 620871 43376 620923
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 43120 620393 43126 620405
rect 42218 620365 43126 620393
rect 42218 620353 42224 620365
rect 43120 620353 43126 620365
rect 43178 620353 43184 620405
rect 672784 619169 672790 619221
rect 672842 619209 672848 619221
rect 673840 619209 673846 619221
rect 672842 619181 673846 619209
rect 672842 619169 672848 619181
rect 673840 619169 673846 619181
rect 673898 619169 673904 619221
rect 42064 617837 42070 617889
rect 42122 617877 42128 617889
rect 42640 617877 42646 617889
rect 42122 617849 42646 617877
rect 42122 617837 42128 617849
rect 42640 617837 42646 617849
rect 42698 617837 42704 617889
rect 42160 617319 42166 617371
rect 42218 617359 42224 617371
rect 42448 617359 42454 617371
rect 42218 617331 42454 617359
rect 42218 617319 42224 617331
rect 42448 617319 42454 617331
rect 42506 617319 42512 617371
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 42352 616693 42358 616705
rect 42218 616665 42358 616693
rect 42218 616653 42224 616665
rect 42352 616653 42358 616665
rect 42410 616653 42416 616705
rect 42160 615839 42166 615891
rect 42218 615879 42224 615891
rect 43120 615879 43126 615891
rect 42218 615851 43126 615879
rect 42218 615839 42224 615851
rect 43120 615839 43126 615851
rect 43178 615839 43184 615891
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 43504 614177 43510 614189
rect 42218 614149 43510 614177
rect 42218 614137 42224 614149
rect 43504 614137 43510 614149
rect 43562 614137 43568 614189
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42352 613659 42358 613671
rect 42218 613631 42358 613659
rect 42218 613619 42224 613631
rect 42352 613619 42358 613631
rect 42410 613619 42416 613671
rect 42352 613471 42358 613523
rect 42410 613511 42416 613523
rect 59536 613511 59542 613523
rect 42410 613483 59542 613511
rect 42410 613471 42416 613483
rect 59536 613471 59542 613483
rect 59594 613471 59600 613523
rect 650032 613471 650038 613523
rect 650090 613511 650096 613523
rect 677104 613511 677110 613523
rect 650090 613483 677110 613511
rect 650090 613471 650096 613483
rect 677104 613471 677110 613483
rect 677162 613471 677168 613523
rect 654352 613397 654358 613449
rect 654410 613437 654416 613449
rect 669520 613437 669526 613449
rect 654410 613409 669526 613437
rect 654410 613397 654416 613409
rect 669520 613397 669526 613409
rect 669578 613397 669584 613449
rect 674224 613397 674230 613449
rect 674282 613437 674288 613449
rect 675184 613437 675190 613449
rect 674282 613409 675190 613437
rect 674282 613397 674288 613409
rect 675184 613397 675190 613409
rect 675242 613397 675248 613449
rect 42064 612953 42070 613005
rect 42122 612993 42128 613005
rect 42448 612993 42454 613005
rect 42122 612965 42454 612993
rect 42122 612953 42128 612965
rect 42448 612953 42454 612965
rect 42506 612953 42512 613005
rect 672112 604073 672118 604125
rect 672170 604113 672176 604125
rect 675472 604113 675478 604125
rect 672170 604085 675478 604113
rect 672170 604073 672176 604085
rect 675472 604073 675478 604085
rect 675530 604073 675536 604125
rect 672016 603259 672022 603311
rect 672074 603299 672080 603311
rect 675376 603299 675382 603311
rect 672074 603271 675382 603299
rect 672074 603259 672080 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 673264 602667 673270 602719
rect 673322 602707 673328 602719
rect 675376 602707 675382 602719
rect 673322 602679 675382 602707
rect 673322 602667 673328 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 672400 602149 672406 602201
rect 672458 602189 672464 602201
rect 675184 602189 675190 602201
rect 672458 602161 675190 602189
rect 672458 602149 672464 602161
rect 675184 602149 675190 602161
rect 675242 602189 675248 602201
rect 675376 602189 675382 602201
rect 675242 602161 675382 602189
rect 675242 602149 675248 602161
rect 675376 602149 675382 602161
rect 675434 602149 675440 602201
rect 673456 602075 673462 602127
rect 673514 602115 673520 602127
rect 674512 602115 674518 602127
rect 673514 602087 674518 602115
rect 673514 602075 673520 602087
rect 674512 602075 674518 602087
rect 674570 602115 674576 602127
rect 675472 602115 675478 602127
rect 674570 602087 675478 602115
rect 674570 602075 674576 602087
rect 675472 602075 675478 602087
rect 675530 602075 675536 602127
rect 43216 601927 43222 601979
rect 43274 601967 43280 601979
rect 46000 601967 46006 601979
rect 43274 601939 46006 601967
rect 43274 601927 43280 601939
rect 46000 601927 46006 601939
rect 46058 601927 46064 601979
rect 663760 601927 663766 601979
rect 663818 601967 663824 601979
rect 675088 601967 675094 601979
rect 663818 601939 675094 601967
rect 663818 601927 663824 601939
rect 675088 601927 675094 601939
rect 675146 601927 675152 601979
rect 42448 601853 42454 601905
rect 42506 601893 42512 601905
rect 59536 601893 59542 601905
rect 42506 601865 59542 601893
rect 42506 601853 42512 601865
rect 59536 601853 59542 601865
rect 59594 601853 59600 601905
rect 673168 601705 673174 601757
rect 673226 601745 673232 601757
rect 673744 601745 673750 601757
rect 673226 601717 673750 601745
rect 673226 601705 673232 601717
rect 673744 601705 673750 601717
rect 673802 601705 673808 601757
rect 674608 600373 674614 600425
rect 674666 600413 674672 600425
rect 675472 600413 675478 600425
rect 674666 600385 675478 600413
rect 674666 600373 674672 600385
rect 675472 600373 675478 600385
rect 675530 600373 675536 600425
rect 673072 599559 673078 599611
rect 673130 599599 673136 599611
rect 675376 599599 675382 599611
rect 673130 599571 675382 599599
rect 673130 599559 673136 599571
rect 675376 599559 675382 599571
rect 675434 599559 675440 599611
rect 654448 599041 654454 599093
rect 654506 599081 654512 599093
rect 669520 599081 669526 599093
rect 654506 599053 669526 599081
rect 654506 599041 654512 599053
rect 669520 599041 669526 599053
rect 669578 599041 669584 599093
rect 671824 599041 671830 599093
rect 671882 599081 671888 599093
rect 675376 599081 675382 599093
rect 671882 599053 675382 599081
rect 671882 599041 671888 599053
rect 675376 599041 675382 599053
rect 675434 599041 675440 599093
rect 672976 598375 672982 598427
rect 673034 598415 673040 598427
rect 675472 598415 675478 598427
rect 673034 598387 675478 598415
rect 673034 598375 673040 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 672784 597117 672790 597169
rect 672842 597157 672848 597169
rect 675472 597157 675478 597169
rect 672842 597129 675478 597157
rect 672842 597117 672848 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 675088 596821 675094 596873
rect 675146 596861 675152 596873
rect 675376 596861 675382 596873
rect 675146 596833 675382 596861
rect 675146 596821 675152 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 675088 590457 675094 590509
rect 675146 590497 675152 590509
rect 675472 590497 675478 590509
rect 675146 590469 675478 590497
rect 675146 590457 675152 590469
rect 675472 590457 675478 590469
rect 675530 590457 675536 590509
rect 673168 590383 673174 590435
rect 673226 590423 673232 590435
rect 673840 590423 673846 590435
rect 673226 590395 673846 590423
rect 673226 590383 673232 590395
rect 673840 590383 673846 590395
rect 673898 590383 673904 590435
rect 671920 588755 671926 588807
rect 671978 588795 671984 588807
rect 676912 588795 676918 588807
rect 671978 588767 676918 588795
rect 671978 588755 671984 588767
rect 676912 588755 676918 588767
rect 676970 588755 676976 588807
rect 654448 587497 654454 587549
rect 654506 587537 654512 587549
rect 666832 587537 666838 587549
rect 654506 587509 666838 587537
rect 654506 587497 654512 587509
rect 666832 587497 666838 587509
rect 666890 587497 666896 587549
rect 673840 587497 673846 587549
rect 673898 587537 673904 587549
rect 676816 587537 676822 587549
rect 673898 587509 676822 587537
rect 673898 587497 673904 587509
rect 676816 587497 676822 587509
rect 676874 587497 676880 587549
rect 46000 584907 46006 584959
rect 46058 584947 46064 584959
rect 58768 584947 58774 584959
rect 46058 584919 58774 584947
rect 46058 584907 46064 584919
rect 58768 584907 58774 584919
rect 58826 584907 58832 584959
rect 43120 584611 43126 584663
rect 43178 584651 43184 584663
rect 43312 584651 43318 584663
rect 43178 584623 43318 584651
rect 43178 584611 43184 584623
rect 43312 584611 43318 584623
rect 43370 584611 43376 584663
rect 43408 584611 43414 584663
rect 43466 584651 43472 584663
rect 43888 584651 43894 584663
rect 43466 584623 43894 584651
rect 43466 584611 43472 584623
rect 43888 584611 43894 584623
rect 43946 584611 43952 584663
rect 41584 584537 41590 584589
rect 41642 584577 41648 584589
rect 43504 584577 43510 584589
rect 41642 584549 43510 584577
rect 41642 584537 41648 584549
rect 43504 584537 43510 584549
rect 43562 584537 43568 584589
rect 41680 584463 41686 584515
rect 41738 584503 41744 584515
rect 43120 584503 43126 584515
rect 41738 584475 43126 584503
rect 41738 584463 41744 584475
rect 43120 584463 43126 584475
rect 43178 584463 43184 584515
rect 42928 584389 42934 584441
rect 42986 584429 42992 584441
rect 43408 584429 43414 584441
rect 42986 584401 43414 584429
rect 42986 584389 42992 584401
rect 43408 584389 43414 584401
rect 43466 584389 43472 584441
rect 43024 584315 43030 584367
rect 43082 584355 43088 584367
rect 43600 584355 43606 584367
rect 43082 584327 43606 584355
rect 43082 584315 43088 584327
rect 43600 584315 43606 584327
rect 43658 584315 43664 584367
rect 41776 584241 41782 584293
rect 41834 584281 41840 584293
rect 42928 584281 42934 584293
rect 41834 584253 42934 584281
rect 41834 584241 41840 584253
rect 42928 584241 42934 584253
rect 42986 584241 42992 584293
rect 41872 584167 41878 584219
rect 41930 584167 41936 584219
rect 42064 584167 42070 584219
rect 42122 584207 42128 584219
rect 43024 584207 43030 584219
rect 42122 584179 43030 584207
rect 42122 584167 42128 584179
rect 43024 584167 43030 584179
rect 43082 584167 43088 584219
rect 41890 583997 41918 584167
rect 42448 584093 42454 584145
rect 42506 584133 42512 584145
rect 50416 584133 50422 584145
rect 42506 584105 50422 584133
rect 42506 584093 42512 584105
rect 50416 584093 50422 584105
rect 50474 584093 50480 584145
rect 41872 583945 41878 583997
rect 41930 583945 41936 583997
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 43312 582135 43318 582147
rect 42218 582107 43318 582135
rect 42218 582095 42224 582107
rect 43312 582095 43318 582107
rect 43370 582095 43376 582147
rect 663952 582021 663958 582073
rect 664010 582061 664016 582073
rect 674416 582061 674422 582073
rect 664010 582033 674422 582061
rect 664010 582021 664016 582033
rect 674416 582021 674422 582033
rect 674474 582021 674480 582073
rect 655216 581947 655222 581999
rect 655274 581987 655280 581999
rect 674608 581987 674614 581999
rect 655274 581959 674614 581987
rect 655274 581947 655280 581959
rect 674608 581947 674614 581959
rect 674666 581947 674672 581999
rect 666928 581577 666934 581629
rect 666986 581617 666992 581629
rect 674608 581617 674614 581629
rect 666986 581589 674614 581617
rect 666986 581577 666992 581589
rect 674608 581577 674614 581589
rect 674666 581577 674672 581629
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 42448 581469 42454 581481
rect 42122 581441 42454 581469
rect 42122 581429 42128 581441
rect 42448 581429 42454 581441
rect 42506 581429 42512 581481
rect 670960 580837 670966 580889
rect 671018 580877 671024 580889
rect 674416 580877 674422 580889
rect 671018 580849 674422 580877
rect 671018 580837 671024 580849
rect 674416 580837 674422 580849
rect 674474 580837 674480 580889
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 43408 580285 43414 580297
rect 42122 580257 43414 580285
rect 42122 580245 42128 580257
rect 43408 580245 43414 580257
rect 43466 580245 43472 580297
rect 671920 580023 671926 580075
rect 671978 580063 671984 580075
rect 674608 580063 674614 580075
rect 671978 580035 674614 580063
rect 671978 580023 671984 580035
rect 674608 580023 674614 580035
rect 674666 580023 674672 580075
rect 42064 578395 42070 578447
rect 42122 578435 42128 578447
rect 43024 578435 43030 578447
rect 42122 578407 43030 578435
rect 42122 578395 42128 578407
rect 43024 578395 43030 578407
rect 43082 578395 43088 578447
rect 43024 578247 43030 578299
rect 43082 578287 43088 578299
rect 43504 578287 43510 578299
rect 43082 578259 43510 578287
rect 43082 578247 43088 578259
rect 43504 578247 43510 578259
rect 43562 578247 43568 578299
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 43600 577695 43606 577707
rect 42218 577667 43606 577695
rect 42218 577655 42224 577667
rect 43600 577655 43606 577667
rect 43658 577655 43664 577707
rect 42064 577137 42070 577189
rect 42122 577177 42128 577189
rect 42928 577177 42934 577189
rect 42122 577149 42934 577177
rect 42122 577137 42128 577149
rect 42928 577137 42934 577149
rect 42986 577137 42992 577189
rect 654448 576027 654454 576079
rect 654506 576067 654512 576079
rect 669712 576067 669718 576079
rect 654506 576039 669718 576067
rect 654506 576027 654512 576039
rect 669712 576027 669718 576039
rect 669770 576027 669776 576079
rect 671728 574473 671734 574525
rect 671786 574513 671792 574525
rect 674608 574513 674614 574525
rect 671786 574485 674614 574513
rect 671786 574473 671792 574485
rect 674608 574473 674614 574485
rect 674666 574473 674672 574525
rect 42160 573955 42166 574007
rect 42218 573995 42224 574007
rect 43120 573995 43126 574007
rect 42218 573967 43126 573995
rect 42218 573955 42224 573967
rect 43120 573955 43126 573967
rect 43178 573955 43184 574007
rect 672592 573437 672598 573489
rect 672650 573477 672656 573489
rect 674608 573477 674614 573489
rect 672650 573449 674614 573477
rect 672650 573437 672656 573449
rect 674608 573437 674614 573449
rect 674666 573437 674672 573489
rect 42064 573215 42070 573267
rect 42122 573255 42128 573267
rect 42448 573255 42454 573267
rect 42122 573227 42454 573255
rect 42122 573215 42128 573227
rect 42448 573215 42454 573227
rect 42506 573215 42512 573267
rect 672208 573067 672214 573119
rect 672266 573107 672272 573119
rect 673744 573107 673750 573119
rect 672266 573079 673750 573107
rect 672266 573067 672272 573079
rect 673744 573067 673750 573079
rect 673802 573067 673808 573119
rect 672304 572845 672310 572897
rect 672362 572885 672368 572897
rect 674608 572885 674614 572897
rect 672362 572857 674614 572885
rect 672362 572845 672368 572857
rect 674608 572845 674614 572857
rect 674666 572845 674672 572897
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 43024 572663 43030 572675
rect 42218 572635 43030 572663
rect 42218 572623 42224 572635
rect 43024 572623 43030 572635
rect 43082 572623 43088 572675
rect 672880 571809 672886 571861
rect 672938 571849 672944 571861
rect 674608 571849 674614 571861
rect 672938 571821 674614 571849
rect 672938 571809 672944 571821
rect 674608 571809 674614 571821
rect 674666 571809 674672 571861
rect 43504 571661 43510 571713
rect 43562 571701 43568 571713
rect 43888 571701 43894 571713
rect 43562 571673 43894 571701
rect 43562 571661 43568 571673
rect 43888 571661 43894 571673
rect 43946 571661 43952 571713
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 42928 571035 42934 571047
rect 42218 571007 42934 571035
rect 42218 570995 42224 571007
rect 42928 570995 42934 571007
rect 42986 570995 42992 571047
rect 42160 570403 42166 570455
rect 42218 570443 42224 570455
rect 42448 570443 42454 570455
rect 42218 570415 42454 570443
rect 42218 570403 42224 570415
rect 42448 570403 42454 570415
rect 42506 570403 42512 570455
rect 42928 570255 42934 570307
rect 42986 570295 42992 570307
rect 59536 570295 59542 570307
rect 42986 570267 59542 570295
rect 42986 570255 42992 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 43024 569703 43030 569715
rect 42122 569675 43030 569703
rect 42122 569663 42128 569675
rect 43024 569663 43030 569675
rect 43082 569663 43088 569715
rect 650128 567369 650134 567421
rect 650186 567409 650192 567421
rect 677008 567409 677014 567421
rect 650186 567381 677014 567409
rect 650186 567369 650192 567381
rect 677008 567369 677014 567381
rect 677066 567369 677072 567421
rect 654448 567295 654454 567347
rect 654506 567335 654512 567347
rect 666640 567335 666646 567347
rect 654506 567307 666646 567335
rect 654506 567295 654512 567307
rect 666640 567295 666646 567307
rect 666698 567295 666704 567347
rect 672400 564261 672406 564313
rect 672458 564301 672464 564313
rect 675088 564301 675094 564313
rect 672458 564273 675094 564301
rect 672458 564261 672464 564273
rect 675088 564261 675094 564273
rect 675146 564261 675152 564313
rect 673456 563891 673462 563943
rect 673514 563931 673520 563943
rect 675184 563931 675190 563943
rect 673514 563903 675190 563931
rect 673514 563891 673520 563903
rect 675184 563891 675190 563903
rect 675242 563891 675248 563943
rect 674608 559377 674614 559429
rect 674666 559417 674672 559429
rect 675376 559417 675382 559429
rect 674666 559389 675382 559417
rect 674666 559377 674672 559389
rect 675376 559377 675382 559389
rect 675434 559377 675440 559429
rect 42448 559007 42454 559059
rect 42506 559047 42512 559059
rect 50224 559047 50230 559059
rect 42506 559019 50230 559047
rect 42506 559007 42512 559019
rect 50224 559007 50230 559019
rect 50282 559007 50288 559059
rect 42544 558859 42550 558911
rect 42602 558899 42608 558911
rect 59536 558899 59542 558911
rect 42602 558871 59542 558899
rect 42602 558859 42608 558871
rect 59536 558859 59542 558871
rect 59594 558859 59600 558911
rect 674896 558045 674902 558097
rect 674954 558085 674960 558097
rect 675376 558085 675382 558097
rect 674954 558057 675382 558085
rect 674954 558045 674960 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 675184 557823 675190 557875
rect 675242 557863 675248 557875
rect 675376 557863 675382 557875
rect 675242 557835 675382 557863
rect 675242 557823 675248 557835
rect 675376 557823 675382 557835
rect 675434 557823 675440 557875
rect 673456 557601 673462 557653
rect 673514 557641 673520 557653
rect 675472 557641 675478 557653
rect 673514 557613 675478 557641
rect 673514 557601 673520 557613
rect 675472 557601 675478 557613
rect 675530 557601 675536 557653
rect 675088 557083 675094 557135
rect 675146 557123 675152 557135
rect 675472 557123 675478 557135
rect 675146 557095 675478 557123
rect 675146 557083 675152 557095
rect 675472 557083 675478 557095
rect 675530 557083 675536 557135
rect 660880 555825 660886 555877
rect 660938 555865 660944 555877
rect 675088 555865 675094 555877
rect 660938 555837 675094 555865
rect 660938 555825 660944 555837
rect 675088 555825 675094 555837
rect 675146 555825 675152 555877
rect 674416 555233 674422 555285
rect 674474 555273 674480 555285
rect 675472 555273 675478 555285
rect 674474 555245 675478 555273
rect 674474 555233 674480 555245
rect 675472 555233 675478 555245
rect 675530 555233 675536 555285
rect 673168 553901 673174 553953
rect 673226 553941 673232 553953
rect 675472 553941 675478 553953
rect 673226 553913 675478 553941
rect 673226 553901 673232 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 673360 553161 673366 553213
rect 673418 553201 673424 553213
rect 675376 553201 675382 553213
rect 673418 553173 675382 553201
rect 673418 553161 673424 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 654448 552939 654454 552991
rect 654506 552979 654512 552991
rect 666640 552979 666646 552991
rect 654506 552951 666646 552979
rect 654506 552939 654512 552951
rect 666640 552939 666646 552951
rect 666698 552939 666704 552991
rect 674320 551903 674326 551955
rect 674378 551943 674384 551955
rect 675472 551943 675478 551955
rect 674378 551915 675478 551943
rect 674378 551903 674384 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 675088 551607 675094 551659
rect 675146 551647 675152 551659
rect 675376 551647 675382 551659
rect 675146 551619 675382 551647
rect 675146 551607 675152 551619
rect 675376 551607 675382 551619
rect 675434 551607 675440 551659
rect 674896 550053 674902 550105
rect 674954 550053 674960 550105
rect 675088 550053 675094 550105
rect 675146 550093 675152 550105
rect 675472 550093 675478 550105
rect 675146 550065 675478 550093
rect 675146 550053 675152 550065
rect 675472 550053 675478 550065
rect 675530 550053 675536 550105
rect 674914 549883 674942 550053
rect 41584 549831 41590 549883
rect 41642 549871 41648 549883
rect 41776 549871 41782 549883
rect 41642 549843 41782 549871
rect 41642 549831 41648 549843
rect 41776 549831 41782 549843
rect 41834 549831 41840 549883
rect 674896 549831 674902 549883
rect 674954 549831 674960 549883
rect 674512 548203 674518 548255
rect 674570 548243 674576 548255
rect 675472 548243 675478 548255
rect 674570 548215 675478 548243
rect 674570 548203 674576 548215
rect 675472 548203 675478 548215
rect 675530 548203 675536 548255
rect 50224 544503 50230 544555
rect 50282 544543 50288 544555
rect 59536 544543 59542 544555
rect 50282 544515 59542 544543
rect 50282 544503 50288 544515
rect 59536 544503 59542 544515
rect 59594 544503 59600 544555
rect 42160 542357 42166 542409
rect 42218 542397 42224 542409
rect 43120 542397 43126 542409
rect 42218 542369 43126 542397
rect 42218 542357 42224 542369
rect 43120 542357 43126 542369
rect 43178 542357 43184 542409
rect 42928 541469 42934 541521
rect 42986 541509 42992 541521
rect 53680 541509 53686 541521
rect 42986 541481 53686 541509
rect 42986 541469 42992 541481
rect 53680 541469 53686 541481
rect 53738 541469 53744 541521
rect 654448 541469 654454 541521
rect 654506 541509 654512 541521
rect 672400 541509 672406 541521
rect 654506 541481 672406 541509
rect 654506 541469 654512 541481
rect 672400 541469 672406 541481
rect 672458 541469 672464 541521
rect 41584 541247 41590 541299
rect 41642 541287 41648 541299
rect 43696 541287 43702 541299
rect 41642 541259 43702 541287
rect 41642 541247 41648 541259
rect 43696 541247 43702 541259
rect 43754 541247 43760 541299
rect 42832 541099 42838 541151
rect 42890 541139 42896 541151
rect 43312 541139 43318 541151
rect 42890 541111 43318 541139
rect 42890 541099 42896 541111
rect 43312 541099 43318 541111
rect 43370 541099 43376 541151
rect 41968 540951 41974 541003
rect 42026 540951 42032 541003
rect 42064 540951 42070 541003
rect 42122 540991 42128 541003
rect 42832 540991 42838 541003
rect 42122 540963 42838 540991
rect 42122 540951 42128 540963
rect 42832 540951 42838 540963
rect 42890 540951 42896 541003
rect 41986 540917 42014 540951
rect 41986 540889 42494 540917
rect 42466 540411 42494 540889
rect 42448 540359 42454 540411
rect 42506 540359 42512 540411
rect 42064 538879 42070 538931
rect 42122 538919 42128 538931
rect 42448 538919 42454 538931
rect 42122 538891 42454 538919
rect 42122 538879 42128 538891
rect 42448 538879 42454 538891
rect 42506 538879 42512 538931
rect 42448 538731 42454 538783
rect 42506 538771 42512 538783
rect 43216 538771 43222 538783
rect 42506 538743 43222 538771
rect 42506 538731 42512 538743
rect 43216 538731 43222 538743
rect 43274 538731 43280 538783
rect 672496 538509 672502 538561
rect 672554 538549 672560 538561
rect 673744 538549 673750 538561
rect 672554 538521 673750 538549
rect 672554 538509 672560 538521
rect 673744 538509 673750 538521
rect 673802 538509 673808 538561
rect 42160 538287 42166 538339
rect 42218 538327 42224 538339
rect 42928 538327 42934 538339
rect 42218 538299 42934 538327
rect 42218 538287 42224 538299
rect 42928 538287 42934 538299
rect 42986 538287 42992 538339
rect 42928 538139 42934 538191
rect 42986 538179 42992 538191
rect 43312 538179 43318 538191
rect 42986 538151 43318 538179
rect 42986 538139 42992 538151
rect 43312 538139 43318 538151
rect 43370 538139 43376 538191
rect 42064 537029 42070 537081
rect 42122 537069 42128 537081
rect 42448 537069 42454 537081
rect 42122 537041 42454 537069
rect 42122 537029 42128 537041
rect 42448 537029 42454 537041
rect 42506 537029 42512 537081
rect 671920 536733 671926 536785
rect 671978 536773 671984 536785
rect 673744 536773 673750 536785
rect 671978 536745 673750 536773
rect 671978 536733 671984 536745
rect 673744 536733 673750 536745
rect 673802 536733 673808 536785
rect 674608 536733 674614 536785
rect 674666 536773 674672 536785
rect 674896 536773 674902 536785
rect 674666 536745 674902 536773
rect 674666 536733 674672 536745
rect 674896 536733 674902 536745
rect 674954 536733 674960 536785
rect 661072 536585 661078 536637
rect 661130 536625 661136 536637
rect 674608 536625 674614 536637
rect 661130 536597 674614 536625
rect 661130 536585 661136 536597
rect 674608 536585 674614 536597
rect 674666 536585 674672 536637
rect 674512 536289 674518 536341
rect 674570 536329 674576 536341
rect 675088 536329 675094 536341
rect 674570 536301 675094 536329
rect 674570 536289 674576 536301
rect 675088 536289 675094 536301
rect 675146 536289 675152 536341
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 43024 535811 43030 535823
rect 42122 535783 43030 535811
rect 42122 535771 42128 535783
rect 43024 535771 43030 535783
rect 43082 535771 43088 535823
rect 655120 535771 655126 535823
rect 655178 535811 655184 535823
rect 676816 535811 676822 535823
rect 655178 535783 676822 535811
rect 655178 535771 655184 535783
rect 676816 535771 676822 535783
rect 676874 535771 676880 535823
rect 42160 535031 42166 535083
rect 42218 535071 42224 535083
rect 43120 535071 43126 535083
rect 42218 535043 43126 535071
rect 42218 535031 42224 535043
rect 43120 535031 43126 535043
rect 43178 535031 43184 535083
rect 43120 534883 43126 534935
rect 43178 534923 43184 534935
rect 43696 534923 43702 534935
rect 43178 534895 43702 534923
rect 43178 534883 43184 534895
rect 43696 534883 43702 534895
rect 43754 534883 43760 534935
rect 42160 534439 42166 534491
rect 42218 534479 42224 534491
rect 42928 534479 42934 534491
rect 42218 534451 42934 534479
rect 42218 534439 42224 534451
rect 42928 534439 42934 534451
rect 42986 534439 42992 534491
rect 42064 533699 42070 533751
rect 42122 533739 42128 533751
rect 43024 533739 43030 533751
rect 42122 533711 43030 533739
rect 42122 533699 42128 533711
rect 43024 533699 43030 533711
rect 43082 533699 43088 533751
rect 42160 531331 42166 531383
rect 42218 531371 42224 531383
rect 42352 531371 42358 531383
rect 42218 531343 42358 531371
rect 42218 531331 42224 531343
rect 42352 531331 42358 531343
rect 42410 531331 42416 531383
rect 42160 530887 42166 530939
rect 42218 530927 42224 530939
rect 42448 530927 42454 530939
rect 42218 530899 42454 530927
rect 42218 530887 42224 530899
rect 42448 530887 42454 530899
rect 42506 530887 42512 530939
rect 42448 530739 42454 530791
rect 42506 530779 42512 530791
rect 42928 530779 42934 530791
rect 42506 530751 42934 530779
rect 42506 530739 42512 530751
rect 42928 530739 42934 530751
rect 42986 530739 42992 530791
rect 42064 530221 42070 530273
rect 42122 530261 42128 530273
rect 42832 530261 42838 530273
rect 42122 530233 42838 530261
rect 42122 530221 42128 530233
rect 42832 530221 42838 530233
rect 42890 530221 42896 530273
rect 42832 529925 42838 529977
rect 42890 529965 42896 529977
rect 59536 529965 59542 529977
rect 42890 529937 59542 529965
rect 42890 529925 42896 529937
rect 59536 529925 59542 529937
rect 59594 529925 59600 529977
rect 654064 529925 654070 529977
rect 654122 529965 654128 529977
rect 672592 529965 672598 529977
rect 654122 529937 672598 529965
rect 654122 529925 654128 529937
rect 672592 529925 672598 529937
rect 672650 529925 672656 529977
rect 672112 529851 672118 529903
rect 672170 529891 672176 529903
rect 673744 529891 673750 529903
rect 672170 529863 673750 529891
rect 672170 529851 672176 529863
rect 673744 529851 673750 529863
rect 673802 529851 673808 529903
rect 674896 529851 674902 529903
rect 674954 529891 674960 529903
rect 675184 529891 675190 529903
rect 674954 529863 675190 529891
rect 674954 529851 674960 529863
rect 675184 529851 675190 529863
rect 675242 529851 675248 529903
rect 672784 529555 672790 529607
rect 672842 529595 672848 529607
rect 673744 529595 673750 529607
rect 672842 529567 673750 529595
rect 672842 529555 672848 529567
rect 673744 529555 673750 529567
rect 673802 529555 673808 529607
rect 672016 529481 672022 529533
rect 672074 529521 672080 529533
rect 674896 529521 674902 529533
rect 672074 529493 674902 529521
rect 672074 529481 672080 529493
rect 674896 529481 674902 529493
rect 674954 529481 674960 529533
rect 42160 529407 42166 529459
rect 42218 529447 42224 529459
rect 43120 529447 43126 529459
rect 42218 529419 43126 529447
rect 42218 529407 42224 529419
rect 43120 529407 43126 529419
rect 43178 529407 43184 529459
rect 671824 528593 671830 528645
rect 671882 528633 671888 528645
rect 673744 528633 673750 528645
rect 671882 528605 673750 528633
rect 671882 528593 671888 528605
rect 673744 528593 673750 528605
rect 673802 528593 673808 528645
rect 42160 527779 42166 527831
rect 42218 527819 42224 527831
rect 42448 527819 42454 527831
rect 42218 527791 42454 527819
rect 42218 527779 42224 527791
rect 42448 527779 42454 527791
rect 42506 527779 42512 527831
rect 42064 527187 42070 527239
rect 42122 527227 42128 527239
rect 42352 527227 42358 527239
rect 42122 527199 42358 527227
rect 42122 527187 42128 527199
rect 42352 527187 42358 527199
rect 42410 527187 42416 527239
rect 42160 526447 42166 526499
rect 42218 526487 42224 526499
rect 42928 526487 42934 526499
rect 42218 526459 42934 526487
rect 42218 526447 42224 526459
rect 42928 526447 42934 526459
rect 42986 526447 42992 526499
rect 650224 524301 650230 524353
rect 650282 524341 650288 524353
rect 677104 524341 677110 524353
rect 650282 524313 677110 524341
rect 650282 524301 650288 524313
rect 677104 524301 677110 524313
rect 677162 524301 677168 524353
rect 42352 524153 42358 524205
rect 42410 524193 42416 524205
rect 42832 524193 42838 524205
rect 42410 524165 42838 524193
rect 42410 524153 42416 524165
rect 42832 524153 42838 524165
rect 42890 524153 42896 524205
rect 654448 519269 654454 519321
rect 654506 519309 654512 519321
rect 663856 519309 663862 519321
rect 654506 519281 663862 519309
rect 654506 519269 654512 519281
rect 663856 519269 663862 519281
rect 663914 519269 663920 519321
rect 50512 515495 50518 515547
rect 50570 515535 50576 515547
rect 59536 515535 59542 515547
rect 50570 515507 59542 515535
rect 50570 515495 50576 515507
rect 59536 515495 59542 515507
rect 59594 515495 59600 515547
rect 674896 514089 674902 514141
rect 674954 514129 674960 514141
rect 675088 514129 675094 514141
rect 674954 514101 675094 514129
rect 674954 514089 674960 514101
rect 675088 514089 675094 514101
rect 675146 514089 675152 514141
rect 654448 506911 654454 506963
rect 654506 506951 654512 506963
rect 663856 506951 663862 506963
rect 654506 506923 663862 506951
rect 654506 506911 654512 506923
rect 663856 506911 663862 506923
rect 663914 506911 663920 506963
rect 53872 501139 53878 501191
rect 53930 501179 53936 501191
rect 59536 501179 59542 501191
rect 53930 501151 59542 501179
rect 53930 501139 53936 501151
rect 59536 501139 59542 501151
rect 59594 501139 59600 501191
rect 674608 499659 674614 499711
rect 674666 499699 674672 499711
rect 674992 499699 674998 499711
rect 674666 499671 674998 499699
rect 674666 499659 674672 499671
rect 674992 499659 674998 499671
rect 675050 499659 675056 499711
rect 675088 495959 675094 496011
rect 675146 495999 675152 496011
rect 675376 495999 675382 496011
rect 675146 495971 675382 495999
rect 675146 495959 675152 495971
rect 675376 495959 675382 495971
rect 675434 495959 675440 496011
rect 654352 495367 654358 495419
rect 654410 495407 654416 495419
rect 661168 495407 661174 495419
rect 654410 495379 661174 495407
rect 654410 495367 654416 495379
rect 661168 495367 661174 495379
rect 661226 495367 661232 495419
rect 664048 492925 664054 492977
rect 664106 492965 664112 492977
rect 674320 492965 674326 492977
rect 664106 492937 674326 492965
rect 664106 492925 664112 492937
rect 674320 492925 674326 492937
rect 674378 492925 674384 492977
rect 655312 492481 655318 492533
rect 655370 492521 655376 492533
rect 674608 492521 674614 492533
rect 655370 492493 674614 492521
rect 655370 492481 655376 492493
rect 674608 492481 674614 492493
rect 674666 492481 674672 492533
rect 672688 492407 672694 492459
rect 672746 492447 672752 492459
rect 673840 492447 673846 492459
rect 672746 492419 673846 492447
rect 672746 492407 672752 492419
rect 673840 492407 673846 492419
rect 673898 492407 673904 492459
rect 50416 486709 50422 486761
rect 50474 486749 50480 486761
rect 58576 486749 58582 486761
rect 50474 486721 58582 486749
rect 50474 486709 50480 486721
rect 58576 486709 58582 486721
rect 58634 486709 58640 486761
rect 654256 483823 654262 483875
rect 654314 483863 654320 483875
rect 666928 483863 666934 483875
rect 654314 483835 666934 483863
rect 654314 483823 654320 483835
rect 666928 483823 666934 483835
rect 666986 483823 666992 483875
rect 650320 479457 650326 479509
rect 650378 479497 650384 479509
rect 677008 479497 677014 479509
rect 650378 479469 677014 479497
rect 650378 479457 650384 479469
rect 677008 479457 677014 479469
rect 677066 479457 677072 479509
rect 44944 472353 44950 472405
rect 45002 472393 45008 472405
rect 59536 472393 59542 472405
rect 45002 472365 59542 472393
rect 45002 472353 45008 472365
rect 59536 472353 59542 472365
rect 59594 472353 59600 472405
rect 654448 472205 654454 472257
rect 654506 472245 654512 472257
rect 660976 472245 660982 472257
rect 654506 472217 660982 472245
rect 654506 472205 654512 472217
rect 660976 472205 660982 472217
rect 661034 472205 661040 472257
rect 47824 457923 47830 457975
rect 47882 457963 47888 457975
rect 59536 457963 59542 457975
rect 47882 457935 59542 457963
rect 47882 457923 47888 457935
rect 59536 457923 59542 457935
rect 59594 457923 59600 457975
rect 654448 457923 654454 457975
rect 654506 457963 654512 457975
rect 660976 457963 660982 457975
rect 654506 457935 660982 457963
rect 654506 457923 654512 457935
rect 660976 457923 660982 457935
rect 661034 457923 661040 457975
rect 654352 446379 654358 446431
rect 654410 446419 654416 446431
rect 672496 446419 672502 446431
rect 654410 446391 672502 446419
rect 654410 446379 654416 446391
rect 672496 446379 672502 446391
rect 672554 446379 672560 446431
rect 53680 443567 53686 443619
rect 53738 443607 53744 443619
rect 59536 443607 59542 443619
rect 53738 443579 59542 443607
rect 53738 443567 53744 443579
rect 59536 443567 59542 443579
rect 59594 443567 59600 443619
rect 654448 434909 654454 434961
rect 654506 434949 654512 434961
rect 663952 434949 663958 434961
rect 654506 434921 663958 434949
rect 654506 434909 654512 434921
rect 663952 434909 663958 434921
rect 664010 434909 664016 434961
rect 42832 432245 42838 432297
rect 42890 432285 42896 432297
rect 50512 432285 50518 432297
rect 42890 432257 50518 432285
rect 42890 432245 42896 432257
rect 50512 432245 50518 432257
rect 50570 432245 50576 432297
rect 42832 431727 42838 431779
rect 42890 431767 42896 431779
rect 53872 431767 53878 431779
rect 42890 431739 53878 431767
rect 42890 431727 42896 431739
rect 53872 431727 53878 431739
rect 53930 431727 53936 431779
rect 42832 429581 42838 429633
rect 42890 429621 42896 429633
rect 43600 429621 43606 429633
rect 42890 429593 43606 429621
rect 42890 429581 42896 429593
rect 43600 429581 43606 429593
rect 43658 429581 43664 429633
rect 47632 429137 47638 429189
rect 47690 429177 47696 429189
rect 59536 429177 59542 429189
rect 47690 429149 59542 429177
rect 47690 429137 47696 429149
rect 59536 429137 59542 429149
rect 59594 429137 59600 429189
rect 654448 426177 654454 426229
rect 654506 426217 654512 426229
rect 669616 426217 669622 426229
rect 654506 426189 669622 426217
rect 654506 426177 654512 426189
rect 669616 426177 669622 426189
rect 669674 426177 669680 426229
rect 42352 417593 42358 417645
rect 42410 417633 42416 417645
rect 56176 417633 56182 417645
rect 42410 417605 56182 417633
rect 42410 417593 42416 417605
rect 56176 417593 56182 417605
rect 56234 417593 56240 417645
rect 40240 416261 40246 416313
rect 40298 416301 40304 416313
rect 42736 416301 42742 416313
rect 40298 416273 42742 416301
rect 40298 416261 40304 416273
rect 42736 416261 42742 416273
rect 42794 416261 42800 416313
rect 40048 415669 40054 415721
rect 40106 415709 40112 415721
rect 43120 415709 43126 415721
rect 40106 415681 43126 415709
rect 40106 415669 40112 415681
rect 43120 415669 43126 415681
rect 43178 415669 43184 415721
rect 40144 415373 40150 415425
rect 40202 415413 40208 415425
rect 43024 415413 43030 415425
rect 40202 415385 43030 415413
rect 40202 415373 40208 415385
rect 43024 415373 43030 415385
rect 43082 415373 43088 415425
rect 39952 414707 39958 414759
rect 40010 414747 40016 414759
rect 43408 414747 43414 414759
rect 40010 414719 43414 414747
rect 40010 414707 40016 414719
rect 43408 414707 43414 414719
rect 43466 414707 43472 414759
rect 50512 414707 50518 414759
rect 50570 414747 50576 414759
rect 58384 414747 58390 414759
rect 50570 414719 58390 414747
rect 50570 414707 50576 414719
rect 58384 414707 58390 414719
rect 58442 414707 58448 414759
rect 41872 413375 41878 413427
rect 41930 413375 41936 413427
rect 41890 413205 41918 413375
rect 41872 413153 41878 413205
rect 41930 413153 41936 413205
rect 653872 411821 653878 411873
rect 653930 411861 653936 411873
rect 669616 411861 669622 411873
rect 653930 411833 669622 411861
rect 653930 411821 653936 411833
rect 669616 411821 669622 411833
rect 669674 411821 669680 411873
rect 42160 411303 42166 411355
rect 42218 411343 42224 411355
rect 42832 411343 42838 411355
rect 42218 411315 42838 411343
rect 42218 411303 42224 411315
rect 42832 411303 42838 411315
rect 42890 411303 42896 411355
rect 42064 410489 42070 410541
rect 42122 410529 42128 410541
rect 47440 410529 47446 410541
rect 42122 410501 47446 410529
rect 42122 410489 42128 410501
rect 47440 410489 47446 410501
rect 47498 410489 47504 410541
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42736 409493 42742 409505
rect 42218 409465 42742 409493
rect 42218 409453 42224 409465
rect 42736 409453 42742 409465
rect 42794 409453 42800 409505
rect 43024 409271 43030 409283
rect 42850 409243 43030 409271
rect 42850 409209 42878 409243
rect 43024 409231 43030 409243
rect 43082 409231 43088 409283
rect 42832 409157 42838 409209
rect 42890 409157 42896 409209
rect 42928 409083 42934 409135
rect 42986 409123 42992 409135
rect 43120 409123 43126 409135
rect 42986 409095 43126 409123
rect 42986 409083 42992 409095
rect 43120 409083 43126 409095
rect 43178 409083 43184 409135
rect 43120 408935 43126 408987
rect 43178 408975 43184 408987
rect 43408 408975 43414 408987
rect 43178 408947 43414 408975
rect 43178 408935 43184 408947
rect 43408 408935 43414 408947
rect 43466 408935 43472 408987
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 42736 408235 42742 408247
rect 42218 408207 42742 408235
rect 42218 408195 42224 408207
rect 42736 408195 42742 408207
rect 42794 408195 42800 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43120 407495 43126 407507
rect 42122 407467 43126 407495
rect 42122 407455 42128 407467
rect 43120 407455 43126 407467
rect 43178 407455 43184 407507
rect 42160 407011 42166 407063
rect 42218 407051 42224 407063
rect 42832 407051 42838 407063
rect 42218 407023 42838 407051
rect 42218 407011 42224 407023
rect 42832 407011 42838 407023
rect 42890 407011 42896 407063
rect 666832 405457 666838 405509
rect 666890 405497 666896 405509
rect 674704 405497 674710 405509
rect 666890 405469 674710 405497
rect 666890 405457 666896 405469
rect 674704 405457 674710 405469
rect 674762 405457 674768 405509
rect 669520 404717 669526 404769
rect 669578 404757 669584 404769
rect 674416 404757 674422 404769
rect 669578 404729 674422 404757
rect 669578 404717 669584 404729
rect 674416 404717 674422 404729
rect 674474 404717 674480 404769
rect 669712 404421 669718 404473
rect 669770 404461 669776 404473
rect 674704 404461 674710 404473
rect 669770 404433 674710 404461
rect 669770 404421 669776 404433
rect 674704 404421 674710 404433
rect 674762 404421 674768 404473
rect 42160 403681 42166 403733
rect 42218 403721 42224 403733
rect 42736 403721 42742 403733
rect 42218 403693 42742 403721
rect 42218 403681 42224 403693
rect 42736 403681 42742 403693
rect 42794 403681 42800 403733
rect 673456 400499 673462 400551
rect 673514 400539 673520 400551
rect 677296 400539 677302 400551
rect 673514 400511 677302 400539
rect 673514 400499 673520 400511
rect 677296 400499 677302 400511
rect 677354 400499 677360 400551
rect 673360 400425 673366 400477
rect 673418 400465 673424 400477
rect 677104 400465 677110 400477
rect 673418 400437 677110 400465
rect 673418 400425 673424 400437
rect 677104 400425 677110 400437
rect 677162 400425 677168 400477
rect 45040 400351 45046 400403
rect 45098 400391 45104 400403
rect 58384 400391 58390 400403
rect 45098 400363 58390 400391
rect 45098 400351 45104 400363
rect 58384 400351 58390 400363
rect 58442 400351 58448 400403
rect 654448 400351 654454 400403
rect 654506 400391 654512 400403
rect 666832 400391 666838 400403
rect 654506 400363 666838 400391
rect 654506 400351 654512 400363
rect 666832 400351 666838 400363
rect 666890 400351 666896 400403
rect 673648 400351 673654 400403
rect 673706 400391 673712 400403
rect 673840 400391 673846 400403
rect 673706 400363 673846 400391
rect 673706 400351 673712 400363
rect 673840 400351 673846 400363
rect 673898 400351 673904 400403
rect 650416 391767 650422 391819
rect 650474 391807 650480 391819
rect 677104 391807 677110 391819
rect 650474 391779 677110 391807
rect 650474 391767 650480 391779
rect 677104 391767 677110 391779
rect 677162 391767 677168 391819
rect 42352 389325 42358 389377
rect 42410 389365 42416 389377
rect 44944 389365 44950 389377
rect 42410 389337 44950 389365
rect 42410 389325 42416 389337
rect 44944 389325 44950 389337
rect 45002 389325 45008 389377
rect 654448 388807 654454 388859
rect 654506 388847 654512 388859
rect 669520 388847 669526 388859
rect 654506 388819 669526 388847
rect 654506 388807 654512 388819
rect 669520 388807 669526 388819
rect 669578 388807 669584 388859
rect 42352 388733 42358 388785
rect 42410 388773 42416 388785
rect 47824 388773 47830 388785
rect 42410 388745 47830 388773
rect 42410 388733 42416 388745
rect 47824 388733 47830 388745
rect 47882 388733 47888 388785
rect 42736 387993 42742 388045
rect 42794 388033 42800 388045
rect 50416 388033 50422 388045
rect 42794 388005 50422 388033
rect 42794 387993 42800 388005
rect 50416 387993 50422 388005
rect 50474 387993 50480 388045
rect 674992 386143 674998 386195
rect 675050 386183 675056 386195
rect 675376 386183 675382 386195
rect 675050 386155 675382 386183
rect 675050 386143 675056 386155
rect 675376 386143 675382 386155
rect 675434 386143 675440 386195
rect 47728 385921 47734 385973
rect 47786 385961 47792 385973
rect 59248 385961 59254 385973
rect 47786 385933 59254 385961
rect 47786 385921 47792 385933
rect 59248 385921 59254 385933
rect 59306 385921 59312 385973
rect 675184 385477 675190 385529
rect 675242 385517 675248 385529
rect 675242 385489 675518 385517
rect 675242 385477 675248 385489
rect 675490 385455 675518 385489
rect 675472 385403 675478 385455
rect 675530 385403 675536 385455
rect 674704 385181 674710 385233
rect 674762 385221 674768 385233
rect 674992 385221 674998 385233
rect 674762 385193 674998 385221
rect 674762 385181 674768 385193
rect 674992 385181 674998 385193
rect 675050 385181 675056 385233
rect 674896 384811 674902 384863
rect 674954 384851 674960 384863
rect 675376 384851 675382 384863
rect 674954 384823 675382 384851
rect 674954 384811 674960 384823
rect 675376 384811 675382 384823
rect 675434 384811 675440 384863
rect 674512 383109 674518 383161
rect 674570 383149 674576 383161
rect 675376 383149 675382 383161
rect 674570 383121 675382 383149
rect 674570 383109 674576 383121
rect 675376 383109 675382 383121
rect 675434 383109 675440 383161
rect 674416 382295 674422 382347
rect 674474 382335 674480 382347
rect 675472 382335 675478 382347
rect 674474 382307 675478 382335
rect 674474 382295 674480 382307
rect 675472 382295 675478 382307
rect 675530 382295 675536 382347
rect 654448 380075 654454 380127
rect 654506 380115 654512 380127
rect 666736 380115 666742 380127
rect 654506 380087 666742 380115
rect 654506 380075 654512 380087
rect 666736 380075 666742 380087
rect 666794 380075 666800 380127
rect 674800 378151 674806 378203
rect 674858 378191 674864 378203
rect 675376 378191 675382 378203
rect 674858 378163 675382 378191
rect 674858 378151 674864 378163
rect 675376 378151 675382 378163
rect 675434 378151 675440 378203
rect 674608 377559 674614 377611
rect 674666 377599 674672 377611
rect 675376 377599 675382 377611
rect 674666 377571 675382 377599
rect 674666 377559 674672 377571
rect 675376 377559 675382 377571
rect 675434 377559 675440 377611
rect 674224 376819 674230 376871
rect 674282 376859 674288 376871
rect 675472 376859 675478 376871
rect 674282 376831 675478 376859
rect 674282 376819 674288 376831
rect 675472 376819 675478 376831
rect 675530 376819 675536 376871
rect 42640 376523 42646 376575
rect 42698 376563 42704 376575
rect 44944 376563 44950 376575
rect 42698 376535 44950 376563
rect 42698 376523 42704 376535
rect 44944 376523 44950 376535
rect 45002 376523 45008 376575
rect 673936 375709 673942 375761
rect 673994 375749 674000 375761
rect 675472 375749 675478 375761
rect 673994 375721 675478 375749
rect 673994 375709 674000 375721
rect 675472 375709 675478 375721
rect 675530 375709 675536 375761
rect 40240 373341 40246 373393
rect 40298 373381 40304 373393
rect 43408 373381 43414 373393
rect 40298 373353 43414 373381
rect 40298 373341 40304 373353
rect 43408 373341 43414 373353
rect 43466 373341 43472 373393
rect 39952 372379 39958 372431
rect 40010 372419 40016 372431
rect 43024 372419 43030 372431
rect 40010 372391 43030 372419
rect 40010 372379 40016 372391
rect 43024 372379 43030 372391
rect 43082 372379 43088 372431
rect 39856 371565 39862 371617
rect 39914 371605 39920 371617
rect 43312 371605 43318 371617
rect 39914 371577 43318 371605
rect 39914 371565 39920 371577
rect 43312 371565 43318 371577
rect 43370 371565 43376 371617
rect 50416 371565 50422 371617
rect 50474 371605 50480 371617
rect 59536 371605 59542 371617
rect 50474 371577 59542 371605
rect 50474 371565 50480 371577
rect 59536 371565 59542 371577
rect 59594 371565 59600 371617
rect 42160 370159 42166 370211
rect 42218 370199 42224 370211
rect 42218 370171 42590 370199
rect 42218 370159 42224 370171
rect 42160 369937 42166 369989
rect 42218 369977 42224 369989
rect 42352 369977 42358 369989
rect 42218 369949 42358 369977
rect 42218 369937 42224 369949
rect 42352 369937 42358 369949
rect 42410 369937 42416 369989
rect 42562 368879 42590 370171
rect 42544 368827 42550 368879
rect 42602 368827 42608 368879
rect 42064 368087 42070 368139
rect 42122 368127 42128 368139
rect 42544 368127 42550 368139
rect 42122 368099 42550 368127
rect 42122 368087 42128 368099
rect 42544 368087 42550 368099
rect 42602 368087 42608 368139
rect 42928 367569 42934 367621
rect 42986 367609 42992 367621
rect 43312 367609 43318 367621
rect 42986 367581 43318 367609
rect 42986 367569 42992 367581
rect 43312 367569 43318 367581
rect 43370 367569 43376 367621
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 50320 367387 50326 367399
rect 42122 367359 50326 367387
rect 42122 367347 42128 367359
rect 50320 367347 50326 367359
rect 50378 367347 50384 367399
rect 42064 366163 42070 366215
rect 42122 366203 42128 366215
rect 43024 366203 43030 366215
rect 42122 366175 43030 366203
rect 42122 366163 42128 366175
rect 43024 366163 43030 366175
rect 43082 366163 43088 366215
rect 654448 365793 654454 365845
rect 654506 365833 654512 365845
rect 661072 365833 661078 365845
rect 654506 365805 661078 365833
rect 654506 365793 654512 365805
rect 661072 365793 661078 365805
rect 661130 365793 661136 365845
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 43120 365019 43126 365031
rect 42218 364991 43126 365019
rect 42218 364979 42224 364991
rect 43120 364979 43126 364991
rect 43178 364979 43184 365031
rect 42064 364387 42070 364439
rect 42122 364427 42128 364439
rect 42640 364427 42646 364439
rect 42122 364399 42646 364427
rect 42122 364387 42128 364399
rect 42640 364387 42646 364399
rect 42698 364387 42704 364439
rect 42160 363795 42166 363847
rect 42218 363835 42224 363847
rect 43408 363835 43414 363847
rect 42218 363807 43414 363835
rect 42218 363795 42224 363807
rect 43408 363795 43414 363807
rect 43466 363795 43472 363847
rect 42160 360613 42166 360665
rect 42218 360653 42224 360665
rect 42928 360653 42934 360665
rect 42218 360625 42934 360653
rect 42218 360613 42224 360625
rect 42928 360613 42934 360625
rect 42986 360613 42992 360665
rect 672400 360021 672406 360073
rect 672458 360061 672464 360073
rect 674416 360061 674422 360073
rect 672458 360033 674422 360061
rect 672458 360021 672464 360033
rect 674416 360021 674422 360033
rect 674474 360021 674480 360073
rect 666640 359725 666646 359777
rect 666698 359765 666704 359777
rect 674704 359765 674710 359777
rect 666698 359737 674710 359765
rect 666698 359725 666704 359737
rect 674704 359725 674710 359737
rect 674762 359725 674768 359777
rect 672592 358985 672598 359037
rect 672650 359025 672656 359037
rect 674416 359025 674422 359037
rect 672650 358997 674422 359025
rect 672650 358985 672656 358997
rect 674416 358985 674422 358997
rect 674474 358985 674480 359037
rect 47440 357135 47446 357187
rect 47498 357175 47504 357187
rect 59536 357175 59542 357187
rect 47498 357147 59542 357175
rect 47498 357135 47504 357147
rect 59536 357135 59542 357147
rect 59594 357135 59600 357187
rect 42448 346109 42454 346161
rect 42506 346149 42512 346161
rect 47632 346149 47638 346161
rect 42506 346121 47638 346149
rect 42506 346109 42512 346121
rect 47632 346109 47638 346121
rect 47690 346109 47696 346161
rect 650512 345591 650518 345643
rect 650570 345631 650576 345643
rect 677104 345631 677110 345643
rect 650570 345603 677110 345631
rect 650570 345591 650576 345603
rect 677104 345591 677110 345603
rect 677162 345591 677168 345643
rect 42448 345517 42454 345569
rect 42506 345557 42512 345569
rect 50512 345557 50518 345569
rect 42506 345529 50518 345557
rect 42506 345517 42512 345529
rect 50512 345517 50518 345529
rect 50570 345517 50576 345569
rect 42928 344777 42934 344829
rect 42986 344817 42992 344829
rect 53680 344817 53686 344829
rect 42986 344789 53686 344817
rect 42986 344777 42992 344789
rect 53680 344777 53686 344789
rect 53738 344777 53744 344829
rect 53872 342779 53878 342831
rect 53930 342819 53936 342831
rect 58384 342819 58390 342831
rect 53930 342791 58390 342819
rect 53930 342779 53936 342791
rect 58384 342779 58390 342791
rect 58442 342779 58448 342831
rect 654448 342705 654454 342757
rect 654506 342745 654512 342757
rect 666640 342745 666646 342757
rect 654506 342717 666646 342745
rect 654506 342705 654512 342717
rect 666640 342705 666646 342717
rect 666698 342705 666704 342757
rect 674800 341595 674806 341647
rect 674858 341635 674864 341647
rect 675184 341635 675190 341647
rect 674858 341607 675190 341635
rect 674858 341595 674864 341607
rect 675184 341595 675190 341607
rect 675242 341595 675248 341647
rect 674896 341299 674902 341351
rect 674954 341339 674960 341351
rect 675088 341339 675094 341351
rect 674954 341311 675094 341339
rect 674954 341299 674960 341311
rect 675088 341299 675094 341311
rect 675146 341299 675152 341351
rect 674608 339745 674614 339797
rect 674666 339785 674672 339797
rect 675088 339785 675094 339797
rect 674666 339757 675094 339785
rect 674666 339745 674672 339757
rect 675088 339745 675094 339757
rect 675146 339745 675152 339797
rect 674416 339523 674422 339575
rect 674474 339563 674480 339575
rect 675376 339563 675382 339575
rect 674474 339535 675382 339563
rect 674474 339523 674480 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 674512 337229 674518 337281
rect 674570 337269 674576 337281
rect 675088 337269 675094 337281
rect 674570 337241 675094 337269
rect 674570 337229 674576 337241
rect 675088 337229 675094 337241
rect 675146 337229 675152 337281
rect 673936 333529 673942 333581
rect 673994 333569 674000 333581
rect 675376 333569 675382 333581
rect 673994 333541 675382 333569
rect 673994 333529 674000 333541
rect 675376 333529 675382 333541
rect 675434 333529 675440 333581
rect 42832 333307 42838 333359
rect 42890 333347 42896 333359
rect 47632 333347 47638 333359
rect 42890 333319 47638 333347
rect 42890 333307 42896 333319
rect 47632 333307 47638 333319
rect 47690 333307 47696 333359
rect 674224 332937 674230 332989
rect 674282 332977 674288 332989
rect 675376 332977 675382 332989
rect 674282 332949 675382 332977
rect 674282 332937 674288 332949
rect 675376 332937 675382 332949
rect 675434 332937 675440 332989
rect 654448 332271 654454 332323
rect 654506 332311 654512 332323
rect 663760 332311 663766 332323
rect 654506 332283 663766 332311
rect 654506 332271 654512 332283
rect 663760 332271 663766 332283
rect 663818 332271 663824 332323
rect 674320 332197 674326 332249
rect 674378 332237 674384 332249
rect 675472 332237 675478 332249
rect 674378 332209 675478 332237
rect 674378 332197 674384 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 674032 331531 674038 331583
rect 674090 331571 674096 331583
rect 675376 331571 675382 331583
rect 674090 331543 675382 331571
rect 674090 331531 674096 331543
rect 675376 331531 675382 331543
rect 675434 331531 675440 331583
rect 39856 329755 39862 329807
rect 39914 329795 39920 329807
rect 43120 329795 43126 329807
rect 39914 329767 43126 329795
rect 39914 329755 39920 329767
rect 43120 329755 43126 329767
rect 43178 329755 43184 329807
rect 40048 329459 40054 329511
rect 40106 329499 40112 329511
rect 42832 329499 42838 329511
rect 40106 329471 42838 329499
rect 40106 329459 40112 329471
rect 42832 329459 42838 329471
rect 42890 329459 42896 329511
rect 39952 329311 39958 329363
rect 40010 329351 40016 329363
rect 42448 329351 42454 329363
rect 40010 329323 42454 329351
rect 40010 329311 40016 329323
rect 42448 329311 42454 329323
rect 42506 329311 42512 329363
rect 40240 329163 40246 329215
rect 40298 329203 40304 329215
rect 42352 329203 42358 329215
rect 40298 329175 42358 329203
rect 40298 329163 40304 329175
rect 42352 329163 42358 329175
rect 42410 329163 42416 329215
rect 50320 328349 50326 328401
rect 50378 328389 50384 328401
rect 57808 328389 57814 328401
rect 50378 328361 57814 328389
rect 50378 328349 50384 328361
rect 57808 328349 57814 328361
rect 57866 328349 57872 328401
rect 41872 327017 41878 327069
rect 41930 327017 41936 327069
rect 41890 326773 41918 327017
rect 41872 326721 41878 326773
rect 41930 326721 41936 326773
rect 42448 325611 42454 325663
rect 42506 325651 42512 325663
rect 42506 325623 42878 325651
rect 42506 325611 42512 325623
rect 42736 325315 42742 325367
rect 42794 325355 42800 325367
rect 42850 325355 42878 325623
rect 42794 325327 42878 325355
rect 42794 325315 42800 325327
rect 42064 324871 42070 324923
rect 42122 324911 42128 324923
rect 42928 324911 42934 324923
rect 42122 324883 42934 324911
rect 42122 324871 42128 324883
rect 42928 324871 42934 324883
rect 42986 324871 42992 324923
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 44656 324171 44662 324183
rect 42218 324143 44662 324171
rect 42218 324131 42224 324143
rect 44656 324131 44662 324143
rect 44714 324131 44720 324183
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 42736 323135 42742 323147
rect 42218 323107 42742 323135
rect 42218 323095 42224 323107
rect 42736 323095 42742 323107
rect 42794 323095 42800 323147
rect 42832 322987 42838 322999
rect 42370 322959 42838 322987
rect 42370 322765 42398 322959
rect 42832 322947 42838 322959
rect 42890 322947 42896 322999
rect 42448 322765 42454 322777
rect 42370 322737 42454 322765
rect 42448 322725 42454 322737
rect 42506 322725 42512 322777
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 43024 321803 43030 321815
rect 42122 321775 43030 321803
rect 42122 321763 42128 321775
rect 43024 321763 43030 321775
rect 43082 321763 43088 321815
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 42448 321063 42454 321075
rect 42218 321035 42454 321063
rect 42218 321023 42224 321035
rect 42448 321023 42454 321035
rect 42506 321023 42512 321075
rect 42160 320579 42166 320631
rect 42218 320619 42224 320631
rect 43120 320619 43126 320631
rect 42218 320591 43126 320619
rect 42218 320579 42224 320591
rect 43120 320579 43126 320591
rect 43178 320579 43184 320631
rect 42160 317471 42166 317523
rect 42218 317511 42224 317523
rect 42448 317511 42454 317523
rect 42218 317483 42454 317511
rect 42218 317471 42224 317483
rect 42448 317471 42454 317483
rect 42506 317471 42512 317523
rect 661168 315029 661174 315081
rect 661226 315069 661232 315081
rect 674416 315069 674422 315081
rect 661226 315041 674422 315069
rect 661226 315029 661232 315041
rect 674416 315029 674422 315041
rect 674474 315029 674480 315081
rect 663856 314733 663862 314785
rect 663914 314773 663920 314785
rect 674704 314773 674710 314785
rect 663914 314745 674710 314773
rect 663914 314733 663920 314745
rect 674704 314733 674710 314745
rect 674762 314733 674768 314785
rect 666928 313993 666934 314045
rect 666986 314033 666992 314045
rect 674416 314033 674422 314045
rect 666986 314005 674422 314033
rect 666986 313993 666992 314005
rect 674416 313993 674422 314005
rect 674474 313993 674480 314045
rect 44656 313919 44662 313971
rect 44714 313959 44720 313971
rect 58000 313959 58006 313971
rect 44714 313931 58006 313959
rect 44714 313919 44720 313931
rect 58000 313919 58006 313931
rect 58058 313919 58064 313971
rect 42544 302893 42550 302945
rect 42602 302933 42608 302945
rect 47728 302933 47734 302945
rect 42602 302905 47734 302933
rect 42602 302893 42608 302905
rect 47728 302893 47734 302905
rect 47786 302893 47792 302945
rect 650608 302597 650614 302649
rect 650666 302637 650672 302649
rect 674416 302637 674422 302649
rect 650666 302609 674422 302637
rect 650666 302597 650672 302609
rect 674416 302597 674422 302609
rect 674474 302597 674480 302649
rect 42544 302301 42550 302353
rect 42602 302341 42608 302353
rect 50416 302341 50422 302353
rect 42602 302313 50422 302341
rect 42602 302301 42608 302313
rect 50416 302301 50422 302313
rect 50474 302301 50480 302353
rect 42544 301857 42550 301909
rect 42602 301897 42608 301909
rect 45040 301897 45046 301909
rect 42602 301869 45046 301897
rect 42602 301857 42608 301869
rect 45040 301857 45046 301869
rect 45098 301857 45104 301909
rect 674512 300525 674518 300577
rect 674570 300565 674576 300577
rect 674704 300565 674710 300577
rect 674570 300537 674710 300565
rect 674570 300525 674576 300537
rect 674704 300525 674710 300537
rect 674762 300525 674768 300577
rect 45136 299563 45142 299615
rect 45194 299603 45200 299615
rect 59440 299603 59446 299615
rect 45194 299575 59446 299603
rect 45194 299563 45200 299575
rect 59440 299563 59446 299575
rect 59498 299563 59504 299615
rect 674512 295937 674518 295989
rect 674570 295977 674576 295989
rect 675376 295977 675382 295989
rect 674570 295949 675382 295977
rect 674570 295937 674576 295949
rect 675376 295937 675382 295949
rect 675434 295937 675440 295989
rect 674896 295345 674902 295397
rect 674954 295385 674960 295397
rect 675472 295385 675478 295397
rect 674954 295357 675478 295385
rect 674954 295345 674960 295357
rect 675472 295345 675478 295357
rect 675530 295345 675536 295397
rect 673936 294531 673942 294583
rect 673994 294571 674000 294583
rect 675376 294571 675382 294583
rect 673994 294543 675382 294571
rect 673994 294531 674000 294543
rect 675376 294531 675382 294543
rect 675434 294531 675440 294583
rect 654544 293791 654550 293843
rect 654602 293831 654608 293843
rect 663760 293831 663766 293843
rect 654602 293803 663766 293831
rect 654602 293791 654608 293803
rect 663760 293791 663766 293803
rect 663818 293791 663824 293843
rect 674320 292903 674326 292955
rect 674378 292943 674384 292955
rect 675376 292943 675382 292955
rect 674378 292915 675382 292943
rect 674378 292903 674384 292915
rect 675376 292903 675382 292915
rect 675434 292903 675440 292955
rect 674800 291719 674806 291771
rect 674858 291759 674864 291771
rect 675088 291759 675094 291771
rect 674858 291731 675094 291759
rect 674858 291719 674864 291731
rect 675088 291719 675094 291731
rect 675146 291719 675152 291771
rect 674608 291053 674614 291105
rect 674666 291093 674672 291105
rect 675088 291093 675094 291105
rect 674666 291065 675094 291093
rect 674666 291053 674672 291065
rect 675088 291053 675094 291065
rect 675146 291053 675152 291105
rect 42544 289795 42550 289847
rect 42602 289835 42608 289847
rect 47728 289835 47734 289847
rect 42602 289807 47734 289835
rect 42602 289795 42608 289807
rect 47728 289795 47734 289807
rect 47786 289795 47792 289847
rect 674992 288537 674998 288589
rect 675050 288577 675056 288589
rect 675472 288577 675478 288589
rect 675050 288549 675478 288577
rect 675050 288537 675056 288549
rect 675472 288537 675478 288549
rect 675530 288537 675536 288589
rect 674416 287723 674422 287775
rect 674474 287763 674480 287775
rect 675376 287763 675382 287775
rect 674474 287735 675382 287763
rect 674474 287723 674480 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 674032 287205 674038 287257
rect 674090 287245 674096 287257
rect 675472 287245 675478 287257
rect 674090 287217 675478 287245
rect 674090 287205 674096 287217
rect 675472 287205 675478 287217
rect 675530 287205 675536 287257
rect 674224 286761 674230 286813
rect 674282 286801 674288 286813
rect 675376 286801 675382 286813
rect 674282 286773 675382 286801
rect 674282 286761 674288 286773
rect 675376 286761 675382 286773
rect 675434 286761 675440 286813
rect 39856 285429 39862 285481
rect 39914 285469 39920 285481
rect 43120 285469 43126 285481
rect 39914 285441 43126 285469
rect 39914 285429 39920 285441
rect 43120 285429 43126 285441
rect 43178 285429 43184 285481
rect 40048 285281 40054 285333
rect 40106 285321 40112 285333
rect 43120 285321 43126 285333
rect 40106 285293 43126 285321
rect 40106 285281 40112 285293
rect 43120 285281 43126 285293
rect 43178 285281 43184 285333
rect 40144 285133 40150 285185
rect 40202 285173 40208 285185
rect 43024 285173 43030 285185
rect 40202 285145 43030 285173
rect 40202 285133 40208 285145
rect 43024 285133 43030 285145
rect 43082 285133 43088 285185
rect 45040 285133 45046 285185
rect 45098 285173 45104 285185
rect 58096 285173 58102 285185
rect 45098 285145 58102 285173
rect 45098 285133 45104 285145
rect 58096 285133 58102 285145
rect 58154 285133 58160 285185
rect 654064 284763 654070 284815
rect 654122 284803 654128 284815
rect 660880 284803 660886 284815
rect 654122 284775 660886 284803
rect 654122 284763 654128 284775
rect 660880 284763 660886 284775
rect 660938 284763 660944 284815
rect 41200 284097 41206 284149
rect 41258 284137 41264 284149
rect 41258 284109 42494 284137
rect 41258 284097 41264 284109
rect 41968 283801 41974 283853
rect 42026 283801 42032 283853
rect 41986 283557 42014 283801
rect 42466 283631 42494 284109
rect 42448 283579 42454 283631
rect 42506 283579 42512 283631
rect 41968 283505 41974 283557
rect 42026 283505 42032 283557
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42448 281769 42454 281781
rect 42218 281741 42454 281769
rect 42218 281729 42224 281741
rect 42448 281729 42454 281741
rect 42506 281729 42512 281781
rect 42160 281063 42166 281115
rect 42218 281103 42224 281115
rect 53488 281103 53494 281115
rect 42218 281075 53494 281103
rect 42218 281063 42224 281075
rect 53488 281063 53494 281075
rect 53546 281063 53552 281115
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 43024 279919 43030 279931
rect 42218 279891 43030 279919
rect 42218 279879 42224 279891
rect 43024 279879 43030 279891
rect 43082 279879 43088 279931
rect 43120 279879 43126 279931
rect 43178 279879 43184 279931
rect 43138 279709 43166 279879
rect 43120 279657 43126 279709
rect 43178 279657 43184 279709
rect 318160 278661 318166 278673
rect 295810 278633 318166 278661
rect 295810 278599 295838 278633
rect 318160 278621 318166 278633
rect 318218 278621 318224 278673
rect 379426 278633 403358 278661
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42928 278587 42934 278599
rect 42218 278559 42934 278587
rect 42218 278547 42224 278559
rect 42928 278547 42934 278559
rect 42986 278547 42992 278599
rect 64720 278547 64726 278599
rect 64778 278587 64784 278599
rect 66640 278587 66646 278599
rect 64778 278559 66646 278587
rect 64778 278547 64784 278559
rect 66640 278547 66646 278559
rect 66698 278547 66704 278599
rect 295792 278547 295798 278599
rect 295850 278547 295856 278599
rect 309040 278547 309046 278599
rect 309098 278587 309104 278599
rect 370480 278587 370486 278599
rect 309098 278559 370486 278587
rect 309098 278547 309104 278559
rect 370480 278547 370486 278559
rect 370538 278547 370544 278599
rect 370960 278547 370966 278599
rect 371018 278587 371024 278599
rect 379024 278587 379030 278599
rect 371018 278559 379030 278587
rect 371018 278547 371024 278559
rect 379024 278547 379030 278559
rect 379082 278547 379088 278599
rect 379120 278547 379126 278599
rect 379178 278587 379184 278599
rect 379426 278587 379454 278633
rect 403330 278599 403358 278633
rect 379178 278559 379454 278587
rect 379178 278547 379184 278559
rect 379696 278547 379702 278599
rect 379754 278587 379760 278599
rect 396208 278587 396214 278599
rect 379754 278559 396214 278587
rect 379754 278547 379760 278559
rect 396208 278547 396214 278559
rect 396266 278547 396272 278599
rect 403312 278547 403318 278599
rect 403370 278547 403376 278599
rect 266032 278473 266038 278525
rect 266090 278513 266096 278525
rect 334384 278513 334390 278525
rect 266090 278485 334390 278513
rect 266090 278473 266096 278485
rect 334384 278473 334390 278485
rect 334442 278473 334448 278525
rect 338320 278473 338326 278525
rect 338378 278513 338384 278525
rect 358576 278513 358582 278525
rect 338378 278485 358582 278513
rect 338378 278473 338384 278485
rect 358576 278473 358582 278485
rect 358634 278473 358640 278525
rect 373168 278473 373174 278525
rect 373226 278513 373232 278525
rect 387760 278513 387766 278525
rect 373226 278485 387766 278513
rect 373226 278473 373232 278485
rect 387760 278473 387766 278485
rect 387818 278473 387824 278525
rect 388336 278473 388342 278525
rect 388394 278513 388400 278525
rect 490192 278513 490198 278525
rect 388394 278485 490198 278513
rect 388394 278473 388400 278485
rect 490192 278473 490198 278485
rect 490250 278473 490256 278525
rect 223120 278399 223126 278451
rect 223178 278439 223184 278451
rect 329104 278439 329110 278451
rect 223178 278411 329110 278439
rect 223178 278399 223184 278411
rect 329104 278399 329110 278411
rect 329162 278399 329168 278451
rect 350320 278399 350326 278451
rect 350378 278439 350384 278451
rect 393808 278439 393814 278451
rect 350378 278411 393814 278439
rect 350378 278399 350384 278411
rect 393808 278399 393814 278411
rect 393866 278399 393872 278451
rect 293776 278325 293782 278377
rect 293834 278365 293840 278377
rect 389008 278365 389014 278377
rect 293834 278337 389014 278365
rect 293834 278325 293840 278337
rect 389008 278325 389014 278337
rect 389066 278325 389072 278377
rect 292048 278251 292054 278303
rect 292106 278291 292112 278303
rect 374800 278291 374806 278303
rect 292106 278263 374806 278291
rect 292106 278251 292112 278263
rect 374800 278251 374806 278263
rect 374858 278251 374864 278303
rect 375472 278251 375478 278303
rect 375530 278291 375536 278303
rect 385072 278291 385078 278303
rect 375530 278263 385078 278291
rect 375530 278251 375536 278263
rect 385072 278251 385078 278263
rect 385130 278251 385136 278303
rect 301840 278177 301846 278229
rect 301898 278217 301904 278229
rect 453232 278217 453238 278229
rect 301898 278189 453238 278217
rect 301898 278177 301904 278189
rect 453232 278177 453238 278189
rect 453290 278177 453296 278229
rect 198160 278103 198166 278155
rect 198218 278143 198224 278155
rect 325264 278143 325270 278155
rect 198218 278115 325270 278143
rect 198218 278103 198224 278115
rect 325264 278103 325270 278115
rect 325322 278103 325328 278155
rect 326608 278103 326614 278155
rect 326666 278143 326672 278155
rect 635248 278143 635254 278155
rect 326666 278115 635254 278143
rect 326666 278103 326672 278115
rect 635248 278103 635254 278115
rect 635306 278103 635312 278155
rect 297520 278029 297526 278081
rect 297578 278069 297584 278081
rect 417616 278069 417622 278081
rect 297578 278041 417622 278069
rect 297578 278029 297584 278041
rect 417616 278029 417622 278041
rect 417674 278029 417680 278081
rect 290800 277955 290806 278007
rect 290858 277995 290864 278007
rect 309424 277995 309430 278007
rect 290858 277967 309430 277995
rect 290858 277955 290864 277967
rect 309424 277955 309430 277967
rect 309482 277955 309488 278007
rect 311824 277955 311830 278007
rect 311882 277995 311888 278007
rect 328144 277995 328150 278007
rect 311882 277967 328150 277995
rect 311882 277955 311888 277967
rect 328144 277955 328150 277967
rect 328202 277955 328208 278007
rect 353488 277955 353494 278007
rect 353546 277995 353552 278007
rect 353546 277967 357374 277995
rect 353546 277955 353552 277967
rect 64816 277881 64822 277933
rect 64874 277921 64880 277933
rect 182224 277921 182230 277933
rect 64874 277893 182230 277921
rect 64874 277881 64880 277893
rect 182224 277881 182230 277893
rect 182282 277881 182288 277933
rect 301552 277881 301558 277933
rect 301610 277921 301616 277933
rect 311920 277921 311926 277933
rect 301610 277893 311926 277921
rect 301610 277881 301616 277893
rect 311920 277881 311926 277893
rect 311978 277881 311984 277933
rect 312400 277881 312406 277933
rect 312458 277921 312464 277933
rect 339952 277921 339958 277933
rect 312458 277893 339958 277921
rect 312458 277881 312464 277893
rect 339952 277881 339958 277893
rect 340010 277881 340016 277933
rect 355504 277881 355510 277933
rect 355562 277921 355568 277933
rect 357346 277921 357374 277967
rect 357424 277955 357430 278007
rect 357482 277995 357488 278007
rect 415312 277995 415318 278007
rect 357482 277967 415318 277995
rect 357482 277955 357488 277967
rect 415312 277955 415318 277967
rect 415370 277955 415376 278007
rect 422320 277921 422326 277933
rect 355562 277893 357278 277921
rect 357346 277893 422326 277921
rect 355562 277881 355568 277893
rect 287248 277807 287254 277859
rect 287306 277847 287312 277859
rect 335536 277847 335542 277859
rect 287306 277819 335542 277847
rect 287306 277807 287312 277819
rect 335536 277807 335542 277819
rect 335594 277807 335600 277859
rect 356848 277807 356854 277859
rect 356906 277847 356912 277859
rect 357250 277847 357278 277893
rect 422320 277881 422326 277893
rect 422378 277881 422384 277933
rect 436624 277847 436630 277859
rect 356906 277819 357182 277847
rect 357250 277819 436630 277847
rect 356906 277807 356912 277819
rect 289936 277733 289942 277785
rect 289994 277773 290000 277785
rect 357040 277773 357046 277785
rect 289994 277745 357046 277773
rect 289994 277733 290000 277745
rect 357040 277733 357046 277745
rect 357098 277733 357104 277785
rect 357154 277773 357182 277819
rect 436624 277807 436630 277819
rect 436682 277807 436688 277859
rect 450832 277773 450838 277785
rect 357154 277745 450838 277773
rect 450832 277733 450838 277745
rect 450890 277733 450896 277785
rect 291472 277659 291478 277711
rect 291530 277699 291536 277711
rect 356944 277699 356950 277711
rect 291530 277671 356950 277699
rect 291530 277659 291536 277671
rect 356944 277659 356950 277671
rect 357002 277659 357008 277711
rect 358864 277659 358870 277711
rect 358922 277699 358928 277711
rect 465520 277699 465526 277711
rect 358922 277671 465526 277699
rect 358922 277659 358928 277671
rect 465520 277659 465526 277671
rect 465578 277659 465584 277711
rect 296464 277585 296470 277637
rect 296522 277625 296528 277637
rect 410800 277625 410806 277637
rect 296522 277597 410806 277625
rect 296522 277585 296528 277597
rect 410800 277585 410806 277597
rect 410858 277585 410864 277637
rect 293200 277511 293206 277563
rect 293258 277551 293264 277563
rect 382288 277551 382294 277563
rect 293258 277523 382294 277551
rect 293258 277511 293264 277523
rect 382288 277511 382294 277523
rect 382346 277511 382352 277563
rect 307984 277437 307990 277489
rect 308042 277477 308048 277489
rect 318064 277477 318070 277489
rect 308042 277449 318070 277477
rect 308042 277437 308048 277449
rect 318064 277437 318070 277449
rect 318122 277437 318128 277489
rect 318352 277437 318358 277489
rect 318410 277477 318416 277489
rect 331312 277477 331318 277489
rect 318410 277449 331318 277477
rect 318410 277437 318416 277449
rect 331312 277437 331318 277449
rect 331370 277437 331376 277489
rect 352912 277437 352918 277489
rect 352970 277477 352976 277489
rect 357424 277477 357430 277489
rect 352970 277449 357430 277477
rect 352970 277437 352976 277449
rect 357424 277437 357430 277449
rect 357482 277437 357488 277489
rect 361552 277437 361558 277489
rect 361610 277477 361616 277489
rect 486832 277477 486838 277489
rect 361610 277449 486838 277477
rect 361610 277437 361616 277449
rect 486832 277437 486838 277449
rect 486890 277437 486896 277489
rect 247888 277363 247894 277415
rect 247946 277403 247952 277415
rect 292240 277403 292246 277415
rect 247946 277375 292246 277403
rect 247946 277363 247952 277375
rect 292240 277363 292246 277375
rect 292298 277363 292304 277415
rect 298192 277363 298198 277415
rect 298250 277403 298256 277415
rect 425008 277403 425014 277415
rect 298250 277375 318110 277403
rect 298250 277363 298256 277375
rect 318082 277329 318110 277375
rect 318274 277375 425014 277403
rect 318274 277329 318302 277375
rect 425008 277363 425014 277375
rect 425066 277363 425072 277415
rect 318082 277301 318302 277329
rect 318448 277289 318454 277341
rect 318506 277329 318512 277341
rect 327376 277329 327382 277341
rect 318506 277301 327382 277329
rect 318506 277289 318512 277301
rect 327376 277289 327382 277301
rect 327434 277289 327440 277341
rect 327664 277289 327670 277341
rect 327722 277329 327728 277341
rect 460720 277329 460726 277341
rect 327722 277301 460726 277329
rect 327722 277289 327728 277301
rect 460720 277289 460726 277301
rect 460778 277289 460784 277341
rect 42064 277215 42070 277267
rect 42122 277255 42128 277267
rect 43120 277255 43126 277267
rect 42122 277227 43126 277255
rect 42122 277215 42128 277227
rect 43120 277215 43126 277227
rect 43178 277215 43184 277267
rect 240688 277215 240694 277267
rect 240746 277255 240752 277267
rect 290800 277255 290806 277267
rect 240746 277227 290806 277255
rect 240746 277215 240752 277227
rect 290800 277215 290806 277227
rect 290858 277215 290864 277267
rect 299056 277215 299062 277267
rect 299114 277255 299120 277267
rect 432208 277255 432214 277267
rect 299114 277227 432214 277255
rect 299114 277215 299120 277227
rect 432208 277215 432214 277227
rect 432266 277215 432272 277267
rect 300208 277141 300214 277193
rect 300266 277181 300272 277193
rect 439312 277181 439318 277193
rect 300266 277153 439318 277181
rect 300266 277141 300272 277153
rect 439312 277141 439318 277153
rect 439370 277141 439376 277193
rect 233488 277067 233494 277119
rect 233546 277107 233552 277119
rect 330160 277107 330166 277119
rect 233546 277079 330166 277107
rect 233546 277067 233552 277079
rect 330160 277067 330166 277079
rect 330218 277067 330224 277119
rect 349072 277067 349078 277119
rect 349130 277107 349136 277119
rect 386992 277107 386998 277119
rect 349130 277079 386998 277107
rect 349130 277067 349136 277079
rect 386992 277067 386998 277079
rect 387050 277067 387056 277119
rect 388432 277067 388438 277119
rect 388490 277107 388496 277119
rect 402448 277107 402454 277119
rect 388490 277079 402454 277107
rect 388490 277067 388496 277079
rect 402448 277067 402454 277079
rect 402506 277067 402512 277119
rect 225232 276993 225238 277045
rect 225290 277033 225296 277045
rect 273616 277033 273622 277045
rect 225290 277005 273622 277033
rect 225290 276993 225296 277005
rect 273616 276993 273622 277005
rect 273674 276993 273680 277045
rect 290800 276993 290806 277045
rect 290858 277033 290864 277045
rect 364432 277033 364438 277045
rect 290858 277005 364438 277033
rect 290858 276993 290864 277005
rect 364432 276993 364438 277005
rect 364490 276993 364496 277045
rect 364816 276993 364822 277045
rect 364874 277033 364880 277045
rect 364874 277005 376766 277033
rect 364874 276993 364880 277005
rect 300784 276919 300790 276971
rect 300842 276959 300848 276971
rect 376624 276959 376630 276971
rect 300842 276931 376630 276959
rect 300842 276919 300848 276931
rect 376624 276919 376630 276931
rect 376682 276919 376688 276971
rect 289264 276845 289270 276897
rect 289322 276885 289328 276897
rect 350032 276885 350038 276897
rect 289322 276857 350038 276885
rect 289322 276845 289328 276857
rect 350032 276845 350038 276857
rect 350090 276845 350096 276897
rect 365296 276845 365302 276897
rect 365354 276885 365360 276897
rect 370960 276885 370966 276897
rect 365354 276857 370966 276885
rect 365354 276845 365360 276857
rect 370960 276845 370966 276857
rect 371018 276845 371024 276897
rect 376738 276885 376766 277005
rect 377008 276993 377014 277045
rect 377066 277033 377072 277045
rect 378544 277033 378550 277045
rect 377066 277005 378550 277033
rect 377066 276993 377072 277005
rect 378544 276993 378550 277005
rect 378602 276993 378608 277045
rect 378640 276993 378646 277045
rect 378698 277033 378704 277045
rect 504688 277033 504694 277045
rect 378698 277005 504694 277033
rect 378698 276993 378704 277005
rect 504688 276993 504694 277005
rect 504746 276993 504752 277045
rect 376912 276919 376918 276971
rect 376970 276959 376976 276971
rect 446512 276959 446518 276971
rect 376970 276931 446518 276959
rect 376970 276919 376976 276931
rect 446512 276919 446518 276931
rect 446570 276919 446576 276971
rect 515440 276885 515446 276897
rect 376738 276857 515446 276885
rect 515440 276845 515446 276857
rect 515498 276845 515504 276897
rect 254896 276771 254902 276823
rect 254954 276811 254960 276823
rect 332752 276811 332758 276823
rect 254954 276783 332758 276811
rect 254954 276771 254960 276783
rect 332752 276771 332758 276783
rect 332810 276771 332816 276823
rect 348880 276771 348886 276823
rect 348938 276811 348944 276823
rect 383344 276811 383350 276823
rect 348938 276783 383350 276811
rect 348938 276771 348944 276783
rect 383344 276771 383350 276783
rect 383402 276771 383408 276823
rect 383728 276771 383734 276823
rect 383786 276811 383792 276823
rect 523792 276811 523798 276823
rect 383786 276783 523798 276811
rect 383786 276771 383792 276783
rect 523792 276771 523798 276783
rect 523850 276771 523856 276823
rect 639376 276771 639382 276823
rect 639434 276811 639440 276823
rect 649552 276811 649558 276823
rect 639434 276783 649558 276811
rect 639434 276771 639440 276783
rect 649552 276771 649558 276783
rect 649610 276771 649616 276823
rect 215728 276697 215734 276749
rect 215786 276737 215792 276749
rect 311824 276737 311830 276749
rect 215786 276709 311830 276737
rect 215786 276697 215792 276709
rect 311824 276697 311830 276709
rect 311882 276697 311888 276749
rect 311920 276697 311926 276749
rect 311978 276737 311984 276749
rect 338704 276737 338710 276749
rect 311978 276709 338710 276737
rect 311978 276697 311984 276709
rect 338704 276697 338710 276709
rect 338762 276697 338768 276749
rect 370960 276697 370966 276749
rect 371018 276737 371024 276749
rect 518992 276737 518998 276749
rect 371018 276709 518998 276737
rect 371018 276697 371024 276709
rect 518992 276697 518998 276709
rect 519050 276697 519056 276749
rect 208528 276623 208534 276675
rect 208586 276663 208592 276675
rect 309616 276663 309622 276675
rect 208586 276635 309622 276663
rect 208586 276623 208592 276635
rect 309616 276623 309622 276635
rect 309674 276623 309680 276675
rect 318160 276623 318166 276675
rect 318218 276663 318224 276675
rect 338320 276663 338326 276675
rect 318218 276635 338326 276663
rect 318218 276623 318224 276635
rect 338320 276623 338326 276635
rect 338378 276623 338384 276675
rect 363760 276623 363766 276675
rect 363818 276663 363824 276675
rect 368560 276663 368566 276675
rect 363818 276635 368566 276663
rect 363818 276623 363824 276635
rect 368560 276623 368566 276635
rect 368618 276623 368624 276675
rect 368752 276623 368758 276675
rect 368810 276663 368816 276675
rect 378640 276663 378646 276675
rect 368810 276635 378646 276663
rect 368810 276623 368816 276635
rect 378640 276623 378646 276635
rect 378698 276623 378704 276675
rect 378736 276623 378742 276675
rect 378794 276663 378800 276675
rect 611824 276663 611830 276675
rect 378794 276635 611830 276663
rect 378794 276623 378800 276635
rect 611824 276623 611830 276635
rect 611882 276623 611888 276675
rect 292240 276549 292246 276601
rect 292298 276589 292304 276601
rect 307984 276589 307990 276601
rect 292298 276561 307990 276589
rect 292298 276549 292304 276561
rect 307984 276549 307990 276561
rect 308042 276549 308048 276601
rect 318064 276549 318070 276601
rect 318122 276589 318128 276601
rect 332176 276589 332182 276601
rect 318122 276561 332182 276589
rect 318122 276549 318128 276561
rect 332176 276549 332182 276561
rect 332234 276549 332240 276601
rect 358576 276549 358582 276601
rect 358634 276589 358640 276601
rect 379120 276589 379126 276601
rect 358634 276561 379126 276589
rect 358634 276549 358640 276561
rect 379120 276549 379126 276561
rect 379178 276549 379184 276601
rect 379792 276549 379798 276601
rect 379850 276589 379856 276601
rect 636688 276589 636694 276601
rect 379850 276561 636694 276589
rect 379850 276549 379856 276561
rect 636688 276549 636694 276561
rect 636746 276549 636752 276601
rect 288400 276475 288406 276527
rect 288458 276515 288464 276527
rect 342928 276515 342934 276527
rect 288458 276487 342934 276515
rect 288458 276475 288464 276487
rect 342928 276475 342934 276487
rect 342986 276475 342992 276527
rect 351088 276475 351094 276527
rect 351146 276515 351152 276527
rect 401200 276515 401206 276527
rect 351146 276487 401206 276515
rect 351146 276475 351152 276487
rect 401200 276475 401206 276487
rect 401258 276475 401264 276527
rect 243760 276401 243766 276453
rect 243818 276441 243824 276453
rect 434512 276441 434518 276453
rect 243818 276413 434518 276441
rect 243818 276401 243824 276413
rect 434512 276401 434518 276413
rect 434570 276401 434576 276453
rect 231952 276327 231958 276379
rect 232010 276367 232016 276379
rect 338224 276367 338230 276379
rect 232010 276339 338230 276367
rect 232010 276327 232016 276339
rect 338224 276327 338230 276339
rect 338282 276327 338288 276379
rect 346768 276327 346774 276379
rect 346826 276367 346832 276379
rect 365584 276367 365590 276379
rect 346826 276339 365590 276367
rect 346826 276327 346832 276339
rect 365584 276327 365590 276339
rect 365642 276327 365648 276379
rect 370960 276327 370966 276379
rect 371018 276367 371024 276379
rect 375472 276367 375478 276379
rect 371018 276339 375478 276367
rect 371018 276327 371024 276339
rect 375472 276327 375478 276339
rect 375530 276327 375536 276379
rect 375568 276327 375574 276379
rect 375626 276367 375632 276379
rect 380464 276367 380470 276379
rect 375626 276339 380470 276367
rect 375626 276327 375632 276339
rect 380464 276327 380470 276339
rect 380522 276327 380528 276379
rect 380560 276327 380566 276379
rect 380618 276367 380624 276379
rect 380618 276339 385022 276367
rect 380618 276327 380624 276339
rect 232336 276253 232342 276305
rect 232394 276293 232400 276305
rect 341776 276293 341782 276305
rect 232394 276265 341782 276293
rect 232394 276253 232400 276265
rect 341776 276253 341782 276265
rect 341834 276253 341840 276305
rect 348400 276253 348406 276305
rect 348458 276293 348464 276305
rect 379504 276293 379510 276305
rect 348458 276265 379510 276293
rect 348458 276253 348464 276265
rect 379504 276253 379510 276265
rect 379562 276253 379568 276305
rect 379984 276253 379990 276305
rect 380042 276293 380048 276305
rect 384880 276293 384886 276305
rect 380042 276265 384886 276293
rect 380042 276253 380048 276265
rect 384880 276253 384886 276265
rect 384938 276253 384944 276305
rect 384994 276293 385022 276339
rect 385072 276327 385078 276379
rect 385130 276367 385136 276379
rect 565456 276367 565462 276379
rect 385130 276339 565462 276367
rect 385130 276327 385136 276339
rect 565456 276327 565462 276339
rect 565514 276327 565520 276379
rect 572464 276293 572470 276305
rect 384994 276265 572470 276293
rect 572464 276253 572470 276265
rect 572522 276253 572528 276305
rect 244720 276179 244726 276231
rect 244778 276219 244784 276231
rect 441712 276219 441718 276231
rect 244778 276191 441718 276219
rect 244778 276179 244784 276191
rect 441712 276179 441718 276191
rect 441770 276179 441776 276231
rect 245392 276105 245398 276157
rect 245450 276145 245456 276157
rect 448816 276145 448822 276157
rect 245450 276117 448822 276145
rect 245450 276105 245456 276117
rect 448816 276105 448822 276117
rect 448874 276105 448880 276157
rect 246352 276031 246358 276083
rect 246410 276071 246416 276083
rect 455920 276071 455926 276083
rect 246410 276043 455926 276071
rect 246410 276031 246416 276043
rect 455920 276031 455926 276043
rect 455978 276031 455984 276083
rect 233488 275957 233494 276009
rect 233546 275997 233552 276009
rect 348976 275997 348982 276009
rect 233546 275969 348982 275997
rect 233546 275957 233552 275969
rect 348976 275957 348982 275969
rect 349034 275957 349040 276009
rect 370384 275957 370390 276009
rect 370442 275997 370448 276009
rect 384784 275997 384790 276009
rect 370442 275969 384790 275997
rect 370442 275957 370448 275969
rect 384784 275957 384790 275969
rect 384842 275957 384848 276009
rect 384880 275957 384886 276009
rect 384938 275997 384944 276009
rect 579664 275997 579670 276009
rect 384938 275969 579670 275997
rect 384938 275957 384944 275969
rect 579664 275957 579670 275969
rect 579722 275957 579728 276009
rect 247408 275883 247414 275935
rect 247466 275923 247472 275935
rect 463120 275923 463126 275935
rect 247466 275895 463126 275923
rect 247466 275883 247472 275895
rect 463120 275883 463126 275895
rect 463178 275883 463184 275935
rect 227440 275809 227446 275861
rect 227498 275849 227504 275861
rect 298960 275849 298966 275861
rect 227498 275821 298966 275849
rect 227498 275809 227504 275821
rect 298960 275809 298966 275821
rect 299018 275809 299024 275861
rect 311536 275809 311542 275861
rect 311594 275849 311600 275861
rect 532144 275849 532150 275861
rect 311594 275821 532150 275849
rect 311594 275809 311600 275821
rect 532144 275809 532150 275821
rect 532202 275809 532208 275861
rect 248080 275735 248086 275787
rect 248138 275775 248144 275787
rect 470224 275775 470230 275787
rect 248138 275747 470230 275775
rect 248138 275735 248144 275747
rect 470224 275735 470230 275747
rect 470282 275735 470288 275787
rect 234064 275661 234070 275713
rect 234122 275701 234128 275713
rect 356080 275701 356086 275713
rect 234122 275673 356086 275701
rect 234122 275661 234128 275673
rect 356080 275661 356086 275673
rect 356138 275661 356144 275713
rect 364240 275661 364246 275713
rect 364298 275701 364304 275713
rect 380272 275701 380278 275713
rect 364298 275673 380278 275701
rect 364298 275661 364304 275673
rect 380272 275661 380278 275673
rect 380330 275661 380336 275713
rect 380464 275661 380470 275713
rect 380522 275701 380528 275713
rect 601072 275701 601078 275713
rect 380522 275673 601078 275701
rect 380522 275661 380528 275673
rect 601072 275661 601078 275673
rect 601130 275661 601136 275713
rect 249136 275587 249142 275639
rect 249194 275627 249200 275639
rect 477424 275627 477430 275639
rect 249194 275599 477430 275627
rect 249194 275587 249200 275599
rect 477424 275587 477430 275599
rect 477482 275587 477488 275639
rect 249808 275513 249814 275565
rect 249866 275553 249872 275565
rect 484432 275553 484438 275565
rect 249866 275525 484438 275553
rect 249866 275513 249872 275525
rect 484432 275513 484438 275525
rect 484490 275513 484496 275565
rect 200176 275439 200182 275491
rect 200234 275479 200240 275491
rect 270736 275479 270742 275491
rect 200234 275451 270742 275479
rect 200234 275439 200240 275451
rect 270736 275439 270742 275451
rect 270794 275439 270800 275491
rect 323248 275439 323254 275491
rect 323306 275479 323312 275491
rect 564208 275479 564214 275491
rect 323306 275451 564214 275479
rect 323306 275439 323312 275451
rect 564208 275439 564214 275451
rect 564266 275439 564272 275491
rect 235024 275365 235030 275417
rect 235082 275405 235088 275417
rect 363184 275405 363190 275417
rect 235082 275377 363190 275405
rect 235082 275365 235088 275377
rect 363184 275365 363190 275377
rect 363242 275365 363248 275417
rect 371824 275365 371830 275417
rect 371882 275405 371888 275417
rect 371882 275377 377726 275405
rect 371882 275365 371888 275377
rect 235984 275291 235990 275343
rect 236042 275331 236048 275343
rect 370288 275331 370294 275343
rect 236042 275303 370294 275331
rect 236042 275291 236048 275303
rect 370288 275291 370294 275303
rect 370346 275291 370352 275343
rect 372880 275291 372886 275343
rect 372938 275331 372944 275343
rect 377584 275331 377590 275343
rect 372938 275303 377590 275331
rect 372938 275291 372944 275303
rect 377584 275291 377590 275303
rect 377642 275291 377648 275343
rect 377698 275331 377726 275377
rect 377872 275365 377878 275417
rect 377930 275405 377936 275417
rect 622480 275405 622486 275417
rect 377930 275377 622486 275405
rect 377930 275365 377936 275377
rect 622480 275365 622486 275377
rect 622538 275365 622544 275417
rect 379408 275331 379414 275343
rect 377698 275303 379414 275331
rect 379408 275291 379414 275303
rect 379466 275291 379472 275343
rect 379504 275291 379510 275343
rect 379562 275331 379568 275343
rect 633136 275331 633142 275343
rect 379562 275303 633142 275331
rect 379562 275291 379568 275303
rect 633136 275291 633142 275303
rect 633194 275291 633200 275343
rect 196720 275217 196726 275269
rect 196778 275257 196784 275269
rect 270544 275257 270550 275269
rect 196778 275229 270550 275257
rect 196778 275217 196784 275229
rect 270544 275217 270550 275229
rect 270602 275217 270608 275269
rect 284944 275217 284950 275269
rect 285002 275257 285008 275269
rect 314416 275257 314422 275269
rect 285002 275229 314422 275257
rect 285002 275217 285008 275229
rect 314416 275217 314422 275229
rect 314474 275217 314480 275269
rect 316048 275217 316054 275269
rect 316106 275257 316112 275269
rect 571312 275257 571318 275269
rect 316106 275229 571318 275257
rect 316106 275217 316112 275229
rect 571312 275217 571318 275229
rect 571370 275217 571376 275269
rect 228016 275143 228022 275195
rect 228074 275183 228080 275195
rect 306064 275183 306070 275195
rect 228074 275155 306070 275183
rect 228074 275143 228080 275155
rect 306064 275143 306070 275155
rect 306122 275143 306128 275195
rect 317296 275143 317302 275195
rect 317354 275183 317360 275195
rect 578512 275183 578518 275195
rect 317354 275155 578518 275183
rect 317354 275143 317360 275155
rect 578512 275143 578518 275155
rect 578570 275143 578576 275195
rect 236752 275069 236758 275121
rect 236810 275109 236816 275121
rect 377488 275109 377494 275121
rect 236810 275081 377494 275109
rect 236810 275069 236816 275081
rect 377488 275069 377494 275081
rect 377546 275069 377552 275121
rect 377584 275069 377590 275121
rect 377642 275109 377648 275121
rect 379984 275109 379990 275121
rect 377642 275081 379990 275109
rect 377642 275069 377648 275081
rect 379984 275069 379990 275081
rect 380042 275069 380048 275121
rect 380080 275069 380086 275121
rect 380138 275109 380144 275121
rect 380560 275109 380566 275121
rect 380138 275081 380566 275109
rect 380138 275069 380144 275081
rect 380560 275069 380566 275081
rect 380618 275069 380624 275121
rect 381424 275069 381430 275121
rect 381482 275109 381488 275121
rect 647536 275109 647542 275121
rect 381482 275081 647542 275109
rect 381482 275069 381488 275081
rect 647536 275069 647542 275081
rect 647594 275069 647600 275121
rect 229072 274995 229078 275047
rect 229130 275035 229136 275047
rect 313264 275035 313270 275047
rect 229130 275007 313270 275035
rect 229130 274995 229136 275007
rect 313264 274995 313270 275007
rect 313322 274995 313328 275047
rect 318064 274995 318070 275047
rect 318122 275035 318128 275047
rect 585616 275035 585622 275047
rect 318122 275007 585622 275035
rect 318122 274995 318128 275007
rect 585616 274995 585622 275007
rect 585674 274995 585680 275047
rect 258544 274921 258550 274973
rect 258602 274961 258608 274973
rect 333136 274961 333142 274973
rect 258602 274933 333142 274961
rect 258602 274921 258608 274933
rect 333136 274921 333142 274933
rect 333194 274921 333200 274973
rect 368080 274921 368086 274973
rect 368138 274961 368144 274973
rect 378640 274961 378646 274973
rect 368138 274933 378646 274961
rect 368138 274921 368144 274933
rect 378640 274921 378646 274933
rect 378698 274921 378704 274973
rect 378736 274921 378742 274973
rect 378794 274961 378800 274973
rect 384688 274961 384694 274973
rect 378794 274933 384694 274961
rect 378794 274921 378800 274933
rect 384688 274921 384694 274933
rect 384746 274921 384752 274973
rect 384784 274921 384790 274973
rect 384842 274961 384848 274973
rect 558256 274961 558262 274973
rect 384842 274933 558262 274961
rect 384842 274921 384848 274933
rect 558256 274921 558262 274933
rect 558314 274921 558320 274973
rect 242992 274847 242998 274899
rect 243050 274887 243056 274899
rect 427408 274887 427414 274899
rect 243050 274859 427414 274887
rect 243050 274847 243056 274859
rect 427408 274847 427414 274859
rect 427466 274847 427472 274899
rect 223024 274773 223030 274825
rect 223082 274813 223088 274825
rect 263344 274813 263350 274825
rect 223082 274785 263350 274813
rect 223082 274773 223088 274785
rect 263344 274773 263350 274785
rect 263402 274773 263408 274825
rect 269200 274773 269206 274825
rect 269258 274813 269264 274825
rect 334480 274813 334486 274825
rect 269258 274785 334486 274813
rect 269258 274773 269264 274785
rect 334480 274773 334486 274785
rect 334538 274773 334544 274825
rect 372304 274773 372310 274825
rect 372362 274813 372368 274825
rect 384592 274813 384598 274825
rect 372362 274785 384598 274813
rect 372362 274773 372368 274785
rect 384592 274773 384598 274785
rect 384650 274773 384656 274825
rect 384688 274773 384694 274825
rect 384746 274813 384752 274825
rect 551056 274813 551062 274825
rect 384746 274785 551062 274813
rect 384746 274773 384752 274785
rect 551056 274773 551062 274785
rect 551114 274773 551120 274825
rect 242224 274699 242230 274751
rect 242282 274739 242288 274751
rect 420208 274739 420214 274751
rect 242282 274711 420214 274739
rect 242282 274699 242288 274711
rect 420208 274699 420214 274711
rect 420266 274699 420272 274751
rect 226288 274625 226294 274677
rect 226346 274665 226352 274677
rect 291856 274665 291862 274677
rect 226346 274637 291862 274665
rect 226346 274625 226352 274637
rect 291856 274625 291862 274637
rect 291914 274625 291920 274677
rect 297808 274625 297814 274677
rect 297866 274665 297872 274677
rect 337936 274665 337942 274677
rect 297866 274637 337942 274665
rect 297866 274625 297872 274637
rect 337936 274625 337942 274637
rect 337994 274625 338000 274677
rect 369520 274625 369526 274677
rect 369578 274665 369584 274677
rect 378544 274665 378550 274677
rect 369578 274637 378550 274665
rect 369578 274625 369584 274637
rect 378544 274625 378550 274637
rect 378602 274625 378608 274677
rect 378640 274625 378646 274677
rect 378698 274665 378704 274677
rect 540400 274665 540406 274677
rect 378698 274637 540406 274665
rect 378698 274625 378704 274637
rect 540400 274625 540406 274637
rect 540458 274625 540464 274677
rect 240496 274551 240502 274603
rect 240554 274591 240560 274603
rect 406000 274591 406006 274603
rect 240554 274563 406006 274591
rect 240554 274551 240560 274563
rect 406000 274551 406006 274563
rect 406058 274551 406064 274603
rect 239344 274477 239350 274529
rect 239402 274517 239408 274529
rect 398896 274517 398902 274529
rect 239402 274489 398902 274517
rect 239402 274477 239408 274489
rect 398896 274477 398902 274489
rect 398954 274477 398960 274529
rect 238480 274403 238486 274455
rect 238538 274443 238544 274455
rect 391696 274443 391702 274455
rect 238538 274415 391702 274443
rect 238538 274403 238544 274415
rect 391696 274403 391702 274415
rect 391754 274403 391760 274455
rect 237808 274329 237814 274381
rect 237866 274369 237872 274381
rect 372304 274369 372310 274381
rect 237866 274341 372310 274369
rect 237866 274329 237872 274341
rect 372304 274329 372310 274341
rect 372362 274329 372368 274381
rect 378736 274369 378742 274381
rect 372418 274341 378742 274369
rect 42160 274255 42166 274307
rect 42218 274295 42224 274307
rect 43024 274295 43030 274307
rect 42218 274267 43030 274295
rect 42218 274255 42224 274267
rect 43024 274255 43030 274267
rect 43082 274255 43088 274307
rect 207376 274255 207382 274307
rect 207434 274295 207440 274307
rect 271312 274295 271318 274307
rect 207434 274267 271318 274295
rect 207434 274255 207440 274267
rect 271312 274255 271318 274267
rect 271370 274255 271376 274307
rect 271408 274255 271414 274307
rect 271466 274295 271472 274307
rect 271466 274267 272606 274295
rect 271466 274255 271472 274267
rect 214576 274181 214582 274233
rect 214634 274221 214640 274233
rect 272464 274221 272470 274233
rect 214634 274193 272470 274221
rect 214634 274181 214640 274193
rect 272464 274181 272470 274193
rect 272522 274181 272528 274233
rect 272578 274221 272606 274267
rect 276400 274255 276406 274307
rect 276458 274295 276464 274307
rect 335632 274295 335638 274307
rect 276458 274267 335638 274295
rect 276458 274255 276464 274267
rect 335632 274255 335638 274267
rect 335690 274255 335696 274307
rect 358768 274255 358774 274307
rect 358826 274295 358832 274307
rect 372418 274295 372446 274341
rect 378736 274329 378742 274341
rect 378794 274329 378800 274381
rect 378832 274329 378838 274381
rect 378890 274369 378896 274381
rect 385552 274369 385558 274381
rect 378890 274341 385558 274369
rect 378890 274329 378896 274341
rect 385552 274329 385558 274341
rect 385610 274329 385616 274381
rect 385840 274329 385846 274381
rect 385898 274369 385904 274381
rect 395344 274369 395350 274381
rect 385898 274341 395350 274369
rect 385898 274329 385904 274341
rect 395344 274329 395350 274341
rect 395402 274329 395408 274381
rect 511888 274295 511894 274307
rect 358826 274267 372446 274295
rect 372514 274267 511894 274295
rect 358826 274255 358832 274267
rect 272578 274193 284894 274221
rect 225424 274107 225430 274159
rect 225482 274147 225488 274159
rect 284656 274147 284662 274159
rect 225482 274119 284662 274147
rect 225482 274107 225488 274119
rect 284656 274107 284662 274119
rect 284714 274107 284720 274159
rect 225232 274033 225238 274085
rect 225290 274073 225296 274085
rect 281104 274073 281110 274085
rect 225290 274045 281110 274073
rect 225290 274033 225296 274045
rect 281104 274033 281110 274045
rect 281162 274033 281168 274085
rect 239440 273959 239446 274011
rect 239498 273999 239504 274011
rect 275248 273999 275254 274011
rect 239498 273971 275254 273999
rect 239498 273959 239504 273971
rect 275248 273959 275254 273971
rect 275306 273959 275312 274011
rect 284866 273999 284894 274193
rect 287056 274181 287062 274233
rect 287114 274221 287120 274233
rect 337552 274221 337558 274233
rect 287114 274193 337558 274221
rect 287114 274181 287120 274193
rect 337552 274181 337558 274193
rect 337610 274181 337616 274233
rect 352240 274181 352246 274233
rect 352298 274221 352304 274233
rect 372400 274221 372406 274233
rect 352298 274193 372406 274221
rect 352298 274181 352304 274193
rect 372400 274181 372406 274193
rect 372458 274181 372464 274233
rect 286768 274107 286774 274159
rect 286826 274147 286832 274159
rect 328720 274147 328726 274159
rect 286826 274119 328726 274147
rect 286826 274107 286832 274119
rect 328720 274107 328726 274119
rect 328778 274107 328784 274159
rect 364336 274107 364342 274159
rect 364394 274147 364400 274159
rect 372514 274147 372542 274267
rect 511888 274255 511894 274267
rect 511946 274255 511952 274307
rect 374128 274181 374134 274233
rect 374186 274221 374192 274233
rect 378448 274221 378454 274233
rect 374186 274193 378454 274221
rect 374186 274181 374192 274193
rect 378448 274181 378454 274193
rect 378506 274181 378512 274233
rect 378544 274181 378550 274233
rect 378602 274221 378608 274233
rect 380176 274221 380182 274233
rect 378602 274193 380182 274221
rect 378602 274181 378608 274193
rect 380176 274181 380182 274193
rect 380234 274181 380240 274233
rect 380272 274181 380278 274233
rect 380330 274221 380336 274233
rect 508336 274221 508342 274233
rect 380330 274193 508342 274221
rect 380330 274181 380336 274193
rect 508336 274181 508342 274193
rect 508394 274181 508400 274233
rect 364394 274119 372542 274147
rect 364394 274107 364400 274119
rect 374320 274107 374326 274159
rect 374378 274147 374384 274159
rect 374378 274119 378782 274147
rect 374378 274107 374384 274119
rect 296656 274033 296662 274085
rect 296714 274073 296720 274085
rect 297136 274073 297142 274085
rect 296714 274045 297142 274073
rect 296714 274033 296720 274045
rect 297136 274033 297142 274045
rect 297194 274033 297200 274085
rect 304912 274033 304918 274085
rect 304970 274073 304976 274085
rect 338896 274073 338902 274085
rect 304970 274045 338902 274073
rect 304970 274033 304976 274045
rect 338896 274033 338902 274045
rect 338954 274033 338960 274085
rect 360496 274033 360502 274085
rect 360554 274073 360560 274085
rect 378640 274073 378646 274085
rect 360554 274045 378646 274073
rect 360554 274033 360560 274045
rect 378640 274033 378646 274045
rect 378698 274033 378704 274085
rect 378754 274073 378782 274119
rect 378832 274107 378838 274159
rect 378890 274147 378896 274159
rect 479728 274147 479734 274159
rect 378890 274119 479734 274147
rect 378890 274107 378896 274119
rect 479728 274107 479734 274119
rect 479786 274107 479792 274159
rect 385744 274073 385750 274085
rect 378754 274045 385750 274073
rect 385744 274033 385750 274045
rect 385802 274033 385808 274085
rect 388912 274033 388918 274085
rect 388970 274073 388976 274085
rect 476176 274073 476182 274085
rect 388970 274045 476182 274073
rect 388970 274033 388976 274045
rect 476176 274033 476182 274045
rect 476234 274033 476240 274085
rect 378544 273999 378550 274011
rect 284866 273971 378550 273999
rect 378544 273959 378550 273971
rect 378602 273959 378608 274011
rect 383056 273999 383062 274011
rect 378658 273971 383062 273999
rect 232432 273885 232438 273937
rect 232490 273925 232496 273937
rect 274672 273925 274678 273937
rect 232490 273897 274678 273925
rect 232490 273885 232496 273897
rect 274672 273885 274678 273897
rect 274730 273885 274736 273937
rect 308848 273885 308854 273937
rect 308906 273925 308912 273937
rect 308906 273897 322718 273925
rect 308906 273885 308912 273897
rect 230608 273811 230614 273863
rect 230666 273851 230672 273863
rect 319696 273851 319702 273863
rect 230666 273823 319702 273851
rect 230666 273811 230672 273823
rect 319696 273811 319702 273823
rect 319754 273811 319760 273863
rect 229744 273737 229750 273789
rect 229802 273777 229808 273789
rect 320080 273777 320086 273789
rect 229802 273749 320086 273777
rect 229802 273737 229808 273749
rect 320080 273737 320086 273749
rect 320138 273737 320144 273789
rect 322690 273777 322718 273897
rect 322768 273885 322774 273937
rect 322826 273925 322832 273937
rect 341296 273925 341302 273937
rect 322826 273897 341302 273925
rect 322826 273885 322832 273897
rect 341296 273885 341302 273897
rect 341354 273885 341360 273937
rect 360016 273885 360022 273937
rect 360074 273925 360080 273937
rect 378658 273925 378686 273971
rect 383056 273959 383062 273971
rect 383114 273959 383120 274011
rect 360074 273897 378686 273925
rect 360074 273885 360080 273897
rect 378736 273885 378742 273937
rect 378794 273925 378800 273937
rect 461968 273925 461974 273937
rect 378794 273897 461974 273925
rect 378794 273885 378800 273897
rect 461968 273885 461974 273897
rect 462026 273885 462032 273937
rect 325264 273811 325270 273863
rect 325322 273851 325328 273863
rect 325936 273851 325942 273863
rect 325322 273823 325942 273851
rect 325322 273811 325328 273823
rect 325936 273811 325942 273823
rect 325994 273811 326000 273863
rect 356176 273811 356182 273863
rect 356234 273851 356240 273863
rect 444112 273851 444118 273863
rect 356234 273823 444118 273851
rect 356234 273811 356240 273823
rect 444112 273811 444118 273823
rect 444170 273811 444176 273863
rect 377488 273777 377494 273789
rect 322690 273749 377494 273777
rect 377488 273737 377494 273749
rect 377546 273737 377552 273789
rect 377584 273737 377590 273789
rect 377642 273777 377648 273789
rect 392944 273777 392950 273789
rect 377642 273749 392950 273777
rect 377642 273737 377648 273749
rect 392944 273737 392950 273749
rect 393002 273737 393008 273789
rect 231760 273663 231766 273715
rect 231818 273703 231824 273715
rect 325456 273703 325462 273715
rect 231818 273675 325462 273703
rect 231818 273663 231824 273675
rect 325456 273663 325462 273675
rect 325514 273663 325520 273715
rect 325648 273663 325654 273715
rect 325706 273703 325712 273715
rect 327664 273703 327670 273715
rect 325706 273675 327670 273703
rect 325706 273663 325712 273675
rect 327664 273663 327670 273675
rect 327722 273663 327728 273715
rect 354448 273663 354454 273715
rect 354506 273703 354512 273715
rect 429808 273703 429814 273715
rect 354506 273675 429814 273703
rect 354506 273663 354512 273675
rect 429808 273663 429814 273675
rect 429866 273663 429872 273715
rect 66640 273589 66646 273641
rect 66698 273629 66704 273641
rect 66698 273601 69182 273629
rect 66698 273589 66704 273601
rect 69154 273555 69182 273601
rect 236272 273589 236278 273641
rect 236330 273629 236336 273641
rect 245488 273629 245494 273641
rect 236330 273601 245494 273629
rect 236330 273589 236336 273601
rect 245488 273589 245494 273601
rect 245546 273589 245552 273641
rect 262672 273589 262678 273641
rect 262730 273629 262736 273641
rect 262730 273601 372350 273629
rect 262730 273589 262736 273601
rect 79216 273555 79222 273567
rect 69154 273527 79222 273555
rect 79216 273515 79222 273527
rect 79274 273515 79280 273567
rect 106288 273515 106294 273567
rect 106346 273555 106352 273567
rect 198736 273555 198742 273567
rect 106346 273527 198742 273555
rect 106346 273515 106352 273527
rect 198736 273515 198742 273527
rect 198794 273515 198800 273567
rect 212368 273555 212374 273567
rect 198850 273527 212374 273555
rect 91984 273441 91990 273493
rect 92042 273481 92048 273493
rect 190576 273481 190582 273493
rect 92042 273453 190582 273481
rect 92042 273441 92048 273453
rect 190576 273441 190582 273453
rect 190634 273441 190640 273493
rect 190672 273441 190678 273493
rect 190730 273481 190736 273493
rect 198850 273481 198878 273527
rect 212368 273515 212374 273527
rect 212426 273515 212432 273567
rect 227536 273515 227542 273567
rect 227594 273555 227600 273567
rect 247600 273555 247606 273567
rect 227594 273527 247606 273555
rect 227594 273515 227600 273527
rect 247600 273515 247606 273527
rect 247658 273515 247664 273567
rect 262384 273515 262390 273567
rect 262442 273555 262448 273567
rect 270352 273555 270358 273567
rect 262442 273527 270358 273555
rect 262442 273515 262448 273527
rect 270352 273515 270358 273527
rect 270410 273515 270416 273567
rect 270448 273515 270454 273567
rect 270506 273555 270512 273567
rect 271408 273555 271414 273567
rect 270506 273527 271414 273555
rect 270506 273515 270512 273527
rect 271408 273515 271414 273527
rect 271466 273515 271472 273567
rect 271600 273515 271606 273567
rect 271658 273555 271664 273567
rect 279472 273555 279478 273567
rect 271658 273527 279478 273555
rect 271658 273515 271664 273527
rect 279472 273515 279478 273527
rect 279530 273515 279536 273567
rect 284464 273515 284470 273567
rect 284522 273555 284528 273567
rect 284522 273527 285950 273555
rect 284522 273515 284528 273527
rect 190730 273453 198878 273481
rect 190730 273441 190736 273453
rect 224080 273441 224086 273493
rect 224138 273481 224144 273493
rect 274000 273481 274006 273493
rect 224138 273453 274006 273481
rect 224138 273441 224144 273453
rect 274000 273441 274006 273453
rect 274058 273441 274064 273493
rect 275152 273441 275158 273493
rect 275210 273481 275216 273493
rect 279664 273481 279670 273493
rect 275210 273453 279670 273481
rect 275210 273441 275216 273453
rect 279664 273441 279670 273453
rect 279722 273441 279728 273493
rect 281200 273441 281206 273493
rect 281258 273481 281264 273493
rect 285808 273481 285814 273493
rect 281258 273453 285814 273481
rect 281258 273441 281264 273453
rect 285808 273441 285814 273453
rect 285866 273441 285872 273493
rect 285922 273481 285950 273527
rect 290896 273515 290902 273567
rect 290954 273555 290960 273567
rect 293008 273555 293014 273567
rect 290954 273527 293014 273555
rect 290954 273515 290960 273527
rect 293008 273515 293014 273527
rect 293066 273515 293072 273567
rect 294736 273515 294742 273567
rect 294794 273555 294800 273567
rect 309040 273555 309046 273567
rect 294794 273527 309046 273555
rect 294794 273515 294800 273527
rect 309040 273515 309046 273527
rect 309098 273515 309104 273567
rect 319792 273515 319798 273567
rect 319850 273555 319856 273567
rect 321520 273555 321526 273567
rect 319850 273527 321526 273555
rect 319850 273515 319856 273527
rect 321520 273515 321526 273527
rect 321578 273515 321584 273567
rect 325456 273515 325462 273567
rect 325514 273555 325520 273567
rect 334576 273555 334582 273567
rect 325514 273527 334582 273555
rect 325514 273515 325520 273527
rect 334576 273515 334582 273527
rect 334634 273515 334640 273567
rect 340624 273515 340630 273567
rect 340682 273555 340688 273567
rect 343504 273555 343510 273567
rect 340682 273527 343510 273555
rect 340682 273515 340688 273527
rect 343504 273515 343510 273527
rect 343562 273515 343568 273567
rect 344656 273515 344662 273567
rect 344714 273555 344720 273567
rect 347728 273555 347734 273567
rect 344714 273527 347734 273555
rect 344714 273515 344720 273527
rect 347728 273515 347734 273527
rect 347786 273515 347792 273567
rect 356944 273515 356950 273567
rect 357002 273555 357008 273567
rect 367888 273555 367894 273567
rect 357002 273527 367894 273555
rect 357002 273515 357008 273527
rect 367888 273515 367894 273527
rect 367946 273515 367952 273567
rect 372322 273555 372350 273601
rect 372400 273589 372406 273641
rect 372458 273629 372464 273641
rect 411952 273629 411958 273641
rect 372458 273601 411958 273629
rect 372458 273589 372464 273601
rect 411952 273589 411958 273601
rect 412010 273589 412016 273641
rect 630736 273589 630742 273641
rect 630794 273629 630800 273641
rect 639376 273629 639382 273641
rect 630794 273601 639382 273629
rect 630794 273589 630800 273601
rect 639376 273589 639382 273601
rect 639434 273589 639440 273641
rect 649456 273629 649462 273641
rect 645154 273601 649462 273629
rect 380272 273555 380278 273567
rect 372322 273527 380278 273555
rect 380272 273515 380278 273527
rect 380330 273515 380336 273567
rect 380368 273515 380374 273567
rect 380426 273555 380432 273567
rect 396208 273555 396214 273567
rect 380426 273527 396214 273555
rect 380426 273515 380432 273527
rect 396208 273515 396214 273527
rect 396266 273515 396272 273567
rect 396304 273515 396310 273567
rect 396362 273555 396368 273567
rect 612976 273555 612982 273567
rect 396362 273527 612982 273555
rect 396362 273515 396368 273527
rect 612976 273515 612982 273527
rect 613034 273515 613040 273567
rect 642256 273515 642262 273567
rect 642314 273555 642320 273567
rect 645154 273555 645182 273601
rect 649456 273589 649462 273601
rect 649514 273589 649520 273641
rect 642314 273527 645182 273555
rect 642314 273515 642320 273527
rect 310864 273481 310870 273493
rect 285922 273453 310870 273481
rect 310864 273441 310870 273453
rect 310922 273441 310928 273493
rect 319696 273441 319702 273493
rect 319754 273481 319760 273493
rect 327472 273481 327478 273493
rect 319754 273453 327478 273481
rect 319754 273441 319760 273453
rect 327472 273441 327478 273453
rect 327530 273441 327536 273493
rect 327568 273441 327574 273493
rect 327626 273481 327632 273493
rect 557008 273481 557014 273493
rect 327626 273453 557014 273481
rect 327626 273441 327632 273453
rect 557008 273441 557014 273453
rect 557066 273441 557072 273493
rect 153808 273367 153814 273419
rect 153866 273407 153872 273419
rect 160912 273407 160918 273419
rect 153866 273379 160918 273407
rect 153866 273367 153872 273379
rect 160912 273367 160918 273379
rect 160970 273367 160976 273419
rect 161008 273367 161014 273419
rect 161066 273407 161072 273419
rect 404944 273407 404950 273419
rect 161066 273379 404950 273407
rect 161066 273367 161072 273379
rect 404944 273367 404950 273379
rect 405002 273367 405008 273419
rect 157456 273293 157462 273345
rect 157514 273333 157520 273345
rect 404080 273333 404086 273345
rect 157514 273305 404086 273333
rect 157514 273293 157520 273305
rect 404080 273293 404086 273305
rect 404138 273293 404144 273345
rect 161296 273219 161302 273271
rect 161354 273259 161360 273271
rect 161354 273231 164222 273259
rect 161354 273219 161360 273231
rect 147952 273145 147958 273197
rect 148010 273185 148016 273197
rect 149680 273185 149686 273197
rect 148010 273157 149686 273185
rect 148010 273145 148016 273157
rect 149680 273145 149686 273157
rect 149738 273145 149744 273197
rect 151408 273145 151414 273197
rect 151466 273185 151472 273197
rect 152560 273185 152566 273197
rect 151466 273157 152566 273185
rect 151466 273145 151472 273157
rect 152560 273145 152566 273157
rect 152618 273145 152624 273197
rect 152656 273145 152662 273197
rect 152714 273185 152720 273197
rect 155344 273185 155350 273197
rect 152714 273157 155350 273185
rect 152714 273145 152720 273157
rect 155344 273145 155350 273157
rect 155402 273145 155408 273197
rect 156208 273145 156214 273197
rect 156266 273185 156272 273197
rect 158320 273185 158326 273197
rect 156266 273157 158326 273185
rect 156266 273145 156272 273157
rect 158320 273145 158326 273157
rect 158378 273145 158384 273197
rect 162160 273145 162166 273197
rect 162218 273185 162224 273197
rect 164080 273185 164086 273197
rect 162218 273157 164086 273185
rect 162218 273145 162224 273157
rect 164080 273145 164086 273157
rect 164138 273145 164144 273197
rect 164194 273185 164222 273231
rect 164272 273219 164278 273271
rect 164330 273259 164336 273271
rect 371536 273259 371542 273271
rect 164330 273231 371542 273259
rect 164330 273219 164336 273231
rect 371536 273219 371542 273231
rect 371594 273219 371600 273271
rect 374320 273219 374326 273271
rect 374378 273259 374384 273271
rect 401296 273259 401302 273271
rect 374378 273231 401302 273259
rect 374378 273219 374384 273231
rect 401296 273219 401302 273231
rect 401354 273219 401360 273271
rect 403216 273185 403222 273197
rect 164194 273157 403222 273185
rect 403216 273145 403222 273157
rect 403274 273145 403280 273197
rect 139600 273071 139606 273123
rect 139658 273111 139664 273123
rect 139658 273083 144062 273111
rect 139658 273071 139664 273083
rect 142000 272997 142006 273049
rect 142058 273037 142064 273049
rect 143920 273037 143926 273049
rect 142058 273009 143926 273037
rect 142058 272997 142064 273009
rect 143920 272997 143926 273009
rect 143978 272997 143984 273049
rect 144034 273037 144062 273083
rect 146704 273071 146710 273123
rect 146762 273111 146768 273123
rect 373840 273111 373846 273123
rect 146762 273083 373846 273111
rect 146762 273071 146768 273083
rect 373840 273071 373846 273083
rect 373898 273071 373904 273123
rect 374608 273071 374614 273123
rect 374666 273111 374672 273123
rect 400624 273111 400630 273123
rect 374666 273083 400630 273111
rect 374666 273071 374672 273083
rect 400624 273071 400630 273083
rect 400682 273071 400688 273123
rect 399664 273037 399670 273049
rect 144034 273009 399670 273037
rect 399664 272997 399670 273009
rect 399722 272997 399728 273049
rect 143152 272923 143158 272975
rect 143210 272963 143216 272975
rect 374416 272963 374422 272975
rect 143210 272935 374422 272963
rect 143210 272923 143216 272935
rect 374416 272923 374422 272935
rect 374474 272923 374480 272975
rect 396976 272963 396982 272975
rect 374530 272935 396982 272963
rect 65872 272849 65878 272901
rect 65930 272889 65936 272901
rect 190672 272889 190678 272901
rect 65930 272861 190678 272889
rect 65930 272849 65936 272861
rect 190672 272849 190678 272861
rect 190730 272849 190736 272901
rect 190768 272849 190774 272901
rect 190826 272889 190832 272901
rect 192880 272889 192886 272901
rect 190826 272861 192886 272889
rect 190826 272849 190832 272861
rect 192880 272849 192886 272861
rect 192938 272849 192944 272901
rect 197104 272849 197110 272901
rect 197162 272889 197168 272901
rect 213232 272889 213238 272901
rect 197162 272861 213238 272889
rect 197162 272849 197168 272861
rect 213232 272849 213238 272861
rect 213290 272849 213296 272901
rect 213328 272849 213334 272901
rect 213386 272889 213392 272901
rect 216688 272889 216694 272901
rect 213386 272861 216694 272889
rect 213386 272849 213392 272861
rect 216688 272849 216694 272861
rect 216746 272849 216752 272901
rect 217552 272849 217558 272901
rect 217610 272889 217616 272901
rect 220432 272889 220438 272901
rect 217610 272861 220438 272889
rect 217610 272849 217616 272861
rect 220432 272849 220438 272861
rect 220490 272849 220496 272901
rect 221008 272849 221014 272901
rect 221066 272889 221072 272901
rect 249040 272889 249046 272901
rect 221066 272861 249046 272889
rect 221066 272849 221072 272861
rect 249040 272849 249046 272861
rect 249098 272849 249104 272901
rect 258352 272849 258358 272901
rect 258410 272889 258416 272901
rect 374320 272889 374326 272901
rect 258410 272861 374326 272889
rect 258410 272849 258416 272861
rect 374320 272849 374326 272861
rect 374378 272849 374384 272901
rect 135952 272775 135958 272827
rect 136010 272815 136016 272827
rect 374530 272815 374558 272935
rect 396976 272923 396982 272935
rect 397034 272923 397040 272975
rect 374608 272849 374614 272901
rect 374666 272889 374672 272901
rect 378448 272889 378454 272901
rect 374666 272861 378454 272889
rect 374666 272849 374672 272861
rect 378448 272849 378454 272861
rect 378506 272849 378512 272901
rect 380368 272889 380374 272901
rect 378562 272861 380374 272889
rect 136010 272787 374558 272815
rect 136010 272775 136016 272787
rect 374800 272775 374806 272827
rect 374858 272815 374864 272827
rect 376240 272815 376246 272827
rect 374858 272787 376246 272815
rect 374858 272775 374864 272787
rect 376240 272775 376246 272787
rect 376298 272775 376304 272827
rect 376336 272775 376342 272827
rect 376394 272815 376400 272827
rect 377392 272815 377398 272827
rect 376394 272787 377398 272815
rect 376394 272775 376400 272787
rect 377392 272775 377398 272787
rect 377450 272775 377456 272827
rect 377488 272775 377494 272827
rect 377546 272815 377552 272827
rect 378160 272815 378166 272827
rect 377546 272787 378166 272815
rect 377546 272775 377552 272787
rect 378160 272775 378166 272787
rect 378218 272775 378224 272827
rect 125296 272701 125302 272753
rect 125354 272741 125360 272753
rect 125354 272713 130334 272741
rect 125354 272701 125360 272713
rect 128944 272627 128950 272679
rect 129002 272667 129008 272679
rect 130306 272667 130334 272713
rect 132496 272701 132502 272753
rect 132554 272741 132560 272753
rect 146896 272741 146902 272753
rect 132554 272713 146902 272741
rect 132554 272701 132560 272713
rect 146896 272701 146902 272713
rect 146954 272701 146960 272753
rect 166960 272701 166966 272753
rect 167018 272741 167024 272753
rect 227536 272741 227542 272753
rect 167018 272713 227542 272741
rect 167018 272701 167024 272713
rect 227536 272701 227542 272713
rect 227594 272701 227600 272753
rect 247600 272701 247606 272753
rect 247658 272741 247664 272753
rect 378448 272741 378454 272753
rect 247658 272713 378454 272741
rect 247658 272701 247664 272713
rect 378448 272701 378454 272713
rect 378506 272701 378512 272753
rect 378562 272667 378590 272861
rect 380368 272849 380374 272861
rect 380426 272849 380432 272901
rect 380560 272849 380566 272901
rect 380618 272889 380624 272901
rect 643888 272889 643894 272901
rect 380618 272861 643894 272889
rect 380618 272849 380624 272861
rect 643888 272849 643894 272861
rect 643946 272849 643952 272901
rect 397072 272815 397078 272827
rect 129002 272639 130142 272667
rect 130306 272639 378590 272667
rect 378658 272787 397078 272815
rect 129002 272627 129008 272639
rect 127696 272553 127702 272605
rect 127754 272593 127760 272605
rect 129520 272593 129526 272605
rect 127754 272565 129526 272593
rect 127754 272553 127760 272565
rect 129520 272553 129526 272565
rect 129578 272553 129584 272605
rect 130114 272593 130142 272639
rect 322576 272593 322582 272605
rect 130114 272565 322582 272593
rect 322576 272553 322582 272565
rect 322634 272553 322640 272605
rect 322960 272553 322966 272605
rect 323018 272593 323024 272605
rect 378658 272593 378686 272787
rect 397072 272775 397078 272787
rect 397130 272775 397136 272827
rect 378832 272701 378838 272753
rect 378890 272741 378896 272753
rect 398320 272741 398326 272753
rect 378890 272713 398326 272741
rect 378890 272701 378896 272713
rect 398320 272701 398326 272713
rect 398378 272701 398384 272753
rect 378736 272627 378742 272679
rect 378794 272667 378800 272679
rect 392464 272667 392470 272679
rect 378794 272639 392470 272667
rect 378794 272627 378800 272639
rect 392464 272627 392470 272639
rect 392522 272627 392528 272679
rect 392560 272627 392566 272679
rect 392618 272667 392624 272679
rect 407248 272667 407254 272679
rect 392618 272639 407254 272667
rect 392618 272627 392624 272639
rect 407248 272627 407254 272639
rect 407306 272627 407312 272679
rect 391696 272593 391702 272605
rect 323018 272565 378686 272593
rect 378850 272565 391702 272593
rect 323018 272553 323024 272565
rect 121744 272479 121750 272531
rect 121802 272519 121808 272531
rect 378736 272519 378742 272531
rect 121802 272491 378742 272519
rect 121802 272479 121808 272491
rect 378736 272479 378742 272491
rect 378794 272479 378800 272531
rect 378850 272457 378878 272565
rect 391696 272553 391702 272565
rect 391754 272553 391760 272605
rect 396784 272593 396790 272605
rect 391810 272565 396790 272593
rect 379216 272479 379222 272531
rect 379274 272519 379280 272531
rect 391810 272519 391838 272565
rect 396784 272553 396790 272565
rect 396842 272553 396848 272605
rect 397360 272553 397366 272605
rect 397418 272593 397424 272605
rect 595120 272593 595126 272605
rect 397418 272565 595126 272593
rect 397418 272553 397424 272565
rect 595120 272553 595126 272565
rect 595178 272553 595184 272605
rect 379274 272491 391838 272519
rect 379274 272479 379280 272491
rect 394576 272479 394582 272531
rect 394634 272519 394640 272531
rect 408112 272519 408118 272531
rect 394634 272491 408118 272519
rect 394634 272479 394640 272491
rect 408112 272479 408118 272491
rect 408170 272479 408176 272531
rect 408226 272491 408446 272519
rect 64912 272405 64918 272457
rect 64970 272445 64976 272457
rect 71920 272445 71926 272457
rect 64970 272417 71926 272445
rect 64970 272405 64976 272417
rect 71920 272405 71926 272417
rect 71978 272405 71984 272457
rect 84880 272405 84886 272457
rect 84938 272445 84944 272457
rect 86320 272445 86326 272457
rect 84938 272417 86326 272445
rect 84938 272405 84944 272417
rect 86320 272405 86326 272417
rect 86378 272405 86384 272457
rect 105040 272405 105046 272457
rect 105098 272445 105104 272457
rect 106480 272445 106486 272457
rect 105098 272417 106486 272445
rect 105098 272405 105104 272417
rect 106480 272405 106486 272417
rect 106538 272405 106544 272457
rect 118096 272405 118102 272457
rect 118154 272445 118160 272457
rect 322576 272445 322582 272457
rect 118154 272417 322582 272445
rect 118154 272405 118160 272417
rect 322576 272405 322582 272417
rect 322634 272405 322640 272457
rect 322768 272405 322774 272457
rect 322826 272445 322832 272457
rect 378448 272445 378454 272457
rect 322826 272417 378454 272445
rect 322826 272405 322832 272417
rect 378448 272405 378454 272417
rect 378506 272405 378512 272457
rect 378832 272405 378838 272457
rect 378890 272405 378896 272457
rect 379120 272405 379126 272457
rect 379178 272445 379184 272457
rect 394192 272445 394198 272457
rect 379178 272417 394198 272445
rect 379178 272405 379184 272417
rect 394192 272405 394198 272417
rect 394250 272405 394256 272457
rect 394480 272405 394486 272457
rect 394538 272445 394544 272457
rect 408226 272445 408254 272491
rect 394538 272417 408254 272445
rect 408418 272445 408446 272491
rect 591568 272445 591574 272457
rect 408418 272417 591574 272445
rect 394538 272405 394544 272417
rect 591568 272405 591574 272417
rect 591626 272405 591632 272457
rect 111088 272331 111094 272383
rect 111146 272371 111152 272383
rect 378064 272371 378070 272383
rect 111146 272343 378070 272371
rect 111146 272331 111152 272343
rect 378064 272331 378070 272343
rect 378122 272331 378128 272383
rect 378928 272331 378934 272383
rect 378986 272371 378992 272383
rect 389488 272371 389494 272383
rect 378986 272343 389494 272371
rect 378986 272331 378992 272343
rect 389488 272331 389494 272343
rect 389546 272331 389552 272383
rect 389584 272331 389590 272383
rect 389642 272371 389648 272383
rect 408208 272371 408214 272383
rect 389642 272343 408214 272371
rect 389642 272331 389648 272343
rect 408208 272331 408214 272343
rect 408266 272331 408272 272383
rect 408304 272331 408310 272383
rect 408362 272371 408368 272383
rect 587920 272371 587926 272383
rect 408362 272343 587926 272371
rect 408362 272331 408368 272343
rect 587920 272331 587926 272343
rect 587978 272331 587984 272383
rect 67024 272257 67030 272309
rect 67082 272297 67088 272309
rect 197104 272297 197110 272309
rect 67082 272269 197110 272297
rect 67082 272257 67088 272269
rect 197104 272257 197110 272269
rect 197162 272257 197168 272309
rect 209776 272257 209782 272309
rect 209834 272297 209840 272309
rect 216112 272297 216118 272309
rect 209834 272269 216118 272297
rect 209834 272257 209840 272269
rect 216112 272257 216118 272269
rect 216170 272257 216176 272309
rect 218224 272257 218230 272309
rect 218282 272297 218288 272309
rect 223984 272297 223990 272309
rect 218282 272269 223990 272297
rect 218282 272257 218288 272269
rect 223984 272257 223990 272269
rect 224042 272257 224048 272309
rect 224560 272257 224566 272309
rect 224618 272297 224624 272309
rect 277552 272297 277558 272309
rect 224618 272269 277558 272297
rect 224618 272257 224624 272269
rect 277552 272257 277558 272269
rect 277610 272257 277616 272309
rect 278800 272257 278806 272309
rect 278858 272297 278864 272309
rect 280048 272297 280054 272309
rect 278858 272269 280054 272297
rect 278858 272257 278864 272269
rect 280048 272257 280054 272269
rect 280106 272257 280112 272309
rect 280720 272257 280726 272309
rect 280778 272297 280784 272309
rect 282352 272297 282358 272309
rect 280778 272269 282358 272297
rect 280778 272257 280784 272269
rect 282352 272257 282358 272269
rect 282410 272257 282416 272309
rect 285520 272257 285526 272309
rect 285578 272297 285584 272309
rect 319792 272297 319798 272309
rect 285578 272269 319798 272297
rect 285578 272257 285584 272269
rect 319792 272257 319798 272269
rect 319850 272257 319856 272309
rect 320368 272257 320374 272309
rect 320426 272297 320432 272309
rect 607024 272297 607030 272309
rect 320426 272269 607030 272297
rect 320426 272257 320432 272269
rect 607024 272257 607030 272269
rect 607082 272257 607088 272309
rect 103888 272183 103894 272235
rect 103946 272223 103952 272235
rect 103946 272195 378686 272223
rect 103946 272183 103952 272195
rect 107440 272109 107446 272161
rect 107498 272149 107504 272161
rect 378352 272149 378358 272161
rect 107498 272121 378358 272149
rect 107498 272109 107504 272121
rect 378352 272109 378358 272121
rect 378410 272109 378416 272161
rect 378658 272149 378686 272195
rect 379024 272183 379030 272235
rect 379082 272223 379088 272235
rect 385264 272223 385270 272235
rect 379082 272195 385270 272223
rect 379082 272183 379088 272195
rect 385264 272183 385270 272195
rect 385322 272183 385328 272235
rect 385552 272183 385558 272235
rect 385610 272223 385616 272235
rect 386800 272223 386806 272235
rect 385610 272195 386806 272223
rect 385610 272183 385616 272195
rect 386800 272183 386806 272195
rect 386858 272183 386864 272235
rect 566512 272223 566518 272235
rect 396514 272195 566518 272223
rect 383056 272149 383062 272161
rect 378658 272121 383062 272149
rect 383056 272109 383062 272121
rect 383114 272109 383120 272161
rect 383248 272109 383254 272161
rect 383306 272149 383312 272161
rect 396400 272149 396406 272161
rect 383306 272121 396406 272149
rect 383306 272109 383312 272121
rect 396400 272109 396406 272121
rect 396458 272109 396464 272161
rect 150256 272035 150262 272087
rect 150314 272075 150320 272087
rect 164272 272075 164278 272087
rect 150314 272047 164278 272075
rect 150314 272035 150320 272047
rect 164272 272035 164278 272047
rect 164330 272035 164336 272087
rect 164560 272035 164566 272087
rect 164618 272075 164624 272087
rect 382960 272075 382966 272087
rect 164618 272047 382966 272075
rect 164618 272035 164624 272047
rect 382960 272035 382966 272047
rect 383018 272035 383024 272087
rect 383344 272035 383350 272087
rect 383402 272075 383408 272087
rect 392560 272075 392566 272087
rect 383402 272047 392566 272075
rect 383402 272035 383408 272047
rect 392560 272035 392566 272047
rect 392618 272035 392624 272087
rect 99184 271961 99190 272013
rect 99242 272001 99248 272013
rect 197200 272001 197206 272013
rect 99242 271973 197206 272001
rect 99242 271961 99248 271973
rect 197200 271961 197206 271973
rect 197258 271961 197264 272013
rect 197296 271961 197302 272013
rect 197354 272001 197360 272013
rect 207856 272001 207862 272013
rect 197354 271973 207862 272001
rect 197354 271961 197360 271973
rect 207856 271961 207862 271973
rect 207914 271961 207920 272013
rect 223696 271961 223702 272013
rect 223754 272001 223760 272013
rect 262384 272001 262390 272013
rect 223754 271973 262390 272001
rect 223754 271961 223760 271973
rect 262384 271961 262390 271973
rect 262442 271961 262448 272013
rect 268048 271961 268054 272013
rect 268106 272001 268112 272013
rect 278992 272001 278998 272013
rect 268106 271973 278998 272001
rect 268106 271961 268112 271973
rect 278992 271961 278998 271973
rect 279050 271961 279056 272013
rect 283792 271961 283798 272013
rect 283850 272001 283856 272013
rect 307312 272001 307318 272013
rect 283850 271973 307318 272001
rect 283850 271961 283856 271973
rect 307312 271961 307318 271973
rect 307370 271961 307376 272013
rect 308464 271961 308470 272013
rect 308522 272001 308528 272013
rect 331408 272001 331414 272013
rect 308522 271973 331414 272001
rect 308522 271961 308528 271973
rect 331408 271961 331414 271973
rect 331466 271961 331472 272013
rect 336976 271961 336982 272013
rect 337034 272001 337040 272013
rect 343024 272001 343030 272013
rect 337034 271973 343030 272001
rect 337034 271961 337040 271973
rect 343024 271961 343030 271973
rect 343082 271961 343088 272013
rect 347920 271961 347926 272013
rect 347978 272001 347984 272013
rect 374512 272001 374518 272013
rect 347978 271973 374518 272001
rect 347978 271961 347984 271973
rect 374512 271961 374518 271973
rect 374570 271961 374576 272013
rect 374704 271961 374710 272013
rect 374762 272001 374768 272013
rect 378544 272001 378550 272013
rect 374762 271973 378550 272001
rect 374762 271961 374768 271973
rect 378544 271961 378550 271973
rect 378602 271961 378608 272013
rect 378640 271961 378646 272013
rect 378698 272001 378704 272013
rect 389584 272001 389590 272013
rect 378698 271973 389590 272001
rect 378698 271961 378704 271973
rect 389584 271961 389590 271973
rect 389642 271961 389648 272013
rect 391600 271961 391606 272013
rect 391658 272001 391664 272013
rect 396514 272001 396542 272195
rect 566512 272183 566518 272195
rect 566570 272183 566576 272235
rect 573712 272149 573718 272161
rect 391658 271973 396542 272001
rect 396610 272121 573718 272149
rect 391658 271961 391664 271973
rect 165808 271887 165814 271939
rect 165866 271927 165872 271939
rect 166960 271927 166966 271939
rect 165866 271899 166966 271927
rect 165866 271887 165872 271899
rect 166960 271887 166966 271899
rect 167018 271887 167024 271939
rect 170512 271887 170518 271939
rect 170570 271927 170576 271939
rect 172720 271927 172726 271939
rect 170570 271899 172726 271927
rect 170570 271887 170576 271899
rect 172720 271887 172726 271899
rect 172778 271887 172784 271939
rect 177616 271887 177622 271939
rect 177674 271927 177680 271939
rect 178384 271927 178390 271939
rect 177674 271899 178390 271927
rect 177674 271887 177680 271899
rect 178384 271887 178390 271899
rect 178442 271887 178448 271939
rect 180016 271887 180022 271939
rect 180074 271927 180080 271939
rect 181360 271927 181366 271939
rect 180074 271899 181366 271927
rect 180074 271887 180080 271899
rect 181360 271887 181366 271899
rect 181418 271887 181424 271939
rect 187024 271887 187030 271939
rect 187082 271927 187088 271939
rect 207280 271927 207286 271939
rect 187082 271899 207286 271927
rect 187082 271887 187088 271899
rect 207280 271887 207286 271899
rect 207338 271887 207344 271939
rect 207376 271887 207382 271939
rect 207434 271927 207440 271939
rect 296848 271927 296854 271939
rect 207434 271899 296854 271927
rect 207434 271887 207440 271899
rect 296848 271887 296854 271899
rect 296906 271887 296912 271939
rect 296944 271887 296950 271939
rect 297002 271927 297008 271939
rect 322576 271927 322582 271939
rect 297002 271899 322582 271927
rect 297002 271887 297008 271899
rect 322576 271887 322582 271899
rect 322634 271887 322640 271939
rect 323056 271887 323062 271939
rect 323114 271927 323120 271939
rect 383248 271927 383254 271939
rect 323114 271899 383254 271927
rect 323114 271887 323120 271899
rect 383248 271887 383254 271899
rect 383306 271887 383312 271939
rect 383440 271887 383446 271939
rect 383498 271927 383504 271939
rect 383498 271899 383582 271927
rect 383498 271887 383504 271899
rect 95632 271813 95638 271865
rect 95690 271853 95696 271865
rect 195856 271853 195862 271865
rect 95690 271825 195862 271853
rect 95690 271813 95696 271825
rect 195856 271813 195862 271825
rect 195914 271813 195920 271865
rect 208048 271813 208054 271865
rect 208106 271853 208112 271865
rect 210256 271853 210262 271865
rect 208106 271825 210262 271853
rect 208106 271813 208112 271825
rect 210256 271813 210262 271825
rect 210314 271813 210320 271865
rect 210352 271813 210358 271865
rect 210410 271853 210416 271865
rect 215440 271853 215446 271865
rect 210410 271825 215446 271853
rect 210410 271813 210416 271825
rect 215440 271813 215446 271825
rect 215498 271813 215504 271865
rect 220816 271813 220822 271865
rect 220874 271853 220880 271865
rect 236176 271853 236182 271865
rect 220874 271825 236182 271853
rect 220874 271813 220880 271825
rect 236176 271813 236182 271825
rect 236234 271813 236240 271865
rect 250192 271813 250198 271865
rect 250250 271853 250256 271865
rect 276784 271853 276790 271865
rect 250250 271825 276790 271853
rect 250250 271813 250256 271825
rect 276784 271813 276790 271825
rect 276842 271813 276848 271865
rect 283408 271813 283414 271865
rect 283466 271853 283472 271865
rect 303664 271853 303670 271865
rect 283466 271825 303670 271853
rect 283466 271813 283472 271825
rect 303664 271813 303670 271825
rect 303722 271813 303728 271865
rect 313648 271813 313654 271865
rect 313706 271853 313712 271865
rect 383344 271853 383350 271865
rect 313706 271825 383350 271853
rect 313706 271813 313712 271825
rect 383344 271813 383350 271825
rect 383402 271813 383408 271865
rect 383554 271853 383582 271899
rect 385264 271887 385270 271939
rect 385322 271927 385328 271939
rect 387472 271927 387478 271939
rect 385322 271899 387478 271927
rect 385322 271887 385328 271899
rect 387472 271887 387478 271899
rect 387530 271887 387536 271939
rect 394384 271887 394390 271939
rect 394442 271927 394448 271939
rect 396610 271927 396638 272121
rect 573712 272109 573718 272121
rect 573770 272109 573776 272161
rect 396784 271961 396790 272013
rect 396842 272001 396848 272013
rect 618832 272001 618838 272013
rect 396842 271973 618838 272001
rect 396842 271961 396848 271973
rect 618832 271961 618838 271973
rect 618890 271961 618896 272013
rect 394442 271899 396638 271927
rect 394442 271887 394448 271899
rect 396688 271887 396694 271939
rect 396746 271927 396752 271939
rect 405712 271927 405718 271939
rect 396746 271899 405718 271927
rect 396746 271887 396752 271899
rect 405712 271887 405718 271899
rect 405770 271887 405776 271939
rect 549904 271853 549910 271865
rect 383554 271825 549910 271853
rect 549904 271813 549910 271825
rect 549962 271813 549968 271865
rect 101488 271739 101494 271791
rect 101546 271779 101552 271791
rect 103600 271779 103606 271791
rect 101546 271751 103606 271779
rect 101546 271739 101552 271751
rect 103600 271739 103606 271751
rect 103658 271739 103664 271791
rect 146896 271739 146902 271791
rect 146954 271779 146960 271791
rect 166768 271779 166774 271791
rect 146954 271751 166774 271779
rect 146954 271739 146960 271751
rect 166768 271739 166774 271751
rect 166826 271739 166832 271791
rect 176464 271739 176470 271791
rect 176522 271779 176528 271791
rect 178480 271779 178486 271791
rect 176522 271751 178486 271779
rect 176522 271739 176528 271751
rect 178480 271739 178486 271751
rect 178538 271739 178544 271791
rect 186832 271779 186838 271791
rect 178786 271751 186838 271779
rect 75376 271665 75382 271717
rect 75434 271705 75440 271717
rect 77680 271705 77686 271717
rect 75434 271677 77686 271705
rect 75434 271665 75440 271677
rect 77680 271665 77686 271677
rect 77738 271665 77744 271717
rect 120976 271665 120982 271717
rect 121034 271705 121040 271717
rect 141040 271705 141046 271717
rect 121034 271677 141046 271705
rect 121034 271665 121040 271677
rect 141040 271665 141046 271677
rect 141098 271665 141104 271717
rect 141328 271665 141334 271717
rect 141386 271705 141392 271717
rect 161104 271705 161110 271717
rect 141386 271677 161110 271705
rect 141386 271665 141392 271677
rect 161104 271665 161110 271677
rect 161162 271665 161168 271717
rect 166576 271665 166582 271717
rect 166634 271705 166640 271717
rect 166864 271705 166870 271717
rect 166634 271677 166870 271705
rect 166634 271665 166640 271677
rect 166864 271665 166870 271677
rect 166922 271665 166928 271717
rect 171664 271665 171670 271717
rect 171722 271705 171728 271717
rect 178786 271705 178814 271751
rect 186832 271739 186838 271751
rect 186890 271739 186896 271791
rect 187024 271739 187030 271791
rect 187082 271779 187088 271791
rect 259312 271779 259318 271791
rect 187082 271751 259318 271779
rect 187082 271739 187088 271751
rect 259312 271739 259318 271751
rect 259370 271739 259376 271791
rect 273520 271739 273526 271791
rect 273578 271779 273584 271791
rect 296656 271779 296662 271791
rect 273578 271751 296662 271779
rect 273578 271739 273584 271751
rect 296656 271739 296662 271751
rect 296714 271739 296720 271791
rect 316720 271739 316726 271791
rect 316778 271779 316784 271791
rect 334096 271779 334102 271791
rect 316778 271751 334102 271779
rect 316778 271739 316784 271751
rect 334096 271739 334102 271751
rect 334154 271739 334160 271791
rect 357040 271739 357046 271791
rect 357098 271779 357104 271791
rect 377488 271779 377494 271791
rect 357098 271751 377494 271779
rect 357098 271739 357104 271751
rect 377488 271739 377494 271751
rect 377546 271739 377552 271791
rect 377776 271739 377782 271791
rect 377834 271779 377840 271791
rect 378736 271779 378742 271791
rect 377834 271751 378742 271779
rect 377834 271739 377840 271751
rect 378736 271739 378742 271751
rect 378794 271739 378800 271791
rect 379024 271739 379030 271791
rect 379082 271779 379088 271791
rect 383728 271779 383734 271791
rect 379082 271751 383734 271779
rect 379082 271739 379088 271751
rect 383728 271739 383734 271751
rect 383786 271739 383792 271791
rect 394096 271739 394102 271791
rect 394154 271779 394160 271791
rect 406576 271779 406582 271791
rect 394154 271751 406582 271779
rect 394154 271739 394160 271751
rect 406576 271739 406582 271751
rect 406634 271739 406640 271791
rect 171722 271677 178814 271705
rect 171722 271665 171728 271677
rect 178864 271665 178870 271717
rect 178922 271705 178928 271717
rect 382960 271705 382966 271717
rect 178922 271677 382966 271705
rect 178922 271665 178928 271677
rect 382960 271665 382966 271677
rect 383018 271665 383024 271717
rect 383248 271665 383254 271717
rect 383306 271705 383312 271717
rect 409264 271705 409270 271717
rect 383306 271677 409270 271705
rect 383306 271665 383312 271677
rect 409264 271665 409270 271677
rect 409322 271665 409328 271717
rect 89584 271591 89590 271643
rect 89642 271631 89648 271643
rect 92080 271631 92086 271643
rect 89642 271603 92086 271631
rect 89642 271591 89648 271603
rect 92080 271591 92086 271603
rect 92138 271591 92144 271643
rect 100816 271591 100822 271643
rect 100874 271631 100880 271643
rect 120784 271631 120790 271643
rect 100874 271603 120790 271631
rect 100874 271591 100880 271603
rect 120784 271591 120790 271603
rect 120842 271591 120848 271643
rect 182416 271591 182422 271643
rect 182474 271631 182480 271643
rect 296848 271631 296854 271643
rect 182474 271603 296854 271631
rect 182474 271591 182480 271603
rect 296848 271591 296854 271603
rect 296906 271591 296912 271643
rect 297040 271591 297046 271643
rect 297098 271631 297104 271643
rect 383056 271631 383062 271643
rect 297098 271603 383062 271631
rect 297098 271591 297104 271603
rect 383056 271591 383062 271603
rect 383114 271591 383120 271643
rect 392752 271591 392758 271643
rect 392810 271631 392816 271643
rect 409936 271631 409942 271643
rect 392810 271603 409942 271631
rect 392810 271591 392816 271603
rect 409936 271591 409942 271603
rect 409994 271591 410000 271643
rect 141136 271517 141142 271569
rect 141194 271557 141200 271569
rect 141616 271557 141622 271569
rect 141194 271529 141622 271557
rect 141194 271517 141200 271529
rect 141616 271517 141622 271529
rect 141674 271517 141680 271569
rect 185968 271517 185974 271569
rect 186026 271557 186032 271569
rect 410992 271557 410998 271569
rect 186026 271529 186974 271557
rect 186026 271517 186032 271529
rect 156880 271443 156886 271495
rect 156938 271483 156944 271495
rect 168112 271483 168118 271495
rect 156938 271455 168118 271483
rect 156938 271443 156944 271455
rect 168112 271443 168118 271455
rect 168170 271443 168176 271495
rect 175312 271443 175318 271495
rect 175370 271483 175376 271495
rect 186832 271483 186838 271495
rect 175370 271455 186838 271483
rect 175370 271443 175376 271455
rect 186832 271443 186838 271455
rect 186890 271443 186896 271495
rect 186946 271483 186974 271529
rect 187138 271529 410998 271557
rect 187138 271483 187166 271529
rect 410992 271517 410998 271529
rect 411050 271517 411056 271569
rect 197296 271483 197302 271495
rect 186946 271455 187166 271483
rect 187234 271455 197302 271483
rect 102640 271369 102646 271421
rect 102698 271409 102704 271421
rect 187234 271409 187262 271455
rect 197296 271443 197302 271455
rect 197354 271443 197360 271495
rect 205840 271443 205846 271495
rect 205898 271483 205904 271495
rect 411952 271483 411958 271495
rect 205898 271455 411958 271483
rect 205898 271443 205904 271455
rect 411952 271443 411958 271455
rect 412010 271443 412016 271495
rect 421840 271443 421846 271495
rect 421898 271483 421904 271495
rect 431920 271483 431926 271495
rect 421898 271455 431926 271483
rect 421898 271443 421904 271455
rect 431920 271443 431926 271455
rect 431978 271443 431984 271495
rect 211888 271409 211894 271421
rect 102698 271381 187262 271409
rect 195298 271381 211894 271409
rect 102698 271369 102704 271381
rect 113488 271295 113494 271347
rect 113546 271335 113552 271347
rect 195298 271335 195326 271381
rect 211888 271369 211894 271381
rect 211946 271369 211952 271421
rect 220336 271369 220342 271421
rect 220394 271409 220400 271421
rect 241840 271409 241846 271421
rect 220394 271381 241846 271409
rect 220394 271369 220400 271381
rect 241840 271369 241846 271381
rect 241898 271369 241904 271421
rect 246640 271369 246646 271421
rect 246698 271409 246704 271421
rect 257680 271409 257686 271421
rect 246698 271381 257686 271409
rect 246698 271369 246704 271381
rect 257680 271369 257686 271381
rect 257738 271369 257744 271421
rect 277264 271409 277270 271421
rect 260770 271381 277270 271409
rect 113546 271307 195326 271335
rect 113546 271295 113552 271307
rect 195952 271295 195958 271347
rect 196010 271335 196016 271347
rect 206608 271335 206614 271347
rect 196010 271307 206614 271335
rect 196010 271295 196016 271307
rect 206608 271295 206614 271307
rect 206666 271295 206672 271347
rect 219760 271295 219766 271347
rect 219818 271335 219824 271347
rect 238288 271335 238294 271347
rect 219818 271307 238294 271335
rect 219818 271295 219824 271307
rect 238288 271295 238294 271307
rect 238346 271295 238352 271347
rect 241552 271295 241558 271347
rect 241610 271335 241616 271347
rect 242032 271335 242038 271347
rect 241610 271307 242038 271335
rect 241610 271295 241616 271307
rect 242032 271295 242038 271307
rect 242090 271295 242096 271347
rect 253744 271295 253750 271347
rect 253802 271335 253808 271347
rect 260770 271335 260798 271381
rect 277264 271369 277270 271381
rect 277322 271369 277328 271421
rect 314320 271369 314326 271421
rect 314378 271409 314384 271421
rect 327568 271409 327574 271421
rect 314378 271381 327574 271409
rect 314378 271369 314384 271381
rect 327568 271369 327574 271381
rect 327626 271369 327632 271421
rect 333424 271369 333430 271421
rect 333482 271409 333488 271421
rect 342640 271409 342646 271421
rect 333482 271381 342646 271409
rect 333482 271369 333488 271381
rect 342640 271369 342646 271381
rect 342698 271369 342704 271421
rect 347440 271369 347446 271421
rect 347498 271409 347504 271421
rect 372688 271409 372694 271421
rect 347498 271381 372694 271409
rect 347498 271369 347504 271381
rect 372688 271369 372694 271381
rect 372746 271369 372752 271421
rect 380176 271409 380182 271421
rect 372802 271381 380182 271409
rect 253802 271307 260798 271335
rect 253802 271295 253808 271307
rect 264496 271295 264502 271347
rect 264554 271335 264560 271347
rect 278512 271335 278518 271347
rect 264554 271307 278518 271335
rect 264554 271295 264560 271307
rect 278512 271295 278518 271307
rect 278570 271295 278576 271347
rect 282928 271295 282934 271347
rect 282986 271335 282992 271347
rect 300112 271335 300118 271347
rect 282986 271307 300118 271335
rect 282986 271295 282992 271307
rect 300112 271295 300118 271307
rect 300170 271295 300176 271347
rect 315376 271295 315382 271347
rect 315434 271335 315440 271347
rect 322672 271335 322678 271347
rect 315434 271307 322678 271335
rect 315434 271295 315440 271307
rect 322672 271295 322678 271307
rect 322730 271295 322736 271347
rect 322768 271295 322774 271347
rect 322826 271335 322832 271347
rect 325648 271335 325654 271347
rect 322826 271307 325654 271335
rect 322826 271295 322832 271307
rect 325648 271295 325654 271307
rect 325706 271295 325712 271347
rect 327472 271335 327478 271347
rect 326242 271307 327478 271335
rect 116944 271221 116950 271273
rect 117002 271261 117008 271273
rect 156880 271261 156886 271273
rect 117002 271233 156886 271261
rect 117002 271221 117008 271233
rect 156880 271221 156886 271233
rect 156938 271221 156944 271273
rect 168112 271221 168118 271273
rect 168170 271261 168176 271273
rect 211792 271261 211798 271273
rect 168170 271233 211798 271261
rect 168170 271221 168176 271233
rect 211792 271221 211798 271233
rect 211850 271221 211856 271273
rect 262192 271221 262198 271273
rect 262250 271261 262256 271273
rect 282160 271261 282166 271273
rect 262250 271233 282166 271261
rect 262250 271221 262256 271233
rect 282160 271221 282166 271233
rect 282218 271221 282224 271273
rect 306256 271221 306262 271273
rect 306314 271261 306320 271273
rect 315184 271261 315190 271273
rect 306314 271233 315190 271261
rect 306314 271221 306320 271233
rect 315184 271221 315190 271233
rect 315242 271221 315248 271273
rect 315664 271221 315670 271273
rect 315722 271261 315728 271273
rect 322000 271261 322006 271273
rect 315722 271233 322006 271261
rect 315722 271221 315728 271233
rect 322000 271221 322006 271233
rect 322058 271221 322064 271273
rect 322096 271221 322102 271273
rect 322154 271261 322160 271273
rect 326242 271261 326270 271307
rect 327472 271295 327478 271307
rect 327530 271295 327536 271347
rect 329968 271295 329974 271347
rect 330026 271335 330032 271347
rect 341968 271335 341974 271347
rect 330026 271307 341974 271335
rect 330026 271295 330032 271307
rect 341968 271295 341974 271307
rect 342026 271295 342032 271347
rect 357328 271295 357334 271347
rect 357386 271335 357392 271347
rect 357386 271307 362174 271335
rect 357386 271295 357392 271307
rect 322154 271233 326270 271261
rect 322154 271221 322160 271233
rect 326320 271221 326326 271273
rect 326378 271261 326384 271273
rect 341488 271261 341494 271273
rect 326378 271233 341494 271261
rect 326378 271221 326384 271233
rect 341488 271221 341494 271233
rect 341546 271221 341552 271273
rect 345712 271221 345718 271273
rect 345770 271261 345776 271273
rect 358096 271261 358102 271273
rect 345770 271233 358102 271261
rect 345770 271221 345776 271233
rect 358096 271221 358102 271233
rect 358154 271221 358160 271273
rect 120496 271147 120502 271199
rect 120554 271187 120560 271199
rect 197104 271187 197110 271199
rect 120554 271159 197110 271187
rect 120554 271147 120560 271159
rect 197104 271147 197110 271159
rect 197162 271147 197168 271199
rect 202576 271147 202582 271199
rect 202634 271187 202640 271199
rect 202634 271159 205214 271187
rect 202634 271147 202640 271159
rect 109840 271073 109846 271125
rect 109898 271113 109904 271125
rect 109898 271085 188318 271113
rect 109898 271073 109904 271085
rect 184720 270999 184726 271051
rect 184778 271039 184784 271051
rect 187024 271039 187030 271051
rect 184778 271011 187030 271039
rect 184778 270999 184784 271011
rect 187024 270999 187030 271011
rect 187082 270999 187088 271051
rect 188290 271039 188318 271085
rect 188368 271073 188374 271125
rect 188426 271113 188432 271125
rect 190000 271113 190006 271125
rect 188426 271085 190006 271113
rect 188426 271073 188432 271085
rect 190000 271073 190006 271085
rect 190058 271073 190064 271125
rect 190576 271073 190582 271125
rect 190634 271113 190640 271125
rect 204496 271113 204502 271125
rect 190634 271085 204502 271113
rect 190634 271073 190640 271085
rect 204496 271073 204502 271085
rect 204554 271073 204560 271125
rect 205186 271113 205214 271159
rect 219280 271147 219286 271199
rect 219338 271187 219344 271199
rect 234640 271187 234646 271199
rect 219338 271159 234646 271187
rect 219338 271147 219344 271159
rect 234640 271147 234646 271159
rect 234698 271147 234704 271199
rect 269392 271147 269398 271199
rect 269450 271187 269456 271199
rect 270448 271187 270454 271199
rect 269450 271159 270454 271187
rect 269450 271147 269456 271159
rect 270448 271147 270454 271159
rect 270506 271147 270512 271199
rect 282736 271147 282742 271199
rect 282794 271187 282800 271199
rect 282794 271159 292286 271187
rect 282794 271147 282800 271159
rect 210352 271113 210358 271125
rect 205186 271085 210358 271113
rect 210352 271073 210358 271085
rect 210410 271073 210416 271125
rect 210448 271073 210454 271125
rect 210506 271113 210512 271125
rect 215536 271113 215542 271125
rect 210506 271085 215542 271113
rect 210506 271073 210512 271085
rect 215536 271073 215542 271085
rect 215594 271073 215600 271125
rect 218896 271073 218902 271125
rect 218954 271113 218960 271125
rect 231184 271113 231190 271125
rect 218954 271085 231190 271113
rect 218954 271073 218960 271085
rect 231184 271073 231190 271085
rect 231242 271073 231248 271125
rect 260944 271073 260950 271125
rect 261002 271113 261008 271125
rect 278128 271113 278134 271125
rect 261002 271085 278134 271113
rect 261002 271073 261008 271085
rect 278128 271073 278134 271085
rect 278186 271073 278192 271125
rect 282160 271073 282166 271125
rect 282218 271113 282224 271125
rect 290896 271113 290902 271125
rect 282218 271085 290902 271113
rect 282218 271073 282224 271085
rect 290896 271073 290902 271085
rect 290954 271073 290960 271125
rect 195856 271039 195862 271051
rect 188290 271011 195862 271039
rect 195856 270999 195862 271011
rect 195914 270999 195920 271051
rect 196240 270999 196246 271051
rect 196298 271039 196304 271051
rect 269872 271039 269878 271051
rect 196298 271011 269878 271039
rect 196298 270999 196304 271011
rect 269872 270999 269878 271011
rect 269930 270999 269936 271051
rect 281680 270999 281686 271051
rect 281738 271039 281744 271051
rect 289456 271039 289462 271051
rect 281738 271011 289462 271039
rect 281738 270999 281744 271011
rect 289456 270999 289462 271011
rect 289514 270999 289520 271051
rect 292258 271039 292286 271159
rect 292528 271147 292534 271199
rect 292586 271187 292592 271199
rect 315280 271187 315286 271199
rect 292586 271159 315286 271187
rect 292586 271147 292592 271159
rect 315280 271147 315286 271159
rect 315338 271147 315344 271199
rect 315472 271147 315478 271199
rect 315530 271187 315536 271199
rect 327088 271187 327094 271199
rect 315530 271159 327094 271187
rect 315530 271147 315536 271159
rect 327088 271147 327094 271159
rect 327146 271147 327152 271199
rect 327952 271187 327958 271199
rect 327202 271159 327958 271187
rect 297136 271113 297142 271125
rect 293122 271085 297142 271113
rect 293122 271039 293150 271085
rect 297136 271073 297142 271085
rect 297194 271073 297200 271125
rect 302800 271073 302806 271125
rect 302858 271113 302864 271125
rect 302858 271085 319262 271113
rect 302858 271073 302864 271085
rect 292258 271011 293150 271039
rect 294256 270999 294262 271051
rect 294314 271039 294320 271051
rect 319024 271039 319030 271051
rect 294314 271011 319030 271039
rect 294314 270999 294320 271011
rect 319024 270999 319030 271011
rect 319082 270999 319088 271051
rect 319234 271039 319262 271085
rect 319312 271073 319318 271125
rect 319370 271113 319376 271125
rect 319370 271085 322718 271113
rect 319370 271073 319376 271085
rect 322288 271039 322294 271051
rect 319234 271011 322294 271039
rect 322288 270999 322294 271011
rect 322346 270999 322352 271051
rect 322690 271039 322718 271085
rect 322768 271073 322774 271125
rect 322826 271113 322832 271125
rect 327202 271113 327230 271159
rect 327952 271147 327958 271159
rect 328010 271147 328016 271199
rect 346384 271147 346390 271199
rect 346442 271187 346448 271199
rect 362032 271187 362038 271199
rect 346442 271159 362038 271187
rect 346442 271147 346448 271159
rect 362032 271147 362038 271159
rect 362090 271147 362096 271199
rect 362146 271187 362174 271307
rect 366448 271295 366454 271347
rect 366506 271335 366512 271347
rect 372802 271335 372830 271381
rect 380176 271369 380182 271381
rect 380234 271369 380240 271421
rect 380368 271369 380374 271421
rect 380426 271409 380432 271421
rect 380426 271381 383294 271409
rect 380426 271369 380432 271381
rect 383152 271335 383158 271347
rect 366506 271307 372830 271335
rect 372898 271307 383158 271335
rect 366506 271295 366512 271307
rect 367120 271221 367126 271273
rect 367178 271261 367184 271273
rect 372898 271261 372926 271307
rect 383152 271295 383158 271307
rect 383210 271295 383216 271347
rect 383266 271335 383294 271381
rect 383440 271369 383446 271421
rect 383498 271409 383504 271421
rect 384112 271409 384118 271421
rect 383498 271381 384118 271409
rect 383498 271369 383504 271381
rect 384112 271369 384118 271381
rect 384170 271369 384176 271421
rect 384208 271369 384214 271421
rect 384266 271409 384272 271421
rect 593968 271409 593974 271421
rect 384266 271381 593974 271409
rect 384266 271369 384272 271381
rect 593968 271369 593974 271381
rect 594026 271369 594032 271421
rect 590320 271335 590326 271347
rect 383266 271307 590326 271335
rect 590320 271295 590326 271307
rect 590378 271295 590384 271347
rect 367178 271233 372926 271261
rect 367178 271221 367184 271233
rect 372976 271221 372982 271273
rect 373034 271261 373040 271273
rect 421840 271261 421846 271273
rect 373034 271233 421846 271261
rect 373034 271221 373040 271233
rect 421840 271221 421846 271233
rect 421898 271221 421904 271273
rect 431920 271221 431926 271273
rect 431978 271261 431984 271273
rect 480976 271261 480982 271273
rect 431978 271233 480982 271261
rect 431978 271221 431984 271233
rect 480976 271221 480982 271233
rect 481034 271221 481040 271273
rect 501040 271221 501046 271273
rect 501098 271261 501104 271273
rect 543952 271261 543958 271273
rect 501098 271233 543958 271261
rect 501098 271221 501104 271233
rect 543952 271221 543958 271233
rect 544010 271221 544016 271273
rect 377104 271187 377110 271199
rect 362146 271159 377110 271187
rect 377104 271147 377110 271159
rect 377162 271147 377168 271199
rect 377200 271147 377206 271199
rect 377258 271187 377264 271199
rect 431632 271187 431638 271199
rect 377258 271159 431638 271187
rect 377258 271147 377264 271159
rect 431632 271147 431638 271159
rect 431690 271147 431696 271199
rect 431824 271147 431830 271199
rect 431882 271187 431888 271199
rect 545200 271187 545206 271199
rect 431882 271159 545206 271187
rect 431882 271147 431888 271159
rect 545200 271147 545206 271159
rect 545258 271147 545264 271199
rect 340912 271113 340918 271125
rect 322826 271085 327230 271113
rect 327298 271085 340918 271113
rect 322826 271073 322832 271085
rect 327298 271039 327326 271085
rect 340912 271073 340918 271085
rect 340970 271073 340976 271125
rect 345232 271073 345238 271125
rect 345290 271113 345296 271125
rect 354832 271113 354838 271125
rect 345290 271085 354838 271113
rect 345290 271073 345296 271085
rect 354832 271073 354838 271085
rect 354890 271073 354896 271125
rect 357712 271073 357718 271125
rect 357770 271113 357776 271125
rect 371440 271113 371446 271125
rect 357770 271085 371446 271113
rect 357770 271073 357776 271085
rect 371440 271073 371446 271085
rect 371498 271073 371504 271125
rect 371536 271073 371542 271125
rect 371594 271113 371600 271125
rect 371594 271085 398942 271113
rect 371594 271073 371600 271085
rect 322690 271011 327326 271039
rect 327472 270999 327478 271051
rect 327530 271039 327536 271051
rect 377008 271039 377014 271051
rect 327530 271011 377014 271039
rect 327530 270999 327536 271011
rect 377008 270999 377014 271011
rect 377066 270999 377072 271051
rect 377104 270999 377110 271051
rect 377162 271039 377168 271051
rect 378640 271039 378646 271051
rect 377162 271011 378646 271039
rect 377162 270999 377168 271011
rect 378640 270999 378646 271011
rect 378698 270999 378704 271051
rect 378736 270999 378742 271051
rect 378794 271039 378800 271051
rect 384208 271039 384214 271051
rect 378794 271011 384214 271039
rect 378794 270999 378800 271011
rect 384208 270999 384214 271011
rect 384266 270999 384272 271051
rect 385648 270999 385654 271051
rect 385706 271039 385712 271051
rect 398800 271039 398806 271051
rect 385706 271011 398806 271039
rect 385706 270999 385712 271011
rect 398800 270999 398806 271011
rect 398858 270999 398864 271051
rect 398914 271039 398942 271085
rect 398992 271073 398998 271125
rect 399050 271113 399056 271125
rect 449296 271113 449302 271125
rect 399050 271085 449302 271113
rect 399050 271073 399056 271085
rect 449296 271073 449302 271085
rect 449354 271073 449360 271125
rect 449584 271073 449590 271125
rect 449642 271113 449648 271125
rect 481072 271113 481078 271125
rect 449642 271085 481078 271113
rect 449642 271073 449648 271085
rect 481072 271073 481078 271085
rect 481130 271073 481136 271125
rect 481168 271073 481174 271125
rect 481226 271113 481232 271125
rect 534448 271113 534454 271125
rect 481226 271085 534454 271113
rect 481226 271073 481232 271085
rect 534448 271073 534454 271085
rect 534506 271073 534512 271125
rect 402352 271039 402358 271051
rect 398914 271011 402358 271039
rect 402352 270999 402358 271011
rect 402410 270999 402416 271051
rect 428176 271039 428182 271051
rect 418978 271011 428182 271039
rect 241840 270965 241846 270977
rect 187330 270937 196094 270965
rect 175600 270851 175606 270903
rect 175658 270891 175664 270903
rect 175658 270863 185822 270891
rect 175658 270851 175664 270863
rect 130096 270777 130102 270829
rect 130154 270817 130160 270829
rect 132400 270817 132406 270829
rect 130154 270789 132406 270817
rect 130154 270777 130160 270789
rect 132400 270777 132406 270789
rect 132458 270777 132464 270829
rect 144400 270777 144406 270829
rect 144458 270817 144464 270829
rect 146800 270817 146806 270829
rect 144458 270789 146806 270817
rect 144458 270777 144464 270789
rect 146800 270777 146806 270789
rect 146858 270777 146864 270829
rect 168400 270777 168406 270829
rect 168458 270817 168464 270829
rect 175504 270817 175510 270829
rect 168458 270789 175510 270817
rect 168458 270777 168464 270789
rect 175504 270777 175510 270789
rect 175562 270777 175568 270829
rect 185794 270817 185822 270863
rect 187330 270817 187358 270937
rect 189520 270851 189526 270903
rect 189578 270891 189584 270903
rect 196066 270891 196094 270937
rect 218626 270937 241846 270965
rect 218626 270891 218654 270937
rect 241840 270925 241846 270937
rect 241898 270925 241904 270977
rect 241936 270925 241942 270977
rect 241994 270965 242000 270977
rect 241994 270937 252062 270965
rect 241994 270925 242000 270937
rect 189578 270863 195998 270891
rect 196066 270863 218654 270891
rect 189578 270851 189584 270863
rect 185794 270789 187358 270817
rect 193072 270777 193078 270829
rect 193130 270817 193136 270829
rect 195856 270817 195862 270829
rect 193130 270789 195862 270817
rect 193130 270777 193136 270789
rect 195856 270777 195862 270789
rect 195914 270777 195920 270829
rect 195970 270817 195998 270863
rect 218704 270851 218710 270903
rect 218762 270891 218768 270903
rect 227632 270891 227638 270903
rect 218762 270863 227638 270891
rect 218762 270851 218768 270863
rect 227632 270851 227638 270863
rect 227690 270851 227696 270903
rect 252034 270891 252062 270937
rect 257680 270925 257686 270977
rect 257738 270965 257744 270977
rect 276208 270965 276214 270977
rect 257738 270937 276214 270965
rect 257738 270925 257744 270937
rect 276208 270925 276214 270937
rect 276266 270925 276272 270977
rect 394096 270965 394102 270977
rect 277762 270937 320030 270965
rect 277762 270891 277790 270937
rect 252034 270863 277790 270891
rect 315184 270851 315190 270903
rect 315242 270891 315248 270903
rect 316912 270891 316918 270903
rect 315242 270863 316918 270891
rect 315242 270851 315248 270863
rect 316912 270851 316918 270863
rect 316970 270851 316976 270903
rect 320002 270891 320030 270937
rect 320194 270937 394102 270965
rect 320194 270891 320222 270937
rect 394096 270925 394102 270937
rect 394154 270925 394160 270977
rect 394288 270925 394294 270977
rect 394346 270965 394352 270977
rect 402832 270965 402838 270977
rect 394346 270937 402838 270965
rect 394346 270925 394352 270937
rect 402832 270925 402838 270937
rect 402890 270925 402896 270977
rect 402928 270925 402934 270977
rect 402986 270965 402992 270977
rect 418978 270965 419006 271011
rect 428176 270999 428182 271011
rect 428234 270999 428240 271051
rect 446320 270999 446326 271051
rect 446378 271039 446384 271051
rect 452176 271039 452182 271051
rect 446378 271011 452182 271039
rect 446378 270999 446384 271011
rect 452176 270999 452182 271011
rect 452234 270999 452240 271051
rect 469456 270999 469462 271051
rect 469514 271039 469520 271051
rect 489520 271039 489526 271051
rect 469514 271011 489526 271039
rect 469514 270999 469520 271011
rect 489520 270999 489526 271011
rect 489578 270999 489584 271051
rect 518416 271039 518422 271051
rect 511138 271011 518422 271039
rect 402986 270937 419006 270965
rect 402986 270925 402992 270937
rect 489616 270925 489622 270977
rect 489674 270965 489680 270977
rect 511138 270965 511166 271011
rect 518416 270999 518422 271011
rect 518474 270999 518480 271051
rect 518512 270999 518518 271051
rect 518570 271039 518576 271051
rect 548560 271039 548566 271051
rect 518570 271011 548566 271039
rect 518570 270999 518576 271011
rect 548560 270999 548566 271011
rect 548618 270999 548624 271051
rect 558640 270999 558646 271051
rect 558698 271039 558704 271051
rect 564496 271039 564502 271051
rect 558698 271011 564502 271039
rect 558698 270999 558704 271011
rect 564496 270999 564502 271011
rect 564554 270999 564560 271051
rect 489674 270937 511166 270965
rect 489674 270925 489680 270937
rect 320002 270863 320222 270891
rect 322000 270851 322006 270903
rect 322058 270891 322064 270903
rect 340432 270891 340438 270903
rect 322058 270863 340438 270891
rect 322058 270851 322064 270863
rect 340432 270851 340438 270863
rect 340490 270851 340496 270903
rect 344752 270851 344758 270903
rect 344810 270891 344816 270903
rect 351280 270891 351286 270903
rect 344810 270863 351286 270891
rect 344810 270851 344816 270863
rect 351280 270851 351286 270863
rect 351338 270851 351344 270903
rect 369136 270891 369142 270903
rect 358498 270863 369142 270891
rect 205840 270817 205846 270829
rect 195970 270789 205846 270817
rect 205840 270777 205846 270789
rect 205898 270777 205904 270829
rect 206146 270789 210590 270817
rect 68176 270703 68182 270755
rect 68234 270743 68240 270755
rect 69040 270743 69046 270755
rect 68234 270715 69046 270743
rect 68234 270703 68240 270715
rect 69040 270703 69046 270715
rect 69098 270703 69104 270755
rect 98032 270703 98038 270755
rect 98090 270743 98096 270755
rect 100720 270743 100726 270755
rect 98090 270715 100726 270743
rect 98090 270703 98096 270715
rect 100720 270703 100726 270715
rect 100778 270703 100784 270755
rect 115792 270703 115798 270755
rect 115850 270743 115856 270755
rect 118000 270743 118006 270755
rect 115850 270715 118006 270743
rect 115850 270703 115856 270715
rect 118000 270703 118006 270715
rect 118058 270703 118064 270755
rect 119344 270703 119350 270755
rect 119402 270743 119408 270755
rect 120880 270743 120886 270755
rect 119402 270715 120886 270743
rect 119402 270703 119408 270715
rect 120880 270703 120886 270715
rect 120938 270703 120944 270755
rect 122896 270703 122902 270755
rect 122954 270743 122960 270755
rect 123760 270743 123766 270755
rect 122954 270715 123766 270743
rect 122954 270703 122960 270715
rect 123760 270703 123766 270715
rect 123818 270703 123824 270755
rect 124144 270703 124150 270755
rect 124202 270743 124208 270755
rect 126544 270743 126550 270755
rect 124202 270715 126550 270743
rect 124202 270703 124208 270715
rect 126544 270703 126550 270715
rect 126602 270703 126608 270755
rect 131248 270703 131254 270755
rect 131306 270743 131312 270755
rect 132304 270743 132310 270755
rect 131306 270715 132310 270743
rect 131306 270703 131312 270715
rect 132304 270703 132310 270715
rect 132362 270703 132368 270755
rect 133552 270703 133558 270755
rect 133610 270743 133616 270755
rect 135280 270743 135286 270755
rect 133610 270715 135286 270743
rect 133610 270703 133616 270715
rect 135280 270703 135286 270715
rect 135338 270703 135344 270755
rect 137200 270703 137206 270755
rect 137258 270743 137264 270755
rect 138160 270743 138166 270755
rect 137258 270715 138166 270743
rect 137258 270703 137264 270715
rect 138160 270703 138166 270715
rect 138218 270703 138224 270755
rect 138352 270703 138358 270755
rect 138410 270743 138416 270755
rect 140944 270743 140950 270755
rect 138410 270715 140950 270743
rect 138410 270703 138416 270715
rect 140944 270703 140950 270715
rect 141002 270703 141008 270755
rect 145552 270703 145558 270755
rect 145610 270743 145616 270755
rect 146704 270743 146710 270755
rect 145610 270715 146710 270743
rect 145610 270703 145616 270715
rect 146704 270703 146710 270715
rect 146762 270703 146768 270755
rect 191920 270703 191926 270755
rect 191978 270743 191984 270755
rect 191978 270715 195422 270743
rect 191978 270703 191984 270715
rect 195394 270669 195422 270715
rect 195472 270703 195478 270755
rect 195530 270743 195536 270755
rect 206146 270743 206174 270789
rect 195530 270715 206174 270743
rect 195530 270703 195536 270715
rect 206224 270703 206230 270755
rect 206282 270743 206288 270755
rect 210448 270743 210454 270755
rect 206282 270715 210454 270743
rect 206282 270703 206288 270715
rect 210448 270703 210454 270715
rect 210506 270703 210512 270755
rect 210562 270743 210590 270789
rect 210640 270777 210646 270829
rect 210698 270817 210704 270829
rect 212176 270817 212182 270829
rect 210698 270789 212182 270817
rect 210698 270777 210704 270789
rect 212176 270777 212182 270789
rect 212234 270777 212240 270829
rect 257296 270777 257302 270829
rect 257354 270817 257360 270829
rect 277456 270817 277462 270829
rect 257354 270789 277462 270817
rect 257354 270777 257360 270789
rect 277456 270777 277462 270789
rect 277514 270777 277520 270829
rect 314800 270777 314806 270829
rect 314858 270817 314864 270829
rect 319696 270817 319702 270829
rect 314858 270789 319702 270817
rect 314858 270777 314864 270789
rect 319696 270777 319702 270789
rect 319754 270777 319760 270829
rect 322960 270777 322966 270829
rect 323018 270817 323024 270829
rect 324880 270817 324886 270829
rect 323018 270789 324886 270817
rect 323018 270777 323024 270789
rect 324880 270777 324886 270789
rect 324938 270777 324944 270829
rect 324976 270777 324982 270829
rect 325034 270817 325040 270829
rect 328240 270817 328246 270829
rect 325034 270789 328246 270817
rect 325034 270777 325040 270789
rect 328240 270777 328246 270789
rect 328298 270777 328304 270829
rect 328336 270777 328342 270829
rect 328394 270817 328400 270829
rect 331216 270817 331222 270829
rect 328394 270789 331222 270817
rect 328394 270777 328400 270789
rect 331216 270777 331222 270789
rect 331274 270777 331280 270829
rect 339856 270777 339862 270829
rect 339914 270817 339920 270829
rect 345328 270817 345334 270829
rect 339914 270789 345334 270817
rect 339914 270777 339920 270789
rect 345328 270777 345334 270789
rect 345386 270777 345392 270829
rect 347824 270777 347830 270829
rect 347882 270817 347888 270829
rect 358498 270817 358526 270863
rect 369136 270851 369142 270863
rect 369194 270851 369200 270903
rect 369232 270851 369238 270903
rect 369290 270891 369296 270903
rect 380272 270891 380278 270903
rect 369290 270863 380278 270891
rect 369290 270851 369296 270863
rect 380272 270851 380278 270863
rect 380330 270851 380336 270903
rect 380944 270851 380950 270903
rect 381002 270891 381008 270903
rect 381424 270891 381430 270903
rect 381002 270863 381430 270891
rect 381002 270851 381008 270863
rect 381424 270851 381430 270863
rect 381482 270851 381488 270903
rect 383056 270851 383062 270903
rect 383114 270891 383120 270903
rect 392752 270891 392758 270903
rect 383114 270863 392758 270891
rect 383114 270851 383120 270863
rect 392752 270851 392758 270863
rect 392810 270851 392816 270903
rect 392848 270851 392854 270903
rect 392906 270891 392912 270903
rect 452176 270891 452182 270903
rect 392906 270863 452182 270891
rect 392906 270851 392912 270863
rect 452176 270851 452182 270863
rect 452234 270851 452240 270903
rect 452464 270851 452470 270903
rect 452522 270891 452528 270903
rect 541552 270891 541558 270903
rect 452522 270863 541558 270891
rect 452522 270851 452528 270863
rect 541552 270851 541558 270863
rect 541610 270851 541616 270903
rect 548560 270851 548566 270903
rect 548618 270891 548624 270903
rect 558640 270891 558646 270903
rect 548618 270863 558646 270891
rect 548618 270851 548624 270863
rect 558640 270851 558646 270863
rect 558698 270851 558704 270903
rect 347882 270789 358526 270817
rect 347882 270777 347888 270789
rect 362032 270777 362038 270829
rect 362090 270817 362096 270829
rect 369424 270817 369430 270829
rect 362090 270789 369430 270817
rect 362090 270777 362096 270789
rect 369424 270777 369430 270789
rect 369482 270777 369488 270829
rect 369904 270777 369910 270829
rect 369962 270817 369968 270829
rect 374416 270817 374422 270829
rect 369962 270789 374422 270817
rect 369962 270777 369968 270789
rect 374416 270777 374422 270789
rect 374474 270777 374480 270829
rect 374512 270777 374518 270829
rect 374570 270817 374576 270829
rect 380368 270817 380374 270829
rect 374570 270789 380374 270817
rect 374570 270777 374576 270789
rect 380368 270777 380374 270789
rect 380426 270777 380432 270829
rect 383152 270777 383158 270829
rect 383210 270817 383216 270829
rect 386320 270817 386326 270829
rect 383210 270789 386326 270817
rect 383210 270777 383216 270789
rect 386320 270777 386326 270789
rect 386378 270777 386384 270829
rect 387472 270777 387478 270829
rect 387530 270817 387536 270829
rect 510640 270817 510646 270829
rect 387530 270789 510646 270817
rect 387530 270777 387536 270789
rect 510640 270777 510646 270789
rect 510698 270777 510704 270829
rect 214480 270743 214486 270755
rect 210562 270715 214486 270743
rect 214480 270703 214486 270715
rect 214538 270703 214544 270755
rect 251248 270703 251254 270755
rect 251306 270743 251312 270755
rect 252208 270743 252214 270755
rect 251306 270715 252214 270743
rect 251306 270703 251312 270715
rect 252208 270703 252214 270715
rect 252266 270703 252272 270755
rect 268720 270703 268726 270755
rect 268778 270743 268784 270755
rect 316720 270743 316726 270755
rect 268778 270715 316726 270743
rect 268778 270703 268784 270715
rect 316720 270703 316726 270715
rect 316778 270703 316784 270755
rect 317104 270703 317110 270755
rect 317162 270743 317168 270755
rect 392080 270743 392086 270755
rect 317162 270715 392086 270743
rect 317162 270703 317168 270715
rect 392080 270703 392086 270715
rect 392138 270703 392144 270755
rect 394480 270703 394486 270755
rect 394538 270743 394544 270755
rect 452176 270743 452182 270755
rect 394538 270715 452182 270743
rect 394538 270703 394544 270715
rect 452176 270703 452182 270715
rect 452234 270703 452240 270755
rect 452656 270703 452662 270755
rect 452714 270743 452720 270755
rect 570160 270743 570166 270755
rect 452714 270715 570166 270743
rect 452714 270703 452720 270715
rect 570160 270703 570166 270715
rect 570218 270703 570224 270755
rect 213808 270669 213814 270681
rect 195394 270641 213814 270669
rect 213808 270629 213814 270641
rect 213866 270629 213872 270681
rect 243280 270629 243286 270681
rect 243338 270669 243344 270681
rect 431056 270669 431062 270681
rect 243338 270641 431062 270669
rect 243338 270629 243344 270641
rect 431056 270629 431062 270641
rect 431114 270629 431120 270681
rect 672496 270629 672502 270681
rect 672554 270669 672560 270681
rect 673840 270669 673846 270681
rect 672554 270641 673846 270669
rect 672554 270629 672560 270641
rect 673840 270629 673846 270641
rect 673898 270629 673904 270681
rect 231280 270555 231286 270607
rect 231338 270595 231344 270607
rect 328432 270595 328438 270607
rect 231338 270567 328438 270595
rect 231338 270555 231344 270567
rect 328432 270555 328438 270567
rect 328490 270555 328496 270607
rect 368464 270555 368470 270607
rect 368522 270595 368528 270607
rect 368752 270595 368758 270607
rect 368522 270567 368758 270595
rect 368522 270555 368528 270567
rect 368752 270555 368758 270567
rect 368810 270555 368816 270607
rect 372496 270555 372502 270607
rect 372554 270595 372560 270607
rect 387280 270595 387286 270607
rect 372554 270567 387286 270595
rect 372554 270555 372560 270567
rect 387280 270555 387286 270567
rect 387338 270555 387344 270607
rect 387376 270555 387382 270607
rect 387434 270595 387440 270607
rect 561808 270595 561814 270607
rect 387434 270567 561814 270595
rect 387434 270555 387440 270567
rect 561808 270555 561814 270567
rect 561866 270555 561872 270607
rect 221968 270481 221974 270533
rect 222026 270521 222032 270533
rect 256144 270521 256150 270533
rect 222026 270493 256150 270521
rect 222026 270481 222032 270493
rect 256144 270481 256150 270493
rect 256202 270481 256208 270533
rect 292144 270481 292150 270533
rect 292202 270521 292208 270533
rect 304912 270521 304918 270533
rect 292202 270493 304918 270521
rect 292202 270481 292208 270493
rect 304912 270481 304918 270493
rect 304970 270481 304976 270533
rect 316720 270481 316726 270533
rect 316778 270521 316784 270533
rect 370000 270521 370006 270533
rect 316778 270493 370006 270521
rect 316778 270481 316784 270493
rect 370000 270481 370006 270493
rect 370058 270481 370064 270533
rect 371440 270481 371446 270533
rect 371498 270521 371504 270533
rect 454768 270521 454774 270533
rect 371498 270493 454774 270521
rect 371498 270481 371504 270493
rect 454768 270481 454774 270493
rect 454826 270481 454832 270533
rect 548560 270481 548566 270533
rect 548618 270521 548624 270533
rect 575824 270521 575830 270533
rect 548618 270493 575830 270521
rect 548618 270481 548624 270493
rect 575824 270481 575830 270493
rect 575882 270481 575888 270533
rect 203824 270407 203830 270459
rect 203882 270447 203888 270459
rect 270928 270447 270934 270459
rect 203882 270419 270934 270447
rect 203882 270407 203888 270419
rect 270928 270407 270934 270419
rect 270986 270407 270992 270459
rect 307792 270407 307798 270459
rect 307850 270447 307856 270459
rect 503536 270447 503542 270459
rect 307850 270419 503542 270447
rect 307850 270407 307856 270419
rect 503536 270407 503542 270419
rect 503594 270407 503600 270459
rect 245296 270333 245302 270385
rect 245354 270373 245360 270385
rect 445264 270373 445270 270385
rect 245354 270345 445270 270373
rect 245354 270333 245360 270345
rect 445264 270333 445270 270345
rect 445322 270333 445328 270385
rect 232816 270259 232822 270311
rect 232874 270299 232880 270311
rect 328336 270299 328342 270311
rect 232874 270271 328342 270299
rect 232874 270259 232880 270271
rect 328336 270259 328342 270271
rect 328394 270259 328400 270311
rect 328432 270259 328438 270311
rect 328490 270299 328496 270311
rect 331120 270299 331126 270311
rect 328490 270271 331126 270299
rect 328490 270259 328496 270271
rect 331120 270259 331126 270271
rect 331178 270259 331184 270311
rect 331216 270259 331222 270311
rect 331274 270299 331280 270311
rect 339856 270299 339862 270311
rect 331274 270271 339862 270299
rect 331274 270259 331280 270271
rect 339856 270259 339862 270271
rect 339914 270259 339920 270311
rect 357616 270259 357622 270311
rect 357674 270299 357680 270311
rect 366736 270299 366742 270311
rect 357674 270271 366742 270299
rect 357674 270259 357680 270271
rect 366736 270259 366742 270271
rect 366794 270259 366800 270311
rect 367024 270259 367030 270311
rect 367082 270299 367088 270311
rect 371632 270299 371638 270311
rect 367082 270271 371638 270299
rect 367082 270259 367088 270271
rect 371632 270259 371638 270271
rect 371690 270259 371696 270311
rect 373360 270259 373366 270311
rect 373418 270299 373424 270311
rect 387184 270299 387190 270311
rect 373418 270271 387190 270299
rect 373418 270259 373424 270271
rect 387184 270259 387190 270271
rect 387242 270259 387248 270311
rect 387376 270259 387382 270311
rect 387434 270299 387440 270311
rect 568912 270299 568918 270311
rect 387434 270271 568918 270299
rect 387434 270259 387440 270271
rect 568912 270259 568918 270271
rect 568970 270259 568976 270311
rect 233968 270185 233974 270237
rect 234026 270225 234032 270237
rect 352432 270225 352438 270237
rect 234026 270197 352438 270225
rect 234026 270185 234032 270197
rect 352432 270185 352438 270197
rect 352490 270185 352496 270237
rect 358480 270185 358486 270237
rect 358538 270225 358544 270237
rect 373456 270225 373462 270237
rect 358538 270197 373462 270225
rect 358538 270185 358544 270197
rect 373456 270185 373462 270197
rect 373514 270185 373520 270237
rect 373552 270185 373558 270237
rect 373610 270225 373616 270237
rect 387088 270225 387094 270237
rect 373610 270197 387094 270225
rect 373610 270185 373616 270197
rect 387088 270185 387094 270197
rect 387146 270185 387152 270237
rect 387280 270185 387286 270237
rect 387338 270225 387344 270237
rect 576112 270225 576118 270237
rect 387338 270197 576118 270225
rect 387338 270185 387344 270197
rect 576112 270185 576118 270197
rect 576170 270185 576176 270237
rect 245872 270111 245878 270163
rect 245930 270151 245936 270163
rect 452368 270151 452374 270163
rect 245930 270123 452374 270151
rect 245930 270111 245936 270123
rect 452368 270111 452374 270123
rect 452426 270111 452432 270163
rect 234544 270037 234550 270089
rect 234602 270077 234608 270089
rect 359632 270077 359638 270089
rect 234602 270049 359638 270077
rect 234602 270037 234608 270049
rect 359632 270037 359638 270049
rect 359690 270037 359696 270089
rect 363088 270037 363094 270089
rect 363146 270077 363152 270089
rect 386992 270077 386998 270089
rect 363146 270049 386998 270077
rect 363146 270037 363152 270049
rect 386992 270037 386998 270049
rect 387050 270037 387056 270089
rect 387184 270037 387190 270089
rect 387242 270077 387248 270089
rect 583216 270077 583222 270089
rect 387242 270049 583222 270077
rect 387242 270037 387248 270049
rect 583216 270037 583222 270049
rect 583274 270037 583280 270089
rect 158608 269963 158614 270015
rect 158666 270003 158672 270015
rect 161200 270003 161206 270015
rect 158666 269975 161206 270003
rect 158666 269963 158672 269975
rect 161200 269963 161206 269975
rect 161258 269963 161264 270015
rect 194320 269963 194326 270015
rect 194378 270003 194384 270015
rect 318448 270003 318454 270015
rect 194378 269975 318454 270003
rect 194378 269963 194384 269975
rect 318448 269963 318454 269975
rect 318506 269963 318512 270015
rect 318544 269963 318550 270015
rect 318602 270003 318608 270015
rect 323344 270003 323350 270015
rect 318602 269975 323350 270003
rect 318602 269963 318608 269975
rect 323344 269963 323350 269975
rect 323402 269963 323408 270015
rect 323440 269963 323446 270015
rect 323498 270003 323504 270015
rect 366640 270003 366646 270015
rect 323498 269975 366646 270003
rect 323498 269963 323504 269975
rect 366640 269963 366646 269975
rect 366698 269963 366704 270015
rect 366736 269963 366742 270015
rect 366794 270003 366800 270015
rect 373744 270003 373750 270015
rect 366794 269975 373750 270003
rect 366794 269963 366800 269975
rect 373744 269963 373750 269975
rect 373802 269963 373808 270015
rect 374032 269963 374038 270015
rect 374090 270003 374096 270015
rect 374512 270003 374518 270015
rect 374090 269975 374518 270003
rect 374090 269963 374096 269975
rect 374512 269963 374518 269975
rect 374570 269963 374576 270015
rect 374896 269963 374902 270015
rect 374954 270003 374960 270015
rect 379120 270003 379126 270015
rect 374954 269975 379126 270003
rect 374954 269963 374960 269975
rect 379120 269963 379126 269975
rect 379178 269963 379184 270015
rect 379216 269963 379222 270015
rect 379274 270003 379280 270015
rect 386896 270003 386902 270015
rect 379274 269975 386902 270003
rect 379274 269963 379280 269975
rect 386896 269963 386902 269975
rect 386954 269963 386960 270015
rect 387088 269963 387094 270015
rect 387146 270003 387152 270015
rect 586768 270003 586774 270015
rect 387146 269975 586774 270003
rect 387146 269963 387152 269975
rect 586768 269963 586774 269975
rect 586826 269963 586832 270015
rect 247024 269889 247030 269941
rect 247082 269929 247088 269941
rect 459568 269929 459574 269941
rect 247082 269901 459574 269929
rect 247082 269889 247088 269901
rect 459568 269889 459574 269901
rect 459626 269889 459632 269941
rect 172912 269815 172918 269867
rect 172970 269855 172976 269867
rect 175600 269855 175606 269867
rect 172970 269827 175606 269855
rect 172970 269815 172976 269827
rect 175600 269815 175606 269827
rect 175658 269815 175664 269867
rect 226960 269815 226966 269867
rect 227018 269855 227024 269867
rect 295408 269855 295414 269867
rect 227018 269827 295414 269855
rect 227018 269815 227024 269827
rect 295408 269815 295414 269827
rect 295466 269815 295472 269867
rect 310384 269815 310390 269867
rect 310442 269855 310448 269867
rect 524944 269855 524950 269867
rect 310442 269827 524950 269855
rect 310442 269815 310448 269827
rect 524944 269815 524950 269827
rect 525002 269815 525008 269867
rect 247600 269741 247606 269793
rect 247658 269781 247664 269793
rect 466576 269781 466582 269793
rect 247658 269753 466582 269781
rect 247658 269741 247664 269753
rect 466576 269741 466582 269753
rect 466634 269741 466640 269793
rect 660976 269741 660982 269793
rect 661034 269781 661040 269793
rect 674704 269781 674710 269793
rect 661034 269753 674710 269781
rect 661034 269741 661040 269753
rect 674704 269741 674710 269753
rect 674762 269741 674768 269793
rect 235696 269667 235702 269719
rect 235754 269707 235760 269719
rect 357616 269707 357622 269719
rect 235754 269679 357622 269707
rect 235754 269667 235760 269679
rect 357616 269667 357622 269679
rect 357674 269667 357680 269719
rect 358576 269667 358582 269719
rect 358634 269707 358640 269719
rect 375664 269707 375670 269719
rect 358634 269679 375670 269707
rect 358634 269667 358640 269679
rect 375664 269667 375670 269679
rect 375722 269667 375728 269719
rect 375760 269667 375766 269719
rect 375818 269707 375824 269719
rect 379024 269707 379030 269719
rect 375818 269679 379030 269707
rect 375818 269667 375824 269679
rect 379024 269667 379030 269679
rect 379082 269667 379088 269719
rect 379120 269667 379126 269719
rect 379178 269707 379184 269719
rect 597520 269707 597526 269719
rect 379178 269679 597526 269707
rect 379178 269667 379184 269679
rect 597520 269667 597526 269679
rect 597578 269667 597584 269719
rect 174064 269593 174070 269645
rect 174122 269633 174128 269645
rect 175504 269633 175510 269645
rect 174122 269605 175510 269633
rect 174122 269593 174128 269605
rect 175504 269593 175510 269605
rect 175562 269593 175568 269645
rect 248560 269593 248566 269645
rect 248618 269633 248624 269645
rect 473776 269633 473782 269645
rect 248618 269605 473782 269633
rect 248618 269593 248624 269605
rect 473776 269593 473782 269605
rect 473834 269593 473840 269645
rect 236272 269519 236278 269571
rect 236330 269559 236336 269571
rect 358480 269559 358486 269571
rect 236330 269531 358486 269559
rect 236330 269519 236336 269531
rect 358480 269519 358486 269531
rect 358538 269519 358544 269571
rect 368464 269519 368470 269571
rect 368522 269559 368528 269571
rect 372976 269559 372982 269571
rect 368522 269531 372982 269559
rect 368522 269519 368528 269531
rect 372976 269519 372982 269531
rect 373034 269519 373040 269571
rect 374416 269519 374422 269571
rect 374474 269559 374480 269571
rect 378928 269559 378934 269571
rect 374474 269531 378934 269559
rect 374474 269519 374480 269531
rect 378928 269519 378934 269531
rect 378986 269519 378992 269571
rect 379024 269519 379030 269571
rect 379082 269559 379088 269571
rect 604624 269559 604630 269571
rect 379082 269531 604630 269559
rect 379082 269519 379088 269531
rect 604624 269519 604630 269531
rect 604682 269519 604688 269571
rect 227536 269445 227542 269497
rect 227594 269485 227600 269497
rect 302512 269485 302518 269497
rect 227594 269457 302518 269485
rect 227594 269445 227600 269457
rect 302512 269445 302518 269457
rect 302570 269445 302576 269497
rect 312592 269445 312598 269497
rect 312650 269485 312656 269497
rect 542800 269485 542806 269497
rect 312650 269457 542806 269485
rect 312650 269445 312656 269457
rect 542800 269445 542806 269457
rect 542858 269445 542864 269497
rect 249616 269371 249622 269423
rect 249674 269411 249680 269423
rect 481360 269411 481366 269423
rect 249674 269383 481366 269411
rect 249674 269371 249680 269383
rect 481360 269371 481366 269383
rect 481418 269371 481424 269423
rect 228496 269297 228502 269349
rect 228554 269337 228560 269349
rect 309712 269337 309718 269349
rect 228554 269309 309718 269337
rect 228554 269297 228560 269309
rect 309712 269297 309718 269309
rect 309770 269297 309776 269349
rect 313840 269297 313846 269349
rect 313898 269337 313904 269349
rect 553456 269337 553462 269349
rect 313898 269309 553462 269337
rect 313898 269297 313904 269309
rect 553456 269297 553462 269309
rect 553514 269297 553520 269349
rect 221488 269223 221494 269275
rect 221546 269263 221552 269275
rect 251248 269263 251254 269275
rect 221546 269235 251254 269263
rect 221546 269223 221552 269235
rect 251248 269223 251254 269235
rect 251306 269223 251312 269275
rect 251344 269223 251350 269275
rect 251402 269263 251408 269275
rect 495184 269263 495190 269275
rect 251402 269235 495190 269263
rect 251402 269223 251408 269235
rect 495184 269223 495190 269235
rect 495242 269223 495248 269275
rect 242608 269149 242614 269201
rect 242666 269189 242672 269201
rect 423856 269189 423862 269201
rect 242666 269161 423862 269189
rect 242666 269149 242672 269161
rect 423856 269149 423862 269161
rect 423914 269149 423920 269201
rect 486640 269189 486646 269201
rect 466594 269161 486646 269189
rect 241552 269075 241558 269127
rect 241610 269115 241616 269127
rect 416656 269115 416662 269127
rect 241610 269087 416662 269115
rect 241610 269075 241616 269087
rect 416656 269075 416662 269087
rect 416714 269075 416720 269127
rect 240880 269001 240886 269053
rect 240938 269041 240944 269053
rect 409552 269041 409558 269053
rect 240938 269013 409558 269041
rect 240938 269001 240944 269013
rect 409552 269001 409558 269013
rect 409610 269001 409616 269053
rect 416272 269001 416278 269053
rect 416330 269041 416336 269053
rect 466594 269041 466622 269161
rect 486640 269149 486646 269161
rect 486698 269149 486704 269201
rect 663952 269149 663958 269201
rect 664010 269189 664016 269201
rect 674704 269189 674710 269201
rect 664010 269161 674710 269189
rect 664010 269149 664016 269161
rect 674704 269149 674710 269161
rect 674762 269149 674768 269201
rect 416330 269013 466622 269041
rect 416330 269001 416336 269013
rect 486640 269001 486646 269053
rect 486698 269041 486704 269053
rect 518320 269041 518326 269053
rect 486698 269013 489662 269041
rect 486698 269001 486704 269013
rect 489634 268979 489662 269013
rect 515554 269013 518326 269041
rect 230224 268927 230230 268979
rect 230282 268967 230288 268979
rect 230282 268939 316478 268967
rect 230282 268927 230288 268939
rect 229552 268853 229558 268905
rect 229610 268893 229616 268905
rect 316336 268893 316342 268905
rect 229610 268865 316342 268893
rect 229610 268853 229616 268865
rect 316336 268853 316342 268865
rect 316394 268853 316400 268905
rect 316450 268893 316478 268939
rect 317968 268927 317974 268979
rect 318026 268967 318032 268979
rect 337264 268967 337270 268979
rect 318026 268939 337270 268967
rect 318026 268927 318032 268939
rect 337264 268927 337270 268939
rect 337322 268927 337328 268979
rect 349072 268927 349078 268979
rect 349130 268967 349136 268979
rect 369808 268967 369814 268979
rect 349130 268939 369814 268967
rect 349130 268927 349136 268939
rect 369808 268927 369814 268939
rect 369866 268927 369872 268979
rect 371344 268927 371350 268979
rect 371402 268967 371408 268979
rect 378448 268967 378454 268979
rect 371402 268939 378454 268967
rect 371402 268927 371408 268939
rect 378448 268927 378454 268939
rect 378506 268927 378512 268979
rect 385552 268967 385558 268979
rect 378562 268939 385558 268967
rect 318256 268893 318262 268905
rect 316450 268865 318262 268893
rect 318256 268853 318262 268865
rect 318314 268853 318320 268905
rect 318352 268853 318358 268905
rect 318410 268893 318416 268905
rect 337840 268893 337846 268905
rect 318410 268865 337846 268893
rect 318410 268853 318416 268865
rect 337840 268853 337846 268865
rect 337898 268853 337904 268905
rect 351760 268853 351766 268905
rect 351818 268893 351824 268905
rect 378562 268893 378590 268939
rect 385552 268927 385558 268939
rect 385610 268927 385616 268979
rect 386992 268927 386998 268979
rect 387050 268967 387056 268979
rect 388528 268967 388534 268979
rect 387050 268939 388534 268967
rect 387050 268927 387056 268939
rect 388528 268927 388534 268939
rect 388586 268927 388592 268979
rect 388720 268927 388726 268979
rect 388778 268927 388784 268979
rect 388816 268927 388822 268979
rect 388874 268927 388880 268979
rect 489616 268927 489622 268979
rect 489674 268927 489680 268979
rect 489712 268927 489718 268979
rect 489770 268967 489776 268979
rect 515554 268967 515582 269013
rect 518320 269001 518326 269013
rect 518378 269001 518384 269053
rect 536848 269041 536854 269053
rect 535618 269013 536854 269041
rect 489770 268939 515582 268967
rect 489770 268927 489776 268939
rect 518416 268927 518422 268979
rect 518474 268967 518480 268979
rect 535618 268967 535646 269013
rect 536848 269001 536854 269013
rect 536906 269001 536912 269053
rect 518474 268939 535646 268967
rect 518474 268927 518480 268939
rect 351818 268865 378590 268893
rect 351818 268853 351824 268865
rect 378640 268853 378646 268905
rect 378698 268893 378704 268905
rect 388738 268893 388766 268927
rect 378698 268865 388766 268893
rect 388834 268893 388862 268927
rect 529744 268893 529750 268905
rect 388834 268865 529750 268893
rect 378698 268853 378704 268865
rect 529744 268853 529750 268865
rect 529802 268853 529808 268905
rect 240016 268779 240022 268831
rect 240074 268819 240080 268831
rect 378544 268819 378550 268831
rect 240074 268791 378550 268819
rect 240074 268779 240080 268791
rect 378544 268779 378550 268791
rect 378602 268779 378608 268831
rect 416272 268819 416278 268831
rect 378658 268791 416278 268819
rect 225808 268705 225814 268757
rect 225866 268745 225872 268757
rect 288208 268745 288214 268757
rect 225866 268717 288214 268745
rect 225866 268705 225872 268717
rect 288208 268705 288214 268717
rect 288266 268705 288272 268757
rect 290608 268705 290614 268757
rect 290666 268745 290672 268757
rect 317968 268745 317974 268757
rect 290666 268717 317974 268745
rect 290666 268705 290672 268717
rect 317968 268705 317974 268717
rect 318026 268705 318032 268757
rect 318256 268705 318262 268757
rect 318314 268745 318320 268757
rect 334960 268745 334966 268757
rect 318314 268717 334966 268745
rect 318314 268705 318320 268717
rect 334960 268705 334966 268717
rect 335018 268705 335024 268757
rect 335056 268705 335062 268757
rect 335114 268745 335120 268757
rect 348016 268745 348022 268757
rect 335114 268717 348022 268745
rect 335114 268705 335120 268717
rect 348016 268705 348022 268717
rect 348074 268705 348080 268757
rect 367504 268705 367510 268757
rect 367562 268745 367568 268757
rect 378658 268745 378686 268791
rect 416272 268779 416278 268791
rect 416330 268779 416336 268831
rect 367562 268717 378686 268745
rect 367562 268705 367568 268717
rect 378736 268705 378742 268757
rect 378794 268745 378800 268757
rect 526096 268745 526102 268757
rect 378794 268717 526102 268745
rect 378794 268705 378800 268717
rect 526096 268705 526102 268717
rect 526154 268705 526160 268757
rect 238864 268631 238870 268683
rect 238922 268671 238928 268683
rect 378352 268671 378358 268683
rect 238922 268643 378358 268671
rect 238922 268631 238928 268643
rect 378352 268631 378358 268643
rect 378410 268631 378416 268683
rect 378466 268643 388862 268671
rect 238288 268557 238294 268609
rect 238346 268597 238352 268609
rect 366736 268597 366742 268609
rect 238346 268569 366742 268597
rect 238346 268557 238352 268569
rect 366736 268557 366742 268569
rect 366794 268557 366800 268609
rect 370768 268557 370774 268609
rect 370826 268597 370832 268609
rect 376816 268597 376822 268609
rect 370826 268569 376822 268597
rect 370826 268557 370832 268569
rect 376816 268557 376822 268569
rect 376874 268557 376880 268609
rect 377008 268557 377014 268609
rect 377066 268597 377072 268609
rect 378466 268597 378494 268643
rect 377066 268569 378494 268597
rect 377066 268557 377072 268569
rect 378544 268557 378550 268609
rect 378602 268597 378608 268609
rect 388432 268597 388438 268609
rect 378602 268569 388438 268597
rect 378602 268557 378608 268569
rect 388432 268557 388438 268569
rect 388490 268557 388496 268609
rect 237136 268483 237142 268535
rect 237194 268523 237200 268535
rect 358576 268523 358582 268535
rect 237194 268495 358582 268523
rect 237194 268483 237200 268495
rect 358576 268483 358582 268495
rect 358634 268483 358640 268535
rect 366544 268483 366550 268535
rect 366602 268523 366608 268535
rect 378640 268523 378646 268535
rect 366602 268495 378646 268523
rect 366602 268483 366608 268495
rect 378640 268483 378646 268495
rect 378698 268483 378704 268535
rect 378832 268483 378838 268535
rect 378890 268523 378896 268535
rect 387280 268523 387286 268535
rect 378890 268495 387286 268523
rect 378890 268483 378896 268495
rect 387280 268483 387286 268495
rect 387338 268483 387344 268535
rect 388528 268483 388534 268535
rect 388586 268523 388592 268535
rect 388834 268523 388862 268643
rect 389200 268631 389206 268683
rect 389258 268671 389264 268683
rect 415120 268671 415126 268683
rect 389258 268643 415126 268671
rect 389258 268631 389264 268643
rect 415120 268631 415126 268643
rect 415178 268631 415184 268683
rect 388912 268557 388918 268609
rect 388970 268597 388976 268609
rect 389392 268597 389398 268609
rect 388970 268569 389398 268597
rect 388970 268557 388976 268569
rect 389392 268557 389398 268569
rect 389450 268557 389456 268609
rect 389488 268557 389494 268609
rect 389546 268597 389552 268609
rect 395344 268597 395350 268609
rect 389546 268569 395350 268597
rect 389546 268557 389552 268569
rect 395344 268557 395350 268569
rect 395402 268557 395408 268609
rect 395440 268557 395446 268609
rect 395498 268597 395504 268609
rect 399568 268597 399574 268609
rect 395498 268569 399574 268597
rect 395498 268557 395504 268569
rect 399568 268557 399574 268569
rect 399626 268557 399632 268609
rect 399280 268523 399286 268535
rect 388586 268495 388670 268523
rect 388834 268495 399286 268523
rect 388586 268483 388592 268495
rect 210928 268409 210934 268461
rect 210986 268449 210992 268461
rect 271984 268449 271990 268461
rect 210986 268421 271990 268449
rect 210986 268409 210992 268421
rect 271984 268409 271990 268421
rect 272042 268409 272048 268461
rect 272752 268409 272758 268461
rect 272810 268449 272816 268461
rect 272810 268421 316766 268449
rect 272810 268409 272816 268421
rect 228784 268335 228790 268387
rect 228842 268375 228848 268387
rect 274192 268375 274198 268387
rect 228842 268347 274198 268375
rect 228842 268335 228848 268347
rect 274192 268335 274198 268347
rect 274250 268335 274256 268387
rect 287056 268335 287062 268387
rect 287114 268375 287120 268387
rect 316738 268375 316766 268421
rect 316912 268409 316918 268461
rect 316970 268449 316976 268461
rect 336496 268449 336502 268461
rect 316970 268421 336502 268449
rect 316970 268409 316976 268421
rect 336496 268409 336502 268421
rect 336554 268409 336560 268461
rect 336592 268409 336598 268461
rect 336650 268449 336656 268461
rect 337360 268449 337366 268461
rect 336650 268421 337366 268449
rect 336650 268409 336656 268421
rect 337360 268409 337366 268421
rect 337418 268409 337424 268461
rect 337744 268409 337750 268461
rect 337802 268449 337808 268461
rect 366448 268449 366454 268461
rect 337802 268421 366454 268449
rect 337802 268409 337808 268421
rect 366448 268409 366454 268421
rect 366506 268409 366512 268461
rect 366640 268409 366646 268461
rect 366698 268449 366704 268461
rect 377872 268449 377878 268461
rect 366698 268421 377878 268449
rect 366698 268409 366704 268421
rect 377872 268409 377878 268421
rect 377930 268409 377936 268461
rect 378928 268409 378934 268461
rect 378986 268449 378992 268461
rect 388432 268449 388438 268461
rect 378986 268421 388438 268449
rect 378986 268409 378992 268421
rect 388432 268409 388438 268421
rect 388490 268409 388496 268461
rect 388642 268449 388670 268495
rect 399280 268483 399286 268495
rect 399338 268483 399344 268535
rect 403696 268483 403702 268535
rect 403754 268523 403760 268535
rect 406096 268523 406102 268535
rect 403754 268495 406102 268523
rect 403754 268483 403760 268495
rect 406096 268483 406102 268495
rect 406154 268483 406160 268535
rect 501136 268449 501142 268461
rect 388642 268421 501142 268449
rect 501136 268409 501142 268421
rect 501194 268409 501200 268461
rect 318256 268375 318262 268387
rect 287114 268347 316670 268375
rect 316738 268347 318262 268375
rect 287114 268335 287120 268347
rect 222544 268261 222550 268313
rect 222602 268301 222608 268313
rect 259696 268301 259702 268313
rect 222602 268273 259702 268301
rect 222602 268261 222608 268273
rect 259696 268261 259702 268273
rect 259754 268261 259760 268313
rect 260080 268261 260086 268313
rect 260138 268301 260144 268313
rect 292144 268301 292150 268313
rect 260138 268273 292150 268301
rect 260138 268261 260144 268273
rect 292144 268261 292150 268273
rect 292202 268261 292208 268313
rect 296656 268261 296662 268313
rect 296714 268301 296720 268313
rect 312688 268301 312694 268313
rect 296714 268273 312694 268301
rect 296714 268261 296720 268273
rect 312688 268261 312694 268273
rect 312746 268261 312752 268313
rect 218032 268187 218038 268239
rect 218090 268227 218096 268239
rect 272656 268227 272662 268239
rect 218090 268199 272662 268227
rect 218090 268187 218096 268199
rect 272656 268187 272662 268199
rect 272714 268187 272720 268239
rect 277648 268187 277654 268239
rect 277706 268227 277712 268239
rect 282256 268227 282262 268239
rect 277706 268199 282262 268227
rect 277706 268187 277712 268199
rect 282256 268187 282262 268199
rect 282314 268187 282320 268239
rect 283504 268187 283510 268239
rect 283562 268227 283568 268239
rect 316528 268227 316534 268239
rect 283562 268199 316534 268227
rect 283562 268187 283568 268199
rect 316528 268187 316534 268199
rect 316586 268187 316592 268239
rect 316642 268227 316670 268347
rect 318256 268335 318262 268347
rect 318314 268335 318320 268387
rect 318544 268335 318550 268387
rect 318602 268375 318608 268387
rect 322960 268375 322966 268387
rect 318602 268347 322966 268375
rect 318602 268335 318608 268347
rect 322960 268335 322966 268347
rect 323018 268335 323024 268387
rect 323056 268335 323062 268387
rect 323114 268375 323120 268387
rect 338320 268375 338326 268387
rect 323114 268347 338326 268375
rect 323114 268335 323120 268347
rect 338320 268335 338326 268347
rect 338378 268335 338384 268387
rect 360976 268335 360982 268387
rect 361034 268375 361040 268387
rect 483280 268375 483286 268387
rect 361034 268347 483286 268375
rect 361034 268335 361040 268347
rect 483280 268335 483286 268347
rect 483338 268335 483344 268387
rect 317104 268261 317110 268313
rect 317162 268301 317168 268313
rect 326704 268301 326710 268313
rect 317162 268273 326710 268301
rect 317162 268261 317168 268273
rect 326704 268261 326710 268273
rect 326762 268261 326768 268313
rect 326800 268261 326806 268313
rect 326858 268301 326864 268313
rect 332272 268301 332278 268313
rect 326858 268273 332278 268301
rect 326858 268261 326864 268273
rect 332272 268261 332278 268273
rect 332330 268261 332336 268313
rect 332560 268261 332566 268313
rect 332618 268301 332624 268313
rect 337456 268301 337462 268313
rect 332618 268273 337462 268301
rect 332618 268261 332624 268273
rect 337456 268261 337462 268273
rect 337514 268261 337520 268313
rect 348496 268261 348502 268313
rect 348554 268301 348560 268313
rect 374320 268301 374326 268313
rect 348554 268273 374326 268301
rect 348554 268261 348560 268273
rect 374320 268261 374326 268273
rect 374378 268261 374384 268313
rect 374416 268261 374422 268313
rect 374474 268301 374480 268313
rect 376336 268301 376342 268313
rect 374474 268273 376342 268301
rect 374474 268261 374480 268273
rect 376336 268261 376342 268273
rect 376394 268261 376400 268313
rect 376816 268261 376822 268313
rect 376874 268301 376880 268313
rect 388720 268301 388726 268313
rect 376874 268273 388726 268301
rect 376874 268261 376880 268273
rect 388720 268261 388726 268273
rect 388778 268261 388784 268313
rect 388816 268261 388822 268313
rect 388874 268301 388880 268313
rect 554704 268301 554710 268313
rect 388874 268273 554710 268301
rect 388874 268261 388880 268273
rect 554704 268261 554710 268273
rect 554762 268261 554768 268313
rect 322576 268227 322582 268239
rect 316642 268199 322582 268227
rect 322576 268187 322582 268199
rect 322634 268187 322640 268239
rect 322864 268187 322870 268239
rect 322922 268227 322928 268239
rect 323920 268227 323926 268239
rect 322922 268199 323926 268227
rect 322922 268187 322928 268199
rect 323920 268187 323926 268199
rect 323978 268187 323984 268239
rect 324016 268187 324022 268239
rect 324074 268227 324080 268239
rect 324496 268227 324502 268239
rect 324074 268199 324502 268227
rect 324074 268187 324080 268199
rect 324496 268187 324502 268199
rect 324554 268187 324560 268239
rect 324592 268187 324598 268239
rect 324650 268227 324656 268239
rect 347536 268227 347542 268239
rect 324650 268199 347542 268227
rect 324650 268187 324656 268199
rect 347536 268187 347542 268199
rect 347594 268187 347600 268239
rect 359440 268187 359446 268239
rect 359498 268227 359504 268239
rect 468976 268227 468982 268239
rect 359498 268199 468982 268227
rect 359498 268187 359504 268199
rect 468976 268187 468982 268199
rect 469034 268187 469040 268239
rect 223216 268113 223222 268165
rect 223274 268153 223280 268165
rect 266800 268153 266806 268165
rect 223274 268125 266806 268153
rect 223274 268113 223280 268125
rect 266800 268113 266806 268125
rect 266858 268113 266864 268165
rect 267376 268113 267382 268165
rect 267434 268153 267440 268165
rect 268048 268153 268054 268165
rect 267434 268125 268054 268153
rect 267434 268113 267440 268125
rect 268048 268113 268054 268125
rect 268106 268113 268112 268165
rect 294544 268113 294550 268165
rect 294602 268153 294608 268165
rect 318352 268153 318358 268165
rect 294602 268125 318358 268153
rect 294602 268113 294608 268125
rect 318352 268113 318358 268125
rect 318410 268113 318416 268165
rect 318448 268113 318454 268165
rect 318506 268153 318512 268165
rect 325648 268153 325654 268165
rect 318506 268125 325654 268153
rect 318506 268113 318512 268125
rect 325648 268113 325654 268125
rect 325706 268113 325712 268165
rect 328432 268113 328438 268165
rect 328490 268153 328496 268165
rect 336976 268153 336982 268165
rect 328490 268125 336982 268153
rect 328490 268113 328496 268125
rect 336976 268113 336982 268125
rect 337034 268113 337040 268165
rect 355696 268113 355702 268165
rect 355754 268153 355760 268165
rect 440464 268153 440470 268165
rect 355754 268125 440470 268153
rect 355754 268113 355760 268125
rect 440464 268113 440470 268125
rect 440522 268113 440528 268165
rect 235888 268039 235894 268091
rect 235946 268079 235952 268091
rect 274864 268079 274870 268091
rect 235946 268051 274870 268079
rect 235946 268039 235952 268051
rect 274864 268039 274870 268051
rect 274922 268039 274928 268091
rect 286000 268039 286006 268091
rect 286058 268079 286064 268091
rect 316240 268079 316246 268091
rect 286058 268051 316246 268079
rect 286058 268039 286064 268051
rect 316240 268039 316246 268051
rect 316298 268039 316304 268091
rect 317104 268039 317110 268091
rect 317162 268079 317168 268091
rect 326992 268079 326998 268091
rect 317162 268051 326998 268079
rect 317162 268039 317168 268051
rect 326992 268039 326998 268051
rect 327050 268039 327056 268091
rect 327760 268039 327766 268091
rect 327818 268079 327824 268091
rect 336400 268079 336406 268091
rect 327818 268051 336406 268079
rect 327818 268039 327824 268051
rect 336400 268039 336406 268051
rect 336458 268039 336464 268091
rect 337360 268039 337366 268091
rect 337418 268079 337424 268091
rect 348592 268079 348598 268091
rect 337418 268051 348598 268079
rect 337418 268039 337424 268051
rect 348592 268039 348598 268051
rect 348650 268039 348656 268091
rect 353968 268039 353974 268091
rect 354026 268079 354032 268091
rect 426256 268079 426262 268091
rect 354026 268051 426262 268079
rect 354026 268039 354032 268051
rect 426256 268039 426262 268051
rect 426314 268039 426320 268091
rect 262000 267965 262006 268017
rect 262058 268005 262064 268017
rect 324016 268005 324022 268017
rect 262058 267977 324022 268005
rect 262058 267965 262064 267977
rect 324016 267965 324022 267977
rect 324074 267965 324080 268017
rect 324112 267965 324118 268017
rect 324170 268005 324176 268017
rect 326608 268005 326614 268017
rect 324170 267977 326614 268005
rect 324170 267965 324176 267977
rect 326608 267965 326614 267977
rect 326666 267965 326672 268017
rect 326704 267965 326710 268017
rect 326762 268005 326768 268017
rect 328240 268005 328246 268017
rect 326762 267977 328246 268005
rect 326762 267965 326768 267977
rect 328240 267965 328246 267977
rect 328298 267965 328304 268017
rect 328336 267965 328342 268017
rect 328394 268005 328400 268017
rect 438064 268005 438070 268017
rect 328394 267977 438070 268005
rect 328394 267965 328400 267977
rect 438064 267965 438070 267977
rect 438122 267965 438128 268017
rect 439120 267965 439126 268017
rect 439178 268005 439184 268017
rect 449104 268005 449110 268017
rect 439178 267977 449110 268005
rect 439178 267965 439184 267977
rect 449104 267965 449110 267977
rect 449162 267965 449168 268017
rect 243088 267891 243094 267943
rect 243146 267931 243152 267943
rect 275728 267931 275734 267943
rect 243146 267903 275734 267931
rect 243146 267891 243152 267903
rect 275728 267891 275734 267903
rect 275786 267891 275792 267943
rect 285040 267891 285046 267943
rect 285098 267931 285104 267943
rect 316144 267931 316150 267943
rect 285098 267903 316150 267931
rect 285098 267891 285104 267903
rect 316144 267891 316150 267903
rect 316202 267891 316208 267943
rect 316240 267891 316246 267943
rect 316298 267931 316304 267943
rect 318544 267931 318550 267943
rect 316298 267903 316862 267931
rect 316298 267891 316304 267903
rect 212272 267817 212278 267869
rect 212330 267857 212336 267869
rect 241072 267857 241078 267869
rect 212330 267829 241078 267857
rect 212330 267817 212336 267829
rect 241072 267817 241078 267829
rect 241130 267817 241136 267869
rect 258544 267817 258550 267869
rect 258602 267857 258608 267869
rect 309616 267857 309622 267869
rect 258602 267829 309622 267857
rect 258602 267817 258608 267829
rect 309616 267817 309622 267829
rect 309674 267817 309680 267869
rect 316834 267857 316862 267903
rect 317794 267903 318550 267931
rect 317794 267857 317822 267903
rect 318544 267891 318550 267903
rect 318602 267891 318608 267943
rect 321328 267891 321334 267943
rect 321386 267931 321392 267943
rect 336592 267931 336598 267943
rect 321386 267903 336598 267931
rect 321386 267891 321392 267903
rect 336592 267891 336598 267903
rect 336650 267891 336656 267943
rect 338320 267891 338326 267943
rect 338378 267931 338384 267943
rect 377008 267931 377014 267943
rect 338378 267903 377014 267931
rect 338378 267891 338384 267903
rect 377008 267891 377014 267903
rect 377066 267891 377072 267943
rect 377872 267891 377878 267943
rect 377930 267931 377936 267943
rect 378256 267931 378262 267943
rect 377930 267903 378262 267931
rect 377930 267891 377936 267903
rect 378256 267891 378262 267903
rect 378314 267891 378320 267943
rect 378544 267891 378550 267943
rect 378602 267931 378608 267943
rect 385456 267931 385462 267943
rect 378602 267903 385462 267931
rect 378602 267891 378608 267903
rect 385456 267891 385462 267903
rect 385514 267891 385520 267943
rect 385552 267891 385558 267943
rect 385610 267931 385616 267943
rect 385610 267903 397502 267931
rect 385610 267891 385616 267903
rect 316834 267829 317822 267857
rect 317872 267817 317878 267869
rect 317930 267857 317936 267869
rect 332560 267857 332566 267869
rect 317930 267829 332566 267857
rect 317930 267817 317936 267829
rect 332560 267817 332566 267829
rect 332618 267817 332624 267869
rect 334096 267817 334102 267869
rect 334154 267857 334160 267869
rect 335056 267857 335062 267869
rect 334154 267829 335062 267857
rect 334154 267817 334160 267829
rect 335056 267817 335062 267829
rect 335114 267817 335120 267869
rect 337456 267817 337462 267869
rect 337514 267857 337520 267869
rect 349072 267857 349078 267869
rect 337514 267829 349078 267857
rect 337514 267817 337520 267829
rect 349072 267817 349078 267829
rect 349130 267817 349136 267869
rect 366352 267817 366358 267869
rect 366410 267857 366416 267869
rect 377968 267857 377974 267869
rect 366410 267829 377974 267857
rect 366410 267817 366416 267829
rect 377968 267817 377974 267829
rect 378026 267817 378032 267869
rect 378352 267817 378358 267869
rect 378410 267857 378416 267869
rect 397264 267857 397270 267869
rect 378410 267829 397270 267857
rect 378410 267817 378416 267829
rect 397264 267817 397270 267829
rect 397322 267817 397328 267869
rect 397474 267857 397502 267903
rect 397552 267891 397558 267943
rect 397610 267931 397616 267943
rect 408784 267931 408790 267943
rect 397610 267903 408790 267931
rect 397610 267891 397616 267903
rect 408784 267891 408790 267903
rect 408842 267891 408848 267943
rect 408400 267857 408406 267869
rect 397474 267829 408406 267857
rect 408400 267817 408406 267829
rect 408458 267817 408464 267869
rect 204976 267743 204982 267795
rect 205034 267783 205040 267795
rect 205034 267755 207422 267783
rect 205034 267743 205040 267755
rect 207394 267635 207422 267755
rect 221776 267743 221782 267795
rect 221834 267783 221840 267795
rect 251920 267783 251926 267795
rect 221834 267755 251926 267783
rect 221834 267743 221840 267755
rect 251920 267743 251926 267755
rect 251978 267743 251984 267795
rect 258640 267743 258646 267795
rect 258698 267783 258704 267795
rect 267472 267783 267478 267795
rect 258698 267755 267478 267783
rect 258698 267743 258704 267755
rect 267472 267743 267478 267755
rect 267530 267743 267536 267795
rect 269296 267743 269302 267795
rect 269354 267783 269360 267795
rect 312016 267783 312022 267795
rect 269354 267755 312022 267783
rect 269354 267743 269360 267755
rect 312016 267743 312022 267755
rect 312074 267743 312080 267795
rect 312112 267743 312118 267795
rect 312170 267783 312176 267795
rect 327760 267783 327766 267795
rect 312170 267755 327766 267783
rect 312170 267743 312176 267755
rect 327760 267743 327766 267755
rect 327818 267743 327824 267795
rect 327856 267743 327862 267795
rect 327914 267783 327920 267795
rect 337744 267783 337750 267795
rect 327914 267755 337750 267783
rect 327914 267743 327920 267755
rect 337744 267743 337750 267755
rect 337802 267743 337808 267795
rect 338032 267743 338038 267795
rect 338090 267783 338096 267795
rect 621232 267783 621238 267795
rect 338090 267755 621238 267783
rect 338090 267743 338096 267755
rect 621232 267743 621238 267755
rect 621290 267743 621296 267795
rect 219568 267669 219574 267721
rect 219626 267709 219632 267721
rect 318256 267709 318262 267721
rect 219626 267681 227246 267709
rect 219626 267669 219632 267681
rect 221776 267635 221782 267647
rect 207394 267607 221782 267635
rect 221776 267595 221782 267607
rect 221834 267595 221840 267647
rect 197200 267521 197206 267573
rect 197258 267561 197264 267573
rect 211504 267561 211510 267573
rect 197258 267533 211510 267561
rect 197258 267521 197264 267533
rect 211504 267521 211510 267533
rect 211562 267521 211568 267573
rect 227218 267413 227246 267681
rect 262114 267681 318262 267709
rect 251920 267595 251926 267647
rect 251978 267635 251984 267647
rect 261808 267635 261814 267647
rect 251978 267607 261814 267635
rect 251978 267595 251984 267607
rect 261808 267595 261814 267607
rect 261866 267595 261872 267647
rect 241840 267521 241846 267573
rect 241898 267561 241904 267573
rect 262114 267561 262142 267681
rect 318256 267669 318262 267681
rect 318314 267669 318320 267721
rect 326896 267709 326902 267721
rect 319138 267681 326902 267709
rect 267472 267595 267478 267647
rect 267530 267635 267536 267647
rect 267760 267635 267766 267647
rect 267530 267607 267766 267635
rect 267530 267595 267536 267607
rect 267760 267595 267766 267607
rect 267818 267595 267824 267647
rect 287728 267595 287734 267647
rect 287786 267635 287792 267647
rect 318448 267635 318454 267647
rect 287786 267607 318454 267635
rect 287786 267595 287792 267607
rect 318448 267595 318454 267607
rect 318506 267595 318512 267647
rect 241898 267533 262142 267561
rect 241898 267521 241904 267533
rect 279952 267521 279958 267573
rect 280010 267561 280016 267573
rect 317104 267561 317110 267573
rect 280010 267533 317110 267561
rect 280010 267521 280016 267533
rect 317104 267521 317110 267533
rect 317162 267521 317168 267573
rect 317200 267521 317206 267573
rect 317258 267561 317264 267573
rect 319138 267561 319166 267681
rect 326896 267669 326902 267681
rect 326954 267669 326960 267721
rect 326992 267669 326998 267721
rect 327050 267709 327056 267721
rect 336112 267709 336118 267721
rect 327050 267681 336118 267709
rect 327050 267669 327056 267681
rect 336112 267669 336118 267681
rect 336170 267669 336176 267721
rect 336208 267669 336214 267721
rect 336266 267709 336272 267721
rect 357328 267709 357334 267721
rect 336266 267681 357334 267709
rect 336266 267669 336272 267681
rect 357328 267669 357334 267681
rect 357386 267669 357392 267721
rect 357424 267669 357430 267721
rect 357482 267709 357488 267721
rect 367792 267709 367798 267721
rect 357482 267681 367798 267709
rect 357482 267669 357488 267681
rect 367792 267669 367798 267681
rect 367850 267669 367856 267721
rect 368560 267669 368566 267721
rect 368618 267709 368624 267721
rect 368618 267681 378686 267709
rect 368618 267669 368624 267681
rect 319216 267595 319222 267647
rect 319274 267635 319280 267647
rect 326800 267635 326806 267647
rect 319274 267607 326806 267635
rect 319274 267595 319280 267607
rect 326800 267595 326806 267607
rect 326858 267595 326864 267647
rect 327088 267595 327094 267647
rect 327146 267635 327152 267647
rect 344848 267635 344854 267647
rect 327146 267607 344854 267635
rect 327146 267595 327152 267607
rect 344848 267595 344854 267607
rect 344906 267595 344912 267647
rect 351280 267595 351286 267647
rect 351338 267635 351344 267647
rect 351338 267607 375134 267635
rect 351338 267595 351344 267607
rect 317258 267533 319166 267561
rect 317258 267521 317264 267533
rect 322480 267521 322486 267573
rect 322538 267561 322544 267573
rect 338032 267561 338038 267573
rect 322538 267533 338038 267561
rect 322538 267521 322544 267533
rect 338032 267521 338038 267533
rect 338090 267521 338096 267573
rect 353296 267521 353302 267573
rect 353354 267561 353360 267573
rect 374992 267561 374998 267573
rect 353354 267533 374998 267561
rect 353354 267521 353360 267533
rect 374992 267521 374998 267533
rect 375050 267521 375056 267573
rect 256144 267447 256150 267499
rect 256202 267487 256208 267499
rect 269008 267487 269014 267499
rect 256202 267459 269014 267487
rect 256202 267447 256208 267459
rect 269008 267447 269014 267459
rect 269066 267447 269072 267499
rect 338320 267487 338326 267499
rect 297058 267459 338326 267487
rect 241840 267413 241846 267425
rect 227218 267385 241846 267413
rect 241840 267373 241846 267385
rect 241898 267373 241904 267425
rect 261808 267373 261814 267425
rect 261866 267413 261872 267425
rect 269296 267413 269302 267425
rect 261866 267385 269302 267413
rect 261866 267373 261872 267385
rect 269296 267373 269302 267385
rect 269354 267373 269360 267425
rect 290320 267373 290326 267425
rect 290378 267413 290384 267425
rect 297058 267413 297086 267459
rect 338320 267447 338326 267459
rect 338378 267447 338384 267499
rect 355024 267447 355030 267499
rect 355082 267487 355088 267499
rect 355082 267459 367166 267487
rect 355082 267447 355088 267459
rect 290378 267385 297086 267413
rect 290378 267373 290384 267385
rect 297136 267373 297142 267425
rect 297194 267413 297200 267425
rect 346576 267413 346582 267425
rect 297194 267385 346582 267413
rect 297194 267373 297200 267385
rect 346576 267373 346582 267385
rect 346634 267373 346640 267425
rect 347248 267373 347254 267425
rect 347306 267413 347312 267425
rect 365200 267413 365206 267425
rect 347306 267385 365206 267413
rect 347306 267373 347312 267385
rect 365200 267373 365206 267385
rect 365258 267373 365264 267425
rect 367138 267413 367166 267459
rect 367792 267447 367798 267499
rect 367850 267487 367856 267499
rect 368752 267487 368758 267499
rect 367850 267459 368758 267487
rect 367850 267447 367856 267459
rect 368752 267447 368758 267459
rect 368810 267447 368816 267499
rect 369136 267447 369142 267499
rect 369194 267487 369200 267499
rect 374800 267487 374806 267499
rect 369194 267459 374806 267487
rect 369194 267447 369200 267459
rect 374800 267447 374806 267459
rect 374858 267447 374864 267499
rect 375106 267487 375134 267607
rect 375184 267595 375190 267647
rect 375242 267635 375248 267647
rect 376816 267635 376822 267647
rect 375242 267607 376822 267635
rect 375242 267595 375248 267607
rect 376816 267595 376822 267607
rect 376874 267595 376880 267647
rect 376912 267595 376918 267647
rect 376970 267635 376976 267647
rect 378352 267635 378358 267647
rect 376970 267607 378358 267635
rect 376970 267595 376976 267607
rect 378352 267595 378358 267607
rect 378410 267595 378416 267647
rect 378658 267635 378686 267681
rect 378832 267669 378838 267721
rect 378890 267709 378896 267721
rect 400048 267709 400054 267721
rect 378890 267681 400054 267709
rect 378890 267669 378896 267681
rect 400048 267669 400054 267681
rect 400106 267669 400112 267721
rect 401680 267669 401686 267721
rect 401738 267709 401744 267721
rect 412816 267709 412822 267721
rect 401738 267681 412822 267709
rect 401738 267669 401744 267681
rect 412816 267669 412822 267681
rect 412874 267669 412880 267721
rect 397456 267635 397462 267647
rect 378658 267607 397462 267635
rect 397456 267595 397462 267607
rect 397514 267595 397520 267647
rect 397552 267595 397558 267647
rect 397610 267635 397616 267647
rect 404656 267635 404662 267647
rect 397610 267607 404662 267635
rect 397610 267595 397616 267607
rect 404656 267595 404662 267607
rect 404714 267595 404720 267647
rect 375376 267521 375382 267573
rect 375434 267561 375440 267573
rect 419056 267561 419062 267573
rect 375434 267533 419062 267561
rect 375434 267521 375440 267533
rect 419056 267521 419062 267533
rect 419114 267521 419120 267573
rect 397552 267487 397558 267499
rect 375106 267459 397558 267487
rect 397552 267447 397558 267459
rect 397610 267447 397616 267499
rect 397648 267447 397654 267499
rect 397706 267487 397712 267499
rect 398800 267487 398806 267499
rect 397706 267459 398806 267487
rect 397706 267447 397712 267459
rect 398800 267447 398806 267459
rect 398858 267447 398864 267499
rect 398896 267447 398902 267499
rect 398954 267487 398960 267499
rect 414352 267487 414358 267499
rect 398954 267459 414358 267487
rect 398954 267447 398960 267459
rect 414352 267447 414358 267459
rect 414410 267447 414416 267499
rect 433360 267413 433366 267425
rect 367138 267385 433366 267413
rect 433360 267373 433366 267385
rect 433418 267373 433424 267425
rect 291664 267299 291670 267351
rect 291722 267339 291728 267351
rect 367024 267339 367030 267351
rect 291722 267311 367030 267339
rect 291722 267299 291728 267311
rect 367024 267299 367030 267311
rect 367082 267299 367088 267351
rect 367120 267299 367126 267351
rect 367178 267339 367184 267351
rect 378352 267339 378358 267351
rect 367178 267311 378358 267339
rect 367178 267299 367184 267311
rect 378352 267299 378358 267311
rect 378410 267299 378416 267351
rect 378448 267299 378454 267351
rect 378506 267339 378512 267351
rect 385840 267339 385846 267351
rect 378506 267311 385846 267339
rect 378506 267299 378512 267311
rect 385840 267299 385846 267311
rect 385898 267299 385904 267351
rect 387472 267299 387478 267351
rect 387530 267339 387536 267351
rect 608176 267339 608182 267351
rect 387530 267311 608182 267339
rect 387530 267299 387536 267311
rect 608176 267299 608182 267311
rect 608234 267299 608240 267351
rect 289456 267225 289462 267277
rect 289514 267265 289520 267277
rect 353680 267265 353686 267277
rect 289514 267237 353686 267265
rect 289514 267225 289520 267237
rect 353680 267225 353686 267237
rect 353738 267225 353744 267277
rect 356560 267225 356566 267277
rect 356618 267265 356624 267277
rect 369040 267265 369046 267277
rect 356618 267237 369046 267265
rect 356618 267225 356624 267237
rect 369040 267225 369046 267237
rect 369098 267225 369104 267277
rect 369328 267225 369334 267277
rect 369386 267265 369392 267277
rect 447664 267265 447670 267277
rect 369386 267237 447670 267265
rect 369386 267225 369392 267237
rect 447664 267225 447670 267237
rect 447722 267225 447728 267277
rect 293584 267151 293590 267203
rect 293642 267191 293648 267203
rect 367120 267191 367126 267203
rect 293642 267163 367126 267191
rect 293642 267151 293648 267163
rect 367120 267151 367126 267163
rect 367178 267151 367184 267203
rect 377008 267191 377014 267203
rect 367234 267163 377014 267191
rect 262096 267077 262102 267129
rect 262154 267117 262160 267129
rect 309424 267117 309430 267129
rect 262154 267089 309430 267117
rect 262154 267077 262160 267089
rect 309424 267077 309430 267089
rect 309482 267077 309488 267129
rect 309616 267077 309622 267129
rect 309674 267117 309680 267129
rect 317872 267117 317878 267129
rect 309674 267089 317878 267117
rect 309674 267077 309680 267089
rect 317872 267077 317878 267089
rect 317930 267077 317936 267129
rect 318256 267077 318262 267129
rect 318314 267117 318320 267129
rect 328528 267117 328534 267129
rect 318314 267089 328534 267117
rect 318314 267077 318320 267089
rect 328528 267077 328534 267089
rect 328586 267077 328592 267129
rect 328624 267077 328630 267129
rect 328682 267117 328688 267129
rect 348496 267117 348502 267129
rect 328682 267089 348502 267117
rect 328682 267077 328688 267089
rect 348496 267077 348502 267089
rect 348554 267077 348560 267129
rect 348592 267077 348598 267129
rect 348650 267117 348656 267129
rect 367234 267117 367262 267163
rect 377008 267151 377014 267163
rect 377066 267151 377072 267203
rect 377200 267151 377206 267203
rect 377258 267191 377264 267203
rect 387472 267191 387478 267203
rect 377258 267163 387478 267191
rect 377258 267151 377264 267163
rect 387472 267151 387478 267163
rect 387530 267151 387536 267203
rect 387568 267151 387574 267203
rect 387626 267191 387632 267203
rect 398512 267191 398518 267203
rect 387626 267163 398518 267191
rect 387626 267151 387632 267163
rect 398512 267151 398518 267163
rect 398570 267151 398576 267203
rect 398800 267151 398806 267203
rect 398858 267191 398864 267203
rect 421456 267191 421462 267203
rect 398858 267163 421462 267191
rect 398858 267151 398864 267163
rect 421456 267151 421462 267163
rect 421514 267151 421520 267203
rect 348650 267089 367262 267117
rect 348650 267077 348656 267089
rect 367312 267077 367318 267129
rect 367370 267117 367376 267129
rect 375184 267117 375190 267129
rect 367370 267089 375190 267117
rect 367370 267077 367376 267089
rect 375184 267077 375190 267089
rect 375242 267077 375248 267129
rect 375952 267077 375958 267129
rect 376010 267117 376016 267129
rect 458320 267117 458326 267129
rect 376010 267089 458326 267117
rect 376010 267077 376016 267089
rect 458320 267077 458326 267089
rect 458378 267077 458384 267129
rect 295312 267003 295318 267055
rect 295370 267043 295376 267055
rect 378832 267043 378838 267055
rect 295370 267015 378838 267043
rect 295370 267003 295376 267015
rect 378832 267003 378838 267015
rect 378890 267003 378896 267055
rect 378928 267003 378934 267055
rect 378986 267043 378992 267055
rect 398224 267043 398230 267055
rect 378986 267015 398230 267043
rect 378986 267003 378992 267015
rect 398224 267003 398230 267015
rect 398282 267003 398288 267055
rect 398434 267015 399422 267043
rect 295984 266929 295990 266981
rect 296042 266969 296048 266981
rect 397168 266969 397174 266981
rect 296042 266941 397174 266969
rect 296042 266929 296048 266941
rect 397168 266929 397174 266941
rect 397226 266929 397232 266981
rect 397264 266929 397270 266981
rect 397322 266969 397328 266981
rect 398434 266969 398462 267015
rect 397322 266941 398462 266969
rect 397322 266929 397328 266941
rect 398512 266929 398518 266981
rect 398570 266969 398576 266981
rect 399184 266969 399190 266981
rect 398570 266941 399190 266969
rect 398570 266929 398576 266941
rect 399184 266929 399190 266941
rect 399242 266929 399248 266981
rect 399394 266969 399422 267015
rect 413680 266969 413686 266981
rect 399394 266941 413686 266969
rect 413680 266929 413686 266941
rect 413738 266929 413744 266981
rect 251632 266855 251638 266907
rect 251690 266895 251696 266907
rect 332368 266895 332374 266907
rect 251690 266867 332374 266895
rect 251690 266855 251696 266867
rect 332368 266855 332374 266867
rect 332426 266855 332432 266907
rect 349552 266855 349558 266907
rect 349610 266895 349616 266907
rect 357424 266895 357430 266907
rect 349610 266867 357430 266895
rect 349610 266855 349616 266867
rect 357424 266855 357430 266867
rect 357482 266855 357488 266907
rect 359824 266855 359830 266907
rect 359882 266895 359888 266907
rect 472624 266895 472630 266907
rect 359882 266867 472630 266895
rect 359882 266855 359888 266867
rect 472624 266855 472630 266867
rect 472682 266855 472688 266907
rect 296848 266781 296854 266833
rect 296906 266821 296912 266833
rect 398896 266821 398902 266833
rect 296906 266793 398902 266821
rect 296906 266781 296912 266793
rect 398896 266781 398902 266793
rect 398954 266781 398960 266833
rect 399088 266781 399094 266833
rect 399146 266821 399152 266833
rect 407152 266821 407158 266833
rect 399146 266793 407158 266821
rect 399146 266781 399152 266793
rect 407152 266781 407158 266793
rect 407210 266781 407216 266833
rect 288784 266707 288790 266759
rect 288842 266747 288848 266759
rect 297136 266747 297142 266759
rect 288842 266719 297142 266747
rect 288842 266707 288848 266719
rect 297136 266707 297142 266719
rect 297194 266707 297200 266759
rect 298000 266707 298006 266759
rect 298058 266747 298064 266759
rect 398800 266747 398806 266759
rect 298058 266719 398806 266747
rect 298058 266707 298064 266719
rect 398800 266707 398806 266719
rect 398858 266707 398864 266759
rect 399280 266707 399286 266759
rect 399338 266747 399344 266759
rect 408784 266747 408790 266759
rect 399338 266719 408790 266747
rect 399338 266707 399344 266719
rect 408784 266707 408790 266719
rect 408842 266707 408848 266759
rect 298576 266633 298582 266685
rect 298634 266673 298640 266685
rect 428656 266673 428662 266685
rect 298634 266645 428662 266673
rect 298634 266633 298640 266645
rect 428656 266633 428662 266645
rect 428714 266633 428720 266685
rect 199120 266559 199126 266611
rect 199178 266599 199184 266611
rect 214960 266599 214966 266611
rect 199178 266571 214966 266599
rect 199178 266559 199184 266571
rect 214960 266559 214966 266571
rect 215018 266559 215024 266611
rect 244240 266559 244246 266611
rect 244298 266599 244304 266611
rect 331696 266599 331702 266611
rect 244298 266571 331702 266599
rect 244298 266559 244304 266571
rect 331696 266559 331702 266571
rect 331754 266559 331760 266611
rect 338320 266559 338326 266611
rect 338378 266599 338384 266611
rect 360784 266599 360790 266611
rect 338378 266571 360790 266599
rect 338378 266559 338384 266571
rect 360784 266559 360790 266571
rect 360842 266559 360848 266611
rect 362224 266559 362230 266611
rect 362282 266599 362288 266611
rect 494032 266599 494038 266611
rect 362282 266571 494038 266599
rect 362282 266559 362288 266571
rect 494032 266559 494038 266571
rect 494090 266559 494096 266611
rect 237424 266485 237430 266537
rect 237482 266525 237488 266537
rect 330640 266525 330646 266537
rect 237482 266497 330646 266525
rect 237482 266485 237488 266497
rect 330640 266485 330646 266497
rect 330698 266485 330704 266537
rect 331408 266485 331414 266537
rect 331466 266525 331472 266537
rect 339376 266525 339382 266537
rect 331466 266497 339382 266525
rect 331466 266485 331472 266497
rect 339376 266485 339382 266497
rect 339434 266485 339440 266537
rect 362704 266485 362710 266537
rect 362762 266525 362768 266537
rect 497584 266525 497590 266537
rect 362762 266497 497590 266525
rect 362762 266485 362768 266497
rect 497584 266485 497590 266497
rect 497642 266485 497648 266537
rect 244144 266411 244150 266463
rect 244202 266451 244208 266463
rect 261904 266451 261910 266463
rect 244202 266423 261910 266451
rect 244202 266411 244208 266423
rect 261904 266411 261910 266423
rect 261962 266411 261968 266463
rect 299728 266411 299734 266463
rect 299786 266451 299792 266463
rect 435664 266451 435670 266463
rect 299786 266423 435670 266451
rect 299786 266411 299792 266423
rect 435664 266411 435670 266423
rect 435722 266411 435728 266463
rect 300304 266337 300310 266389
rect 300362 266377 300368 266389
rect 442864 266377 442870 266389
rect 300362 266349 442870 266377
rect 300362 266337 300368 266349
rect 442864 266337 442870 266349
rect 442922 266337 442928 266389
rect 301264 266263 301270 266315
rect 301322 266303 301328 266315
rect 449968 266303 449974 266315
rect 301322 266275 449974 266303
rect 301322 266263 301328 266275
rect 449968 266263 449974 266275
rect 450026 266263 450032 266315
rect 230032 266189 230038 266241
rect 230090 266229 230096 266241
rect 329968 266229 329974 266241
rect 230090 266201 329974 266229
rect 230090 266189 230096 266201
rect 329968 266189 329974 266201
rect 330026 266189 330032 266241
rect 347248 266189 347254 266241
rect 347306 266229 347312 266241
rect 347824 266229 347830 266241
rect 347306 266201 347830 266229
rect 347306 266189 347312 266201
rect 347824 266189 347830 266201
rect 347882 266189 347888 266241
rect 357808 266189 357814 266241
rect 357866 266229 357872 266241
rect 375952 266229 375958 266241
rect 357866 266201 375958 266229
rect 357866 266189 357872 266201
rect 375952 266189 375958 266201
rect 376010 266189 376016 266241
rect 376912 266189 376918 266241
rect 376970 266229 376976 266241
rect 522544 266229 522550 266241
rect 376970 266201 522550 266229
rect 376970 266189 376976 266201
rect 522544 266189 522550 266201
rect 522602 266189 522608 266241
rect 302320 266115 302326 266167
rect 302378 266155 302384 266167
rect 457168 266155 457174 266167
rect 302378 266127 457174 266155
rect 302378 266115 302384 266127
rect 457168 266115 457174 266127
rect 457226 266115 457232 266167
rect 255088 266041 255094 266093
rect 255146 266081 255152 266093
rect 258640 266081 258646 266093
rect 255146 266053 258646 266081
rect 255146 266041 255152 266053
rect 258640 266041 258646 266053
rect 258698 266041 258704 266093
rect 302992 266041 302998 266093
rect 303050 266081 303056 266093
rect 464272 266081 464278 266093
rect 303050 266053 464278 266081
rect 303050 266041 303056 266053
rect 464272 266041 464278 266053
rect 464330 266041 464336 266093
rect 304048 265967 304054 266019
rect 304106 266007 304112 266019
rect 471376 266007 471382 266019
rect 304106 265979 471382 266007
rect 304106 265967 304112 265979
rect 471376 265967 471382 265979
rect 471434 265967 471440 266019
rect 226384 265893 226390 265945
rect 226442 265933 226448 265945
rect 318352 265933 318358 265945
rect 226442 265905 318358 265933
rect 226442 265893 226448 265905
rect 318352 265893 318358 265905
rect 318410 265893 318416 265945
rect 318448 265893 318454 265945
rect 318506 265933 318512 265945
rect 339088 265933 339094 265945
rect 318506 265905 339094 265933
rect 318506 265893 318512 265905
rect 339088 265893 339094 265905
rect 339146 265893 339152 265945
rect 367024 265893 367030 265945
rect 367082 265933 367088 265945
rect 378352 265933 378358 265945
rect 367082 265905 378358 265933
rect 367082 265893 367088 265905
rect 378352 265893 378358 265905
rect 378410 265893 378416 265945
rect 378448 265893 378454 265945
rect 378506 265933 378512 265945
rect 397840 265933 397846 265945
rect 378506 265905 397846 265933
rect 378506 265893 378512 265905
rect 397840 265893 397846 265905
rect 397898 265893 397904 265945
rect 398224 265893 398230 265945
rect 398282 265933 398288 265945
rect 533200 265933 533206 265945
rect 398282 265905 533206 265933
rect 398282 265893 398288 265905
rect 533200 265893 533206 265905
rect 533258 265893 533264 265945
rect 304720 265819 304726 265871
rect 304778 265859 304784 265871
rect 478576 265859 478582 265871
rect 304778 265831 478582 265859
rect 304778 265819 304784 265831
rect 478576 265819 478582 265831
rect 478634 265819 478640 265871
rect 212464 265745 212470 265797
rect 212522 265785 212528 265797
rect 318832 265785 318838 265797
rect 212522 265757 318838 265785
rect 212522 265745 212528 265757
rect 318832 265745 318838 265757
rect 318890 265745 318896 265797
rect 318928 265745 318934 265797
rect 318986 265785 318992 265797
rect 327856 265785 327862 265797
rect 318986 265757 327862 265785
rect 318986 265745 318992 265757
rect 327856 265745 327862 265757
rect 327914 265745 327920 265797
rect 327952 265745 327958 265797
rect 328010 265785 328016 265797
rect 348496 265785 348502 265797
rect 328010 265757 348502 265785
rect 328010 265745 328016 265757
rect 348496 265745 348502 265757
rect 348554 265745 348560 265797
rect 350704 265745 350710 265797
rect 350762 265785 350768 265797
rect 368560 265785 368566 265797
rect 350762 265757 368566 265785
rect 350762 265745 350768 265757
rect 368560 265745 368566 265757
rect 368618 265745 368624 265797
rect 368752 265745 368758 265797
rect 368810 265785 368816 265797
rect 378736 265785 378742 265797
rect 368810 265757 378742 265785
rect 368810 265745 368816 265757
rect 378736 265745 378742 265757
rect 378794 265745 378800 265797
rect 378832 265745 378838 265797
rect 378890 265785 378896 265797
rect 399088 265785 399094 265797
rect 378890 265757 399094 265785
rect 378890 265745 378896 265757
rect 399088 265745 399094 265757
rect 399146 265745 399152 265797
rect 399184 265745 399190 265797
rect 399242 265785 399248 265797
rect 547600 265785 547606 265797
rect 399242 265757 547606 265785
rect 399242 265745 399248 265757
rect 547600 265745 547606 265757
rect 547658 265745 547664 265797
rect 305584 265671 305590 265723
rect 305642 265711 305648 265723
rect 485680 265711 485686 265723
rect 305642 265683 485686 265711
rect 305642 265671 305648 265683
rect 485680 265671 485686 265683
rect 485738 265671 485744 265723
rect 306736 265597 306742 265649
rect 306794 265637 306800 265649
rect 318736 265637 318742 265649
rect 306794 265609 318742 265637
rect 306794 265597 306800 265609
rect 318736 265597 318742 265609
rect 318794 265597 318800 265649
rect 319024 265597 319030 265649
rect 319082 265637 319088 265649
rect 492880 265637 492886 265649
rect 319082 265609 492886 265637
rect 319082 265597 319088 265609
rect 492880 265597 492886 265609
rect 492938 265597 492944 265649
rect 307312 265523 307318 265575
rect 307370 265563 307376 265575
rect 499888 265563 499894 265575
rect 307370 265535 499894 265563
rect 307370 265523 307376 265535
rect 499888 265523 499894 265535
rect 499946 265523 499952 265575
rect 269008 265449 269014 265501
rect 269066 265489 269072 265501
rect 288496 265489 288502 265501
rect 269066 265461 288502 265489
rect 269066 265449 269072 265461
rect 288496 265449 288502 265461
rect 288554 265449 288560 265501
rect 309328 265449 309334 265501
rect 309386 265489 309392 265501
rect 309386 265461 379070 265489
rect 309386 265449 309392 265461
rect 309904 265375 309910 265427
rect 309962 265415 309968 265427
rect 318544 265415 318550 265427
rect 309962 265387 318550 265415
rect 309962 265375 309968 265387
rect 318544 265375 318550 265387
rect 318602 265375 318608 265427
rect 319216 265375 319222 265427
rect 319274 265415 319280 265427
rect 319696 265415 319702 265427
rect 319274 265387 319702 265415
rect 319274 265375 319280 265387
rect 319696 265375 319702 265387
rect 319754 265375 319760 265427
rect 321040 265375 321046 265427
rect 321098 265415 321104 265427
rect 321098 265387 374654 265415
rect 321098 265375 321104 265387
rect 311632 265301 311638 265353
rect 311690 265341 311696 265353
rect 318928 265341 318934 265353
rect 311690 265313 318934 265341
rect 311690 265301 311696 265313
rect 318928 265301 318934 265313
rect 318986 265301 318992 265353
rect 326464 265341 326470 265353
rect 319138 265313 326470 265341
rect 221680 265227 221686 265279
rect 221738 265267 221744 265279
rect 273136 265267 273142 265279
rect 221738 265239 273142 265267
rect 221738 265227 221744 265239
rect 273136 265227 273142 265239
rect 273194 265227 273200 265279
rect 313264 265227 313270 265279
rect 313322 265267 313328 265279
rect 318832 265267 318838 265279
rect 313322 265239 318838 265267
rect 313322 265227 313328 265239
rect 318832 265227 318838 265239
rect 318890 265227 318896 265279
rect 319138 265267 319166 265313
rect 326464 265301 326470 265313
rect 326522 265301 326528 265353
rect 326608 265301 326614 265353
rect 326666 265341 326672 265353
rect 326666 265313 374558 265341
rect 326666 265301 326672 265313
rect 318946 265239 319166 265267
rect 201424 265153 201430 265205
rect 201482 265193 201488 265205
rect 262096 265193 262102 265205
rect 201482 265165 227486 265193
rect 201482 265153 201488 265165
rect 79216 265005 79222 265057
rect 79274 265045 79280 265057
rect 227458 265045 227486 265165
rect 252034 265165 262102 265193
rect 252034 265119 252062 265165
rect 262096 265153 262102 265165
rect 262154 265153 262160 265205
rect 282256 265153 282262 265205
rect 282314 265193 282320 265205
rect 282314 265165 309374 265193
rect 282314 265153 282320 265165
rect 227554 265091 252062 265119
rect 227554 265045 227582 265091
rect 255664 265079 255670 265131
rect 255722 265119 255728 265131
rect 267568 265119 267574 265131
rect 255722 265091 267574 265119
rect 255722 265079 255728 265091
rect 267568 265079 267574 265091
rect 267626 265079 267632 265131
rect 79274 265017 83582 265045
rect 227458 265017 227582 265045
rect 79274 265005 79280 265017
rect 83554 264971 83582 265017
rect 262096 265005 262102 265057
rect 262154 265045 262160 265057
rect 282256 265045 282262 265057
rect 262154 265017 282262 265045
rect 262154 265005 262160 265017
rect 282256 265005 282262 265017
rect 282314 265005 282320 265057
rect 86416 264971 86422 264983
rect 83554 264943 86422 264971
rect 86416 264931 86422 264943
rect 86474 264931 86480 264983
rect 211216 264931 211222 264983
rect 211274 264971 211280 264983
rect 212272 264971 212278 264983
rect 211274 264943 212278 264971
rect 211274 264931 211280 264943
rect 212272 264931 212278 264943
rect 212330 264931 212336 264983
rect 256624 264931 256630 264983
rect 256682 264971 256688 264983
rect 268240 264971 268246 264983
rect 256682 264943 268246 264971
rect 256682 264931 256688 264943
rect 268240 264931 268246 264943
rect 268298 264931 268304 264983
rect 287536 264931 287542 264983
rect 287594 264971 287600 264983
rect 309346 264971 309374 265165
rect 312016 265153 312022 265205
rect 312074 265193 312080 265205
rect 316624 265193 316630 265205
rect 312074 265165 316630 265193
rect 312074 265153 312080 265165
rect 316624 265153 316630 265165
rect 316682 265153 316688 265205
rect 317680 265193 317686 265205
rect 317122 265165 317686 265193
rect 316528 265079 316534 265131
rect 316586 265119 316592 265131
rect 317122 265119 317150 265165
rect 317680 265153 317686 265165
rect 317738 265153 317744 265205
rect 318736 265153 318742 265205
rect 318794 265193 318800 265205
rect 318946 265193 318974 265239
rect 319696 265227 319702 265279
rect 319754 265267 319760 265279
rect 319754 265239 374462 265267
rect 319754 265227 319760 265239
rect 318794 265165 318974 265193
rect 318794 265153 318800 265165
rect 319312 265153 319318 265205
rect 319370 265193 319376 265205
rect 329296 265193 329302 265205
rect 319370 265165 329302 265193
rect 319370 265153 319376 265165
rect 329296 265153 329302 265165
rect 329354 265153 329360 265205
rect 332272 265153 332278 265205
rect 332330 265193 332336 265205
rect 367312 265193 367318 265205
rect 332330 265165 367318 265193
rect 332330 265153 332336 265165
rect 367312 265153 367318 265165
rect 367370 265153 367376 265205
rect 316586 265091 317150 265119
rect 316586 265079 316592 265091
rect 318544 265079 318550 265131
rect 318602 265119 318608 265131
rect 318928 265119 318934 265131
rect 318602 265091 318934 265119
rect 318602 265079 318608 265091
rect 318928 265079 318934 265091
rect 318986 265079 318992 265131
rect 319216 265079 319222 265131
rect 319274 265119 319280 265131
rect 326608 265119 326614 265131
rect 319274 265091 326614 265119
rect 319274 265079 319280 265091
rect 326608 265079 326614 265091
rect 326666 265079 326672 265131
rect 337072 265079 337078 265131
rect 337130 265119 337136 265131
rect 337552 265119 337558 265131
rect 337130 265091 337558 265119
rect 337130 265079 337136 265091
rect 337552 265079 337558 265091
rect 337610 265079 337616 265131
rect 344848 265079 344854 265131
rect 344906 265119 344912 265131
rect 374224 265119 374230 265131
rect 344906 265091 374230 265119
rect 344906 265079 344912 265091
rect 374224 265079 374230 265091
rect 374282 265079 374288 265131
rect 374434 265119 374462 265239
rect 374530 265193 374558 265313
rect 374626 265267 374654 265387
rect 374800 265375 374806 265427
rect 374858 265415 374864 265427
rect 374858 265387 376190 265415
rect 374858 265375 374864 265387
rect 376162 265341 376190 265387
rect 376432 265375 376438 265427
rect 376490 265415 376496 265427
rect 377200 265415 377206 265427
rect 376490 265387 377206 265415
rect 376490 265375 376496 265387
rect 377200 265375 377206 265387
rect 377258 265375 377264 265427
rect 378928 265415 378934 265427
rect 378370 265387 378934 265415
rect 378370 265341 378398 265387
rect 378928 265375 378934 265387
rect 378986 265375 378992 265427
rect 379042 265415 379070 265461
rect 379120 265449 379126 265501
rect 379178 265489 379184 265501
rect 387184 265489 387190 265501
rect 379178 265461 387190 265489
rect 379178 265449 379184 265461
rect 387184 265449 387190 265461
rect 387242 265449 387248 265501
rect 514288 265489 514294 265501
rect 398866 265461 514294 265489
rect 398866 265415 398894 265461
rect 514288 265449 514294 265461
rect 514346 265449 514352 265501
rect 379042 265387 398894 265415
rect 399856 265375 399862 265427
rect 399914 265415 399920 265427
rect 521392 265415 521398 265427
rect 399914 265387 521398 265415
rect 399914 265375 399920 265387
rect 521392 265375 521398 265387
rect 521450 265375 521456 265427
rect 376162 265313 378398 265341
rect 378736 265301 378742 265353
rect 378794 265341 378800 265353
rect 390544 265341 390550 265353
rect 378794 265313 390550 265341
rect 378794 265301 378800 265313
rect 390544 265301 390550 265313
rect 390602 265301 390608 265353
rect 392848 265301 392854 265353
rect 392906 265341 392912 265353
rect 393616 265341 393622 265353
rect 392906 265313 393622 265341
rect 392906 265301 392912 265313
rect 393616 265301 393622 265313
rect 393674 265301 393680 265353
rect 398704 265301 398710 265353
rect 398762 265341 398768 265353
rect 535600 265341 535606 265353
rect 398762 265313 535606 265341
rect 398762 265301 398768 265313
rect 535600 265301 535606 265313
rect 535658 265301 535664 265353
rect 374626 265239 398846 265267
rect 398512 265193 398518 265205
rect 374530 265165 398518 265193
rect 398512 265153 398518 265165
rect 398570 265153 398576 265205
rect 398818 265193 398846 265239
rect 398992 265227 398998 265279
rect 399050 265267 399056 265279
rect 546352 265267 546358 265279
rect 399050 265239 546358 265267
rect 399050 265227 399056 265239
rect 546352 265227 546358 265239
rect 546410 265227 546416 265279
rect 399856 265193 399862 265205
rect 398818 265165 399862 265193
rect 399856 265153 399862 265165
rect 399914 265153 399920 265205
rect 406480 265153 406486 265205
rect 406538 265193 406544 265205
rect 408112 265193 408118 265205
rect 406538 265165 408118 265193
rect 406538 265153 406544 265165
rect 408112 265153 408118 265165
rect 408170 265153 408176 265205
rect 411760 265153 411766 265205
rect 411818 265193 411824 265205
rect 412048 265193 412054 265205
rect 411818 265165 412054 265193
rect 411818 265153 411824 265165
rect 412048 265153 412054 265165
rect 412106 265153 412112 265205
rect 374434 265091 393182 265119
rect 309424 265005 309430 265057
rect 309482 265045 309488 265057
rect 333616 265045 333622 265057
rect 309482 265017 333622 265045
rect 309482 265005 309488 265017
rect 333616 265005 333622 265017
rect 333674 265005 333680 265057
rect 365968 265005 365974 265057
rect 366026 265045 366032 265057
rect 376720 265045 376726 265057
rect 366026 265017 376726 265045
rect 366026 265005 366032 265017
rect 376720 265005 376726 265017
rect 376778 265005 376784 265057
rect 377200 265005 377206 265057
rect 377258 265045 377264 265057
rect 393154 265045 393182 265091
rect 393328 265079 393334 265131
rect 393386 265119 393392 265131
rect 615376 265119 615382 265131
rect 393386 265091 615382 265119
rect 393386 265079 393392 265091
rect 615376 265079 615382 265091
rect 615434 265079 615440 265131
rect 398992 265045 398998 265057
rect 377258 265017 393086 265045
rect 393154 265017 398998 265045
rect 377258 265005 377264 265017
rect 318736 264971 318742 264983
rect 287594 264943 309278 264971
rect 309346 264943 318742 264971
rect 287594 264931 287600 264943
rect 210640 264857 210646 264909
rect 210698 264897 210704 264909
rect 212464 264897 212470 264909
rect 210698 264869 212470 264897
rect 210698 264857 210704 264869
rect 212464 264857 212470 264869
rect 212522 264857 212528 264909
rect 309250 264897 309278 264943
rect 318736 264931 318742 264943
rect 318794 264931 318800 264983
rect 318928 264931 318934 264983
rect 318986 264971 318992 264983
rect 321040 264971 321046 264983
rect 318986 264943 321046 264971
rect 318986 264931 318992 264943
rect 321040 264931 321046 264943
rect 321098 264931 321104 264983
rect 348592 264971 348598 264983
rect 325186 264943 348598 264971
rect 325186 264897 325214 264943
rect 348592 264931 348598 264943
rect 348650 264931 348656 264983
rect 365200 264931 365206 264983
rect 365258 264971 365264 264983
rect 385648 264971 385654 264983
rect 365258 264943 385654 264971
rect 365258 264931 365264 264943
rect 385648 264931 385654 264943
rect 385706 264931 385712 264983
rect 392848 264971 392854 264983
rect 385762 264943 392854 264971
rect 309250 264869 325214 264897
rect 348496 264857 348502 264909
rect 348554 264897 348560 264909
rect 382384 264897 382390 264909
rect 348554 264869 382390 264897
rect 348554 264857 348560 264869
rect 382384 264857 382390 264869
rect 382442 264857 382448 264909
rect 383440 264857 383446 264909
rect 383498 264897 383504 264909
rect 385762 264897 385790 264943
rect 392848 264931 392854 264943
rect 392906 264931 392912 264983
rect 393058 264971 393086 265017
rect 398992 265005 398998 265017
rect 399050 265005 399056 265057
rect 399088 265005 399094 265057
rect 399146 265045 399152 265057
rect 629680 265045 629686 265057
rect 399146 265017 629686 265045
rect 399146 265005 399152 265017
rect 629680 265005 629686 265017
rect 629738 265005 629744 265057
rect 393328 264971 393334 264983
rect 393058 264943 393334 264971
rect 393328 264931 393334 264943
rect 393386 264931 393392 264983
rect 396976 264931 396982 264983
rect 397034 264971 397040 264983
rect 398608 264971 398614 264983
rect 397034 264943 398614 264971
rect 397034 264931 397040 264943
rect 398608 264931 398614 264943
rect 398666 264931 398672 264983
rect 399568 264931 399574 264983
rect 399626 264971 399632 264983
rect 412624 264971 412630 264983
rect 399626 264943 412630 264971
rect 399626 264931 399632 264943
rect 412624 264931 412630 264943
rect 412682 264931 412688 264983
rect 383498 264869 385790 264897
rect 388983 264909 389035 264915
rect 383498 264857 383504 264869
rect 412720 264897 412726 264909
rect 389035 264869 412726 264897
rect 412720 264857 412726 264869
rect 412778 264857 412784 264909
rect 388983 264851 389035 264857
rect 449392 264709 449398 264761
rect 449450 264749 449456 264761
rect 469360 264749 469366 264761
rect 449450 264721 469366 264749
rect 449450 264709 449456 264721
rect 469360 264709 469366 264721
rect 469418 264709 469424 264761
rect 475792 264709 475798 264761
rect 475850 264749 475856 264761
rect 489520 264749 489526 264761
rect 475850 264721 489526 264749
rect 475850 264709 475856 264721
rect 489520 264709 489526 264721
rect 489578 264709 489584 264761
rect 159856 263451 159862 263503
rect 159914 263491 159920 263503
rect 161104 263491 161110 263503
rect 159914 263463 161110 263491
rect 159914 263451 159920 263463
rect 161104 263451 161110 263463
rect 161162 263451 161168 263503
rect 182224 262119 182230 262171
rect 182282 262159 182288 262171
rect 182282 262131 192926 262159
rect 182282 262119 182288 262131
rect 192898 262085 192926 262131
rect 192976 262085 192982 262097
rect 192898 262057 192982 262085
rect 192976 262045 192982 262057
rect 193034 262045 193040 262097
rect 72016 260639 72022 260691
rect 72074 260679 72080 260691
rect 84688 260679 84694 260691
rect 72074 260651 84694 260679
rect 72074 260639 72080 260651
rect 84688 260639 84694 260651
rect 84746 260639 84752 260691
rect 42448 259677 42454 259729
rect 42506 259717 42512 259729
rect 53872 259717 53878 259729
rect 42506 259689 53878 259717
rect 42506 259677 42512 259689
rect 53872 259677 53878 259689
rect 53930 259677 53936 259729
rect 86416 259233 86422 259285
rect 86474 259273 86480 259285
rect 86474 259245 89342 259273
rect 86474 259233 86480 259245
rect 89314 259199 89342 259245
rect 632464 259233 632470 259285
rect 632522 259273 632528 259285
rect 642160 259273 642166 259285
rect 632522 259245 642166 259273
rect 632522 259233 632528 259245
rect 642160 259233 642166 259245
rect 642218 259233 642224 259285
rect 92272 259199 92278 259211
rect 89314 259171 92278 259199
rect 92272 259159 92278 259171
rect 92330 259159 92336 259211
rect 42832 258937 42838 258989
rect 42890 258977 42896 258989
rect 50320 258977 50326 258989
rect 42890 258949 50326 258977
rect 42890 258937 42896 258949
rect 50320 258937 50326 258949
rect 50378 258937 50384 258989
rect 42448 258641 42454 258693
rect 42506 258681 42512 258693
rect 47440 258681 47446 258693
rect 42506 258653 47446 258681
rect 42506 258641 42512 258653
rect 47440 258641 47446 258653
rect 47498 258641 47504 258693
rect 42448 257827 42454 257879
rect 42506 257867 42512 257879
rect 43216 257867 43222 257879
rect 42506 257839 43222 257867
rect 42506 257827 42512 257839
rect 43216 257827 43222 257839
rect 43274 257827 43280 257879
rect 616336 257753 616342 257805
rect 616394 257793 616400 257805
rect 630736 257793 630742 257805
rect 616394 257765 630742 257793
rect 616394 257753 616400 257765
rect 630736 257753 630742 257765
rect 630794 257753 630800 257805
rect 197104 257605 197110 257657
rect 197162 257645 197168 257657
rect 212080 257645 212086 257657
rect 197162 257617 212086 257645
rect 197162 257605 197168 257617
rect 212080 257605 212086 257617
rect 212138 257605 212144 257657
rect 674608 256421 674614 256473
rect 674666 256461 674672 256473
rect 674896 256461 674902 256473
rect 674666 256433 674902 256461
rect 674666 256421 674672 256433
rect 674896 256421 674902 256433
rect 674954 256421 674960 256473
rect 639280 256347 639286 256399
rect 639338 256387 639344 256399
rect 677104 256387 677110 256399
rect 639338 256359 677110 256387
rect 639338 256347 639344 256359
rect 677104 256347 677110 256359
rect 677162 256347 677168 256399
rect 92272 254867 92278 254919
rect 92330 254907 92336 254919
rect 104368 254907 104374 254919
rect 92330 254879 104374 254907
rect 92330 254867 92336 254879
rect 104368 254867 104374 254879
rect 104426 254867 104432 254919
rect 84688 253461 84694 253513
rect 84746 253501 84752 253513
rect 84746 253473 86462 253501
rect 84746 253461 84752 253473
rect 86434 253427 86462 253473
rect 92176 253427 92182 253439
rect 86434 253399 92182 253427
rect 92176 253387 92182 253399
rect 92234 253387 92240 253439
rect 192976 253387 192982 253439
rect 193034 253427 193040 253439
rect 198736 253427 198742 253439
rect 193034 253399 198742 253427
rect 193034 253387 193040 253399
rect 198736 253387 198742 253399
rect 198794 253387 198800 253439
rect 674608 253387 674614 253439
rect 674666 253427 674672 253439
rect 675280 253427 675286 253439
rect 674666 253399 675286 253427
rect 674666 253387 674672 253399
rect 675280 253387 675286 253399
rect 675338 253387 675344 253439
rect 674512 252721 674518 252773
rect 674570 252761 674576 252773
rect 675088 252761 675094 252773
rect 674570 252733 675094 252761
rect 674570 252721 674576 252733
rect 675088 252721 675094 252733
rect 675146 252721 675152 252773
rect 616336 250615 616342 250627
rect 610594 250587 616342 250615
rect 92176 250501 92182 250553
rect 92234 250541 92240 250553
rect 97168 250541 97174 250553
rect 92234 250513 97174 250541
rect 92234 250501 92240 250513
rect 97168 250501 97174 250513
rect 97226 250501 97232 250553
rect 607696 250501 607702 250553
rect 607754 250541 607760 250553
rect 610594 250541 610622 250587
rect 616336 250575 616342 250587
rect 616394 250575 616400 250627
rect 607754 250513 610622 250541
rect 607754 250501 607760 250513
rect 104368 250057 104374 250109
rect 104426 250097 104432 250109
rect 106576 250097 106582 250109
rect 104426 250069 106582 250097
rect 104426 250057 104432 250069
rect 106576 250057 106582 250069
rect 106634 250057 106640 250109
rect 56176 249243 56182 249295
rect 56234 249283 56240 249295
rect 205648 249283 205654 249295
rect 56234 249255 205654 249283
rect 56234 249243 56240 249255
rect 205648 249243 205654 249255
rect 205706 249243 205712 249295
rect 53776 249169 53782 249221
rect 53834 249209 53840 249221
rect 210736 249209 210742 249221
rect 53834 249181 210742 249209
rect 53834 249169 53840 249181
rect 210736 249169 210742 249181
rect 210794 249169 210800 249221
rect 47632 249095 47638 249147
rect 47690 249135 47696 249147
rect 206896 249135 206902 249147
rect 47690 249107 206902 249135
rect 47690 249095 47696 249107
rect 206896 249095 206902 249107
rect 206954 249095 206960 249147
rect 627856 248059 627862 248111
rect 627914 248099 627920 248111
rect 632464 248099 632470 248111
rect 627914 248071 632470 248099
rect 627914 248059 627920 248071
rect 632464 248059 632470 248071
rect 632522 248059 632528 248111
rect 674416 247911 674422 247963
rect 674474 247951 674480 247963
rect 675472 247951 675478 247963
rect 674474 247923 675478 247951
rect 674474 247911 674480 247923
rect 675472 247911 675478 247923
rect 675530 247911 675536 247963
rect 198736 247689 198742 247741
rect 198794 247729 198800 247741
rect 198794 247701 207326 247729
rect 198794 247689 198800 247701
rect 207298 247655 207326 247701
rect 211024 247689 211030 247741
rect 211082 247729 211088 247741
rect 211312 247729 211318 247741
rect 211082 247701 211318 247729
rect 211082 247689 211088 247701
rect 211312 247689 211318 247701
rect 211370 247689 211376 247741
rect 209392 247655 209398 247667
rect 207298 247627 209398 247655
rect 209392 247615 209398 247627
rect 209450 247615 209456 247667
rect 126544 247319 126550 247371
rect 126602 247359 126608 247371
rect 126602 247331 409406 247359
rect 126602 247319 126608 247331
rect 129520 247245 129526 247297
rect 129578 247285 129584 247297
rect 129578 247257 406334 247285
rect 129578 247245 129584 247257
rect 135184 247171 135190 247223
rect 135242 247211 135248 247223
rect 135242 247183 398894 247211
rect 135242 247171 135248 247183
rect 132304 247097 132310 247149
rect 132362 247137 132368 247149
rect 132362 247109 398750 247137
rect 132362 247097 132368 247109
rect 140944 247023 140950 247075
rect 141002 247063 141008 247075
rect 141002 247035 398078 247063
rect 141002 247023 141008 247035
rect 81136 246989 81142 247001
rect 80674 246961 81142 246989
rect 65200 246727 65206 246779
rect 65258 246767 65264 246779
rect 80674 246767 80702 246961
rect 81136 246949 81142 246961
rect 81194 246949 81200 247001
rect 143920 246949 143926 247001
rect 143978 246989 143984 247001
rect 143978 246961 397694 246989
rect 143978 246949 143984 246961
rect 146704 246875 146710 246927
rect 146762 246915 146768 246927
rect 146762 246887 388094 246915
rect 146762 246875 146768 246887
rect 181456 246801 181462 246853
rect 181514 246841 181520 246853
rect 197584 246841 197590 246853
rect 181514 246813 197590 246841
rect 181514 246801 181520 246813
rect 197584 246801 197590 246813
rect 197642 246801 197648 246853
rect 211792 246801 211798 246853
rect 211850 246841 211856 246853
rect 211850 246813 387038 246841
rect 211850 246801 211856 246813
rect 387010 246779 387038 246813
rect 388066 246779 388094 246887
rect 65258 246739 80702 246767
rect 65258 246727 65264 246739
rect 81136 246727 81142 246779
rect 81194 246767 81200 246779
rect 205072 246767 205078 246779
rect 81194 246739 205078 246767
rect 81194 246727 81200 246739
rect 205072 246727 205078 246739
rect 205130 246727 205136 246779
rect 212272 246727 212278 246779
rect 212330 246767 212336 246779
rect 227056 246767 227062 246779
rect 212330 246739 227062 246767
rect 212330 246727 212336 246739
rect 227056 246727 227062 246739
rect 227114 246727 227120 246779
rect 385072 246767 385078 246779
rect 227218 246739 385078 246767
rect 65008 246653 65014 246705
rect 65066 246693 65072 246705
rect 80656 246693 80662 246705
rect 65066 246665 80662 246693
rect 65066 246653 65072 246665
rect 80656 246653 80662 246665
rect 80714 246653 80720 246705
rect 80944 246653 80950 246705
rect 81002 246693 81008 246705
rect 210928 246693 210934 246705
rect 81002 246665 210934 246693
rect 81002 246653 81008 246665
rect 210928 246653 210934 246665
rect 210986 246653 210992 246705
rect 211888 246653 211894 246705
rect 211946 246693 211952 246705
rect 227218 246693 227246 246739
rect 385072 246727 385078 246739
rect 385130 246727 385136 246779
rect 386992 246727 386998 246779
rect 387050 246727 387056 246779
rect 388048 246727 388054 246779
rect 388106 246727 388112 246779
rect 390256 246727 390262 246779
rect 390314 246767 390320 246779
rect 397666 246767 397694 246961
rect 398050 246767 398078 247035
rect 398722 246989 398750 247109
rect 398866 247063 398894 247183
rect 398866 247035 406238 247063
rect 398722 246961 406142 246989
rect 406114 246779 406142 246961
rect 402160 246767 402166 246779
rect 390314 246739 397598 246767
rect 397666 246739 397790 246767
rect 398050 246739 402166 246767
rect 390314 246727 390320 246739
rect 211946 246665 227246 246693
rect 211946 246653 211952 246665
rect 237808 246653 237814 246705
rect 237866 246693 237872 246705
rect 267472 246693 267478 246705
rect 237866 246665 267478 246693
rect 237866 246653 237872 246665
rect 267472 246653 267478 246665
rect 267530 246653 267536 246705
rect 267568 246653 267574 246705
rect 267626 246693 267632 246705
rect 268624 246693 268630 246705
rect 267626 246665 268630 246693
rect 267626 246653 267632 246665
rect 268624 246653 268630 246665
rect 268682 246653 268688 246705
rect 276688 246693 276694 246705
rect 269218 246665 276694 246693
rect 56080 246579 56086 246631
rect 56138 246619 56144 246631
rect 80752 246619 80758 246631
rect 56138 246591 80758 246619
rect 56138 246579 56144 246591
rect 80752 246579 80758 246591
rect 80810 246579 80816 246631
rect 81232 246579 81238 246631
rect 81290 246619 81296 246631
rect 204880 246619 204886 246631
rect 81290 246591 204886 246619
rect 81290 246579 81296 246591
rect 204880 246579 204886 246591
rect 204938 246579 204944 246631
rect 269218 246619 269246 246665
rect 276688 246653 276694 246665
rect 276746 246653 276752 246705
rect 276802 246665 278750 246693
rect 231778 246591 269246 246619
rect 53200 246505 53206 246557
rect 53258 246545 53264 246557
rect 204688 246545 204694 246557
rect 53258 246517 204694 246545
rect 53258 246505 53264 246517
rect 204688 246505 204694 246517
rect 204746 246505 204752 246557
rect 212176 246505 212182 246557
rect 212234 246545 212240 246557
rect 231778 246545 231806 246591
rect 269296 246579 269302 246631
rect 269354 246619 269360 246631
rect 276802 246619 276830 246665
rect 269354 246591 276830 246619
rect 269354 246579 269360 246591
rect 276880 246579 276886 246631
rect 276938 246619 276944 246631
rect 276938 246591 277118 246619
rect 276938 246579 276944 246591
rect 212234 246517 231806 246545
rect 212234 246505 212240 246517
rect 232144 246505 232150 246557
rect 232202 246545 232208 246557
rect 266608 246545 266614 246557
rect 232202 246517 266614 246545
rect 232202 246505 232208 246517
rect 266608 246505 266614 246517
rect 266666 246505 266672 246557
rect 266704 246505 266710 246557
rect 266762 246545 266768 246557
rect 267568 246545 267574 246557
rect 266762 246517 267574 246545
rect 266762 246505 266768 246517
rect 267568 246505 267574 246517
rect 267626 246505 267632 246557
rect 267952 246505 267958 246557
rect 268010 246545 268016 246557
rect 276592 246545 276598 246557
rect 268010 246517 276598 246545
rect 268010 246505 268016 246517
rect 276592 246505 276598 246517
rect 276650 246505 276656 246557
rect 276688 246505 276694 246557
rect 276746 246545 276752 246557
rect 277090 246545 277118 246591
rect 277360 246579 277366 246631
rect 277418 246619 277424 246631
rect 278608 246619 278614 246631
rect 277418 246591 278614 246619
rect 277418 246579 277424 246591
rect 278608 246579 278614 246591
rect 278666 246579 278672 246631
rect 278722 246619 278750 246665
rect 278800 246653 278806 246705
rect 278858 246693 278864 246705
rect 288016 246693 288022 246705
rect 278858 246665 288022 246693
rect 278858 246653 278864 246665
rect 288016 246653 288022 246665
rect 288074 246653 288080 246705
rect 288130 246665 308414 246693
rect 288130 246619 288158 246665
rect 278722 246591 288158 246619
rect 288880 246579 288886 246631
rect 288938 246619 288944 246631
rect 297904 246619 297910 246631
rect 288938 246591 297910 246619
rect 288938 246579 288944 246591
rect 297904 246579 297910 246591
rect 297962 246579 297968 246631
rect 298000 246579 298006 246631
rect 298058 246619 298064 246631
rect 302416 246619 302422 246631
rect 298058 246591 302422 246619
rect 298058 246579 298064 246591
rect 302416 246579 302422 246591
rect 302474 246579 302480 246631
rect 308080 246619 308086 246631
rect 304258 246591 308086 246619
rect 276746 246517 277022 246545
rect 277090 246517 278654 246545
rect 276746 246505 276752 246517
rect 53392 246431 53398 246483
rect 53450 246471 53456 246483
rect 204784 246471 204790 246483
rect 53450 246443 204790 246471
rect 53450 246431 53456 246443
rect 204784 246431 204790 246443
rect 204842 246431 204848 246483
rect 211696 246431 211702 246483
rect 211754 246471 211760 246483
rect 226960 246471 226966 246483
rect 211754 246443 226966 246471
rect 211754 246431 211760 246443
rect 226960 246431 226966 246443
rect 227018 246431 227024 246483
rect 276880 246471 276886 246483
rect 227458 246443 276886 246471
rect 47728 246357 47734 246409
rect 47786 246397 47792 246409
rect 210160 246397 210166 246409
rect 47786 246369 210166 246397
rect 47786 246357 47792 246369
rect 210160 246357 210166 246369
rect 210218 246357 210224 246409
rect 212080 246357 212086 246409
rect 212138 246397 212144 246409
rect 221776 246397 221782 246409
rect 212138 246369 221782 246397
rect 212138 246357 212144 246369
rect 221776 246357 221782 246369
rect 221834 246357 221840 246409
rect 221872 246357 221878 246409
rect 221930 246397 221936 246409
rect 227458 246397 227486 246443
rect 276880 246431 276886 246443
rect 276938 246431 276944 246483
rect 276994 246471 277022 246517
rect 278626 246471 278654 246517
rect 278704 246505 278710 246557
rect 278762 246545 278768 246557
rect 304258 246545 304286 246591
rect 308080 246579 308086 246591
rect 308138 246579 308144 246631
rect 308386 246619 308414 246665
rect 308464 246653 308470 246705
rect 308522 246693 308528 246705
rect 350128 246693 350134 246705
rect 308522 246665 350134 246693
rect 308522 246653 308528 246665
rect 350128 246653 350134 246665
rect 350186 246653 350192 246705
rect 352336 246653 352342 246705
rect 352394 246693 352400 246705
rect 362608 246693 362614 246705
rect 352394 246665 362614 246693
rect 352394 246653 352400 246665
rect 362608 246653 362614 246665
rect 362666 246653 362672 246705
rect 362722 246665 369086 246693
rect 334864 246619 334870 246631
rect 308386 246591 334870 246619
rect 334864 246579 334870 246591
rect 334922 246579 334928 246631
rect 334960 246579 334966 246631
rect 335018 246619 335024 246631
rect 353200 246619 353206 246631
rect 335018 246591 353206 246619
rect 335018 246579 335024 246591
rect 353200 246579 353206 246591
rect 353258 246579 353264 246631
rect 353296 246579 353302 246631
rect 353354 246619 353360 246631
rect 362722 246619 362750 246665
rect 353354 246591 362750 246619
rect 353354 246579 353360 246591
rect 362800 246579 362806 246631
rect 362858 246619 362864 246631
rect 368944 246619 368950 246631
rect 362858 246591 368950 246619
rect 362858 246579 362864 246591
rect 368944 246579 368950 246591
rect 369002 246579 369008 246631
rect 369058 246619 369086 246665
rect 369136 246653 369142 246705
rect 369194 246693 369200 246705
rect 389488 246693 389494 246705
rect 369194 246665 389494 246693
rect 369194 246653 369200 246665
rect 389488 246653 389494 246665
rect 389546 246653 389552 246705
rect 397570 246693 397598 246739
rect 397648 246693 397654 246705
rect 397570 246665 397654 246693
rect 397648 246653 397654 246665
rect 397706 246653 397712 246705
rect 397762 246693 397790 246739
rect 402160 246727 402166 246739
rect 402218 246727 402224 246779
rect 406096 246727 406102 246779
rect 406154 246727 406160 246779
rect 406210 246767 406238 247035
rect 406306 246841 406334 247257
rect 406306 246836 406564 246841
rect 406306 246830 406576 246836
rect 406306 246813 406524 246830
rect 409378 246779 409406 247331
rect 674320 247023 674326 247075
rect 674378 247063 674384 247075
rect 675472 247063 675478 247075
rect 674378 247035 675478 247063
rect 674378 247023 674384 247035
rect 675472 247023 675478 247035
rect 675530 247023 675536 247075
rect 406524 246772 406576 246778
rect 408976 246767 408982 246779
rect 406210 246739 406490 246767
rect 406462 246734 406490 246739
rect 406614 246739 408982 246767
rect 406614 246734 406642 246739
rect 406462 246706 406642 246734
rect 408976 246727 408982 246739
rect 409034 246727 409040 246779
rect 409360 246727 409366 246779
rect 409418 246727 409424 246779
rect 409456 246727 409462 246779
rect 409514 246767 409520 246779
rect 412144 246767 412150 246779
rect 409514 246739 412150 246767
rect 409514 246727 409520 246739
rect 412144 246727 412150 246739
rect 412202 246727 412208 246779
rect 674704 246727 674710 246779
rect 674762 246767 674768 246779
rect 675376 246767 675382 246779
rect 674762 246739 675382 246767
rect 674762 246727 674768 246739
rect 675376 246727 675382 246739
rect 675434 246727 675440 246779
rect 408784 246693 408790 246705
rect 397762 246678 406424 246693
rect 406672 246678 408790 246693
rect 397762 246665 408790 246678
rect 406396 246650 406700 246665
rect 408784 246653 408790 246665
rect 408842 246653 408848 246705
rect 402064 246619 402070 246631
rect 369058 246591 402070 246619
rect 402064 246579 402070 246591
rect 402122 246579 402128 246631
rect 402160 246579 402166 246631
rect 402218 246619 402224 246631
rect 406768 246619 406774 246631
rect 402218 246591 406774 246619
rect 402218 246579 402224 246591
rect 406768 246579 406774 246591
rect 406826 246579 406832 246631
rect 278762 246517 304286 246545
rect 304354 246517 335102 246545
rect 278762 246505 278768 246517
rect 304354 246471 304382 246517
rect 276994 246443 278078 246471
rect 278626 246443 304382 246471
rect 221930 246369 227486 246397
rect 221930 246357 221936 246369
rect 231856 246357 231862 246409
rect 231914 246397 231920 246409
rect 278050 246397 278078 246443
rect 304432 246431 304438 246483
rect 304490 246471 304496 246483
rect 312400 246471 312406 246483
rect 304490 246443 312406 246471
rect 304490 246431 304496 246443
rect 312400 246431 312406 246443
rect 312458 246431 312464 246483
rect 334960 246471 334966 246483
rect 312514 246443 334966 246471
rect 298000 246397 298006 246409
rect 231914 246369 277982 246397
rect 278050 246369 298006 246397
rect 231914 246357 231920 246369
rect 44848 246283 44854 246335
rect 44906 246323 44912 246335
rect 209680 246323 209686 246335
rect 44906 246295 209686 246323
rect 44906 246283 44912 246295
rect 209680 246283 209686 246295
rect 209738 246283 209744 246335
rect 209968 246283 209974 246335
rect 210026 246323 210032 246335
rect 247216 246323 247222 246335
rect 210026 246295 247222 246323
rect 210026 246283 210032 246295
rect 247216 246283 247222 246295
rect 247274 246283 247280 246335
rect 267760 246283 267766 246335
rect 267818 246323 267824 246335
rect 277954 246323 277982 246369
rect 298000 246357 298006 246369
rect 298058 246357 298064 246409
rect 298096 246357 298102 246409
rect 298154 246397 298160 246409
rect 299248 246397 299254 246409
rect 298154 246369 299254 246397
rect 298154 246357 298160 246369
rect 299248 246357 299254 246369
rect 299306 246357 299312 246409
rect 302416 246357 302422 246409
rect 302474 246397 302480 246409
rect 312514 246397 312542 246443
rect 334960 246431 334966 246443
rect 335018 246431 335024 246483
rect 335074 246471 335102 246517
rect 335344 246505 335350 246557
rect 335402 246545 335408 246557
rect 396784 246545 396790 246557
rect 335402 246517 396790 246545
rect 335402 246505 335408 246517
rect 396784 246505 396790 246517
rect 396842 246505 396848 246557
rect 397648 246505 397654 246557
rect 397706 246545 397712 246557
rect 412048 246545 412054 246557
rect 397706 246517 412054 246545
rect 397706 246505 397712 246517
rect 412048 246505 412054 246517
rect 412106 246505 412112 246557
rect 335074 246443 397310 246471
rect 302474 246369 312542 246397
rect 302474 246357 302480 246369
rect 322000 246357 322006 246409
rect 322058 246397 322064 246409
rect 322058 246369 352766 246397
rect 322058 246357 322064 246369
rect 307984 246323 307990 246335
rect 267818 246295 277886 246323
rect 277954 246295 307990 246323
rect 267818 246283 267824 246295
rect 44944 246209 44950 246261
rect 45002 246249 45008 246261
rect 80752 246249 80758 246261
rect 45002 246221 80758 246249
rect 45002 246209 45008 246221
rect 80752 246209 80758 246221
rect 80810 246209 80816 246261
rect 80944 246209 80950 246261
rect 81002 246249 81008 246261
rect 209584 246249 209590 246261
rect 81002 246221 209590 246249
rect 81002 246209 81008 246221
rect 209584 246209 209590 246221
rect 209642 246209 209648 246261
rect 209872 246209 209878 246261
rect 209930 246249 209936 246261
rect 237808 246249 237814 246261
rect 209930 246221 237814 246249
rect 209930 246209 209936 246221
rect 237808 246209 237814 246221
rect 237866 246209 237872 246261
rect 240496 246209 240502 246261
rect 240554 246249 240560 246261
rect 277360 246249 277366 246261
rect 240554 246221 277366 246249
rect 240554 246209 240560 246221
rect 277360 246209 277366 246221
rect 277418 246209 277424 246261
rect 277858 246249 277886 246295
rect 307984 246283 307990 246295
rect 308042 246283 308048 246335
rect 308080 246283 308086 246335
rect 308138 246323 308144 246335
rect 308138 246295 329630 246323
rect 308138 246283 308144 246295
rect 287632 246249 287638 246261
rect 277858 246221 287638 246249
rect 287632 246209 287638 246221
rect 287690 246209 287696 246261
rect 292240 246249 292246 246261
rect 288034 246221 292246 246249
rect 118096 246135 118102 246187
rect 118154 246175 118160 246187
rect 128080 246175 128086 246187
rect 118154 246147 128086 246175
rect 118154 246135 118160 246147
rect 128080 246135 128086 246147
rect 128138 246135 128144 246187
rect 170896 246175 170902 246187
rect 161218 246147 170902 246175
rect 46192 246061 46198 246113
rect 46250 246101 46256 246113
rect 60496 246101 60502 246113
rect 46250 246073 60502 246101
rect 46250 246061 46256 246073
rect 60496 246061 60502 246073
rect 60554 246061 60560 246113
rect 66256 246061 66262 246113
rect 66314 246101 66320 246113
rect 77776 246101 77782 246113
rect 66314 246073 77782 246101
rect 66314 246061 66320 246073
rect 77776 246061 77782 246073
rect 77834 246061 77840 246113
rect 97840 245987 97846 246039
rect 97898 246027 97904 246039
rect 118096 246027 118102 246039
rect 97898 245999 118102 246027
rect 97898 245987 97904 245999
rect 118096 245987 118102 245999
rect 118154 245987 118160 246039
rect 128080 245987 128086 246039
rect 128138 246027 128144 246039
rect 141136 246027 141142 246039
rect 128138 245999 141142 246027
rect 128138 245987 128144 245999
rect 141136 245987 141142 245999
rect 141194 245987 141200 246039
rect 151120 245987 151126 246039
rect 151178 246027 151184 246039
rect 161218 246027 161246 246147
rect 170896 246135 170902 246147
rect 170954 246135 170960 246187
rect 211984 246135 211990 246187
rect 212042 246175 212048 246187
rect 267760 246175 267766 246187
rect 212042 246147 267766 246175
rect 212042 246135 212048 246147
rect 267760 246135 267766 246147
rect 267818 246135 267824 246187
rect 267856 246135 267862 246187
rect 267914 246175 267920 246187
rect 269296 246175 269302 246187
rect 267914 246147 269302 246175
rect 267914 246135 267920 246147
rect 269296 246135 269302 246147
rect 269354 246135 269360 246187
rect 272848 246135 272854 246187
rect 272906 246175 272912 246187
rect 278032 246175 278038 246187
rect 272906 246147 278038 246175
rect 272906 246135 272912 246147
rect 278032 246135 278038 246147
rect 278090 246135 278096 246187
rect 278128 246135 278134 246187
rect 278186 246175 278192 246187
rect 288034 246175 288062 246221
rect 292240 246209 292246 246221
rect 292298 246209 292304 246261
rect 292336 246209 292342 246261
rect 292394 246249 292400 246261
rect 294160 246249 294166 246261
rect 292394 246221 294166 246249
rect 292394 246209 292400 246221
rect 294160 246209 294166 246221
rect 294218 246209 294224 246261
rect 294544 246209 294550 246261
rect 294602 246249 294608 246261
rect 301264 246249 301270 246261
rect 294602 246221 301270 246249
rect 294602 246209 294608 246221
rect 301264 246209 301270 246221
rect 301322 246209 301328 246261
rect 301360 246209 301366 246261
rect 301418 246249 301424 246261
rect 329602 246249 329630 246295
rect 329680 246283 329686 246335
rect 329738 246323 329744 246335
rect 329738 246295 335102 246323
rect 329738 246283 329744 246295
rect 334768 246249 334774 246261
rect 301418 246221 322238 246249
rect 329602 246221 334774 246249
rect 301418 246209 301424 246221
rect 278186 246147 288062 246175
rect 278186 246135 278192 246147
rect 288112 246135 288118 246187
rect 288170 246175 288176 246187
rect 308464 246175 308470 246187
rect 288170 246147 308470 246175
rect 288170 246135 288176 246147
rect 308464 246135 308470 246147
rect 308522 246135 308528 246187
rect 308560 246135 308566 246187
rect 308618 246175 308624 246187
rect 322000 246175 322006 246187
rect 308618 246147 322006 246175
rect 308618 246135 308624 246147
rect 322000 246135 322006 246147
rect 322058 246135 322064 246187
rect 322210 246175 322238 246221
rect 334768 246209 334774 246221
rect 334826 246209 334832 246261
rect 335074 246249 335102 246295
rect 335152 246283 335158 246335
rect 335210 246323 335216 246335
rect 352336 246323 352342 246335
rect 335210 246295 352342 246323
rect 335210 246283 335216 246295
rect 352336 246283 352342 246295
rect 352394 246283 352400 246335
rect 352738 246323 352766 246369
rect 353200 246357 353206 246409
rect 353258 246397 353264 246409
rect 378640 246397 378646 246409
rect 353258 246369 378646 246397
rect 353258 246357 353264 246369
rect 378640 246357 378646 246369
rect 378698 246357 378704 246409
rect 388528 246357 388534 246409
rect 388586 246397 388592 246409
rect 389776 246397 389782 246409
rect 388586 246369 389782 246397
rect 388586 246357 388592 246369
rect 389776 246357 389782 246369
rect 389834 246357 389840 246409
rect 397282 246397 397310 246443
rect 397360 246431 397366 246483
rect 397418 246471 397424 246483
rect 407248 246471 407254 246483
rect 397418 246443 407254 246471
rect 397418 246431 397424 246443
rect 407248 246431 407254 246443
rect 407306 246431 407312 246483
rect 408592 246397 408598 246409
rect 397282 246369 408598 246397
rect 408592 246357 408598 246369
rect 408650 246357 408656 246409
rect 387280 246323 387286 246335
rect 352738 246295 387286 246323
rect 387280 246283 387286 246295
rect 387338 246283 387344 246335
rect 388912 246283 388918 246335
rect 388970 246323 388976 246335
rect 407632 246323 407638 246335
rect 388970 246295 407638 246323
rect 388970 246283 388976 246295
rect 407632 246283 407638 246295
rect 407690 246283 407696 246335
rect 335074 246221 372734 246249
rect 329680 246175 329686 246187
rect 322210 246147 329686 246175
rect 329680 246135 329686 246147
rect 329738 246135 329744 246187
rect 330736 246135 330742 246187
rect 330794 246175 330800 246187
rect 358000 246175 358006 246187
rect 330794 246147 358006 246175
rect 330794 246135 330800 246147
rect 358000 246135 358006 246147
rect 358058 246135 358064 246187
rect 181552 246061 181558 246113
rect 181610 246101 181616 246113
rect 205840 246101 205846 246113
rect 181610 246073 205846 246101
rect 181610 246061 181616 246073
rect 205840 246061 205846 246073
rect 205898 246061 205904 246113
rect 216016 246101 216022 246113
rect 215938 246073 216022 246101
rect 151178 245999 161246 246027
rect 151178 245987 151184 245999
rect 170896 245987 170902 246039
rect 170954 246027 170960 246039
rect 181456 246027 181462 246039
rect 170954 245999 181462 246027
rect 170954 245987 170960 245999
rect 181456 245987 181462 245999
rect 181514 245987 181520 246039
rect 205840 245913 205846 245965
rect 205898 245953 205904 245965
rect 215938 245953 215966 246073
rect 216016 246061 216022 246073
rect 216074 246061 216080 246113
rect 237712 246061 237718 246113
rect 237770 246101 237776 246113
rect 242512 246101 242518 246113
rect 237770 246073 242518 246101
rect 237770 246061 237776 246073
rect 242512 246061 242518 246073
rect 242570 246061 242576 246113
rect 266512 246101 266518 246113
rect 243298 246073 266518 246101
rect 227056 245987 227062 246039
rect 227114 246027 227120 246039
rect 231856 246027 231862 246039
rect 227114 245999 231862 246027
rect 227114 245987 227120 245999
rect 231856 245987 231862 245999
rect 231914 245987 231920 246039
rect 240016 245987 240022 246039
rect 240074 246027 240080 246039
rect 241744 246027 241750 246039
rect 240074 245999 241750 246027
rect 240074 245987 240080 245999
rect 241744 245987 241750 245999
rect 241802 245987 241808 246039
rect 205898 245925 215966 245953
rect 205898 245913 205904 245925
rect 236080 245913 236086 245965
rect 236138 245953 236144 245965
rect 243298 245953 243326 246073
rect 266512 246061 266518 246073
rect 266570 246061 266576 246113
rect 266608 246061 266614 246113
rect 266666 246101 266672 246113
rect 278608 246101 278614 246113
rect 266666 246073 278614 246101
rect 266666 246061 266672 246073
rect 278608 246061 278614 246073
rect 278666 246061 278672 246113
rect 278704 246061 278710 246113
rect 278762 246101 278768 246113
rect 285904 246101 285910 246113
rect 278762 246073 285910 246101
rect 278762 246061 278768 246073
rect 285904 246061 285910 246073
rect 285962 246061 285968 246113
rect 286096 246061 286102 246113
rect 286154 246101 286160 246113
rect 292624 246101 292630 246113
rect 286154 246073 292630 246101
rect 286154 246061 286160 246073
rect 292624 246061 292630 246073
rect 292682 246061 292688 246113
rect 292720 246061 292726 246113
rect 292778 246101 292784 246113
rect 304432 246101 304438 246113
rect 292778 246073 304438 246101
rect 292778 246061 292784 246073
rect 304432 246061 304438 246073
rect 304490 246061 304496 246113
rect 304528 246061 304534 246113
rect 304586 246101 304592 246113
rect 308944 246101 308950 246113
rect 304586 246073 308950 246101
rect 304586 246061 304592 246073
rect 308944 246061 308950 246073
rect 309002 246061 309008 246113
rect 312400 246061 312406 246113
rect 312458 246101 312464 246113
rect 342736 246101 342742 246113
rect 312458 246073 342742 246101
rect 312458 246061 312464 246073
rect 342736 246061 342742 246073
rect 342794 246061 342800 246113
rect 350128 246061 350134 246113
rect 350186 246101 350192 246113
rect 353296 246101 353302 246113
rect 350186 246073 353302 246101
rect 350186 246061 350192 246073
rect 353296 246061 353302 246073
rect 353354 246061 353360 246113
rect 372706 246101 372734 246221
rect 378640 246209 378646 246261
rect 378698 246249 378704 246261
rect 412240 246249 412246 246261
rect 378698 246221 412246 246249
rect 378698 246209 378704 246221
rect 412240 246209 412246 246221
rect 412298 246209 412304 246261
rect 389296 246175 389302 246187
rect 373186 246147 389302 246175
rect 373186 246101 373214 246147
rect 389296 246135 389302 246147
rect 389354 246135 389360 246187
rect 396784 246135 396790 246187
rect 396842 246175 396848 246187
rect 406192 246175 406198 246187
rect 396842 246147 406198 246175
rect 396842 246135 396848 246147
rect 406192 246135 406198 246147
rect 406250 246135 406256 246187
rect 372706 246073 373214 246101
rect 387376 246061 387382 246113
rect 387434 246101 387440 246113
rect 388912 246101 388918 246113
rect 387434 246073 388918 246101
rect 387434 246061 387440 246073
rect 388912 246061 388918 246073
rect 388970 246061 388976 246113
rect 505360 246101 505366 246113
rect 389026 246073 505366 246101
rect 247216 245987 247222 246039
rect 247274 246027 247280 246039
rect 252496 246027 252502 246039
rect 247274 245999 252502 246027
rect 247274 245987 247280 245999
rect 252496 245987 252502 245999
rect 252554 245987 252560 246039
rect 262576 245987 262582 246039
rect 262634 246027 262640 246039
rect 277744 246027 277750 246039
rect 262634 245999 277750 246027
rect 262634 245987 262640 245999
rect 277744 245987 277750 245999
rect 277802 245987 277808 246039
rect 367504 246027 367510 246039
rect 277858 245999 367510 246027
rect 236138 245925 243326 245953
rect 236138 245913 236144 245925
rect 263824 245913 263830 245965
rect 263882 245953 263888 245965
rect 277858 245953 277886 245999
rect 367504 245987 367510 245999
rect 367562 245987 367568 246039
rect 367696 245987 367702 246039
rect 367754 246027 367760 246039
rect 389026 246027 389054 246073
rect 505360 246061 505366 246073
rect 505418 246061 505424 246113
rect 674800 246061 674806 246113
rect 674858 246101 674864 246113
rect 675376 246101 675382 246113
rect 674858 246073 675382 246101
rect 674858 246061 674864 246073
rect 675376 246061 675382 246073
rect 675434 246061 675440 246113
rect 367754 245999 389054 246027
rect 367754 245987 367760 245999
rect 389296 245987 389302 246039
rect 389354 246027 389360 246039
rect 409840 246027 409846 246039
rect 389354 245999 409846 246027
rect 389354 245987 389360 245999
rect 409840 245987 409846 245999
rect 409898 245987 409904 246039
rect 263882 245925 277886 245953
rect 263882 245913 263888 245925
rect 278032 245913 278038 245965
rect 278090 245953 278096 245965
rect 368080 245953 368086 245965
rect 278090 245925 368086 245953
rect 278090 245913 278096 245925
rect 368080 245913 368086 245925
rect 368138 245913 368144 245965
rect 385072 245913 385078 245965
rect 385130 245953 385136 245965
rect 409168 245953 409174 245965
rect 385130 245925 409174 245953
rect 385130 245913 385136 245925
rect 409168 245913 409174 245925
rect 409226 245913 409232 245965
rect 77776 245839 77782 245891
rect 77834 245879 77840 245891
rect 97840 245879 97846 245891
rect 77834 245851 97846 245879
rect 77834 245839 77840 245851
rect 97840 245839 97846 245851
rect 97898 245839 97904 245891
rect 141136 245839 141142 245891
rect 141194 245879 141200 245891
rect 151120 245879 151126 245891
rect 141194 245851 151126 245879
rect 141194 245839 141200 245851
rect 151120 245839 151126 245851
rect 151178 245839 151184 245891
rect 237040 245839 237046 245891
rect 237098 245879 237104 245891
rect 252688 245879 252694 245891
rect 237098 245851 252694 245879
rect 237098 245839 237104 245851
rect 252688 245839 252694 245851
rect 252746 245839 252752 245891
rect 255088 245839 255094 245891
rect 255146 245879 255152 245891
rect 338128 245879 338134 245891
rect 255146 245851 338134 245879
rect 255146 245839 255152 245851
rect 338128 245839 338134 245851
rect 338186 245839 338192 245891
rect 338224 245839 338230 245891
rect 338282 245879 338288 245891
rect 357424 245879 357430 245891
rect 338282 245851 357430 245879
rect 338282 245839 338288 245851
rect 357424 245839 357430 245851
rect 357482 245839 357488 245891
rect 387280 245839 387286 245891
rect 387338 245879 387344 245891
rect 409456 245879 409462 245891
rect 387338 245851 409462 245879
rect 387338 245839 387344 245851
rect 409456 245839 409462 245851
rect 409514 245839 409520 245891
rect 210832 245765 210838 245817
rect 210890 245805 210896 245817
rect 227344 245805 227350 245817
rect 210890 245777 227350 245805
rect 210890 245765 210896 245777
rect 227344 245765 227350 245777
rect 227402 245765 227408 245817
rect 251344 245765 251350 245817
rect 251402 245805 251408 245817
rect 356272 245805 356278 245817
rect 251402 245777 356278 245805
rect 251402 245765 251408 245777
rect 356272 245765 356278 245777
rect 356330 245765 356336 245817
rect 388048 245765 388054 245817
rect 388106 245805 388112 245817
rect 397360 245805 397366 245817
rect 388106 245777 397366 245805
rect 388106 245765 388112 245777
rect 397360 245765 397366 245777
rect 397418 245765 397424 245817
rect 226960 245691 226966 245743
rect 227018 245731 227024 245743
rect 232144 245731 232150 245743
rect 227018 245703 232150 245731
rect 227018 245691 227024 245703
rect 232144 245691 232150 245703
rect 232202 245691 232208 245743
rect 254128 245691 254134 245743
rect 254186 245731 254192 245743
rect 330736 245731 330742 245743
rect 254186 245703 330742 245731
rect 254186 245691 254192 245703
rect 330736 245691 330742 245703
rect 330794 245691 330800 245743
rect 330832 245691 330838 245743
rect 330890 245731 330896 245743
rect 357136 245731 357142 245743
rect 330890 245703 357142 245731
rect 330890 245691 330896 245703
rect 357136 245691 357142 245703
rect 357194 245691 357200 245743
rect 386992 245691 386998 245743
rect 387050 245731 387056 245743
rect 390256 245731 390262 245743
rect 387050 245703 390262 245731
rect 387050 245691 387056 245703
rect 390256 245691 390262 245703
rect 390314 245691 390320 245743
rect 402064 245691 402070 245743
rect 402122 245731 402128 245743
rect 407056 245731 407062 245743
rect 402122 245703 407062 245731
rect 402122 245691 402128 245703
rect 407056 245691 407062 245703
rect 407114 245691 407120 245743
rect 216016 245617 216022 245669
rect 216074 245657 216080 245669
rect 236080 245657 236086 245669
rect 216074 245629 236086 245657
rect 216074 245617 216080 245629
rect 236080 245617 236086 245629
rect 236138 245617 236144 245669
rect 263056 245617 263062 245669
rect 263114 245657 263120 245669
rect 263114 245629 277886 245657
rect 263114 245617 263120 245629
rect 210544 245543 210550 245595
rect 210602 245583 210608 245595
rect 277744 245583 277750 245595
rect 210602 245555 277750 245583
rect 210602 245543 210608 245555
rect 277744 245543 277750 245555
rect 277802 245543 277808 245595
rect 277858 245583 277886 245629
rect 277936 245617 277942 245669
rect 277994 245657 278000 245669
rect 370960 245657 370966 245669
rect 277994 245629 370966 245657
rect 277994 245617 278000 245629
rect 370960 245617 370966 245629
rect 371018 245617 371024 245669
rect 369232 245583 369238 245595
rect 277858 245555 369238 245583
rect 369232 245543 369238 245555
rect 369290 245543 369296 245595
rect 250288 245469 250294 245521
rect 250346 245509 250352 245521
rect 338512 245509 338518 245521
rect 250346 245481 338518 245509
rect 250346 245469 250352 245481
rect 338512 245469 338518 245481
rect 338570 245469 338576 245521
rect 253360 245395 253366 245447
rect 253418 245435 253424 245447
rect 338224 245435 338230 245447
rect 253418 245407 338230 245435
rect 253418 245395 253424 245407
rect 338224 245395 338230 245407
rect 338282 245395 338288 245447
rect 355792 245435 355798 245447
rect 338338 245407 355798 245435
rect 249616 245321 249622 245373
rect 249674 245361 249680 245373
rect 338338 245361 338366 245407
rect 355792 245395 355798 245407
rect 355850 245395 355856 245447
rect 358576 245435 358582 245447
rect 358210 245407 358582 245435
rect 249674 245333 338366 245361
rect 249674 245321 249680 245333
rect 338416 245321 338422 245373
rect 338474 245361 338480 245373
rect 358096 245361 358102 245373
rect 338474 245333 358102 245361
rect 338474 245321 338480 245333
rect 358096 245321 358102 245333
rect 358154 245321 358160 245373
rect 252400 245247 252406 245299
rect 252458 245287 252464 245299
rect 330832 245287 330838 245299
rect 252458 245259 330838 245287
rect 252458 245247 252464 245259
rect 330832 245247 330838 245259
rect 330890 245247 330896 245299
rect 330928 245247 330934 245299
rect 330986 245287 330992 245299
rect 358210 245287 358238 245407
rect 358576 245395 358582 245407
rect 358634 245395 358640 245447
rect 405904 245395 405910 245447
rect 405962 245435 405968 245447
rect 412432 245435 412438 245447
rect 405962 245407 412438 245435
rect 405962 245395 405968 245407
rect 412432 245395 412438 245407
rect 412490 245395 412496 245447
rect 358480 245321 358486 245373
rect 358538 245361 358544 245373
rect 362896 245361 362902 245373
rect 358538 245333 362902 245361
rect 358538 245321 358544 245333
rect 362896 245321 362902 245333
rect 362954 245321 362960 245373
rect 364258 245333 383678 245361
rect 364258 245287 364286 245333
rect 330986 245259 358238 245287
rect 358498 245259 364286 245287
rect 368674 245259 372158 245287
rect 330986 245247 330992 245259
rect 210160 245173 210166 245225
rect 210218 245213 210224 245225
rect 214000 245213 214006 245225
rect 210218 245185 214006 245213
rect 210218 245173 210224 245185
rect 214000 245173 214006 245185
rect 214058 245173 214064 245225
rect 216592 245173 216598 245225
rect 216650 245213 216656 245225
rect 358498 245213 358526 245259
rect 216650 245185 358526 245213
rect 216650 245173 216656 245185
rect 358576 245173 358582 245225
rect 358634 245213 358640 245225
rect 368674 245213 368702 245259
rect 372016 245213 372022 245225
rect 358634 245185 368702 245213
rect 368770 245185 372022 245213
rect 358634 245173 358640 245185
rect 209584 245099 209590 245151
rect 209642 245139 209648 245151
rect 213520 245139 213526 245151
rect 209642 245111 213526 245139
rect 209642 245099 209648 245111
rect 213520 245099 213526 245111
rect 213578 245099 213584 245151
rect 226384 245099 226390 245151
rect 226442 245139 226448 245151
rect 251920 245139 251926 245151
rect 226442 245111 251926 245139
rect 226442 245099 226448 245111
rect 251920 245099 251926 245111
rect 251978 245099 251984 245151
rect 261808 245099 261814 245151
rect 261866 245139 261872 245151
rect 368770 245139 368798 245185
rect 372016 245173 372022 245185
rect 372074 245173 372080 245225
rect 261866 245111 368798 245139
rect 372130 245139 372158 245259
rect 383650 245213 383678 245333
rect 411472 245213 411478 245225
rect 383650 245185 411478 245213
rect 411472 245173 411478 245185
rect 411530 245173 411536 245225
rect 405712 245139 405718 245151
rect 372130 245111 405718 245139
rect 261866 245099 261872 245111
rect 405712 245099 405718 245111
rect 405770 245099 405776 245151
rect 42448 245025 42454 245077
rect 42506 245065 42512 245077
rect 214288 245065 214294 245077
rect 42506 245037 214294 245065
rect 42506 245025 42512 245037
rect 214288 245025 214294 245037
rect 214346 245025 214352 245077
rect 260848 245025 260854 245077
rect 260906 245065 260912 245077
rect 374032 245065 374038 245077
rect 260906 245037 374038 245065
rect 260906 245025 260912 245037
rect 374032 245025 374038 245037
rect 374090 245025 374096 245077
rect 210064 244951 210070 245003
rect 210122 244991 210128 245003
rect 252112 244991 252118 245003
rect 210122 244963 252118 244991
rect 210122 244951 210128 244963
rect 252112 244951 252118 244963
rect 252170 244951 252176 245003
rect 260752 244951 260758 245003
rect 260810 244991 260816 245003
rect 374608 244991 374614 245003
rect 260810 244963 374614 244991
rect 260810 244951 260816 244963
rect 374608 244951 374614 244963
rect 374666 244951 374672 245003
rect 209680 244877 209686 244929
rect 209738 244917 209744 244929
rect 213136 244917 213142 244929
rect 209738 244889 213142 244917
rect 209738 244877 209744 244889
rect 213136 244877 213142 244889
rect 213194 244877 213200 244929
rect 216496 244877 216502 244929
rect 216554 244917 216560 244929
rect 216554 244889 331070 244917
rect 216554 244877 216560 244889
rect 106576 244803 106582 244855
rect 106634 244843 106640 244855
rect 106634 244815 109502 244843
rect 106634 244803 106640 244815
rect 109474 244769 109502 244815
rect 210064 244803 210070 244855
rect 210122 244843 210128 244855
rect 210122 244815 251870 244843
rect 210122 244803 210128 244815
rect 149584 244769 149590 244781
rect 109474 244741 149590 244769
rect 149584 244729 149590 244741
rect 149642 244729 149648 244781
rect 97168 244655 97174 244707
rect 97226 244695 97232 244707
rect 142480 244695 142486 244707
rect 97226 244667 142486 244695
rect 97226 244655 97232 244667
rect 142480 244655 142486 244667
rect 142538 244655 142544 244707
rect 251842 244695 251870 244815
rect 251920 244803 251926 244855
rect 251978 244843 251984 244855
rect 319792 244843 319798 244855
rect 251978 244815 319798 244843
rect 251978 244803 251984 244815
rect 319792 244803 319798 244815
rect 319850 244803 319856 244855
rect 319984 244803 319990 244855
rect 320042 244843 320048 244855
rect 330928 244843 330934 244855
rect 320042 244815 330934 244843
rect 320042 244803 320048 244815
rect 330928 244803 330934 244815
rect 330986 244803 330992 244855
rect 331042 244843 331070 244889
rect 338512 244877 338518 244929
rect 338570 244917 338576 244929
rect 355888 244917 355894 244929
rect 338570 244889 355894 244917
rect 338570 244877 338576 244889
rect 355888 244877 355894 244889
rect 355946 244877 355952 244929
rect 389296 244917 389302 244929
rect 367234 244889 389302 244917
rect 353584 244843 353590 244855
rect 331042 244815 353590 244843
rect 353584 244803 353590 244815
rect 353642 244803 353648 244855
rect 252112 244729 252118 244781
rect 252170 244769 252176 244781
rect 285712 244769 285718 244781
rect 252170 244741 285718 244769
rect 252170 244729 252176 244741
rect 285712 244729 285718 244741
rect 285770 244729 285776 244781
rect 285904 244729 285910 244781
rect 285962 244769 285968 244781
rect 292720 244769 292726 244781
rect 285962 244741 292726 244769
rect 285962 244729 285968 244741
rect 292720 244729 292726 244741
rect 292778 244729 292784 244781
rect 292816 244729 292822 244781
rect 292874 244769 292880 244781
rect 367234 244769 367262 244889
rect 389296 244877 389302 244889
rect 389354 244877 389360 244929
rect 408112 244843 408118 244855
rect 292874 244741 367262 244769
rect 379282 244815 408118 244843
rect 292874 244729 292880 244741
rect 268240 244695 268246 244707
rect 251842 244667 268246 244695
rect 268240 244655 268246 244667
rect 268298 244655 268304 244707
rect 277936 244695 277942 244707
rect 268354 244667 277942 244695
rect 138160 244581 138166 244633
rect 138218 244621 138224 244633
rect 206800 244621 206806 244633
rect 138218 244593 206806 244621
rect 138218 244581 138224 244593
rect 206800 244581 206806 244593
rect 206858 244581 206864 244633
rect 266512 244581 266518 244633
rect 266570 244621 266576 244633
rect 268354 244621 268382 244667
rect 277936 244655 277942 244667
rect 277994 244655 278000 244707
rect 278032 244655 278038 244707
rect 278090 244695 278096 244707
rect 278090 244667 288158 244695
rect 278090 244655 278096 244667
rect 266570 244593 268382 244621
rect 266570 244581 266576 244593
rect 277744 244581 277750 244633
rect 277802 244621 277808 244633
rect 277802 244593 282398 244621
rect 277802 244581 277808 244593
rect 135280 244507 135286 244559
rect 135338 244547 135344 244559
rect 204976 244547 204982 244559
rect 135338 244519 204982 244547
rect 135338 244507 135344 244519
rect 204976 244507 204982 244519
rect 205034 244507 205040 244559
rect 277360 244507 277366 244559
rect 277418 244547 277424 244559
rect 282256 244547 282262 244559
rect 277418 244519 282262 244547
rect 277418 244507 277424 244519
rect 282256 244507 282262 244519
rect 282314 244507 282320 244559
rect 282370 244547 282398 244593
rect 282448 244581 282454 244633
rect 282506 244621 282512 244633
rect 288016 244621 288022 244633
rect 282506 244593 288022 244621
rect 282506 244581 282512 244593
rect 288016 244581 288022 244593
rect 288074 244581 288080 244633
rect 288130 244621 288158 244667
rect 288208 244655 288214 244707
rect 288266 244695 288272 244707
rect 379282 244695 379310 244815
rect 408112 244803 408118 244815
rect 408170 244803 408176 244855
rect 607696 244843 607702 244855
rect 604834 244815 607702 244843
rect 603088 244729 603094 244781
rect 603146 244769 603152 244781
rect 604834 244769 604862 244815
rect 607696 244803 607702 244815
rect 607754 244803 607760 244855
rect 603146 244741 604862 244769
rect 603146 244729 603152 244741
rect 288266 244667 379310 244695
rect 288266 244655 288272 244667
rect 306640 244621 306646 244633
rect 288130 244593 306646 244621
rect 306640 244581 306646 244593
rect 306698 244581 306704 244633
rect 306736 244581 306742 244633
rect 306794 244621 306800 244633
rect 319696 244621 319702 244633
rect 306794 244593 319702 244621
rect 306794 244581 306800 244593
rect 319696 244581 319702 244593
rect 319754 244581 319760 244633
rect 342736 244581 342742 244633
rect 342794 244621 342800 244633
rect 367696 244621 367702 244633
rect 342794 244593 367702 244621
rect 342794 244581 342800 244593
rect 367696 244581 367702 244593
rect 367754 244581 367760 244633
rect 291856 244547 291862 244559
rect 282370 244519 291862 244547
rect 291856 244507 291862 244519
rect 291914 244507 291920 244559
rect 291952 244507 291958 244559
rect 292010 244547 292016 244559
rect 301360 244547 301366 244559
rect 292010 244519 301366 244547
rect 292010 244507 292016 244519
rect 301360 244507 301366 244519
rect 301418 244507 301424 244559
rect 302320 244507 302326 244559
rect 302378 244547 302384 244559
rect 304528 244547 304534 244559
rect 302378 244519 304534 244547
rect 302378 244507 302384 244519
rect 304528 244507 304534 244519
rect 304586 244507 304592 244559
rect 310768 244547 310774 244559
rect 304642 244519 310774 244547
rect 132400 244433 132406 244485
rect 132458 244473 132464 244485
rect 205552 244473 205558 244485
rect 132458 244445 205558 244473
rect 132458 244433 132464 244445
rect 205552 244433 205558 244445
rect 205610 244433 205616 244485
rect 263440 244433 263446 244485
rect 263498 244473 263504 244485
rect 272848 244473 272854 244485
rect 263498 244445 272854 244473
rect 263498 244433 263504 244445
rect 272848 244433 272854 244445
rect 272906 244433 272912 244485
rect 304642 244473 304670 244519
rect 310768 244507 310774 244519
rect 310826 244507 310832 244559
rect 312016 244507 312022 244559
rect 312074 244547 312080 244559
rect 367600 244547 367606 244559
rect 312074 244519 367606 244547
rect 312074 244507 312080 244519
rect 367600 244507 367606 244519
rect 367658 244507 367664 244559
rect 277570 244445 304670 244473
rect 126640 244359 126646 244411
rect 126698 244399 126704 244411
rect 205360 244399 205366 244411
rect 126698 244371 205366 244399
rect 126698 244359 126704 244371
rect 205360 244359 205366 244371
rect 205418 244359 205424 244411
rect 264784 244359 264790 244411
rect 264842 244399 264848 244411
rect 277570 244399 277598 244445
rect 307888 244433 307894 244485
rect 307946 244473 307952 244485
rect 308272 244473 308278 244485
rect 307946 244445 308278 244473
rect 307946 244433 307952 244445
rect 308272 244433 308278 244445
rect 308330 244433 308336 244485
rect 312208 244433 312214 244485
rect 312266 244473 312272 244485
rect 319792 244473 319798 244485
rect 312266 244445 319798 244473
rect 312266 244433 312272 244445
rect 319792 244433 319798 244445
rect 319850 244433 319856 244485
rect 319888 244433 319894 244485
rect 319946 244473 319952 244485
rect 321328 244473 321334 244485
rect 319946 244445 321334 244473
rect 319946 244433 319952 244445
rect 321328 244433 321334 244445
rect 321386 244433 321392 244485
rect 368752 244473 368758 244485
rect 339970 244445 368758 244473
rect 264842 244371 277598 244399
rect 264842 244359 264848 244371
rect 277840 244359 277846 244411
rect 277898 244399 277904 244411
rect 310480 244399 310486 244411
rect 277898 244371 310486 244399
rect 277898 244359 277904 244371
rect 310480 244359 310486 244371
rect 310538 244359 310544 244411
rect 339856 244359 339862 244411
rect 339914 244399 339920 244411
rect 339970 244399 339998 244445
rect 368752 244433 368758 244445
rect 368810 244433 368816 244485
rect 339914 244371 339998 244399
rect 339914 244359 339920 244371
rect 123760 244285 123766 244337
rect 123818 244325 123824 244337
rect 205168 244325 205174 244337
rect 123818 244297 205174 244325
rect 123818 244285 123824 244297
rect 205168 244285 205174 244297
rect 205226 244285 205232 244337
rect 256528 244285 256534 244337
rect 256586 244325 256592 244337
rect 276304 244325 276310 244337
rect 256586 244297 276310 244325
rect 256586 244285 256592 244297
rect 276304 244285 276310 244297
rect 276362 244285 276368 244337
rect 277936 244285 277942 244337
rect 277994 244325 278000 244337
rect 306736 244325 306742 244337
rect 277994 244297 306742 244325
rect 277994 244285 278000 244297
rect 306736 244285 306742 244297
rect 306794 244285 306800 244337
rect 312400 244285 312406 244337
rect 312458 244325 312464 244337
rect 339760 244325 339766 244337
rect 312458 244297 339766 244325
rect 312458 244285 312464 244297
rect 339760 244285 339766 244297
rect 339818 244285 339824 244337
rect 120880 244211 120886 244263
rect 120938 244251 120944 244263
rect 205648 244251 205654 244263
rect 120938 244223 205654 244251
rect 120938 244211 120944 244223
rect 205648 244211 205654 244223
rect 205706 244211 205712 244263
rect 235120 244211 235126 244263
rect 235178 244251 235184 244263
rect 267184 244251 267190 244263
rect 235178 244223 267190 244251
rect 235178 244211 235184 244223
rect 267184 244211 267190 244223
rect 267242 244211 267248 244263
rect 275920 244211 275926 244263
rect 275978 244251 275984 244263
rect 276400 244251 276406 244263
rect 275978 244223 276406 244251
rect 275978 244211 275984 244223
rect 276400 244211 276406 244223
rect 276458 244211 276464 244263
rect 276592 244211 276598 244263
rect 276650 244251 276656 244263
rect 318256 244251 318262 244263
rect 276650 244223 318262 244251
rect 276650 244211 276656 244223
rect 318256 244211 318262 244223
rect 318314 244211 318320 244263
rect 118000 244137 118006 244189
rect 118058 244177 118064 244189
rect 204496 244177 204502 244189
rect 118058 244149 204502 244177
rect 118058 244137 118064 244149
rect 204496 244137 204502 244149
rect 204554 244137 204560 244189
rect 260080 244137 260086 244189
rect 260138 244177 260144 244189
rect 318064 244177 318070 244189
rect 260138 244149 318070 244177
rect 260138 244137 260144 244149
rect 318064 244137 318070 244149
rect 318122 244137 318128 244189
rect 112240 244063 112246 244115
rect 112298 244103 112304 244115
rect 206320 244103 206326 244115
rect 112298 244075 206326 244103
rect 112298 244063 112304 244075
rect 206320 244063 206326 244075
rect 206378 244063 206384 244115
rect 256336 244063 256342 244115
rect 256394 244103 256400 244115
rect 335344 244103 335350 244115
rect 256394 244075 335350 244103
rect 256394 244063 256400 244075
rect 335344 244063 335350 244075
rect 335402 244063 335408 244115
rect 109360 243989 109366 244041
rect 109418 244029 109424 244041
rect 206512 244029 206518 244041
rect 109418 244001 206518 244029
rect 109418 243989 109424 244001
rect 206512 243989 206518 244001
rect 206570 243989 206576 244041
rect 258352 243989 258358 244041
rect 258410 244029 258416 244041
rect 336304 244029 336310 244041
rect 258410 244001 336310 244029
rect 258410 243989 258416 244001
rect 336304 243989 336310 244001
rect 336362 243989 336368 244041
rect 106480 243915 106486 243967
rect 106538 243955 106544 243967
rect 205744 243955 205750 243967
rect 106538 243927 205750 243955
rect 106538 243915 106544 243927
rect 205744 243915 205750 243927
rect 205802 243915 205808 243967
rect 261136 243915 261142 243967
rect 261194 243955 261200 243967
rect 318160 243955 318166 243967
rect 261194 243927 318166 243955
rect 261194 243915 261200 243927
rect 318160 243915 318166 243927
rect 318218 243915 318224 243967
rect 103600 243841 103606 243893
rect 103658 243881 103664 243893
rect 206128 243881 206134 243893
rect 103658 243853 206134 243881
rect 103658 243841 103664 243853
rect 206128 243841 206134 243853
rect 206186 243841 206192 243893
rect 207184 243841 207190 243893
rect 207242 243881 207248 243893
rect 268144 243881 268150 243893
rect 207242 243853 268150 243881
rect 207242 243841 207248 243853
rect 268144 243841 268150 243853
rect 268202 243841 268208 243893
rect 268240 243841 268246 243893
rect 268298 243881 268304 243893
rect 287920 243881 287926 243893
rect 268298 243853 287926 243881
rect 268298 243841 268304 243853
rect 287920 243841 287926 243853
rect 287978 243841 287984 243893
rect 288016 243841 288022 243893
rect 288074 243881 288080 243893
rect 292144 243881 292150 243893
rect 288074 243853 292150 243881
rect 288074 243841 288080 243853
rect 292144 243841 292150 243853
rect 292202 243841 292208 243893
rect 292240 243841 292246 243893
rect 292298 243881 292304 243893
rect 307312 243881 307318 243893
rect 292298 243853 307318 243881
rect 292298 243841 292304 243853
rect 307312 243841 307318 243853
rect 307370 243841 307376 243893
rect 313360 243841 313366 243893
rect 313418 243881 313424 243893
rect 370288 243881 370294 243893
rect 313418 243853 370294 243881
rect 313418 243841 313424 243853
rect 370288 243841 370294 243853
rect 370346 243841 370352 243893
rect 100720 243767 100726 243819
rect 100778 243807 100784 243819
rect 206224 243807 206230 243819
rect 100778 243779 206230 243807
rect 100778 243767 100784 243779
rect 206224 243767 206230 243779
rect 206282 243767 206288 243819
rect 245392 243767 245398 243819
rect 245450 243807 245456 243819
rect 353680 243807 353686 243819
rect 245450 243779 353686 243807
rect 245450 243767 245456 243779
rect 353680 243767 353686 243779
rect 353738 243767 353744 243819
rect 94960 243693 94966 243745
rect 95018 243733 95024 243745
rect 205936 243733 205942 243745
rect 95018 243705 205942 243733
rect 95018 243693 95024 243705
rect 205936 243693 205942 243705
rect 205994 243693 206000 243745
rect 239344 243693 239350 243745
rect 239402 243733 239408 243745
rect 350800 243733 350806 243745
rect 239402 243705 350806 243733
rect 239402 243693 239408 243705
rect 350800 243693 350806 243705
rect 350858 243693 350864 243745
rect 92080 243619 92086 243671
rect 92138 243659 92144 243671
rect 206416 243659 206422 243671
rect 92138 243631 206422 243659
rect 92138 243619 92144 243631
rect 206416 243619 206422 243631
rect 206474 243619 206480 243671
rect 231760 243619 231766 243671
rect 231818 243659 231824 243671
rect 347344 243659 347350 243671
rect 231818 243631 347350 243659
rect 231818 243619 231824 243631
rect 347344 243619 347350 243631
rect 347402 243619 347408 243671
rect 86320 243545 86326 243597
rect 86378 243585 86384 243597
rect 206704 243585 206710 243597
rect 86378 243557 206710 243585
rect 86378 243545 86384 243557
rect 206704 243545 206710 243557
rect 206762 243545 206768 243597
rect 236272 243545 236278 243597
rect 236330 243585 236336 243597
rect 349264 243585 349270 243597
rect 236330 243557 349270 243585
rect 236330 243545 236336 243557
rect 349264 243545 349270 243557
rect 349322 243545 349328 243597
rect 80560 243471 80566 243523
rect 80618 243511 80624 243523
rect 206992 243511 206998 243523
rect 80618 243483 206998 243511
rect 80618 243471 80624 243483
rect 206992 243471 206998 243483
rect 207050 243471 207056 243523
rect 221200 243471 221206 243523
rect 221258 243511 221264 243523
rect 227440 243511 227446 243523
rect 221258 243483 227446 243511
rect 221258 243471 221264 243483
rect 227440 243471 227446 243483
rect 227498 243471 227504 243523
rect 229744 243471 229750 243523
rect 229802 243511 229808 243523
rect 346384 243511 346390 243523
rect 229802 243483 346390 243511
rect 229802 243471 229808 243483
rect 346384 243471 346390 243483
rect 346442 243471 346448 243523
rect 77680 243397 77686 243449
rect 77738 243437 77744 243449
rect 204592 243437 204598 243449
rect 77738 243409 204598 243437
rect 77738 243397 77744 243409
rect 204592 243397 204598 243409
rect 204650 243397 204656 243449
rect 226768 243397 226774 243449
rect 226826 243437 226832 243449
rect 345136 243437 345142 243449
rect 226826 243409 345142 243437
rect 226826 243397 226832 243409
rect 345136 243397 345142 243409
rect 345194 243397 345200 243449
rect 69040 243323 69046 243375
rect 69098 243363 69104 243375
rect 206032 243363 206038 243375
rect 69098 243335 206038 243363
rect 69098 243323 69104 243335
rect 206032 243323 206038 243335
rect 206090 243323 206096 243375
rect 228496 243323 228502 243375
rect 228554 243363 228560 243375
rect 345616 243363 345622 243375
rect 228554 243335 345622 243363
rect 228554 243323 228560 243335
rect 345616 243323 345622 243335
rect 345674 243323 345680 243375
rect 265936 243249 265942 243301
rect 265994 243289 266000 243301
rect 277840 243289 277846 243301
rect 265994 243261 277846 243289
rect 265994 243249 266000 243261
rect 277840 243249 277846 243261
rect 277898 243249 277904 243301
rect 283696 243249 283702 243301
rect 283754 243289 283760 243301
rect 298096 243289 298102 243301
rect 283754 243261 298102 243289
rect 283754 243249 283760 243261
rect 298096 243249 298102 243261
rect 298154 243249 298160 243301
rect 298288 243249 298294 243301
rect 298346 243289 298352 243301
rect 299632 243289 299638 243301
rect 298346 243261 299638 243289
rect 298346 243249 298352 243261
rect 299632 243249 299638 243261
rect 299690 243249 299696 243301
rect 302416 243249 302422 243301
rect 302474 243289 302480 243301
rect 312208 243289 312214 243301
rect 302474 243261 312214 243289
rect 302474 243249 302480 243261
rect 312208 243249 312214 243261
rect 312266 243249 312272 243301
rect 318256 243249 318262 243301
rect 318314 243289 318320 243301
rect 340720 243289 340726 243301
rect 318314 243261 340726 243289
rect 318314 243249 318320 243261
rect 340720 243249 340726 243261
rect 340778 243249 340784 243301
rect 226000 243175 226006 243227
rect 226058 243215 226064 243227
rect 236176 243215 236182 243227
rect 226058 243187 236182 243215
rect 226058 243175 226064 243187
rect 236176 243175 236182 243187
rect 236234 243175 236240 243227
rect 253360 243175 253366 243227
rect 253418 243215 253424 243227
rect 256240 243215 256246 243227
rect 253418 243187 256246 243215
rect 253418 243175 253424 243187
rect 256240 243175 256246 243187
rect 256298 243175 256304 243227
rect 267376 243175 267382 243227
rect 267434 243215 267440 243227
rect 267434 243187 298142 243215
rect 267434 243175 267440 243187
rect 262864 243101 262870 243153
rect 262922 243141 262928 243153
rect 277936 243141 277942 243153
rect 262922 243113 277942 243141
rect 262922 243101 262928 243113
rect 277936 243101 277942 243113
rect 277994 243101 278000 243153
rect 284944 243101 284950 243153
rect 285002 243141 285008 243153
rect 298000 243141 298006 243153
rect 285002 243113 298006 243141
rect 285002 243101 285008 243113
rect 298000 243101 298006 243113
rect 298058 243101 298064 243153
rect 298114 243141 298142 243187
rect 318160 243175 318166 243227
rect 318218 243215 318224 243227
rect 337552 243215 337558 243227
rect 318218 243187 337558 243215
rect 318218 243175 318224 243187
rect 337552 243175 337558 243187
rect 337610 243175 337616 243227
rect 305104 243141 305110 243153
rect 298114 243113 305110 243141
rect 305104 243101 305110 243113
rect 305162 243101 305168 243153
rect 310480 243101 310486 243153
rect 310538 243141 310544 243153
rect 339856 243141 339862 243153
rect 310538 243113 339862 243141
rect 310538 243101 310544 243113
rect 339856 243101 339862 243113
rect 339914 243101 339920 243153
rect 236176 243027 236182 243079
rect 236234 243067 236240 243079
rect 253360 243067 253366 243079
rect 236234 243039 253366 243067
rect 236234 243027 236240 243039
rect 253360 243027 253366 243039
rect 253418 243027 253424 243079
rect 270832 243027 270838 243079
rect 270890 243067 270896 243079
rect 291568 243067 291574 243079
rect 270890 243039 291574 243067
rect 270890 243027 270896 243039
rect 291568 243027 291574 243039
rect 291626 243027 291632 243079
rect 291760 243027 291766 243079
rect 291818 243067 291824 243079
rect 294736 243067 294742 243079
rect 291818 243039 294742 243067
rect 291818 243027 291824 243039
rect 294736 243027 294742 243039
rect 294794 243027 294800 243079
rect 295312 243027 295318 243079
rect 295370 243067 295376 243079
rect 303376 243067 303382 243079
rect 295370 243039 303382 243067
rect 295370 243027 295376 243039
rect 303376 243027 303382 243039
rect 303434 243027 303440 243079
rect 303472 243027 303478 243079
rect 303530 243067 303536 243079
rect 320368 243067 320374 243079
rect 303530 243039 320374 243067
rect 303530 243027 303536 243039
rect 320368 243027 320374 243039
rect 320426 243027 320432 243079
rect 266032 242953 266038 243005
rect 266090 242993 266096 243005
rect 277744 242993 277750 243005
rect 266090 242965 277750 242993
rect 266090 242953 266096 242965
rect 277744 242953 277750 242965
rect 277802 242953 277808 243005
rect 277840 242953 277846 243005
rect 277898 242993 277904 243005
rect 279376 242993 279382 243005
rect 277898 242965 279382 242993
rect 277898 242953 277904 242965
rect 279376 242953 279382 242965
rect 279434 242953 279440 243005
rect 283216 242953 283222 243005
rect 283274 242993 283280 243005
rect 302416 242993 302422 243005
rect 283274 242965 302422 242993
rect 283274 242953 283280 242965
rect 302416 242953 302422 242965
rect 302474 242953 302480 243005
rect 306448 242953 306454 243005
rect 306506 242993 306512 243005
rect 316720 242993 316726 243005
rect 306506 242965 316726 242993
rect 306506 242953 306512 242965
rect 316720 242953 316726 242965
rect 316778 242953 316784 243005
rect 318064 242953 318070 243005
rect 318122 242993 318128 243005
rect 337072 242993 337078 243005
rect 318122 242965 337078 242993
rect 318122 242953 318128 242965
rect 337072 242953 337078 242965
rect 337130 242953 337136 243005
rect 674992 242953 674998 243005
rect 675050 242993 675056 243005
rect 675376 242993 675382 243005
rect 675050 242965 675382 242993
rect 675050 242953 675056 242965
rect 675376 242953 675382 242965
rect 675434 242953 675440 243005
rect 268144 242879 268150 242931
rect 268202 242919 268208 242931
rect 287536 242919 287542 242931
rect 268202 242891 287542 242919
rect 268202 242879 268208 242891
rect 287536 242879 287542 242891
rect 287594 242879 287600 242931
rect 291376 242879 291382 242931
rect 291434 242919 291440 242931
rect 292816 242919 292822 242931
rect 291434 242891 292822 242919
rect 291434 242879 291440 242891
rect 292816 242879 292822 242891
rect 292874 242879 292880 242931
rect 292912 242879 292918 242931
rect 292970 242919 292976 242931
rect 302320 242919 302326 242931
rect 292970 242891 302326 242919
rect 292970 242879 292976 242891
rect 302320 242879 302326 242891
rect 302378 242879 302384 242931
rect 303088 242879 303094 242931
rect 303146 242919 303152 242931
rect 312592 242919 312598 242931
rect 303146 242891 312598 242919
rect 303146 242879 303152 242891
rect 312592 242879 312598 242891
rect 312650 242879 312656 242931
rect 316528 242879 316534 242931
rect 316586 242919 316592 242931
rect 316586 242891 317246 242919
rect 316586 242879 316592 242891
rect 266608 242805 266614 242857
rect 266666 242845 266672 242857
rect 278032 242845 278038 242857
rect 266666 242817 278038 242845
rect 266666 242805 266672 242817
rect 278032 242805 278038 242817
rect 278090 242805 278096 242857
rect 285904 242805 285910 242857
rect 285962 242845 285968 242857
rect 285962 242817 294782 242845
rect 285962 242805 285968 242817
rect 43408 242731 43414 242783
rect 43466 242771 43472 242783
rect 46192 242771 46198 242783
rect 43466 242743 46198 242771
rect 43466 242731 43472 242743
rect 46192 242731 46198 242743
rect 46250 242731 46256 242783
rect 269200 242731 269206 242783
rect 269258 242771 269264 242783
rect 294544 242771 294550 242783
rect 269258 242743 294550 242771
rect 269258 242731 269264 242743
rect 294544 242731 294550 242743
rect 294602 242731 294608 242783
rect 269680 242657 269686 242709
rect 269738 242697 269744 242709
rect 285520 242697 285526 242709
rect 269738 242669 285526 242697
rect 269738 242657 269744 242669
rect 285520 242657 285526 242669
rect 285578 242657 285584 242709
rect 285712 242657 285718 242709
rect 285770 242697 285776 242709
rect 291376 242697 291382 242709
rect 285770 242669 291382 242697
rect 285770 242657 285776 242669
rect 291376 242657 291382 242669
rect 291434 242657 291440 242709
rect 291568 242657 291574 242709
rect 291626 242697 291632 242709
rect 293392 242697 293398 242709
rect 291626 242669 293398 242697
rect 291626 242657 291632 242669
rect 293392 242657 293398 242669
rect 293450 242657 293456 242709
rect 293488 242657 293494 242709
rect 293546 242697 293552 242709
rect 294640 242697 294646 242709
rect 293546 242669 294646 242697
rect 293546 242657 293552 242669
rect 294640 242657 294646 242669
rect 294698 242657 294704 242709
rect 294754 242697 294782 242817
rect 295120 242805 295126 242857
rect 295178 242845 295184 242857
rect 297616 242845 297622 242857
rect 295178 242817 297622 242845
rect 295178 242805 295184 242817
rect 297616 242805 297622 242817
rect 297674 242805 297680 242857
rect 298000 242805 298006 242857
rect 298058 242845 298064 242857
rect 317104 242845 317110 242857
rect 298058 242817 317110 242845
rect 298058 242805 298064 242817
rect 317104 242805 317110 242817
rect 317162 242805 317168 242857
rect 317218 242845 317246 242891
rect 325072 242879 325078 242931
rect 325130 242919 325136 242931
rect 339568 242919 339574 242931
rect 325130 242891 339574 242919
rect 325130 242879 325136 242891
rect 339568 242879 339574 242891
rect 339626 242879 339632 242931
rect 331120 242845 331126 242857
rect 317218 242817 331126 242845
rect 331120 242805 331126 242817
rect 331178 242805 331184 242857
rect 295024 242731 295030 242783
rect 295082 242771 295088 242783
rect 297808 242771 297814 242783
rect 295082 242743 297814 242771
rect 295082 242731 295088 242743
rect 297808 242731 297814 242743
rect 297866 242731 297872 242783
rect 298096 242731 298102 242783
rect 298154 242771 298160 242783
rect 320080 242771 320086 242783
rect 298154 242743 320086 242771
rect 298154 242731 298160 242743
rect 320080 242731 320086 242743
rect 320138 242731 320144 242783
rect 314896 242697 314902 242709
rect 294754 242669 314902 242697
rect 314896 242657 314902 242669
rect 314954 242657 314960 242709
rect 314992 242657 314998 242709
rect 315050 242697 315056 242709
rect 316720 242697 316726 242709
rect 315050 242669 316726 242697
rect 315050 242657 315056 242669
rect 316720 242657 316726 242669
rect 316778 242657 316784 242709
rect 319696 242657 319702 242709
rect 319754 242697 319760 242709
rect 338512 242697 338518 242709
rect 319754 242669 338518 242697
rect 319754 242657 319760 242669
rect 338512 242657 338518 242669
rect 338570 242657 338576 242709
rect 463696 242657 463702 242709
rect 463754 242697 463760 242709
rect 483760 242697 483766 242709
rect 463754 242669 483766 242697
rect 463754 242657 463760 242669
rect 483760 242657 483766 242669
rect 483818 242657 483824 242709
rect 265264 242583 265270 242635
rect 265322 242623 265328 242635
rect 277360 242623 277366 242635
rect 265322 242595 277366 242623
rect 265322 242583 265328 242595
rect 277360 242583 277366 242595
rect 277418 242583 277424 242635
rect 295312 242623 295318 242635
rect 277666 242595 295318 242623
rect 269872 242509 269878 242561
rect 269930 242549 269936 242561
rect 277552 242549 277558 242561
rect 269930 242521 277558 242549
rect 269930 242509 269936 242521
rect 277552 242509 277558 242521
rect 277610 242509 277616 242561
rect 247504 242435 247510 242487
rect 247562 242475 247568 242487
rect 247562 242447 247742 242475
rect 247562 242435 247568 242447
rect 221968 242361 221974 242413
rect 222026 242401 222032 242413
rect 247600 242401 247606 242413
rect 222026 242373 247606 242401
rect 222026 242361 222032 242373
rect 247600 242361 247606 242373
rect 247658 242361 247664 242413
rect 247714 242327 247742 242447
rect 267856 242435 267862 242487
rect 267914 242475 267920 242487
rect 277666 242475 277694 242595
rect 295312 242583 295318 242595
rect 295370 242583 295376 242635
rect 299632 242583 299638 242635
rect 299690 242623 299696 242635
rect 322576 242623 322582 242635
rect 299690 242595 322582 242623
rect 299690 242583 299696 242595
rect 322576 242583 322582 242595
rect 322634 242583 322640 242635
rect 277840 242509 277846 242561
rect 277898 242549 277904 242561
rect 291760 242549 291766 242561
rect 277898 242521 291766 242549
rect 277898 242509 277904 242521
rect 291760 242509 291766 242521
rect 291818 242509 291824 242561
rect 314320 242549 314326 242561
rect 291874 242521 314326 242549
rect 267914 242447 277694 242475
rect 267914 242435 267920 242447
rect 285520 242435 285526 242487
rect 285578 242475 285584 242487
rect 286288 242475 286294 242487
rect 285578 242447 286294 242475
rect 285578 242435 285584 242447
rect 286288 242435 286294 242447
rect 286346 242435 286352 242487
rect 286480 242435 286486 242487
rect 286538 242475 286544 242487
rect 291874 242475 291902 242521
rect 314320 242509 314326 242521
rect 314378 242509 314384 242561
rect 317488 242509 317494 242561
rect 317546 242549 317552 242561
rect 317968 242549 317974 242561
rect 317546 242521 317974 242549
rect 317546 242509 317552 242521
rect 317968 242509 317974 242521
rect 318026 242509 318032 242561
rect 328144 242509 328150 242561
rect 328202 242549 328208 242561
rect 328528 242549 328534 242561
rect 328202 242521 328534 242549
rect 328202 242509 328208 242521
rect 328528 242509 328534 242521
rect 328586 242509 328592 242561
rect 443632 242509 443638 242561
rect 443690 242549 443696 242561
rect 453616 242549 453622 242561
rect 443690 242521 453622 242549
rect 443690 242509 443696 242521
rect 453616 242509 453622 242521
rect 453674 242509 453680 242561
rect 286538 242447 291902 242475
rect 286538 242435 286544 242447
rect 292144 242435 292150 242487
rect 292202 242475 292208 242487
rect 292912 242475 292918 242487
rect 292202 242447 292918 242475
rect 292202 242435 292208 242447
rect 292912 242435 292918 242447
rect 292970 242435 292976 242487
rect 293584 242435 293590 242487
rect 293642 242475 293648 242487
rect 323440 242475 323446 242487
rect 293642 242447 323446 242475
rect 293642 242435 293648 242447
rect 323440 242435 323446 242447
rect 323498 242435 323504 242487
rect 273520 242361 273526 242413
rect 273578 242401 273584 242413
rect 273578 242373 287870 242401
rect 273578 242361 273584 242373
rect 287728 242327 287734 242339
rect 247714 242299 287734 242327
rect 287728 242287 287734 242299
rect 287786 242287 287792 242339
rect 287842 242327 287870 242373
rect 287920 242361 287926 242413
rect 287978 242401 287984 242413
rect 303472 242401 303478 242413
rect 287978 242373 303478 242401
rect 287978 242361 287984 242373
rect 303472 242361 303478 242373
rect 303530 242361 303536 242413
rect 308944 242361 308950 242413
rect 309002 242401 309008 242413
rect 339760 242401 339766 242413
rect 309002 242373 339766 242401
rect 309002 242361 309008 242373
rect 339760 242361 339766 242373
rect 339818 242361 339824 242413
rect 430480 242361 430486 242413
rect 430538 242401 430544 242413
rect 443440 242401 443446 242413
rect 430538 242373 443446 242401
rect 430538 242361 430544 242373
rect 443440 242361 443446 242373
rect 443498 242361 443504 242413
rect 504016 242361 504022 242413
rect 504074 242401 504080 242413
rect 511120 242401 511126 242413
rect 504074 242373 511126 242401
rect 504074 242361 504080 242373
rect 511120 242361 511126 242373
rect 511178 242361 511184 242413
rect 355216 242327 355222 242339
rect 287842 242299 355222 242327
rect 355216 242287 355222 242299
rect 355274 242287 355280 242339
rect 39952 242213 39958 242265
rect 40010 242253 40016 242265
rect 42544 242253 42550 242265
rect 40010 242225 42550 242253
rect 40010 242213 40016 242225
rect 42544 242213 42550 242225
rect 42602 242213 42608 242265
rect 227344 242213 227350 242265
rect 227402 242253 227408 242265
rect 227728 242253 227734 242265
rect 227402 242225 227734 242253
rect 227402 242213 227408 242225
rect 227728 242213 227734 242225
rect 227786 242213 227792 242265
rect 244144 242213 244150 242265
rect 244202 242253 244208 242265
rect 353008 242253 353014 242265
rect 244202 242225 353014 242253
rect 244202 242213 244208 242225
rect 353008 242213 353014 242225
rect 353066 242213 353072 242265
rect 238288 242139 238294 242191
rect 238346 242179 238352 242191
rect 350032 242179 350038 242191
rect 238346 242151 350038 242179
rect 238346 242139 238352 242151
rect 350032 242139 350038 242151
rect 350090 242139 350096 242191
rect 39856 242065 39862 242117
rect 39914 242105 39920 242117
rect 42352 242105 42358 242117
rect 39914 242077 42358 242105
rect 39914 242065 39920 242077
rect 42352 242065 42358 242077
rect 42410 242065 42416 242117
rect 348688 242105 348694 242117
rect 241090 242077 348694 242105
rect 40048 241991 40054 242043
rect 40106 242031 40112 242043
rect 42544 242031 42550 242043
rect 40106 242003 42550 242031
rect 40106 241991 40112 242003
rect 42544 241991 42550 242003
rect 42602 241991 42608 242043
rect 241090 242031 241118 242077
rect 348688 242065 348694 242077
rect 348746 242065 348752 242117
rect 238882 242003 241118 242031
rect 40240 241917 40246 241969
rect 40298 241957 40304 241969
rect 43120 241957 43126 241969
rect 40298 241929 43126 241957
rect 40298 241917 40304 241929
rect 43120 241917 43126 241929
rect 43178 241917 43184 241969
rect 50320 241917 50326 241969
rect 50378 241957 50384 241969
rect 205840 241957 205846 241969
rect 50378 241929 205846 241957
rect 50378 241917 50384 241929
rect 205840 241917 205846 241929
rect 205898 241917 205904 241969
rect 218704 241843 218710 241895
rect 218762 241883 218768 241895
rect 234352 241883 234358 241895
rect 218762 241855 234358 241883
rect 218762 241843 218768 241855
rect 234352 241843 234358 241855
rect 234410 241843 234416 241895
rect 234544 241843 234550 241895
rect 234602 241883 234608 241895
rect 238882 241883 238910 242003
rect 241456 241991 241462 242043
rect 241514 242031 241520 242043
rect 351760 242031 351766 242043
rect 241514 242003 351766 242031
rect 241514 241991 241520 242003
rect 351760 241991 351766 242003
rect 351818 241991 351824 242043
rect 238960 241917 238966 241969
rect 239018 241957 239024 241969
rect 347824 241957 347830 241969
rect 239018 241929 347830 241957
rect 239018 241917 239024 241929
rect 347824 241917 347830 241929
rect 347882 241917 347888 241969
rect 234602 241855 238910 241883
rect 234602 241843 234608 241855
rect 248560 241843 248566 241895
rect 248618 241883 248624 241895
rect 273520 241883 273526 241895
rect 248618 241855 273526 241883
rect 248618 241843 248624 241855
rect 273520 241843 273526 241855
rect 273578 241843 273584 241895
rect 274000 241843 274006 241895
rect 274058 241883 274064 241895
rect 281968 241883 281974 241895
rect 274058 241855 281974 241883
rect 274058 241843 274064 241855
rect 281968 241843 281974 241855
rect 282026 241843 282032 241895
rect 286864 241843 286870 241895
rect 286922 241883 286928 241895
rect 297712 241883 297718 241895
rect 286922 241855 297718 241883
rect 286922 241843 286928 241855
rect 297712 241843 297718 241855
rect 297770 241843 297776 241895
rect 297808 241843 297814 241895
rect 297866 241883 297872 241895
rect 305008 241883 305014 241895
rect 297866 241855 305014 241883
rect 297866 241843 297872 241855
rect 305008 241843 305014 241855
rect 305066 241843 305072 241895
rect 317872 241843 317878 241895
rect 317930 241883 317936 241895
rect 327856 241883 327862 241895
rect 317930 241855 327862 241883
rect 317930 241843 317936 241855
rect 327856 241843 327862 241855
rect 327914 241843 327920 241895
rect 328048 241843 328054 241895
rect 328106 241883 328112 241895
rect 375088 241883 375094 241895
rect 328106 241855 375094 241883
rect 328106 241843 328112 241855
rect 375088 241843 375094 241855
rect 375146 241843 375152 241895
rect 378160 241843 378166 241895
rect 378218 241883 378224 241895
rect 378218 241855 398174 241883
rect 378218 241843 378224 241855
rect 215440 241769 215446 241821
rect 215498 241809 215504 241821
rect 221392 241809 221398 241821
rect 215498 241781 221398 241809
rect 215498 241769 215504 241781
rect 221392 241769 221398 241781
rect 221450 241769 221456 241821
rect 233488 241769 233494 241821
rect 233546 241809 233552 241821
rect 238960 241809 238966 241821
rect 233546 241781 238966 241809
rect 233546 241769 233552 241781
rect 238960 241769 238966 241781
rect 239018 241769 239024 241821
rect 239056 241769 239062 241821
rect 239114 241809 239120 241821
rect 260656 241809 260662 241821
rect 239114 241781 260662 241809
rect 239114 241769 239120 241781
rect 260656 241769 260662 241781
rect 260714 241769 260720 241821
rect 327952 241809 327958 241821
rect 262018 241781 327958 241809
rect 262018 241747 262046 241781
rect 327952 241769 327958 241781
rect 328010 241769 328016 241821
rect 328720 241769 328726 241821
rect 328778 241809 328784 241821
rect 333904 241809 333910 241821
rect 328778 241781 333910 241809
rect 328778 241769 328784 241781
rect 333904 241769 333910 241781
rect 333962 241769 333968 241821
rect 334480 241769 334486 241821
rect 334538 241809 334544 241821
rect 365872 241809 365878 241821
rect 334538 241781 365878 241809
rect 334538 241769 334544 241781
rect 365872 241769 365878 241781
rect 365930 241769 365936 241821
rect 377200 241769 377206 241821
rect 377258 241809 377264 241821
rect 395920 241809 395926 241821
rect 377258 241781 395926 241809
rect 377258 241769 377264 241781
rect 395920 241769 395926 241781
rect 395978 241769 395984 241821
rect 398146 241809 398174 241855
rect 407536 241809 407542 241821
rect 398146 241781 407542 241809
rect 407536 241769 407542 241781
rect 407594 241769 407600 241821
rect 219280 241695 219286 241747
rect 219338 241735 219344 241747
rect 233776 241735 233782 241747
rect 219338 241707 233782 241735
rect 219338 241695 219344 241707
rect 233776 241695 233782 241707
rect 233834 241695 233840 241747
rect 262000 241695 262006 241747
rect 262058 241695 262064 241747
rect 264304 241695 264310 241747
rect 264362 241735 264368 241747
rect 271984 241735 271990 241747
rect 264362 241707 271990 241735
rect 264362 241695 264368 241707
rect 271984 241695 271990 241707
rect 272042 241695 272048 241747
rect 278128 241695 278134 241747
rect 278186 241735 278192 241747
rect 329968 241735 329974 241747
rect 278186 241707 327998 241735
rect 278186 241695 278192 241707
rect 221488 241621 221494 241673
rect 221546 241661 221552 241673
rect 232912 241661 232918 241673
rect 221546 241633 232918 241661
rect 221546 241621 221552 241633
rect 232912 241621 232918 241633
rect 232970 241621 232976 241673
rect 236464 241621 236470 241673
rect 236522 241661 236528 241673
rect 264400 241661 264406 241673
rect 236522 241633 264406 241661
rect 236522 241621 236528 241633
rect 264400 241621 264406 241633
rect 264458 241621 264464 241673
rect 325168 241661 325174 241673
rect 269218 241633 325174 241661
rect 213904 241547 213910 241599
rect 213962 241587 213968 241599
rect 229168 241587 229174 241599
rect 213962 241559 229174 241587
rect 213962 241547 213968 241559
rect 229168 241547 229174 241559
rect 229226 241547 229232 241599
rect 252784 241547 252790 241599
rect 252842 241587 252848 241599
rect 269218 241587 269246 241633
rect 325168 241621 325174 241633
rect 325226 241621 325232 241673
rect 325264 241621 325270 241673
rect 325322 241661 325328 241673
rect 327856 241661 327862 241673
rect 325322 241633 327862 241661
rect 325322 241621 325328 241633
rect 327856 241621 327862 241633
rect 327914 241621 327920 241673
rect 327970 241661 327998 241707
rect 328162 241707 329974 241735
rect 328162 241661 328190 241707
rect 329968 241695 329974 241707
rect 330026 241695 330032 241747
rect 331024 241695 331030 241747
rect 331082 241735 331088 241747
rect 358288 241735 358294 241747
rect 331082 241707 358294 241735
rect 331082 241695 331088 241707
rect 358288 241695 358294 241707
rect 358346 241695 358352 241747
rect 361552 241695 361558 241747
rect 361610 241735 361616 241747
rect 396400 241735 396406 241747
rect 361610 241707 396406 241735
rect 361610 241695 361616 241707
rect 396400 241695 396406 241707
rect 396458 241695 396464 241747
rect 396514 241707 397406 241735
rect 327970 241633 328190 241661
rect 330064 241621 330070 241673
rect 330122 241661 330128 241673
rect 348400 241661 348406 241673
rect 330122 241633 348406 241661
rect 330122 241621 330128 241633
rect 348400 241621 348406 241633
rect 348458 241621 348464 241673
rect 363184 241621 363190 241673
rect 363242 241661 363248 241673
rect 396514 241661 396542 241707
rect 363242 241633 396542 241661
rect 397378 241661 397406 241707
rect 400144 241661 400150 241673
rect 397378 241633 400150 241661
rect 363242 241621 363248 241633
rect 400144 241621 400150 241633
rect 400202 241621 400208 241673
rect 252842 241559 269246 241587
rect 252842 241547 252848 241559
rect 269296 241547 269302 241599
rect 269354 241587 269360 241599
rect 317968 241587 317974 241599
rect 269354 241559 317974 241587
rect 269354 241547 269360 241559
rect 317968 241547 317974 241559
rect 318026 241547 318032 241599
rect 320464 241547 320470 241599
rect 320522 241587 320528 241599
rect 336112 241587 336118 241599
rect 320522 241559 336118 241587
rect 320522 241547 320528 241559
rect 336112 241547 336118 241559
rect 336170 241547 336176 241599
rect 348496 241547 348502 241599
rect 348554 241587 348560 241599
rect 356560 241587 356566 241599
rect 348554 241559 356566 241587
rect 348554 241547 348560 241559
rect 356560 241547 356566 241559
rect 356618 241547 356624 241599
rect 360976 241547 360982 241599
rect 361034 241587 361040 241599
rect 395824 241587 395830 241599
rect 361034 241559 395830 241587
rect 361034 241547 361040 241559
rect 395824 241547 395830 241559
rect 395882 241547 395888 241599
rect 395920 241547 395926 241599
rect 395978 241587 395984 241599
rect 405520 241587 405526 241599
rect 395978 241559 405526 241587
rect 395978 241547 395984 241559
rect 405520 241547 405526 241559
rect 405578 241547 405584 241599
rect 674032 241547 674038 241599
rect 674090 241587 674096 241599
rect 675472 241587 675478 241599
rect 674090 241559 675478 241587
rect 674090 241547 674096 241559
rect 675472 241547 675478 241559
rect 675530 241547 675536 241599
rect 223216 241473 223222 241525
rect 223274 241513 223280 241525
rect 232144 241513 232150 241525
rect 223274 241485 232150 241513
rect 223274 241473 223280 241485
rect 232144 241473 232150 241485
rect 232202 241473 232208 241525
rect 239152 241473 239158 241525
rect 239210 241513 239216 241525
rect 258544 241513 258550 241525
rect 239210 241485 258550 241513
rect 239210 241473 239216 241485
rect 258544 241473 258550 241485
rect 258602 241473 258608 241525
rect 278224 241473 278230 241525
rect 278282 241513 278288 241525
rect 318160 241513 318166 241525
rect 278282 241485 318166 241513
rect 278282 241473 278288 241485
rect 318160 241473 318166 241485
rect 318218 241473 318224 241525
rect 319504 241473 319510 241525
rect 319562 241513 319568 241525
rect 329584 241513 329590 241525
rect 319562 241485 329590 241513
rect 319562 241473 319568 241485
rect 329584 241473 329590 241485
rect 329642 241473 329648 241525
rect 331504 241473 331510 241525
rect 331562 241513 331568 241525
rect 359344 241513 359350 241525
rect 331562 241485 359350 241513
rect 331562 241473 331568 241485
rect 359344 241473 359350 241485
rect 359402 241473 359408 241525
rect 361936 241473 361942 241525
rect 361994 241513 362000 241525
rect 397456 241513 397462 241525
rect 361994 241485 397462 241513
rect 361994 241473 362000 241485
rect 397456 241473 397462 241485
rect 397514 241473 397520 241525
rect 255952 241399 255958 241451
rect 256010 241439 256016 241451
rect 318064 241439 318070 241451
rect 256010 241411 318070 241439
rect 256010 241399 256016 241411
rect 318064 241399 318070 241411
rect 318122 241399 318128 241451
rect 327376 241399 327382 241451
rect 327434 241439 327440 241451
rect 332944 241439 332950 241451
rect 327434 241411 332950 241439
rect 327434 241399 327440 241411
rect 332944 241399 332950 241411
rect 333002 241399 333008 241451
rect 364528 241399 364534 241451
rect 364586 241439 364592 241451
rect 402736 241439 402742 241451
rect 364586 241411 402742 241439
rect 364586 241399 364592 241411
rect 402736 241399 402742 241411
rect 402794 241399 402800 241451
rect 247408 241325 247414 241377
rect 247466 241365 247472 241377
rect 250384 241365 250390 241377
rect 247466 241337 250390 241365
rect 247466 241325 247472 241337
rect 250384 241325 250390 241337
rect 250442 241325 250448 241377
rect 254992 241325 254998 241377
rect 255050 241365 255056 241377
rect 318352 241365 318358 241377
rect 255050 241337 318358 241365
rect 255050 241325 255056 241337
rect 318352 241325 318358 241337
rect 318410 241325 318416 241377
rect 326704 241325 326710 241377
rect 326762 241365 326768 241377
rect 328912 241365 328918 241377
rect 326762 241337 328918 241365
rect 326762 241325 326768 241337
rect 328912 241325 328918 241337
rect 328970 241325 328976 241377
rect 329008 241325 329014 241377
rect 329066 241365 329072 241377
rect 347920 241365 347926 241377
rect 329066 241337 347926 241365
rect 329066 241325 329072 241337
rect 347920 241325 347926 241337
rect 347978 241325 347984 241377
rect 362320 241325 362326 241377
rect 362378 241365 362384 241377
rect 398416 241365 398422 241377
rect 362378 241337 398422 241365
rect 362378 241325 362384 241337
rect 398416 241325 398422 241337
rect 398474 241325 398480 241377
rect 226288 241251 226294 241303
rect 226346 241291 226352 241303
rect 230704 241291 230710 241303
rect 226346 241263 230710 241291
rect 226346 241251 226352 241263
rect 230704 241251 230710 241263
rect 230762 241251 230768 241303
rect 254224 241251 254230 241303
rect 254282 241291 254288 241303
rect 337840 241291 337846 241303
rect 254282 241263 337846 241291
rect 254282 241251 254288 241263
rect 337840 241251 337846 241263
rect 337898 241251 337904 241303
rect 363760 241251 363766 241303
rect 363818 241291 363824 241303
rect 400720 241291 400726 241303
rect 363818 241263 400726 241291
rect 363818 241251 363824 241263
rect 400720 241251 400726 241263
rect 400778 241251 400784 241303
rect 225424 241177 225430 241229
rect 225482 241217 225488 241229
rect 230896 241217 230902 241229
rect 225482 241189 230902 241217
rect 225482 241177 225488 241189
rect 230896 241177 230902 241189
rect 230954 241177 230960 241229
rect 253744 241177 253750 241229
rect 253802 241217 253808 241229
rect 339376 241217 339382 241229
rect 253802 241189 339382 241217
rect 253802 241177 253808 241189
rect 339376 241177 339382 241189
rect 339434 241177 339440 241229
rect 339472 241177 339478 241229
rect 339530 241217 339536 241229
rect 360496 241217 360502 241229
rect 339530 241189 360502 241217
rect 339530 241177 339536 241189
rect 360496 241177 360502 241189
rect 360554 241177 360560 241229
rect 364144 241177 364150 241229
rect 364202 241217 364208 241229
rect 401872 241217 401878 241229
rect 364202 241189 401878 241217
rect 364202 241177 364208 241189
rect 401872 241177 401878 241189
rect 401930 241177 401936 241229
rect 244720 241103 244726 241155
rect 244778 241143 244784 241155
rect 326896 241143 326902 241155
rect 244778 241115 326902 241143
rect 244778 241103 244784 241115
rect 326896 241103 326902 241115
rect 326954 241103 326960 241155
rect 326992 241103 326998 241155
rect 327050 241143 327056 241155
rect 330160 241143 330166 241155
rect 327050 241115 330166 241143
rect 327050 241103 327056 241115
rect 330160 241103 330166 241115
rect 330218 241103 330224 241155
rect 332272 241103 332278 241155
rect 332330 241143 332336 241155
rect 361072 241143 361078 241155
rect 332330 241115 361078 241143
rect 332330 241103 332336 241115
rect 361072 241103 361078 241115
rect 361130 241103 361136 241155
rect 362416 241103 362422 241155
rect 362474 241143 362480 241155
rect 398992 241143 398998 241155
rect 362474 241115 398998 241143
rect 362474 241103 362480 241115
rect 398992 241103 398998 241115
rect 399050 241103 399056 241155
rect 225232 241029 225238 241081
rect 225290 241069 225296 241081
rect 231184 241069 231190 241081
rect 225290 241041 231190 241069
rect 225290 241029 225296 241041
rect 231184 241029 231190 241041
rect 231242 241029 231248 241081
rect 237520 241029 237526 241081
rect 237578 241069 237584 241081
rect 254608 241069 254614 241081
rect 237578 241041 254614 241069
rect 237578 241029 237584 241041
rect 254608 241029 254614 241041
rect 254666 241029 254672 241081
rect 273136 241029 273142 241081
rect 273194 241069 273200 241081
rect 280432 241069 280438 241081
rect 273194 241041 280438 241069
rect 273194 241029 273200 241041
rect 280432 241029 280438 241041
rect 280490 241029 280496 241081
rect 280528 241029 280534 241081
rect 280586 241069 280592 241081
rect 290608 241069 290614 241081
rect 280586 241041 290614 241069
rect 280586 241029 280592 241041
rect 290608 241029 290614 241041
rect 290666 241029 290672 241081
rect 291952 241029 291958 241081
rect 292010 241069 292016 241081
rect 376144 241069 376150 241081
rect 292010 241041 376150 241069
rect 292010 241029 292016 241041
rect 376144 241029 376150 241041
rect 376202 241029 376208 241081
rect 379600 241029 379606 241081
rect 379658 241069 379664 241081
rect 409936 241069 409942 241081
rect 379658 241041 409942 241069
rect 379658 241029 379664 241041
rect 409936 241029 409942 241041
rect 409994 241029 410000 241081
rect 220432 240955 220438 241007
rect 220490 240995 220496 241007
rect 233392 240995 233398 241007
rect 220490 240967 233398 240995
rect 220490 240955 220496 240967
rect 233392 240955 233398 240967
rect 233450 240955 233456 241007
rect 237616 240955 237622 241007
rect 237674 240995 237680 241007
rect 252880 240995 252886 241007
rect 237674 240967 252886 240995
rect 237674 240955 237680 240967
rect 252880 240955 252886 240967
rect 252938 240955 252944 241007
rect 255088 240955 255094 241007
rect 255146 240995 255152 241007
rect 317872 240995 317878 241007
rect 255146 240967 317878 240995
rect 255146 240955 255152 240967
rect 317872 240955 317878 240967
rect 317930 240955 317936 241007
rect 318160 240955 318166 241007
rect 318218 240995 318224 241007
rect 331696 240995 331702 241007
rect 318218 240967 331702 240995
rect 318218 240955 318224 240967
rect 331696 240955 331702 240967
rect 331754 240955 331760 241007
rect 333712 240955 333718 241007
rect 333770 240995 333776 241007
rect 364336 240995 364342 241007
rect 333770 240967 364342 240995
rect 333770 240955 333776 240967
rect 364336 240955 364342 240967
rect 364394 240955 364400 241007
rect 367216 240955 367222 241007
rect 367274 240995 367280 241007
rect 408880 240995 408886 241007
rect 367274 240967 408886 240995
rect 367274 240955 367280 240967
rect 408880 240955 408886 240967
rect 408938 240955 408944 241007
rect 216688 240881 216694 240933
rect 216746 240921 216752 240933
rect 236176 240921 236182 240933
rect 216746 240893 236182 240921
rect 216746 240881 216752 240893
rect 236176 240881 236182 240893
rect 236234 240881 236240 240933
rect 237424 240881 237430 240933
rect 237482 240921 237488 240933
rect 248080 240921 248086 240933
rect 237482 240893 248086 240921
rect 237482 240881 237488 240893
rect 248080 240881 248086 240893
rect 248138 240881 248144 240933
rect 252304 240881 252310 240933
rect 252362 240921 252368 240933
rect 342640 240921 342646 240933
rect 252362 240893 342646 240921
rect 252362 240881 252368 240893
rect 342640 240881 342646 240893
rect 342698 240881 342704 240933
rect 365392 240881 365398 240933
rect 365450 240921 365456 240933
rect 405136 240921 405142 240933
rect 365450 240893 405142 240921
rect 365450 240881 365456 240893
rect 405136 240881 405142 240893
rect 405194 240881 405200 240933
rect 219280 240807 219286 240859
rect 219338 240847 219344 240859
rect 250672 240847 250678 240859
rect 219338 240819 250678 240847
rect 219338 240807 219344 240819
rect 250672 240807 250678 240819
rect 250730 240807 250736 240859
rect 251536 240807 251542 240859
rect 251594 240847 251600 240859
rect 344176 240847 344182 240859
rect 251594 240819 344182 240847
rect 251594 240807 251600 240819
rect 344176 240807 344182 240819
rect 344234 240807 344240 240859
rect 365968 240807 365974 240859
rect 366026 240847 366032 240859
rect 406096 240847 406102 240859
rect 366026 240819 406102 240847
rect 366026 240807 366032 240819
rect 406096 240807 406102 240819
rect 406154 240807 406160 240859
rect 232336 240733 232342 240785
rect 232394 240773 232400 240785
rect 238672 240773 238678 240785
rect 232394 240745 238678 240773
rect 232394 240733 232400 240745
rect 238672 240733 238678 240745
rect 238730 240733 238736 240785
rect 251824 240733 251830 240785
rect 251882 240773 251888 240785
rect 274384 240773 274390 240785
rect 251882 240745 274390 240773
rect 251882 240733 251888 240745
rect 274384 240733 274390 240745
rect 274442 240733 274448 240785
rect 274480 240733 274486 240785
rect 274538 240773 274544 240785
rect 281872 240773 281878 240785
rect 274538 240745 281878 240773
rect 274538 240733 274544 240745
rect 281872 240733 281878 240745
rect 281930 240733 281936 240785
rect 282256 240733 282262 240785
rect 282314 240773 282320 240785
rect 375760 240773 375766 240785
rect 282314 240745 375766 240773
rect 282314 240733 282320 240745
rect 375760 240733 375766 240745
rect 375818 240733 375824 240785
rect 379216 240733 379222 240785
rect 379274 240773 379280 240785
rect 409264 240773 409270 240785
rect 379274 240745 409270 240773
rect 379274 240733 379280 240745
rect 409264 240733 409270 240745
rect 409322 240733 409328 240785
rect 218800 240659 218806 240711
rect 218858 240699 218864 240711
rect 252016 240699 252022 240711
rect 218858 240671 252022 240699
rect 218858 240659 218864 240671
rect 252016 240659 252022 240671
rect 252074 240659 252080 240711
rect 345712 240699 345718 240711
rect 252130 240671 345718 240699
rect 41872 240585 41878 240637
rect 41930 240585 41936 240637
rect 212752 240585 212758 240637
rect 212810 240625 212816 240637
rect 233296 240625 233302 240637
rect 212810 240597 233302 240625
rect 212810 240585 212816 240597
rect 233296 240585 233302 240597
rect 233354 240585 233360 240637
rect 250576 240585 250582 240637
rect 250634 240625 250640 240637
rect 252130 240625 252158 240671
rect 345712 240659 345718 240671
rect 345770 240659 345776 240711
rect 366736 240659 366742 240711
rect 366794 240699 366800 240711
rect 407728 240699 407734 240711
rect 366794 240671 407734 240699
rect 366794 240659 366800 240671
rect 407728 240659 407734 240671
rect 407786 240659 407792 240711
rect 250634 240597 252158 240625
rect 250634 240585 250640 240597
rect 257872 240585 257878 240637
rect 257930 240625 257936 240637
rect 348016 240625 348022 240637
rect 257930 240597 348022 240625
rect 257930 240585 257936 240597
rect 348016 240585 348022 240597
rect 348074 240585 348080 240637
rect 365008 240585 365014 240637
rect 365066 240625 365072 240637
rect 404464 240625 404470 240637
rect 365066 240597 404470 240625
rect 365066 240585 365072 240597
rect 404464 240585 404470 240597
rect 404522 240585 404528 240637
rect 41890 240415 41918 240585
rect 221776 240511 221782 240563
rect 221834 240551 221840 240563
rect 237520 240551 237526 240563
rect 221834 240523 237526 240551
rect 221834 240511 221840 240523
rect 237520 240511 237526 240523
rect 237578 240511 237584 240563
rect 250192 240511 250198 240563
rect 250250 240551 250256 240563
rect 346288 240551 346294 240563
rect 250250 240523 346294 240551
rect 250250 240511 250256 240523
rect 346288 240511 346294 240523
rect 346346 240511 346352 240563
rect 364624 240511 364630 240563
rect 364682 240551 364688 240563
rect 403408 240551 403414 240563
rect 364682 240523 403414 240551
rect 364682 240511 364688 240523
rect 403408 240511 403414 240523
rect 403466 240511 403472 240563
rect 674128 240511 674134 240563
rect 674186 240551 674192 240563
rect 675472 240551 675478 240563
rect 674186 240523 675478 240551
rect 674186 240511 674192 240523
rect 675472 240511 675478 240523
rect 675530 240511 675536 240563
rect 220240 240437 220246 240489
rect 220298 240477 220304 240489
rect 248656 240477 248662 240489
rect 220298 240449 248662 240477
rect 220298 240437 220304 240449
rect 248656 240437 248662 240449
rect 248714 240437 248720 240489
rect 249712 240437 249718 240489
rect 249770 240477 249776 240489
rect 257680 240477 257686 240489
rect 249770 240449 257686 240477
rect 249770 240437 249776 240449
rect 257680 240437 257686 240449
rect 257738 240437 257744 240489
rect 257872 240437 257878 240489
rect 257930 240477 257936 240489
rect 350224 240477 350230 240489
rect 257930 240449 350230 240477
rect 257930 240437 257936 240449
rect 350224 240437 350230 240449
rect 350282 240437 350288 240489
rect 366352 240437 366358 240489
rect 366410 240477 366416 240489
rect 407152 240477 407158 240489
rect 366410 240449 407158 240477
rect 366410 240437 366416 240449
rect 407152 240437 407158 240449
rect 407210 240437 407216 240489
rect 607600 240437 607606 240489
rect 607658 240477 607664 240489
rect 627856 240477 627862 240489
rect 607658 240449 627862 240477
rect 607658 240437 607664 240449
rect 627856 240437 627862 240449
rect 627914 240437 627920 240489
rect 41872 240363 41878 240415
rect 41930 240363 41936 240415
rect 219664 240363 219670 240415
rect 219722 240403 219728 240415
rect 249808 240403 249814 240415
rect 219722 240375 249814 240403
rect 219722 240363 219728 240375
rect 249808 240363 249814 240375
rect 249866 240363 249872 240415
rect 274672 240363 274678 240415
rect 274730 240403 274736 240415
rect 283888 240403 283894 240415
rect 274730 240375 283894 240403
rect 274730 240363 274736 240375
rect 283888 240363 283894 240375
rect 283946 240363 283952 240415
rect 284080 240363 284086 240415
rect 284138 240403 284144 240415
rect 297328 240403 297334 240415
rect 284138 240375 297334 240403
rect 284138 240363 284144 240375
rect 297328 240363 297334 240375
rect 297386 240363 297392 240415
rect 297712 240363 297718 240415
rect 297770 240403 297776 240415
rect 313168 240403 313174 240415
rect 297770 240375 313174 240403
rect 297770 240363 297776 240375
rect 313168 240363 313174 240375
rect 313226 240363 313232 240415
rect 315184 240363 315190 240415
rect 315242 240403 315248 240415
rect 374416 240403 374422 240415
rect 315242 240375 374422 240403
rect 315242 240363 315248 240375
rect 374416 240363 374422 240375
rect 374474 240363 374480 240415
rect 377008 240363 377014 240415
rect 377066 240403 377072 240415
rect 404944 240403 404950 240415
rect 377066 240375 404950 240403
rect 377066 240363 377072 240375
rect 404944 240363 404950 240375
rect 405002 240363 405008 240415
rect 218416 240289 218422 240341
rect 218474 240329 218480 240341
rect 237616 240329 237622 240341
rect 218474 240301 237622 240329
rect 218474 240289 218480 240301
rect 237616 240289 237622 240301
rect 237674 240289 237680 240341
rect 240880 240289 240886 240341
rect 240938 240329 240944 240341
rect 255088 240329 255094 240341
rect 240938 240301 255094 240329
rect 240938 240289 240944 240301
rect 255088 240289 255094 240301
rect 255146 240289 255152 240341
rect 262096 240289 262102 240341
rect 262154 240329 262160 240341
rect 278128 240329 278134 240341
rect 262154 240301 278134 240329
rect 262154 240289 262160 240301
rect 278128 240289 278134 240301
rect 278186 240289 278192 240341
rect 278320 240289 278326 240341
rect 278378 240329 278384 240341
rect 283984 240329 283990 240341
rect 278378 240301 283990 240329
rect 278378 240289 278384 240301
rect 283984 240289 283990 240301
rect 284042 240289 284048 240341
rect 287248 240289 287254 240341
rect 287306 240329 287312 240341
rect 303088 240329 303094 240341
rect 287306 240301 303094 240329
rect 287306 240289 287312 240301
rect 303088 240289 303094 240301
rect 303146 240289 303152 240341
rect 306544 240289 306550 240341
rect 306602 240329 306608 240341
rect 308944 240329 308950 240341
rect 306602 240301 308950 240329
rect 306602 240289 306608 240301
rect 308944 240289 308950 240301
rect 309002 240289 309008 240341
rect 313648 240289 313654 240341
rect 313706 240329 313712 240341
rect 371824 240329 371830 240341
rect 313706 240301 371830 240329
rect 313706 240289 313712 240301
rect 371824 240289 371830 240301
rect 371882 240289 371888 240341
rect 378256 240289 378262 240341
rect 378314 240329 378320 240341
rect 408304 240329 408310 240341
rect 378314 240301 408310 240329
rect 378314 240289 378320 240301
rect 408304 240289 408310 240301
rect 408362 240289 408368 240341
rect 237904 240215 237910 240267
rect 237962 240255 237968 240267
rect 261616 240255 261622 240267
rect 237962 240227 261622 240255
rect 237962 240215 237968 240227
rect 261616 240215 261622 240227
rect 261674 240215 261680 240267
rect 269296 240255 269302 240267
rect 264034 240227 269302 240255
rect 217552 240141 217558 240193
rect 217610 240181 217616 240193
rect 234736 240181 234742 240193
rect 217610 240153 234742 240181
rect 217610 240141 217616 240153
rect 234736 240141 234742 240153
rect 234794 240141 234800 240193
rect 236944 240141 236950 240193
rect 237002 240181 237008 240193
rect 263344 240181 263350 240193
rect 237002 240153 263350 240181
rect 237002 240141 237008 240153
rect 263344 240141 263350 240153
rect 263402 240141 263408 240193
rect 42352 240067 42358 240119
rect 42410 240107 42416 240119
rect 43312 240107 43318 240119
rect 42410 240079 43318 240107
rect 42410 240067 42416 240079
rect 43312 240067 43318 240079
rect 43370 240067 43376 240119
rect 222544 240067 222550 240119
rect 222602 240107 222608 240119
rect 232528 240107 232534 240119
rect 222602 240079 232534 240107
rect 222602 240067 222608 240079
rect 232528 240067 232534 240079
rect 232586 240067 232592 240119
rect 237328 240067 237334 240119
rect 237386 240107 237392 240119
rect 262192 240107 262198 240119
rect 237386 240079 262198 240107
rect 237386 240067 237392 240079
rect 262192 240067 262198 240079
rect 262250 240067 262256 240119
rect 220624 239993 220630 240045
rect 220682 240033 220688 240045
rect 237424 240033 237430 240045
rect 220682 240005 237430 240033
rect 220682 239993 220688 240005
rect 237424 239993 237430 240005
rect 237482 239993 237488 240045
rect 263920 240033 263926 240045
rect 248866 240005 263926 240033
rect 236560 239919 236566 239971
rect 236618 239959 236624 239971
rect 236618 239931 247646 239959
rect 236618 239919 236624 239931
rect 247618 239885 247646 239931
rect 248866 239885 248894 240005
rect 263920 239993 263926 240005
rect 263978 239993 263984 240045
rect 247618 239857 248894 239885
rect 256432 239845 256438 239897
rect 256490 239885 256496 239897
rect 264034 239885 264062 240227
rect 269296 240215 269302 240227
rect 269354 240215 269360 240267
rect 277456 240215 277462 240267
rect 277514 240255 277520 240267
rect 295600 240255 295606 240267
rect 277514 240227 295606 240255
rect 277514 240215 277520 240227
rect 295600 240215 295606 240227
rect 295658 240215 295664 240267
rect 312112 240255 312118 240267
rect 295714 240227 312118 240255
rect 275728 240141 275734 240193
rect 275786 240181 275792 240193
rect 281680 240181 281686 240193
rect 275786 240153 281686 240181
rect 275786 240141 275792 240153
rect 281680 240141 281686 240153
rect 281738 240141 281744 240193
rect 281872 240141 281878 240193
rect 281930 240181 281936 240193
rect 289456 240181 289462 240193
rect 281930 240153 289462 240181
rect 281930 240141 281936 240153
rect 289456 240141 289462 240153
rect 289514 240141 289520 240193
rect 291088 240141 291094 240193
rect 291146 240181 291152 240193
rect 293296 240181 293302 240193
rect 291146 240153 293302 240181
rect 291146 240141 291152 240153
rect 293296 240141 293302 240153
rect 293354 240141 293360 240193
rect 293776 240141 293782 240193
rect 293834 240181 293840 240193
rect 295714 240181 295742 240227
rect 312112 240215 312118 240227
rect 312170 240215 312176 240267
rect 314608 240215 314614 240267
rect 314666 240255 314672 240267
rect 373552 240255 373558 240267
rect 314666 240227 373558 240255
rect 314666 240215 314672 240227
rect 373552 240215 373558 240227
rect 373610 240215 373616 240267
rect 376432 240215 376438 240267
rect 376490 240255 376496 240267
rect 404080 240255 404086 240267
rect 376490 240227 404086 240255
rect 376490 240215 376496 240227
rect 404080 240215 404086 240227
rect 404138 240215 404144 240267
rect 293834 240153 295742 240181
rect 293834 240141 293840 240153
rect 297136 240141 297142 240193
rect 297194 240181 297200 240193
rect 304432 240181 304438 240193
rect 297194 240153 304438 240181
rect 297194 240141 297200 240153
rect 304432 240141 304438 240153
rect 304490 240141 304496 240193
rect 313744 240141 313750 240193
rect 313802 240181 313808 240193
rect 371344 240181 371350 240193
rect 313802 240153 371350 240181
rect 313802 240141 313808 240153
rect 371344 240141 371350 240153
rect 371402 240141 371408 240193
rect 381808 240141 381814 240193
rect 381866 240181 381872 240193
rect 389872 240181 389878 240193
rect 381866 240153 389878 240181
rect 381866 240141 381872 240153
rect 389872 240141 389878 240153
rect 389930 240141 389936 240193
rect 272464 240067 272470 240119
rect 272522 240107 272528 240119
rect 285520 240107 285526 240119
rect 272522 240079 285526 240107
rect 272522 240067 272528 240079
rect 285520 240067 285526 240079
rect 285578 240067 285584 240119
rect 289552 240067 289558 240119
rect 289610 240107 289616 240119
rect 289610 240079 295358 240107
rect 289610 240067 289616 240079
rect 275440 239993 275446 240045
rect 275498 240033 275504 240045
rect 287440 240033 287446 240045
rect 275498 240005 287446 240033
rect 275498 239993 275504 240005
rect 287440 239993 287446 240005
rect 287498 239993 287504 240045
rect 288688 239993 288694 240045
rect 288746 240033 288752 240045
rect 291856 240033 291862 240045
rect 288746 240005 291862 240033
rect 288746 239993 288752 240005
rect 291856 239993 291862 240005
rect 291914 239993 291920 240045
rect 279472 239919 279478 239971
rect 279530 239959 279536 239971
rect 282160 239959 282166 239971
rect 279530 239931 282166 239959
rect 279530 239919 279536 239931
rect 282160 239919 282166 239931
rect 282218 239919 282224 239971
rect 284848 239919 284854 239971
rect 284906 239959 284912 239971
rect 287824 239959 287830 239971
rect 284906 239931 287830 239959
rect 284906 239919 284912 239931
rect 287824 239919 287830 239931
rect 287882 239919 287888 239971
rect 290416 239919 290422 239971
rect 290474 239959 290480 239971
rect 295216 239959 295222 239971
rect 290474 239931 295222 239959
rect 290474 239919 290480 239931
rect 295216 239919 295222 239931
rect 295274 239919 295280 239971
rect 295330 239959 295358 240079
rect 314224 240067 314230 240119
rect 314282 240107 314288 240119
rect 372400 240107 372406 240119
rect 314282 240079 372406 240107
rect 314282 240067 314288 240079
rect 372400 240067 372406 240079
rect 372458 240067 372464 240119
rect 376048 240067 376054 240119
rect 376106 240107 376112 240119
rect 403216 240107 403222 240119
rect 376106 240079 403222 240107
rect 376106 240067 376112 240079
rect 403216 240067 403222 240079
rect 403274 240067 403280 240119
rect 296272 239993 296278 240045
rect 296330 240033 296336 240045
rect 329104 240033 329110 240045
rect 296330 240005 329110 240033
rect 296330 239993 296336 240005
rect 329104 239993 329110 240005
rect 329162 239993 329168 240045
rect 329680 239993 329686 240045
rect 329738 240033 329744 240045
rect 355696 240033 355702 240045
rect 329738 240005 355702 240033
rect 329738 239993 329744 240005
rect 355696 239993 355702 240005
rect 355754 239993 355760 240045
rect 360208 239993 360214 240045
rect 360266 240033 360272 240045
rect 360266 240005 368750 240033
rect 360266 239993 360272 240005
rect 314800 239959 314806 239971
rect 295330 239931 314806 239959
rect 314800 239919 314806 239931
rect 314858 239919 314864 239971
rect 317872 239919 317878 239971
rect 317930 239959 317936 239971
rect 326992 239959 326998 239971
rect 317930 239931 326998 239959
rect 317930 239919 317936 239931
rect 326992 239919 326998 239931
rect 327050 239919 327056 239971
rect 328240 239919 328246 239971
rect 328298 239959 328304 239971
rect 352432 239959 352438 239971
rect 328298 239931 352438 239959
rect 328298 239919 328304 239931
rect 352432 239919 352438 239931
rect 352490 239919 352496 239971
rect 256490 239857 264062 239885
rect 256490 239845 256496 239857
rect 268720 239845 268726 239897
rect 268778 239885 268784 239897
rect 280144 239885 280150 239897
rect 268778 239857 280150 239885
rect 268778 239845 268784 239857
rect 280144 239845 280150 239857
rect 280202 239845 280208 239897
rect 280432 239845 280438 239897
rect 280490 239885 280496 239897
rect 283024 239885 283030 239897
rect 280490 239857 283030 239885
rect 280490 239845 280496 239857
rect 283024 239845 283030 239857
rect 283082 239845 283088 239897
rect 283984 239845 283990 239897
rect 284042 239885 284048 239897
rect 291664 239885 291670 239897
rect 284042 239857 291670 239885
rect 284042 239845 284048 239857
rect 291664 239845 291670 239857
rect 291722 239845 291728 239897
rect 313840 239885 313846 239897
rect 291778 239857 313846 239885
rect 149584 239771 149590 239823
rect 149642 239811 149648 239823
rect 157744 239811 157750 239823
rect 149642 239783 157750 239811
rect 149642 239771 149648 239783
rect 157744 239771 157750 239783
rect 157802 239771 157808 239823
rect 248368 239771 248374 239823
rect 248426 239811 248432 239823
rect 257872 239811 257878 239823
rect 248426 239783 257878 239811
rect 248426 239771 248432 239783
rect 257872 239771 257878 239783
rect 257930 239771 257936 239823
rect 274192 239771 274198 239823
rect 274250 239811 274256 239823
rect 281488 239811 281494 239823
rect 274250 239783 281494 239811
rect 274250 239771 274256 239783
rect 281488 239771 281494 239783
rect 281546 239771 281552 239823
rect 284080 239811 284086 239823
rect 281602 239783 284086 239811
rect 214480 239697 214486 239749
rect 214538 239737 214544 239749
rect 225136 239737 225142 239749
rect 214538 239709 225142 239737
rect 214538 239697 214544 239709
rect 225136 239697 225142 239709
rect 225194 239697 225200 239749
rect 228016 239697 228022 239749
rect 228074 239737 228080 239749
rect 229936 239737 229942 239749
rect 228074 239709 229942 239737
rect 228074 239697 228080 239709
rect 229936 239697 229942 239709
rect 229994 239697 230000 239749
rect 268240 239697 268246 239749
rect 268298 239737 268304 239749
rect 270928 239737 270934 239749
rect 268298 239709 270934 239737
rect 268298 239697 268304 239709
rect 270928 239697 270934 239709
rect 270986 239697 270992 239749
rect 275824 239697 275830 239749
rect 275882 239737 275888 239749
rect 280528 239737 280534 239749
rect 275882 239709 280534 239737
rect 275882 239697 275888 239709
rect 280528 239697 280534 239709
rect 280586 239697 280592 239749
rect 215920 239623 215926 239675
rect 215978 239663 215984 239675
rect 218896 239663 218902 239675
rect 215978 239635 218902 239663
rect 215978 239623 215984 239635
rect 218896 239623 218902 239635
rect 218954 239623 218960 239675
rect 229072 239623 229078 239675
rect 229130 239663 229136 239675
rect 230224 239663 230230 239675
rect 229130 239635 230230 239663
rect 229130 239623 229136 239635
rect 230224 239623 230230 239635
rect 230282 239623 230288 239675
rect 257200 239623 257206 239675
rect 257258 239663 257264 239675
rect 269296 239663 269302 239675
rect 257258 239635 269302 239663
rect 257258 239623 257264 239635
rect 269296 239623 269302 239635
rect 269354 239623 269360 239675
rect 270256 239623 270262 239675
rect 270314 239663 270320 239675
rect 272272 239663 272278 239675
rect 270314 239635 272278 239663
rect 270314 239623 270320 239635
rect 272272 239623 272278 239635
rect 272330 239623 272336 239675
rect 273520 239623 273526 239675
rect 273578 239663 273584 239675
rect 278320 239663 278326 239675
rect 273578 239635 278326 239663
rect 273578 239623 273584 239635
rect 278320 239623 278326 239635
rect 278378 239623 278384 239675
rect 278896 239623 278902 239675
rect 278954 239663 278960 239675
rect 279664 239663 279670 239675
rect 278954 239635 279670 239663
rect 278954 239623 278960 239635
rect 279664 239623 279670 239635
rect 279722 239623 279728 239675
rect 279760 239623 279766 239675
rect 279818 239663 279824 239675
rect 281602 239663 281630 239783
rect 284080 239771 284086 239783
rect 284138 239771 284144 239823
rect 289456 239771 289462 239823
rect 289514 239811 289520 239823
rect 291778 239811 291806 239857
rect 313840 239845 313846 239857
rect 313898 239845 313904 239897
rect 324400 239845 324406 239897
rect 324458 239885 324464 239897
rect 324458 239857 329246 239885
rect 324458 239845 324464 239857
rect 289514 239783 291806 239811
rect 289514 239771 289520 239783
rect 291856 239771 291862 239823
rect 291914 239811 291920 239823
rect 293776 239811 293782 239823
rect 291914 239783 293782 239811
rect 291914 239771 291920 239783
rect 293776 239771 293782 239783
rect 293834 239771 293840 239823
rect 294256 239771 294262 239823
rect 294314 239811 294320 239823
rect 303568 239811 303574 239823
rect 294314 239783 303574 239811
rect 294314 239771 294320 239783
rect 303568 239771 303574 239783
rect 303626 239771 303632 239823
rect 315568 239771 315574 239823
rect 315626 239811 315632 239823
rect 325264 239811 325270 239823
rect 315626 239783 325270 239811
rect 315626 239771 315632 239783
rect 325264 239771 325270 239783
rect 325322 239771 325328 239823
rect 326224 239771 326230 239823
rect 326282 239811 326288 239823
rect 329008 239811 329014 239823
rect 326282 239783 329014 239811
rect 326282 239771 326288 239783
rect 329008 239771 329014 239783
rect 329066 239771 329072 239823
rect 329218 239811 329246 239857
rect 329296 239845 329302 239897
rect 329354 239885 329360 239897
rect 354544 239885 354550 239897
rect 329354 239857 354550 239885
rect 329354 239845 329360 239857
rect 354544 239845 354550 239857
rect 354602 239845 354608 239897
rect 343696 239811 343702 239823
rect 329218 239783 343702 239811
rect 343696 239771 343702 239783
rect 343754 239771 343760 239823
rect 282160 239697 282166 239749
rect 282218 239737 282224 239749
rect 296560 239737 296566 239749
rect 282218 239709 296566 239737
rect 282218 239697 282224 239709
rect 296560 239697 296566 239709
rect 296618 239697 296624 239749
rect 297616 239697 297622 239749
rect 297674 239737 297680 239749
rect 301072 239737 301078 239749
rect 297674 239709 301078 239737
rect 297674 239697 297680 239709
rect 301072 239697 301078 239709
rect 301130 239697 301136 239749
rect 301840 239697 301846 239749
rect 301898 239737 301904 239749
rect 306640 239737 306646 239749
rect 301898 239709 306646 239737
rect 301898 239697 301904 239709
rect 306640 239697 306646 239709
rect 306698 239697 306704 239749
rect 312784 239737 312790 239749
rect 309442 239709 312790 239737
rect 279818 239635 281630 239663
rect 279818 239623 279824 239635
rect 281680 239623 281686 239675
rect 281738 239663 281744 239675
rect 281738 239635 293150 239663
rect 281738 239623 281744 239635
rect 227248 239549 227254 239601
rect 227306 239589 227312 239601
rect 230320 239589 230326 239601
rect 227306 239561 230326 239589
rect 227306 239549 227312 239561
rect 230320 239549 230326 239561
rect 230378 239549 230384 239601
rect 269392 239549 269398 239601
rect 269450 239589 269456 239601
rect 276304 239589 276310 239601
rect 269450 239561 276310 239589
rect 269450 239549 269456 239561
rect 276304 239549 276310 239561
rect 276362 239549 276368 239601
rect 277648 239549 277654 239601
rect 277706 239589 277712 239601
rect 282928 239589 282934 239601
rect 277706 239561 282934 239589
rect 277706 239549 277712 239561
rect 282928 239549 282934 239561
rect 282986 239549 282992 239601
rect 283024 239549 283030 239601
rect 283082 239589 283088 239601
rect 292144 239589 292150 239601
rect 283082 239561 292150 239589
rect 283082 239549 283088 239561
rect 292144 239549 292150 239561
rect 292202 239549 292208 239601
rect 293122 239589 293150 239635
rect 293200 239623 293206 239675
rect 293258 239663 293264 239675
rect 302800 239663 302806 239675
rect 293258 239635 302806 239663
rect 293258 239623 293264 239635
rect 302800 239623 302806 239635
rect 302858 239623 302864 239675
rect 302992 239623 302998 239675
rect 303050 239663 303056 239675
rect 307600 239663 307606 239675
rect 303050 239635 307606 239663
rect 303050 239623 303056 239635
rect 307600 239623 307606 239635
rect 307658 239623 307664 239675
rect 307888 239623 307894 239675
rect 307946 239663 307952 239675
rect 309442 239663 309470 239709
rect 312784 239697 312790 239709
rect 312842 239697 312848 239749
rect 322672 239697 322678 239749
rect 322730 239737 322736 239749
rect 322730 239709 324830 239737
rect 322730 239697 322736 239709
rect 307946 239635 309470 239663
rect 307946 239623 307952 239635
rect 309520 239623 309526 239675
rect 309578 239663 309584 239675
rect 310288 239663 310294 239675
rect 309578 239635 310294 239663
rect 309578 239623 309584 239635
rect 310288 239623 310294 239635
rect 310346 239623 310352 239675
rect 320848 239623 320854 239675
rect 320906 239663 320912 239675
rect 324688 239663 324694 239675
rect 320906 239635 324694 239663
rect 320906 239623 320912 239635
rect 324688 239623 324694 239635
rect 324746 239623 324752 239675
rect 324802 239663 324830 239709
rect 326992 239697 326998 239749
rect 327050 239737 327056 239749
rect 349552 239737 349558 239749
rect 327050 239709 349558 239737
rect 327050 239697 327056 239709
rect 349552 239697 349558 239709
rect 349610 239697 349616 239749
rect 340912 239663 340918 239675
rect 324802 239635 340918 239663
rect 340912 239623 340918 239635
rect 340970 239623 340976 239675
rect 294736 239589 294742 239601
rect 293122 239561 294742 239589
rect 294736 239549 294742 239561
rect 294794 239549 294800 239601
rect 295984 239549 295990 239601
rect 296042 239589 296048 239601
rect 304144 239589 304150 239601
rect 296042 239561 304150 239589
rect 296042 239549 296048 239561
rect 304144 239549 304150 239561
rect 304202 239549 304208 239601
rect 308848 239549 308854 239601
rect 308906 239589 308912 239601
rect 310192 239589 310198 239601
rect 308906 239561 310198 239589
rect 308906 239549 308912 239561
rect 310192 239549 310198 239561
rect 310250 239549 310256 239601
rect 323056 239549 323062 239601
rect 323114 239589 323120 239601
rect 341296 239589 341302 239601
rect 323114 239561 341302 239589
rect 323114 239549 323120 239561
rect 341296 239549 341302 239561
rect 341354 239549 341360 239601
rect 277072 239475 277078 239527
rect 277130 239515 277136 239527
rect 283792 239515 283798 239527
rect 277130 239487 283798 239515
rect 277130 239475 277136 239487
rect 283792 239475 283798 239487
rect 283850 239475 283856 239527
rect 283888 239475 283894 239527
rect 283946 239515 283952 239527
rect 294352 239515 294358 239527
rect 283946 239487 294358 239515
rect 283946 239475 283952 239487
rect 294352 239475 294358 239487
rect 294410 239475 294416 239527
rect 322192 239475 322198 239527
rect 322250 239515 322256 239527
rect 338896 239515 338902 239527
rect 322250 239487 338902 239515
rect 322250 239475 322256 239487
rect 338896 239475 338902 239487
rect 338954 239475 338960 239527
rect 271024 239401 271030 239453
rect 271082 239441 271088 239453
rect 277936 239441 277942 239453
rect 271082 239413 277942 239441
rect 271082 239401 271088 239413
rect 277936 239401 277942 239413
rect 277994 239401 278000 239453
rect 278032 239401 278038 239453
rect 278090 239441 278096 239453
rect 281776 239441 281782 239453
rect 278090 239413 281782 239441
rect 278090 239401 278096 239413
rect 281776 239401 281782 239413
rect 281834 239401 281840 239453
rect 281968 239401 281974 239453
rect 282026 239441 282032 239453
rect 290800 239441 290806 239453
rect 282026 239413 290806 239441
rect 282026 239401 282032 239413
rect 290800 239401 290806 239413
rect 290858 239401 290864 239453
rect 290992 239401 290998 239453
rect 291050 239441 291056 239453
rect 307888 239441 307894 239453
rect 291050 239413 307894 239441
rect 291050 239401 291056 239413
rect 307888 239401 307894 239413
rect 307946 239401 307952 239453
rect 323440 239401 323446 239453
rect 323498 239441 323504 239453
rect 341968 239441 341974 239453
rect 323498 239413 341974 239441
rect 323498 239401 323504 239413
rect 341968 239401 341974 239413
rect 342026 239401 342032 239453
rect 240304 239327 240310 239379
rect 240362 239367 240368 239379
rect 244144 239367 244150 239379
rect 240362 239339 244150 239367
rect 240362 239327 240368 239339
rect 244144 239327 244150 239339
rect 244202 239327 244208 239379
rect 276688 239327 276694 239379
rect 276746 239367 276752 239379
rect 284464 239367 284470 239379
rect 276746 239339 284470 239367
rect 276746 239327 276752 239339
rect 284464 239327 284470 239339
rect 284522 239327 284528 239379
rect 285040 239327 285046 239379
rect 285098 239367 285104 239379
rect 298864 239367 298870 239379
rect 285098 239339 298870 239367
rect 285098 239327 285104 239339
rect 298864 239327 298870 239339
rect 298922 239327 298928 239379
rect 307792 239327 307798 239379
rect 307850 239367 307856 239379
rect 309808 239367 309814 239379
rect 307850 239339 309814 239367
rect 307850 239327 307856 239339
rect 309808 239327 309814 239339
rect 309866 239327 309872 239379
rect 321232 239327 321238 239379
rect 321290 239367 321296 239379
rect 337168 239367 337174 239379
rect 321290 239339 337174 239367
rect 321290 239327 321296 239339
rect 337168 239327 337174 239339
rect 337226 239327 337232 239379
rect 368722 239367 368750 240005
rect 377776 239993 377782 240045
rect 377834 240033 377840 240045
rect 406672 240033 406678 240045
rect 377834 240005 406678 240033
rect 377834 239993 377840 240005
rect 406672 239993 406678 240005
rect 406730 239993 406736 240045
rect 375664 239919 375670 239971
rect 375722 239959 375728 239971
rect 375722 239931 383966 239959
rect 375722 239919 375728 239931
rect 378640 239845 378646 239897
rect 378698 239885 378704 239897
rect 383824 239885 383830 239897
rect 378698 239857 383830 239885
rect 378698 239845 378704 239857
rect 383824 239845 383830 239857
rect 383882 239845 383888 239897
rect 383938 239885 383966 239931
rect 384016 239919 384022 239971
rect 384074 239959 384080 239971
rect 398608 239959 398614 239971
rect 384074 239931 398614 239959
rect 384074 239919 384080 239931
rect 398608 239919 398614 239931
rect 398666 239919 398672 239971
rect 402352 239885 402358 239897
rect 383938 239857 402358 239885
rect 402352 239845 402358 239857
rect 402410 239845 402416 239897
rect 380560 239771 380566 239823
rect 380618 239811 380624 239823
rect 384880 239811 384886 239823
rect 380618 239783 384886 239811
rect 380618 239771 380624 239783
rect 384880 239771 384886 239783
rect 384938 239771 384944 239823
rect 383248 239697 383254 239749
rect 383306 239737 383312 239749
rect 384400 239737 384406 239749
rect 383306 239709 384406 239737
rect 383306 239697 383312 239709
rect 384400 239697 384406 239709
rect 384458 239697 384464 239749
rect 387280 239697 387286 239749
rect 387338 239737 387344 239749
rect 400624 239737 400630 239749
rect 387338 239709 400630 239737
rect 387338 239697 387344 239709
rect 400624 239697 400630 239709
rect 400682 239697 400688 239749
rect 374800 239623 374806 239675
rect 374858 239663 374864 239675
rect 382672 239663 382678 239675
rect 374858 239635 382678 239663
rect 374858 239623 374864 239635
rect 382672 239623 382678 239635
rect 382730 239623 382736 239675
rect 383632 239623 383638 239675
rect 383690 239663 383696 239675
rect 385552 239663 385558 239675
rect 383690 239635 385558 239663
rect 383690 239623 383696 239635
rect 385552 239623 385558 239635
rect 385610 239623 385616 239675
rect 380080 239549 380086 239601
rect 380138 239589 380144 239601
rect 383728 239589 383734 239601
rect 380138 239561 383734 239589
rect 380138 239549 380144 239561
rect 383728 239549 383734 239561
rect 383786 239549 383792 239601
rect 380848 239475 380854 239527
rect 380906 239515 380912 239527
rect 388144 239515 388150 239527
rect 380906 239487 388150 239515
rect 380906 239475 380912 239487
rect 388144 239475 388150 239487
rect 388202 239475 388208 239527
rect 375184 239401 375190 239453
rect 375242 239441 375248 239453
rect 387280 239441 387286 239453
rect 375242 239413 387286 239441
rect 375242 239401 375248 239413
rect 387280 239401 387286 239413
rect 387338 239401 387344 239453
rect 392080 239367 392086 239379
rect 368722 239339 392086 239367
rect 392080 239327 392086 239339
rect 392138 239327 392144 239379
rect 224080 239253 224086 239305
rect 224138 239293 224144 239305
rect 231568 239293 231574 239305
rect 224138 239265 231574 239293
rect 224138 239253 224144 239265
rect 231568 239253 231574 239265
rect 231626 239253 231632 239305
rect 276208 239253 276214 239305
rect 276266 239293 276272 239305
rect 286000 239293 286006 239305
rect 276266 239265 286006 239293
rect 276266 239253 276272 239265
rect 286000 239253 286006 239265
rect 286058 239253 286064 239305
rect 290416 239293 290422 239305
rect 286114 239265 290422 239293
rect 235504 239179 235510 239231
rect 235562 239219 235568 239231
rect 238960 239219 238966 239231
rect 235562 239191 238966 239219
rect 235562 239179 235568 239191
rect 238960 239179 238966 239191
rect 239018 239179 239024 239231
rect 271792 239179 271798 239231
rect 271850 239219 271856 239231
rect 286114 239219 286142 239265
rect 290416 239253 290422 239265
rect 290474 239253 290480 239305
rect 290512 239253 290518 239305
rect 290570 239293 290576 239305
rect 316048 239293 316054 239305
rect 290570 239265 316054 239293
rect 290570 239253 290576 239265
rect 316048 239253 316054 239265
rect 316106 239253 316112 239305
rect 317968 239253 317974 239305
rect 318026 239293 318032 239305
rect 332752 239293 332758 239305
rect 318026 239265 332758 239293
rect 318026 239253 318032 239265
rect 332752 239253 332758 239265
rect 332810 239253 332816 239305
rect 360592 239253 360598 239305
rect 360650 239293 360656 239305
rect 394096 239293 394102 239305
rect 360650 239265 394102 239293
rect 360650 239253 360656 239265
rect 394096 239253 394102 239265
rect 394154 239253 394160 239305
rect 271850 239191 286142 239219
rect 271850 239179 271856 239191
rect 287344 239179 287350 239231
rect 287402 239219 287408 239231
rect 287402 239191 291422 239219
rect 287402 239179 287408 239191
rect 237136 239105 237142 239157
rect 237194 239145 237200 239157
rect 241648 239145 241654 239157
rect 237194 239117 241654 239145
rect 237194 239105 237200 239117
rect 241648 239105 241654 239117
rect 241706 239105 241712 239157
rect 244624 239105 244630 239157
rect 244682 239145 244688 239157
rect 246256 239145 246262 239157
rect 244682 239117 246262 239145
rect 244682 239105 244688 239117
rect 246256 239105 246262 239117
rect 246314 239105 246320 239157
rect 272656 239105 272662 239157
rect 272714 239145 272720 239157
rect 291088 239145 291094 239157
rect 272714 239117 291094 239145
rect 272714 239105 272720 239117
rect 291088 239105 291094 239117
rect 291146 239105 291152 239157
rect 291394 239145 291422 239191
rect 291472 239179 291478 239231
rect 291530 239219 291536 239231
rect 301840 239219 301846 239231
rect 291530 239191 301846 239219
rect 291530 239179 291536 239191
rect 301840 239179 301846 239191
rect 301898 239179 301904 239231
rect 302512 239179 302518 239231
rect 302570 239219 302576 239231
rect 307216 239219 307222 239231
rect 302570 239191 307222 239219
rect 302570 239179 302576 239191
rect 307216 239179 307222 239191
rect 307274 239179 307280 239231
rect 326608 239179 326614 239231
rect 326666 239219 326672 239231
rect 348592 239219 348598 239231
rect 326666 239191 348598 239219
rect 326666 239179 326672 239191
rect 348592 239179 348598 239191
rect 348650 239179 348656 239231
rect 380080 239179 380086 239231
rect 380138 239219 380144 239231
rect 386608 239219 386614 239231
rect 380138 239191 386614 239219
rect 380138 239179 380144 239191
rect 386608 239179 386614 239191
rect 386666 239179 386672 239231
rect 596176 239179 596182 239231
rect 596234 239219 596240 239231
rect 603088 239219 603094 239231
rect 596234 239191 603094 239219
rect 596234 239179 596240 239191
rect 603088 239179 603094 239191
rect 603146 239179 603152 239231
rect 300016 239145 300022 239157
rect 291394 239117 300022 239145
rect 300016 239105 300022 239117
rect 300074 239105 300080 239157
rect 318064 239105 318070 239157
rect 318122 239145 318128 239157
rect 334576 239145 334582 239157
rect 318122 239117 334582 239145
rect 318122 239105 318128 239117
rect 334576 239105 334582 239117
rect 334634 239105 334640 239157
rect 373360 239105 373366 239157
rect 373418 239145 373424 239157
rect 396880 239145 396886 239157
rect 373418 239117 396886 239145
rect 373418 239105 373424 239117
rect 396880 239105 396886 239117
rect 396938 239105 396944 239157
rect 146608 239031 146614 239083
rect 146666 239071 146672 239083
rect 174160 239071 174166 239083
rect 146666 239043 174166 239071
rect 146666 239031 146672 239043
rect 174160 239031 174166 239043
rect 174218 239031 174224 239083
rect 236176 239031 236182 239083
rect 236234 239071 236240 239083
rect 238192 239071 238198 239083
rect 236234 239043 238198 239071
rect 236234 239031 236240 239043
rect 238192 239031 238198 239043
rect 238250 239031 238256 239083
rect 238480 239031 238486 239083
rect 238538 239071 238544 239083
rect 241840 239071 241846 239083
rect 238538 239043 241846 239071
rect 238538 239031 238544 239043
rect 241840 239031 241846 239043
rect 241898 239031 241904 239083
rect 278338 239043 280862 239071
rect 228496 238957 228502 239009
rect 228554 238997 228560 239009
rect 230800 238997 230806 239009
rect 228554 238969 230806 238997
rect 228554 238957 228560 238969
rect 230800 238957 230806 238969
rect 230858 238957 230864 239009
rect 240496 238957 240502 239009
rect 240554 238997 240560 239009
rect 255664 238997 255670 239009
rect 240554 238969 255670 238997
rect 240554 238957 240560 238969
rect 255664 238957 255670 238969
rect 255722 238957 255728 239009
rect 260368 238957 260374 239009
rect 260426 238997 260432 239009
rect 278338 238997 278366 239043
rect 260426 238969 278366 238997
rect 260426 238957 260432 238969
rect 228112 238883 228118 238935
rect 228170 238923 228176 238935
rect 231952 238923 231958 238935
rect 228170 238895 231958 238923
rect 228170 238883 228176 238895
rect 231952 238883 231958 238895
rect 232010 238883 232016 238935
rect 239536 238883 239542 238935
rect 239594 238923 239600 238935
rect 257392 238923 257398 238935
rect 239594 238895 257398 238923
rect 239594 238883 239600 238895
rect 257392 238883 257398 238895
rect 257450 238883 257456 238935
rect 259984 238883 259990 238935
rect 260042 238923 260048 238935
rect 277840 238923 277846 238935
rect 260042 238895 277846 238923
rect 260042 238883 260048 238895
rect 277840 238883 277846 238895
rect 277898 238883 277904 238935
rect 278512 238883 278518 238935
rect 278570 238923 278576 238935
rect 280720 238923 280726 238935
rect 278570 238895 280726 238923
rect 278570 238883 278576 238895
rect 280720 238883 280726 238895
rect 280778 238883 280784 238935
rect 280834 238923 280862 239043
rect 283408 239031 283414 239083
rect 283466 239071 283472 239083
rect 298384 239071 298390 239083
rect 283466 239043 298390 239071
rect 283466 239031 283472 239043
rect 298384 239031 298390 239043
rect 298442 239031 298448 239083
rect 318352 239031 318358 239083
rect 318410 239071 318416 239083
rect 336496 239071 336502 239083
rect 318410 239043 336502 239071
rect 318410 239031 318416 239043
rect 336496 239031 336502 239043
rect 336554 239031 336560 239083
rect 373840 239031 373846 239083
rect 373898 239071 373904 239083
rect 384016 239071 384022 239083
rect 373898 239043 384022 239071
rect 373898 239031 373904 239043
rect 384016 239031 384022 239043
rect 384074 239031 384080 239083
rect 280912 238957 280918 239009
rect 280970 238997 280976 239009
rect 293968 238997 293974 239009
rect 280970 238969 293974 238997
rect 280970 238957 280976 238969
rect 293968 238957 293974 238969
rect 294026 238957 294032 239009
rect 294064 238957 294070 239009
rect 294122 238997 294128 239009
rect 303184 238997 303190 239009
rect 294122 238969 303190 238997
rect 294122 238957 294128 238969
rect 303184 238957 303190 238969
rect 303242 238957 303248 239009
rect 304720 238957 304726 239009
rect 304778 238997 304784 239009
rect 308176 238997 308182 239009
rect 304778 238969 308182 238997
rect 304778 238957 304784 238969
rect 308176 238957 308182 238969
rect 308234 238957 308240 239009
rect 311632 238957 311638 239009
rect 311690 238997 311696 239009
rect 323632 238997 323638 239009
rect 311690 238969 323638 238997
rect 311690 238957 311696 238969
rect 323632 238957 323638 238969
rect 323690 238957 323696 239009
rect 323728 238957 323734 239009
rect 323786 238997 323792 239009
rect 376624 238997 376630 239009
rect 323786 238969 376630 238997
rect 323786 238957 323792 238969
rect 376624 238957 376630 238969
rect 376682 238957 376688 239009
rect 380464 238957 380470 239009
rect 380522 238997 380528 239009
rect 387568 238997 387574 239009
rect 380522 238969 387574 238997
rect 380522 238957 380528 238969
rect 387568 238957 387574 238969
rect 387626 238957 387632 239009
rect 282256 238923 282262 238935
rect 280834 238895 282262 238923
rect 282256 238883 282262 238895
rect 282314 238883 282320 238935
rect 284368 238883 284374 238935
rect 284426 238923 284432 238935
rect 288304 238923 288310 238935
rect 284426 238895 288310 238923
rect 284426 238883 284432 238895
rect 288304 238883 288310 238895
rect 288362 238883 288368 238935
rect 288400 238883 288406 238935
rect 288458 238923 288464 238935
rect 300592 238923 300598 238935
rect 288458 238895 300598 238923
rect 288458 238883 288464 238895
rect 300592 238883 300598 238895
rect 300650 238883 300656 238935
rect 300784 238883 300790 238935
rect 300842 238923 300848 238935
rect 306256 238923 306262 238935
rect 300842 238895 306262 238923
rect 300842 238883 300848 238895
rect 306256 238883 306262 238895
rect 306314 238883 306320 238935
rect 316432 238883 316438 238935
rect 316490 238923 316496 238935
rect 377296 238923 377302 238935
rect 316490 238895 377302 238923
rect 316490 238883 316496 238895
rect 377296 238883 377302 238895
rect 377354 238883 377360 238935
rect 381424 238883 381430 238935
rect 381482 238923 381488 238935
rect 389200 238923 389206 238935
rect 381482 238895 389206 238923
rect 381482 238883 381488 238895
rect 389200 238883 389206 238895
rect 389258 238883 389264 238935
rect 240112 238809 240118 238861
rect 240170 238849 240176 238861
rect 256816 238849 256822 238861
rect 240170 238821 256822 238849
rect 240170 238809 240176 238821
rect 256816 238809 256822 238821
rect 256874 238809 256880 238861
rect 257104 238809 257110 238861
rect 257162 238849 257168 238861
rect 318352 238849 318358 238861
rect 257162 238821 318358 238849
rect 257162 238809 257168 238821
rect 318352 238809 318358 238821
rect 318410 238809 318416 238861
rect 318640 238809 318646 238861
rect 318698 238849 318704 238861
rect 332176 238849 332182 238861
rect 318698 238821 332182 238849
rect 318698 238809 318704 238821
rect 332176 238809 332182 238821
rect 332234 238809 332240 238861
rect 332464 238809 332470 238861
rect 332522 238849 332528 238861
rect 347440 238849 347446 238861
rect 332522 238821 347446 238849
rect 332522 238809 332528 238821
rect 347440 238809 347446 238821
rect 347498 238809 347504 238861
rect 351376 238809 351382 238861
rect 351434 238849 351440 238861
rect 358864 238849 358870 238861
rect 351434 238821 358870 238849
rect 351434 238809 351440 238821
rect 358864 238809 358870 238821
rect 358922 238809 358928 238861
rect 368176 238809 368182 238861
rect 368234 238849 368240 238861
rect 384592 238849 384598 238861
rect 368234 238821 384598 238849
rect 368234 238809 368240 238821
rect 384592 238809 384598 238821
rect 384650 238809 384656 238861
rect 227248 238735 227254 238787
rect 227306 238775 227312 238787
rect 234064 238775 234070 238787
rect 227306 238747 234070 238775
rect 227306 238735 227312 238747
rect 234064 238735 234070 238747
rect 234122 238735 234128 238787
rect 257776 238735 257782 238787
rect 257834 238775 257840 238787
rect 318160 238775 318166 238787
rect 257834 238747 318166 238775
rect 257834 238735 257840 238747
rect 318160 238735 318166 238747
rect 318218 238735 318224 238787
rect 323728 238775 323734 238787
rect 318370 238747 323734 238775
rect 226288 238661 226294 238713
rect 226346 238701 226352 238713
rect 235600 238701 235606 238713
rect 226346 238673 235606 238701
rect 226346 238661 226352 238673
rect 235600 238661 235606 238673
rect 235658 238661 235664 238713
rect 256240 238661 256246 238713
rect 256298 238701 256304 238713
rect 318256 238701 318262 238713
rect 256298 238673 318262 238701
rect 256298 238661 256304 238673
rect 318256 238661 318262 238673
rect 318314 238661 318320 238713
rect 248944 238587 248950 238639
rect 249002 238627 249008 238639
rect 315952 238627 315958 238639
rect 249002 238599 315958 238627
rect 249002 238587 249008 238599
rect 315952 238587 315958 238599
rect 316010 238587 316016 238639
rect 316048 238587 316054 238639
rect 316106 238627 316112 238639
rect 318370 238627 318398 238747
rect 323728 238735 323734 238747
rect 323786 238735 323792 238787
rect 331216 238735 331222 238787
rect 331274 238775 331280 238787
rect 358768 238775 358774 238787
rect 331274 238747 358774 238775
rect 331274 238735 331280 238747
rect 358768 238735 358774 238747
rect 358826 238735 358832 238787
rect 368656 238735 368662 238787
rect 368714 238775 368720 238787
rect 381040 238775 381046 238787
rect 368714 238747 381046 238775
rect 368714 238735 368720 238747
rect 381040 238735 381046 238747
rect 381098 238735 381104 238787
rect 319024 238661 319030 238713
rect 319082 238701 319088 238713
rect 332368 238701 332374 238713
rect 319082 238673 332374 238701
rect 319082 238661 319088 238673
rect 332368 238661 332374 238673
rect 332426 238661 332432 238713
rect 334096 238661 334102 238713
rect 334154 238701 334160 238713
rect 365296 238701 365302 238713
rect 334154 238673 365302 238701
rect 334154 238661 334160 238673
rect 365296 238661 365302 238673
rect 365354 238661 365360 238713
rect 383344 238701 383350 238713
rect 368722 238673 383350 238701
rect 316106 238599 318398 238627
rect 316106 238587 316112 238599
rect 319600 238587 319606 238639
rect 319658 238627 319664 238639
rect 333424 238627 333430 238639
rect 319658 238599 333430 238627
rect 319658 238587 319664 238599
rect 333424 238587 333430 238599
rect 333482 238587 333488 238639
rect 333616 238587 333622 238639
rect 333674 238627 333680 238639
rect 363280 238627 363286 238639
rect 333674 238599 363286 238627
rect 333674 238587 333680 238599
rect 363280 238587 363286 238599
rect 363338 238587 363344 238639
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 43024 238553 43030 238565
rect 42218 238525 43030 238553
rect 42218 238513 42224 238525
rect 43024 238513 43030 238525
rect 43082 238513 43088 238565
rect 227728 238513 227734 238565
rect 227786 238553 227792 238565
rect 232816 238553 232822 238565
rect 227786 238525 232822 238553
rect 227786 238513 227792 238525
rect 232816 238513 232822 238525
rect 232874 238513 232880 238565
rect 255568 238513 255574 238565
rect 255626 238553 255632 238565
rect 318064 238553 318070 238565
rect 255626 238525 318070 238553
rect 255626 238513 255632 238525
rect 318064 238513 318070 238525
rect 318122 238513 318128 238565
rect 318352 238513 318358 238565
rect 318410 238553 318416 238565
rect 324112 238553 324118 238565
rect 318410 238525 324118 238553
rect 318410 238513 318416 238525
rect 324112 238513 324118 238525
rect 324170 238513 324176 238565
rect 329776 238513 329782 238565
rect 329834 238553 329840 238565
rect 332464 238553 332470 238565
rect 329834 238525 332470 238553
rect 329834 238513 329840 238525
rect 332464 238513 332470 238525
rect 332522 238513 332528 238565
rect 334864 238513 334870 238565
rect 334922 238553 334928 238565
rect 367024 238553 367030 238565
rect 334922 238525 367030 238553
rect 334922 238513 334928 238525
rect 367024 238513 367030 238525
rect 367082 238513 367088 238565
rect 254608 238439 254614 238491
rect 254666 238479 254672 238491
rect 254666 238451 332798 238479
rect 254666 238439 254672 238451
rect 42448 238365 42454 238417
rect 42506 238405 42512 238417
rect 43024 238405 43030 238417
rect 42506 238377 43030 238405
rect 42506 238365 42512 238377
rect 43024 238365 43030 238377
rect 43082 238365 43088 238417
rect 221104 238365 221110 238417
rect 221162 238405 221168 238417
rect 246544 238405 246550 238417
rect 221162 238377 246550 238405
rect 221162 238365 221168 238377
rect 246544 238365 246550 238377
rect 246602 238365 246608 238417
rect 254128 238365 254134 238417
rect 254186 238405 254192 238417
rect 332770 238405 332798 238451
rect 332848 238439 332854 238491
rect 332906 238479 332912 238491
rect 362224 238479 362230 238491
rect 332906 238451 362230 238479
rect 332906 238439 332912 238451
rect 362224 238439 362230 238451
rect 362282 238439 362288 238491
rect 366832 238439 366838 238491
rect 366890 238479 366896 238491
rect 368722 238479 368750 238673
rect 383344 238661 383350 238673
rect 383402 238661 383408 238713
rect 370480 238587 370486 238639
rect 370538 238627 370544 238639
rect 382288 238627 382294 238639
rect 370538 238599 382294 238627
rect 370538 238587 370544 238599
rect 382288 238587 382294 238599
rect 382346 238587 382352 238639
rect 370000 238513 370006 238565
rect 370058 238553 370064 238565
rect 380944 238553 380950 238565
rect 370058 238525 380950 238553
rect 370058 238513 370064 238525
rect 380944 238513 380950 238525
rect 381002 238513 381008 238565
rect 381040 238513 381046 238565
rect 381098 238553 381104 238565
rect 385936 238553 385942 238565
rect 381098 238525 385942 238553
rect 381098 238513 381104 238525
rect 385936 238513 385942 238525
rect 385994 238513 386000 238565
rect 366890 238451 368750 238479
rect 366890 238439 366896 238451
rect 369424 238439 369430 238491
rect 369482 238479 369488 238491
rect 388816 238479 388822 238491
rect 369482 238451 388822 238479
rect 369482 238439 369488 238451
rect 388816 238439 388822 238451
rect 388874 238439 388880 238491
rect 336976 238405 336982 238417
rect 254186 238377 332654 238405
rect 332770 238377 336982 238405
rect 254186 238365 254192 238377
rect 218032 238291 218038 238343
rect 218090 238331 218096 238343
rect 253456 238331 253462 238343
rect 218090 238303 253462 238331
rect 218090 238291 218096 238303
rect 253456 238291 253462 238303
rect 253514 238291 253520 238343
rect 258544 238291 258550 238343
rect 258602 238331 258608 238343
rect 280912 238331 280918 238343
rect 258602 238303 280918 238331
rect 258602 238291 258608 238303
rect 280912 238291 280918 238303
rect 280970 238291 280976 238343
rect 283312 238291 283318 238343
rect 283370 238331 283376 238343
rect 284848 238331 284854 238343
rect 283370 238303 284854 238331
rect 283370 238291 283376 238303
rect 284848 238291 284854 238303
rect 284906 238291 284912 238343
rect 285808 238291 285814 238343
rect 285866 238331 285872 238343
rect 298960 238331 298966 238343
rect 285866 238303 298966 238331
rect 285866 238291 285872 238303
rect 298960 238291 298966 238303
rect 299018 238291 299024 238343
rect 299056 238291 299062 238343
rect 299114 238331 299120 238343
rect 305776 238331 305782 238343
rect 299114 238303 305782 238331
rect 299114 238291 299120 238303
rect 305776 238291 305782 238303
rect 305834 238291 305840 238343
rect 305872 238291 305878 238343
rect 305930 238331 305936 238343
rect 332464 238331 332470 238343
rect 305930 238303 332470 238331
rect 305930 238291 305936 238303
rect 332464 238291 332470 238303
rect 332522 238291 332528 238343
rect 221872 238217 221878 238269
rect 221930 238257 221936 238269
rect 244816 238257 244822 238269
rect 221930 238229 244822 238257
rect 221930 238217 221936 238229
rect 244816 238217 244822 238229
rect 244874 238217 244880 238269
rect 252400 238217 252406 238269
rect 252458 238257 252464 238269
rect 332626 238257 332654 238377
rect 336976 238365 336982 238377
rect 337034 238365 337040 238417
rect 369808 238365 369814 238417
rect 369866 238405 369872 238417
rect 389680 238405 389686 238417
rect 369866 238377 389686 238405
rect 369866 238365 369872 238377
rect 389680 238365 389686 238377
rect 389738 238365 389744 238417
rect 332752 238291 332758 238343
rect 332810 238331 332816 238343
rect 385264 238331 385270 238343
rect 332810 238303 385270 238331
rect 332810 238291 332816 238303
rect 385264 238291 385270 238303
rect 385322 238291 385328 238343
rect 338704 238257 338710 238269
rect 252458 238229 332510 238257
rect 332626 238229 338710 238257
rect 252458 238217 252464 238229
rect 222832 238143 222838 238195
rect 222890 238183 222896 238195
rect 243760 238183 243766 238195
rect 222890 238155 243766 238183
rect 222890 238143 222896 238155
rect 243760 238143 243766 238155
rect 243818 238143 243824 238195
rect 253360 238143 253366 238195
rect 253418 238183 253424 238195
rect 332080 238183 332086 238195
rect 253418 238155 332086 238183
rect 253418 238143 253424 238155
rect 332080 238143 332086 238155
rect 332138 238143 332144 238195
rect 223216 238069 223222 238121
rect 223274 238109 223280 238121
rect 242608 238109 242614 238121
rect 223274 238081 242614 238109
rect 223274 238069 223280 238081
rect 242608 238069 242614 238081
rect 242666 238069 242672 238121
rect 251152 238069 251158 238121
rect 251210 238109 251216 238121
rect 332482 238109 332510 238229
rect 338704 238217 338710 238229
rect 338762 238217 338768 238269
rect 370384 238217 370390 238269
rect 370442 238257 370448 238269
rect 390352 238257 390358 238269
rect 370442 238229 390358 238257
rect 370442 238217 370448 238229
rect 390352 238217 390358 238229
rect 390410 238217 390416 238269
rect 332560 238143 332566 238195
rect 332618 238183 332624 238195
rect 340432 238183 340438 238195
rect 332618 238155 340438 238183
rect 332618 238143 332624 238155
rect 340432 238143 340438 238155
rect 340490 238143 340496 238195
rect 372016 238143 372022 238195
rect 372074 238183 372080 238195
rect 394192 238183 394198 238195
rect 372074 238155 394198 238183
rect 372074 238143 372080 238155
rect 394192 238143 394198 238155
rect 394250 238143 394256 238195
rect 341488 238109 341494 238121
rect 251210 238081 332414 238109
rect 332482 238081 341494 238109
rect 251210 238069 251216 238081
rect 251920 237995 251926 238047
rect 251978 238035 251984 238047
rect 332386 238035 332414 238081
rect 341488 238069 341494 238081
rect 341546 238069 341552 238121
rect 371632 238069 371638 238121
rect 371690 238109 371696 238121
rect 393616 238109 393622 238121
rect 371690 238081 393622 238109
rect 371690 238069 371696 238081
rect 393616 238069 393622 238081
rect 393674 238069 393680 238121
rect 251978 238007 329918 238035
rect 332386 238007 332606 238035
rect 251978 237995 251984 238007
rect 42928 237921 42934 237973
rect 42986 237961 42992 237973
rect 43312 237961 43318 237973
rect 42986 237933 43318 237961
rect 42986 237921 42992 237933
rect 43312 237921 43318 237933
rect 43370 237921 43376 237973
rect 181456 237921 181462 237973
rect 181514 237961 181520 237973
rect 201520 237961 201526 237973
rect 181514 237933 201526 237961
rect 181514 237921 181520 237933
rect 201520 237921 201526 237933
rect 201578 237921 201584 237973
rect 223312 237921 223318 237973
rect 223370 237961 223376 237973
rect 242128 237961 242134 237973
rect 223370 237933 242134 237961
rect 223370 237921 223376 237933
rect 242128 237921 242134 237933
rect 242186 237921 242192 237973
rect 249808 237921 249814 237973
rect 249866 237961 249872 237973
rect 329776 237961 329782 237973
rect 249866 237933 329782 237961
rect 249866 237921 249872 237933
rect 329776 237921 329782 237933
rect 329834 237921 329840 237973
rect 329890 237961 329918 238007
rect 332272 237961 332278 237973
rect 329890 237933 332278 237961
rect 332272 237921 332278 237933
rect 332330 237921 332336 237973
rect 332578 237961 332606 238007
rect 332656 237995 332662 238047
rect 332714 238035 332720 238047
rect 343504 238035 343510 238047
rect 332714 238007 343510 238035
rect 332714 237995 332720 238007
rect 343504 237995 343510 238007
rect 343562 237995 343568 238047
rect 371248 237995 371254 238047
rect 371306 238035 371312 238047
rect 392464 238035 392470 238047
rect 371306 238007 392470 238035
rect 371306 237995 371312 238007
rect 392464 237995 392470 238007
rect 392522 237995 392528 238047
rect 345232 237961 345238 237973
rect 332578 237933 345238 237961
rect 345232 237921 345238 237933
rect 345290 237921 345296 237973
rect 371152 237921 371158 237973
rect 371210 237961 371216 237973
rect 391888 237961 391894 237973
rect 371210 237933 391894 237961
rect 371210 237921 371216 237933
rect 391888 237921 391894 237933
rect 391946 237921 391952 237973
rect 42160 237847 42166 237899
rect 42218 237887 42224 237899
rect 47536 237887 47542 237899
rect 42218 237859 47542 237887
rect 42218 237847 42224 237859
rect 47536 237847 47542 237859
rect 47594 237847 47600 237899
rect 224080 237847 224086 237899
rect 224138 237887 224144 237899
rect 240592 237887 240598 237899
rect 224138 237859 240598 237887
rect 224138 237847 224144 237859
rect 240592 237847 240598 237859
rect 240650 237847 240656 237899
rect 249328 237847 249334 237899
rect 249386 237887 249392 237899
rect 349168 237887 349174 237899
rect 249386 237859 349174 237887
rect 249386 237847 249392 237859
rect 349168 237847 349174 237859
rect 349226 237847 349232 237899
rect 362800 237847 362806 237899
rect 362858 237887 362864 237899
rect 370480 237887 370486 237899
rect 362858 237859 370486 237887
rect 362858 237847 362864 237859
rect 370480 237847 370486 237859
rect 370538 237847 370544 237899
rect 370576 237847 370582 237899
rect 370634 237887 370640 237899
rect 379024 237887 379030 237899
rect 370634 237859 379030 237887
rect 370634 237847 370640 237859
rect 379024 237847 379030 237859
rect 379082 237847 379088 237899
rect 384400 237847 384406 237899
rect 384458 237887 384464 237899
rect 410416 237887 410422 237899
rect 384458 237859 410422 237887
rect 384458 237847 384464 237859
rect 410416 237847 410422 237859
rect 410474 237847 410480 237899
rect 43312 237773 43318 237825
rect 43370 237813 43376 237825
rect 43504 237813 43510 237825
rect 43370 237785 43510 237813
rect 43370 237773 43376 237785
rect 43504 237773 43510 237785
rect 43562 237773 43568 237825
rect 171280 237773 171286 237825
rect 171338 237813 171344 237825
rect 181456 237813 181462 237825
rect 171338 237785 181462 237813
rect 171338 237773 171344 237785
rect 181456 237773 181462 237785
rect 181514 237773 181520 237825
rect 201520 237773 201526 237825
rect 201578 237813 201584 237825
rect 207088 237813 207094 237825
rect 201578 237785 207094 237813
rect 201578 237773 201584 237785
rect 207088 237773 207094 237785
rect 207146 237813 207152 237825
rect 221968 237813 221974 237825
rect 207146 237785 221974 237813
rect 207146 237773 207152 237785
rect 221968 237773 221974 237785
rect 222026 237773 222032 237825
rect 225040 237773 225046 237825
rect 225098 237813 225104 237825
rect 238864 237813 238870 237825
rect 225098 237785 238870 237813
rect 225098 237773 225104 237785
rect 238864 237773 238870 237785
rect 238922 237773 238928 237825
rect 247120 237773 247126 237825
rect 247178 237813 247184 237825
rect 353968 237813 353974 237825
rect 247178 237785 353974 237813
rect 247178 237773 247184 237785
rect 353968 237773 353974 237785
rect 354026 237773 354032 237825
rect 375568 237773 375574 237825
rect 375626 237813 375632 237825
rect 401200 237813 401206 237825
rect 375626 237785 401206 237813
rect 375626 237773 375632 237785
rect 401200 237773 401206 237785
rect 401258 237773 401264 237825
rect 221008 237699 221014 237751
rect 221066 237739 221072 237751
rect 246928 237739 246934 237751
rect 221066 237711 246934 237739
rect 221066 237699 221072 237711
rect 246928 237699 246934 237711
rect 246986 237699 246992 237751
rect 247600 237699 247606 237751
rect 247658 237739 247664 237751
rect 351952 237739 351958 237751
rect 247658 237711 351958 237739
rect 247658 237699 247664 237711
rect 351952 237699 351958 237711
rect 352010 237699 352016 237751
rect 359824 237699 359830 237751
rect 359882 237739 359888 237751
rect 370000 237739 370006 237751
rect 359882 237711 370006 237739
rect 359882 237699 359888 237711
rect 370000 237699 370006 237711
rect 370058 237699 370064 237751
rect 370768 237699 370774 237751
rect 370826 237739 370832 237751
rect 381136 237739 381142 237751
rect 370826 237711 381142 237739
rect 370826 237699 370832 237711
rect 381136 237699 381142 237711
rect 381194 237699 381200 237751
rect 384496 237699 384502 237751
rect 384554 237739 384560 237751
rect 410992 237739 410998 237751
rect 384554 237711 410998 237739
rect 384554 237699 384560 237711
rect 410992 237699 410998 237711
rect 411050 237699 411056 237751
rect 549232 237699 549238 237751
rect 549290 237739 549296 237751
rect 649360 237739 649366 237751
rect 549290 237711 649366 237739
rect 549290 237699 549296 237711
rect 649360 237699 649366 237711
rect 649418 237699 649424 237751
rect 245776 237625 245782 237677
rect 245834 237665 245840 237677
rect 356176 237665 356182 237677
rect 245834 237637 356182 237665
rect 245834 237625 245840 237637
rect 356176 237625 356182 237637
rect 356234 237625 356240 237677
rect 373456 237625 373462 237677
rect 373514 237665 373520 237677
rect 397936 237665 397942 237677
rect 373514 237637 397942 237665
rect 373514 237625 373520 237637
rect 397936 237625 397942 237637
rect 397994 237625 398000 237677
rect 497488 237625 497494 237677
rect 497546 237665 497552 237677
rect 596176 237665 596182 237677
rect 497546 237637 596182 237665
rect 497546 237625 497552 237637
rect 596176 237625 596182 237637
rect 596234 237625 596240 237677
rect 148336 237551 148342 237603
rect 148394 237591 148400 237603
rect 161296 237591 161302 237603
rect 148394 237563 161302 237591
rect 148394 237551 148400 237563
rect 161296 237551 161302 237563
rect 161354 237551 161360 237603
rect 246160 237551 246166 237603
rect 246218 237591 246224 237603
rect 355024 237591 355030 237603
rect 246218 237563 355030 237591
rect 246218 237551 246224 237563
rect 355024 237551 355030 237563
rect 355082 237551 355088 237603
rect 355120 237551 355126 237603
rect 355178 237591 355184 237603
rect 370576 237591 370582 237603
rect 355178 237563 370582 237591
rect 355178 237551 355184 237563
rect 370576 237551 370582 237563
rect 370634 237551 370640 237603
rect 374224 237551 374230 237603
rect 374282 237591 374288 237603
rect 399664 237591 399670 237603
rect 374282 237563 399670 237591
rect 374282 237551 374288 237563
rect 399664 237551 399670 237563
rect 399722 237551 399728 237603
rect 420592 237551 420598 237603
rect 420650 237591 420656 237603
rect 607600 237591 607606 237603
rect 420650 237563 607606 237591
rect 420650 237551 420656 237563
rect 607600 237551 607606 237563
rect 607658 237551 607664 237603
rect 275344 237477 275350 237529
rect 275402 237517 275408 237529
rect 281104 237517 281110 237529
rect 275402 237489 281110 237517
rect 275402 237477 275408 237489
rect 281104 237477 281110 237489
rect 281162 237477 281168 237529
rect 288112 237477 288118 237529
rect 288170 237517 288176 237529
rect 292336 237517 292342 237529
rect 288170 237489 292342 237517
rect 288170 237477 288176 237489
rect 292336 237477 292342 237489
rect 292394 237477 292400 237529
rect 293776 237477 293782 237529
rect 293834 237517 293840 237529
rect 305872 237517 305878 237529
rect 293834 237489 305878 237517
rect 293834 237477 293840 237489
rect 305872 237477 305878 237489
rect 305930 237477 305936 237529
rect 305968 237477 305974 237529
rect 306026 237517 306032 237529
rect 317584 237517 317590 237529
rect 306026 237489 317590 237517
rect 306026 237477 306032 237489
rect 317584 237477 317590 237489
rect 317642 237477 317648 237529
rect 317680 237477 317686 237529
rect 317738 237517 317744 237529
rect 318448 237517 318454 237529
rect 317738 237489 318454 237517
rect 317738 237477 317744 237489
rect 318448 237477 318454 237489
rect 318506 237477 318512 237529
rect 318544 237477 318550 237529
rect 318602 237517 318608 237529
rect 319696 237517 319702 237529
rect 318602 237489 319702 237517
rect 318602 237477 318608 237489
rect 319696 237477 319702 237489
rect 319754 237477 319760 237529
rect 329776 237517 329782 237529
rect 319906 237489 329782 237517
rect 161296 237403 161302 237455
rect 161354 237443 161360 237455
rect 171280 237443 171286 237455
rect 161354 237415 171286 237443
rect 161354 237403 161360 237415
rect 171280 237403 171286 237415
rect 171338 237403 171344 237455
rect 227344 237403 227350 237455
rect 227402 237443 227408 237455
rect 233584 237443 233590 237455
rect 227402 237415 233590 237443
rect 227402 237403 227408 237415
rect 233584 237403 233590 237415
rect 233642 237403 233648 237455
rect 238768 237403 238774 237455
rect 238826 237443 238832 237455
rect 259408 237443 259414 237455
rect 238826 237415 259414 237443
rect 238826 237403 238832 237415
rect 259408 237403 259414 237415
rect 259466 237403 259472 237455
rect 275824 237403 275830 237455
rect 275882 237443 275888 237455
rect 286576 237443 286582 237455
rect 275882 237415 286582 237443
rect 275882 237403 275888 237415
rect 286576 237403 286582 237415
rect 286634 237403 286640 237455
rect 288016 237403 288022 237455
rect 288074 237443 288080 237455
rect 291952 237443 291958 237455
rect 288074 237415 291958 237443
rect 288074 237403 288080 237415
rect 291952 237403 291958 237415
rect 292010 237403 292016 237455
rect 294160 237403 294166 237455
rect 294218 237443 294224 237455
rect 302224 237443 302230 237455
rect 294218 237415 302230 237443
rect 294218 237403 294224 237415
rect 302224 237403 302230 237415
rect 302282 237403 302288 237455
rect 316816 237403 316822 237455
rect 316874 237443 316880 237455
rect 319906 237443 319934 237489
rect 329776 237477 329782 237489
rect 329834 237477 329840 237529
rect 331792 237477 331798 237529
rect 331850 237517 331856 237529
rect 337936 237517 337942 237529
rect 331850 237489 337942 237517
rect 331850 237477 331856 237489
rect 337936 237477 337942 237489
rect 337994 237477 338000 237529
rect 372592 237477 372598 237529
rect 372650 237517 372656 237529
rect 395344 237517 395350 237529
rect 372650 237489 395350 237517
rect 372650 237477 372656 237489
rect 395344 237477 395350 237489
rect 395402 237477 395408 237529
rect 316874 237415 319934 237443
rect 316874 237403 316880 237415
rect 319984 237403 319990 237455
rect 320042 237443 320048 237455
rect 331312 237443 331318 237455
rect 320042 237415 331318 237443
rect 320042 237403 320048 237415
rect 331312 237403 331318 237415
rect 331370 237403 331376 237455
rect 339760 237403 339766 237455
rect 339818 237443 339824 237455
rect 348400 237443 348406 237455
rect 339818 237415 348406 237443
rect 339818 237403 339824 237415
rect 348400 237403 348406 237415
rect 348458 237403 348464 237455
rect 348496 237403 348502 237455
rect 348554 237443 348560 237455
rect 348554 237415 368990 237443
rect 348554 237403 348560 237415
rect 221488 237329 221494 237381
rect 221546 237369 221552 237381
rect 245872 237369 245878 237381
rect 221546 237341 245878 237369
rect 221546 237329 221552 237341
rect 245872 237329 245878 237341
rect 245930 237329 245936 237381
rect 277840 237329 277846 237381
rect 277898 237369 277904 237381
rect 287920 237369 287926 237381
rect 277898 237341 287926 237369
rect 277898 237329 277904 237341
rect 287920 237329 287926 237341
rect 287978 237329 287984 237381
rect 289360 237329 289366 237381
rect 289418 237369 289424 237381
rect 300976 237369 300982 237381
rect 289418 237341 300982 237369
rect 289418 237329 289424 237341
rect 300976 237329 300982 237341
rect 301034 237329 301040 237381
rect 317392 237329 317398 237381
rect 317450 237369 317456 237381
rect 317450 237341 319934 237369
rect 317450 237329 317456 237341
rect 319906 237307 319934 237341
rect 338128 237329 338134 237381
rect 338186 237369 338192 237381
rect 338186 237341 348350 237369
rect 338186 237329 338192 237341
rect 217072 237255 217078 237307
rect 217130 237295 217136 237307
rect 255184 237295 255190 237307
rect 217130 237267 255190 237295
rect 217130 237255 217136 237267
rect 255184 237255 255190 237267
rect 255242 237255 255248 237307
rect 273232 237255 273238 237307
rect 273290 237295 273296 237307
rect 287824 237295 287830 237307
rect 273290 237267 287830 237295
rect 273290 237255 273296 237267
rect 287824 237255 287830 237267
rect 287882 237255 287888 237307
rect 290128 237255 290134 237307
rect 290186 237295 290192 237307
rect 301456 237295 301462 237307
rect 290186 237267 301462 237295
rect 290186 237255 290192 237267
rect 301456 237255 301462 237267
rect 301514 237255 301520 237307
rect 317776 237255 317782 237307
rect 317834 237295 317840 237307
rect 319504 237295 319510 237307
rect 317834 237267 319510 237295
rect 317834 237255 317840 237267
rect 319504 237255 319510 237267
rect 319562 237255 319568 237307
rect 319888 237255 319894 237307
rect 319946 237255 319952 237307
rect 321808 237255 321814 237307
rect 321866 237295 321872 237307
rect 331792 237295 331798 237307
rect 321866 237267 331798 237295
rect 321866 237255 321872 237267
rect 331792 237255 331798 237267
rect 331850 237255 331856 237307
rect 331888 237255 331894 237307
rect 331946 237295 331952 237307
rect 339472 237295 339478 237307
rect 331946 237267 339478 237295
rect 331946 237255 331952 237267
rect 339472 237255 339478 237267
rect 339530 237255 339536 237307
rect 348322 237295 348350 237341
rect 353584 237329 353590 237381
rect 353642 237369 353648 237381
rect 358768 237369 358774 237381
rect 353642 237341 358774 237369
rect 353642 237329 353648 237341
rect 358768 237329 358774 237341
rect 358826 237329 358832 237381
rect 355120 237295 355126 237307
rect 348322 237267 355126 237295
rect 355120 237255 355126 237267
rect 355178 237255 355184 237307
rect 368962 237295 368990 237415
rect 372976 237403 372982 237455
rect 373034 237443 373040 237455
rect 396208 237443 396214 237455
rect 373034 237415 396214 237443
rect 373034 237403 373040 237415
rect 396208 237403 396214 237415
rect 396266 237403 396272 237455
rect 369040 237329 369046 237381
rect 369098 237369 369104 237381
rect 387664 237369 387670 237381
rect 369098 237341 387670 237369
rect 369098 237329 369104 237341
rect 387664 237329 387670 237341
rect 387722 237329 387728 237381
rect 378352 237295 378358 237307
rect 368962 237267 378358 237295
rect 378352 237255 378358 237267
rect 378410 237255 378416 237307
rect 379984 237255 379990 237307
rect 380042 237295 380048 237307
rect 385360 237295 385366 237307
rect 380042 237267 385366 237295
rect 380042 237255 380048 237267
rect 385360 237255 385366 237267
rect 385418 237255 385424 237307
rect 274000 237181 274006 237233
rect 274058 237221 274064 237233
rect 290224 237221 290230 237233
rect 274058 237193 290230 237221
rect 274058 237181 274064 237193
rect 290224 237181 290230 237193
rect 290282 237181 290288 237233
rect 291664 237181 291670 237233
rect 291722 237221 291728 237233
rect 317680 237221 317686 237233
rect 291722 237193 317686 237221
rect 291722 237181 291728 237193
rect 317680 237181 317686 237193
rect 317738 237181 317744 237233
rect 318160 237181 318166 237233
rect 318218 237221 318224 237233
rect 330544 237221 330550 237233
rect 318218 237193 330550 237221
rect 318218 237181 318224 237193
rect 330544 237181 330550 237193
rect 330602 237181 330608 237233
rect 330640 237181 330646 237233
rect 330698 237221 330704 237233
rect 357232 237221 357238 237233
rect 330698 237193 357238 237221
rect 330698 237181 330704 237193
rect 357232 237181 357238 237193
rect 357290 237181 357296 237233
rect 288304 237107 288310 237159
rect 288362 237147 288368 237159
rect 290416 237147 290422 237159
rect 288362 237119 290422 237147
rect 288362 237107 288368 237119
rect 290416 237107 290422 237119
rect 290474 237107 290480 237159
rect 290608 237107 290614 237159
rect 290666 237147 290672 237159
rect 290666 237119 295262 237147
rect 290666 237107 290672 237119
rect 225904 237033 225910 237085
rect 225962 237073 225968 237085
rect 236752 237073 236758 237085
rect 225962 237045 236758 237073
rect 225962 237033 225968 237045
rect 236752 237033 236758 237045
rect 236810 237033 236816 237085
rect 278800 237033 278806 237085
rect 278858 237073 278864 237085
rect 295024 237073 295030 237085
rect 278858 237045 295030 237073
rect 278858 237033 278864 237045
rect 295024 237033 295030 237045
rect 295082 237033 295088 237085
rect 295234 237073 295262 237119
rect 318256 237107 318262 237159
rect 318314 237147 318320 237159
rect 328720 237147 328726 237159
rect 318314 237119 328726 237147
rect 318314 237107 318320 237119
rect 328720 237107 328726 237119
rect 328778 237107 328784 237159
rect 328816 237107 328822 237159
rect 328874 237147 328880 237159
rect 353488 237147 353494 237159
rect 328874 237119 353494 237147
rect 328874 237107 328880 237119
rect 353488 237107 353494 237119
rect 353546 237107 353552 237159
rect 296944 237073 296950 237085
rect 295234 237045 296950 237073
rect 296944 237033 296950 237045
rect 297002 237033 297008 237085
rect 315952 237033 315958 237085
rect 316010 237073 316016 237085
rect 325840 237073 325846 237085
rect 316010 237045 325846 237073
rect 316010 237033 316016 237045
rect 325840 237033 325846 237045
rect 325898 237033 325904 237085
rect 327472 237033 327478 237085
rect 327530 237073 327536 237085
rect 350704 237073 350710 237085
rect 327530 237045 350710 237073
rect 327530 237033 327536 237045
rect 350704 237033 350710 237045
rect 350762 237033 350768 237085
rect 224560 236959 224566 237011
rect 224618 236999 224624 237011
rect 239632 236999 239638 237011
rect 224618 236971 239638 236999
rect 224618 236959 224624 236971
rect 239632 236959 239638 236971
rect 239690 236959 239696 237011
rect 276784 236959 276790 237011
rect 276842 236999 276848 237011
rect 295120 236999 295126 237011
rect 276842 236971 295126 236999
rect 276842 236959 276848 236971
rect 295120 236959 295126 236971
rect 295178 236959 295184 237011
rect 295216 236959 295222 237011
rect 295274 236999 295280 237011
rect 303664 236999 303670 237011
rect 295274 236971 303670 236999
rect 295274 236959 295280 236971
rect 303664 236959 303670 236971
rect 303722 236959 303728 237011
rect 327088 236959 327094 237011
rect 327146 236999 327152 237011
rect 349744 236999 349750 237011
rect 327146 236971 349750 236999
rect 327146 236959 327152 236971
rect 349744 236959 349750 236971
rect 349802 236959 349808 237011
rect 223696 236885 223702 236937
rect 223754 236925 223760 236937
rect 241552 236925 241558 236937
rect 223754 236897 241558 236925
rect 223754 236885 223760 236897
rect 241552 236885 241558 236897
rect 241610 236885 241616 236937
rect 286384 236885 286390 236937
rect 286442 236925 286448 236937
rect 299632 236925 299638 236937
rect 286442 236897 299638 236925
rect 286442 236885 286448 236897
rect 299632 236885 299638 236897
rect 299690 236885 299696 236937
rect 327856 236885 327862 236937
rect 327914 236925 327920 236937
rect 351472 236925 351478 236937
rect 327914 236897 351478 236925
rect 327914 236885 327920 236897
rect 351472 236885 351478 236897
rect 351530 236885 351536 236937
rect 277264 236811 277270 236863
rect 277322 236851 277328 236863
rect 279760 236851 279766 236863
rect 277322 236823 279766 236851
rect 277322 236811 277328 236823
rect 279760 236811 279766 236823
rect 279818 236811 279824 236863
rect 288208 236811 288214 236863
rect 288266 236851 288272 236863
rect 289936 236851 289942 236863
rect 288266 236823 289942 236851
rect 288266 236811 288272 236823
rect 289936 236811 289942 236823
rect 289994 236811 290000 236863
rect 291760 236811 291766 236863
rect 291818 236851 291824 236863
rect 291818 236823 308030 236851
rect 291818 236811 291824 236823
rect 288610 236749 290174 236777
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 43120 236703 43126 236715
rect 42218 236675 43126 236703
rect 42218 236663 42224 236675
rect 43120 236663 43126 236675
rect 43178 236663 43184 236715
rect 226864 236663 226870 236715
rect 226922 236703 226928 236715
rect 235024 236703 235030 236715
rect 226922 236675 235030 236703
rect 226922 236663 226928 236675
rect 235024 236663 235030 236675
rect 235082 236663 235088 236715
rect 274096 236663 274102 236715
rect 274154 236703 274160 236715
rect 288208 236703 288214 236715
rect 274154 236675 288214 236703
rect 274154 236663 274160 236675
rect 288208 236663 288214 236675
rect 288266 236663 288272 236715
rect 288610 236703 288638 236749
rect 288322 236675 288638 236703
rect 258160 236589 258166 236641
rect 258218 236629 258224 236641
rect 262096 236629 262102 236641
rect 258218 236601 262102 236629
rect 258218 236589 258224 236601
rect 262096 236589 262102 236601
rect 262154 236589 262160 236641
rect 271888 236589 271894 236641
rect 271946 236629 271952 236641
rect 288322 236629 288350 236675
rect 271946 236601 288350 236629
rect 290146 236629 290174 236749
rect 291280 236737 291286 236789
rect 291338 236777 291344 236789
rect 305968 236777 305974 236789
rect 291338 236749 305974 236777
rect 291338 236737 291344 236749
rect 305968 236737 305974 236749
rect 306026 236737 306032 236789
rect 308002 236777 308030 236823
rect 324016 236811 324022 236863
rect 324074 236851 324080 236863
rect 343024 236851 343030 236863
rect 324074 236823 343030 236851
rect 324074 236811 324080 236823
rect 343024 236811 343030 236823
rect 343082 236811 343088 236863
rect 319312 236777 319318 236789
rect 308002 236749 319318 236777
rect 319312 236737 319318 236749
rect 319370 236737 319376 236789
rect 324784 236737 324790 236789
rect 324842 236777 324848 236789
rect 344752 236777 344758 236789
rect 324842 236749 344758 236777
rect 324842 236737 324848 236749
rect 344752 236737 344758 236749
rect 344810 236737 344816 236789
rect 368944 236737 368950 236789
rect 369002 236777 369008 236789
rect 387088 236777 387094 236789
rect 369002 236749 387094 236777
rect 369002 236737 369008 236749
rect 387088 236737 387094 236749
rect 387146 236737 387152 236789
rect 290416 236663 290422 236715
rect 290474 236703 290480 236715
rect 298768 236703 298774 236715
rect 290474 236675 298774 236703
rect 290474 236663 290480 236675
rect 298768 236663 298774 236675
rect 298826 236663 298832 236715
rect 304048 236663 304054 236715
rect 304106 236703 304112 236715
rect 307984 236703 307990 236715
rect 304106 236675 307990 236703
rect 304106 236663 304112 236675
rect 307984 236663 307990 236675
rect 308042 236663 308048 236715
rect 325648 236663 325654 236715
rect 325706 236703 325712 236715
rect 346960 236703 346966 236715
rect 325706 236675 346966 236703
rect 325706 236663 325712 236675
rect 346960 236663 346966 236675
rect 347018 236663 347024 236715
rect 400336 236663 400342 236715
rect 400394 236703 400400 236715
rect 420400 236703 420406 236715
rect 400394 236675 420406 236703
rect 400394 236663 400400 236675
rect 420400 236663 420406 236675
rect 420458 236663 420464 236715
rect 440656 236663 440662 236715
rect 440714 236703 440720 236715
rect 460720 236703 460726 236715
rect 440714 236675 460726 236703
rect 440714 236663 440720 236675
rect 460720 236663 460726 236675
rect 460778 236663 460784 236715
rect 290146 236601 291998 236629
rect 271946 236589 271952 236601
rect 278416 236515 278422 236567
rect 278474 236555 278480 236567
rect 281200 236555 281206 236567
rect 278474 236527 281206 236555
rect 278474 236515 278480 236527
rect 281200 236515 281206 236527
rect 281258 236515 281264 236567
rect 287344 236515 287350 236567
rect 287402 236555 287408 236567
rect 291856 236555 291862 236567
rect 287402 236527 291862 236555
rect 287402 236515 287408 236527
rect 291856 236515 291862 236527
rect 291914 236515 291920 236567
rect 291970 236555 291998 236601
rect 292048 236589 292054 236641
rect 292106 236629 292112 236641
rect 311440 236629 311446 236641
rect 292106 236601 311446 236629
rect 292106 236589 292112 236601
rect 311440 236589 311446 236601
rect 311498 236589 311504 236641
rect 313648 236589 313654 236641
rect 313706 236629 313712 236641
rect 313840 236629 313846 236641
rect 313706 236601 313846 236629
rect 313706 236589 313712 236601
rect 313840 236589 313846 236601
rect 313898 236589 313904 236641
rect 325264 236589 325270 236641
rect 325322 236629 325328 236641
rect 345904 236629 345910 236641
rect 325322 236601 345910 236629
rect 325322 236589 325328 236601
rect 345904 236589 345910 236601
rect 345962 236589 345968 236641
rect 294448 236555 294454 236567
rect 291970 236527 294454 236555
rect 294448 236515 294454 236527
rect 294506 236515 294512 236567
rect 300208 236515 300214 236567
rect 300266 236555 300272 236567
rect 305872 236555 305878 236567
rect 300266 236527 305878 236555
rect 300266 236515 300272 236527
rect 305872 236515 305878 236527
rect 305930 236515 305936 236567
rect 322480 236515 322486 236567
rect 322538 236555 322544 236567
rect 339952 236555 339958 236567
rect 322538 236527 339958 236555
rect 322538 236515 322544 236527
rect 339952 236515 339958 236527
rect 340010 236515 340016 236567
rect 638032 236515 638038 236567
rect 638090 236555 638096 236567
rect 650512 236555 650518 236567
rect 638090 236527 650518 236555
rect 638090 236515 638096 236527
rect 650512 236515 650518 236527
rect 650570 236515 650576 236567
rect 275920 236441 275926 236493
rect 275978 236481 275984 236493
rect 294832 236481 294838 236493
rect 275978 236453 294838 236481
rect 275978 236441 275984 236453
rect 294832 236441 294838 236453
rect 294890 236441 294896 236493
rect 295024 236441 295030 236493
rect 295082 236481 295088 236493
rect 296176 236481 296182 236493
rect 295082 236453 296182 236481
rect 295082 236441 295088 236453
rect 296176 236441 296182 236453
rect 296234 236441 296240 236493
rect 320368 236441 320374 236493
rect 320426 236481 320432 236493
rect 335248 236481 335254 236493
rect 320426 236453 335254 236481
rect 320426 236441 320432 236453
rect 335248 236441 335254 236453
rect 335306 236441 335312 236493
rect 637360 236441 637366 236493
rect 637418 236481 637424 236493
rect 650224 236481 650230 236493
rect 637418 236453 650230 236481
rect 637418 236441 637424 236453
rect 650224 236441 650230 236453
rect 650282 236441 650288 236493
rect 225520 236367 225526 236419
rect 225578 236407 225584 236419
rect 237232 236407 237238 236419
rect 225578 236379 237238 236407
rect 225578 236367 225584 236379
rect 237232 236367 237238 236379
rect 237290 236367 237296 236419
rect 273424 236367 273430 236419
rect 273482 236407 273488 236419
rect 281584 236407 281590 236419
rect 273482 236379 281590 236407
rect 273482 236367 273488 236379
rect 281584 236367 281590 236379
rect 281642 236367 281648 236419
rect 288112 236407 288118 236419
rect 281698 236379 288118 236407
rect 268336 236293 268342 236345
rect 268394 236333 268400 236345
rect 281698 236333 281726 236379
rect 288112 236367 288118 236379
rect 288170 236367 288176 236419
rect 289936 236367 289942 236419
rect 289994 236407 290000 236419
rect 289994 236379 307454 236407
rect 289994 236367 290000 236379
rect 268394 236305 281726 236333
rect 268394 236293 268400 236305
rect 282736 236293 282742 236345
rect 282794 236333 282800 236345
rect 297808 236333 297814 236345
rect 282794 236305 297814 236333
rect 282794 236293 282800 236305
rect 297808 236293 297814 236305
rect 297866 236293 297872 236345
rect 144112 236219 144118 236271
rect 144170 236259 144176 236271
rect 168400 236259 168406 236271
rect 144170 236231 168406 236259
rect 144170 236219 144176 236231
rect 168400 236219 168406 236231
rect 168458 236219 168464 236271
rect 271408 236219 271414 236271
rect 271466 236259 271472 236271
rect 288976 236259 288982 236271
rect 271466 236231 288982 236259
rect 271466 236219 271472 236231
rect 288976 236219 288982 236231
rect 289034 236219 289040 236271
rect 289072 236219 289078 236271
rect 289130 236259 289136 236271
rect 290704 236259 290710 236271
rect 289130 236231 290710 236259
rect 289130 236219 289136 236231
rect 290704 236219 290710 236231
rect 290762 236219 290768 236271
rect 290800 236219 290806 236271
rect 290858 236259 290864 236271
rect 293968 236259 293974 236271
rect 290858 236231 293974 236259
rect 290858 236219 290864 236231
rect 293968 236219 293974 236231
rect 294026 236219 294032 236271
rect 294064 236219 294070 236271
rect 294122 236259 294128 236271
rect 296464 236259 296470 236271
rect 294122 236231 296470 236259
rect 294122 236219 294128 236231
rect 296464 236219 296470 236231
rect 296522 236219 296528 236271
rect 307426 236259 307454 236379
rect 319984 236367 319990 236419
rect 320042 236407 320048 236419
rect 334384 236407 334390 236419
rect 320042 236379 334390 236407
rect 320042 236367 320048 236379
rect 334384 236367 334390 236379
rect 334442 236367 334448 236419
rect 637936 236367 637942 236419
rect 637994 236407 638000 236419
rect 650320 236407 650326 236419
rect 637994 236379 650326 236407
rect 637994 236367 638000 236379
rect 650320 236367 650326 236379
rect 650378 236367 650384 236419
rect 318064 236293 318070 236345
rect 318122 236333 318128 236345
rect 335632 236333 335638 236345
rect 318122 236305 335638 236333
rect 318122 236293 318128 236305
rect 335632 236293 335638 236305
rect 335690 236293 335696 236345
rect 639184 236293 639190 236345
rect 639242 236333 639248 236345
rect 649840 236333 649846 236345
rect 639242 236305 649846 236333
rect 639242 236293 639248 236305
rect 649840 236293 649846 236305
rect 649898 236293 649904 236345
rect 315376 236259 315382 236271
rect 307426 236231 315382 236259
rect 315376 236219 315382 236231
rect 315434 236219 315440 236271
rect 315952 236219 315958 236271
rect 316010 236259 316016 236271
rect 328432 236259 328438 236271
rect 316010 236231 328438 236259
rect 316010 236219 316016 236231
rect 328432 236219 328438 236231
rect 328490 236219 328496 236271
rect 638800 236219 638806 236271
rect 638858 236259 638864 236271
rect 649648 236259 649654 236271
rect 638858 236231 649654 236259
rect 638858 236219 638864 236231
rect 649648 236219 649654 236231
rect 649706 236219 649712 236271
rect 144016 236145 144022 236197
rect 144074 236185 144080 236197
rect 171280 236185 171286 236197
rect 144074 236157 171286 236185
rect 144074 236145 144080 236157
rect 171280 236145 171286 236157
rect 171338 236145 171344 236197
rect 210352 236145 210358 236197
rect 210410 236185 210416 236197
rect 210736 236185 210742 236197
rect 210410 236157 210742 236185
rect 210410 236145 210416 236157
rect 210736 236145 210742 236157
rect 210794 236185 210800 236197
rect 213040 236185 213046 236197
rect 210794 236157 213046 236185
rect 210794 236145 210800 236157
rect 213040 236145 213046 236157
rect 213098 236145 213104 236197
rect 217456 236145 217462 236197
rect 217514 236185 217520 236197
rect 221776 236185 221782 236197
rect 217514 236157 221782 236185
rect 217514 236145 217520 236157
rect 221776 236145 221782 236157
rect 221834 236145 221840 236197
rect 281680 236145 281686 236197
rect 281738 236185 281744 236197
rect 297424 236185 297430 236197
rect 281738 236157 297430 236185
rect 281738 236145 281744 236157
rect 297424 236145 297430 236157
rect 297482 236145 297488 236197
rect 547120 236145 547126 236197
rect 547178 236185 547184 236197
rect 549232 236185 549238 236197
rect 547178 236157 549238 236185
rect 547178 236145 547184 236157
rect 549232 236145 549238 236157
rect 549290 236145 549296 236197
rect 639760 236145 639766 236197
rect 639818 236185 639824 236197
rect 650032 236185 650038 236197
rect 639818 236157 650038 236185
rect 639818 236145 639824 236157
rect 650032 236145 650038 236157
rect 650090 236145 650096 236197
rect 265648 236071 265654 236123
rect 265706 236111 265712 236123
rect 308272 236111 308278 236123
rect 265706 236083 308278 236111
rect 265706 236071 265712 236083
rect 308272 236071 308278 236083
rect 308330 236071 308336 236123
rect 264880 235997 264886 236049
rect 264938 236037 264944 236049
rect 309904 236037 309910 236049
rect 264938 236009 309910 236037
rect 264938 235997 264944 236009
rect 309904 235997 309910 236009
rect 309962 235997 309968 236049
rect 312976 235997 312982 236049
rect 313034 236037 313040 236049
rect 369616 236037 369622 236049
rect 313034 236009 369622 236037
rect 313034 235997 313040 236009
rect 369616 235997 369622 236009
rect 369674 235997 369680 236049
rect 265072 235923 265078 235975
rect 265130 235963 265136 235975
rect 339376 235963 339382 235975
rect 265130 235935 339382 235963
rect 265130 235923 265136 235935
rect 339376 235923 339382 235935
rect 339434 235923 339440 235975
rect 381904 235923 381910 235975
rect 381962 235963 381968 235975
rect 390928 235963 390934 235975
rect 381962 235935 390934 235963
rect 381962 235923 381968 235935
rect 390928 235923 390934 235935
rect 390986 235923 390992 235975
rect 235696 235849 235702 235901
rect 235754 235889 235760 235901
rect 266128 235889 266134 235901
rect 235754 235861 266134 235889
rect 235754 235849 235760 235861
rect 266128 235849 266134 235861
rect 266186 235849 266192 235901
rect 267088 235849 267094 235901
rect 267146 235889 267152 235901
rect 340336 235889 340342 235901
rect 267146 235861 340342 235889
rect 267146 235849 267152 235861
rect 340336 235849 340342 235861
rect 340394 235849 340400 235901
rect 263728 235775 263734 235827
rect 263786 235815 263792 235827
rect 338896 235815 338902 235827
rect 263786 235787 338902 235815
rect 263786 235775 263792 235787
rect 338896 235775 338902 235787
rect 338954 235775 338960 235827
rect 258928 235701 258934 235753
rect 258986 235741 258992 235753
rect 336688 235741 336694 235753
rect 258986 235713 336694 235741
rect 258986 235701 258992 235713
rect 336688 235701 336694 235713
rect 336746 235701 336752 235753
rect 480976 235701 480982 235753
rect 481034 235741 481040 235753
rect 497488 235741 497494 235753
rect 481034 235713 497494 235741
rect 481034 235701 481040 235713
rect 497488 235701 497494 235713
rect 497546 235701 497552 235753
rect 261904 235627 261910 235679
rect 261962 235667 261968 235679
rect 338128 235667 338134 235679
rect 261962 235639 338134 235667
rect 261962 235627 261968 235639
rect 338128 235627 338134 235639
rect 338186 235627 338192 235679
rect 257296 235553 257302 235605
rect 257354 235593 257360 235605
rect 335920 235593 335926 235605
rect 257354 235565 335926 235593
rect 257354 235553 257360 235565
rect 335920 235553 335926 235565
rect 335978 235553 335984 235605
rect 260560 235479 260566 235531
rect 260618 235519 260624 235531
rect 337168 235519 337174 235531
rect 260618 235491 337174 235519
rect 260618 235479 260624 235491
rect 337168 235479 337174 235491
rect 337226 235479 337232 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 43024 235445 43030 235457
rect 42218 235417 43030 235445
rect 42218 235405 42224 235417
rect 43024 235405 43030 235417
rect 43082 235405 43088 235457
rect 236080 235405 236086 235457
rect 236138 235445 236144 235457
rect 265456 235445 265462 235457
rect 236138 235417 265462 235445
rect 236138 235405 236144 235417
rect 265456 235405 265462 235417
rect 265514 235405 265520 235457
rect 274384 235405 274390 235457
rect 274442 235445 274448 235457
rect 356656 235445 356662 235457
rect 274442 235417 356662 235445
rect 274442 235405 274448 235417
rect 356656 235405 356662 235417
rect 356714 235405 356720 235457
rect 246256 235331 246262 235383
rect 246314 235371 246320 235383
rect 353584 235371 353590 235383
rect 246314 235343 353590 235371
rect 246314 235331 246320 235343
rect 353584 235331 353590 235343
rect 353642 235331 353648 235383
rect 250384 235257 250390 235309
rect 250442 235297 250448 235309
rect 354832 235297 354838 235309
rect 250442 235269 354838 235297
rect 250442 235257 250448 235269
rect 354832 235257 354838 235269
rect 354890 235257 354896 235309
rect 241648 235183 241654 235235
rect 241706 235223 241712 235235
rect 349936 235223 349942 235235
rect 241706 235195 349942 235223
rect 241706 235183 241712 235195
rect 349936 235183 349942 235195
rect 349994 235183 350000 235235
rect 242032 235109 242038 235161
rect 242090 235149 242096 235161
rect 352144 235149 352150 235161
rect 242090 235121 352150 235149
rect 242090 235109 242096 235121
rect 352144 235109 352150 235121
rect 352202 235109 352208 235161
rect 241840 235035 241846 235087
rect 241898 235075 241904 235087
rect 350416 235075 350422 235087
rect 241898 235047 350422 235075
rect 241898 235035 241904 235047
rect 350416 235035 350422 235047
rect 350474 235035 350480 235087
rect 246448 234961 246454 235013
rect 246506 235001 246512 235013
rect 354352 235001 354358 235013
rect 246506 234973 354358 235001
rect 246506 234961 246512 234973
rect 354352 234961 354358 234973
rect 354410 234961 354416 235013
rect 243280 234887 243286 234939
rect 243338 234927 243344 234939
rect 352624 234927 352630 234939
rect 243338 234899 352630 234927
rect 243338 234887 243344 234899
rect 352624 234887 352630 234899
rect 352682 234887 352688 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42448 234853 42454 234865
rect 42218 234825 42454 234853
rect 42218 234813 42224 234825
rect 42448 234813 42454 234825
rect 42506 234813 42512 234865
rect 244144 234813 244150 234865
rect 244202 234853 244208 234865
rect 351376 234853 351382 234865
rect 244202 234825 351382 234853
rect 244202 234813 244208 234825
rect 351376 234813 351382 234825
rect 351434 234813 351440 234865
rect 230608 234739 230614 234791
rect 230666 234779 230672 234791
rect 346960 234779 346966 234791
rect 230666 234751 346966 234779
rect 230666 234739 230672 234751
rect 346960 234739 346966 234751
rect 347018 234739 347024 234791
rect 227824 234665 227830 234717
rect 227882 234705 227888 234717
rect 345520 234705 345526 234717
rect 227882 234677 345526 234705
rect 227882 234665 227888 234677
rect 345520 234665 345526 234677
rect 345578 234665 345584 234717
rect 282448 234591 282454 234643
rect 282506 234631 282512 234643
rect 322768 234631 322774 234643
rect 282506 234603 322774 234631
rect 282506 234591 282512 234603
rect 322768 234591 322774 234603
rect 322826 234591 322832 234643
rect 266992 234517 266998 234569
rect 267050 234557 267056 234569
rect 305680 234557 305686 234569
rect 267050 234529 305686 234557
rect 267050 234517 267056 234529
rect 305680 234517 305686 234529
rect 305738 234517 305744 234569
rect 282832 234443 282838 234495
rect 282890 234483 282896 234495
rect 321904 234483 321910 234495
rect 282890 234455 321910 234483
rect 282890 234443 282896 234455
rect 321904 234443 321910 234455
rect 321962 234443 321968 234495
rect 267472 234369 267478 234421
rect 267530 234409 267536 234421
rect 304240 234409 304246 234421
rect 267530 234381 304246 234409
rect 267530 234369 267536 234381
rect 304240 234369 304246 234381
rect 304298 234369 304304 234421
rect 271600 234295 271606 234347
rect 271658 234335 271664 234347
rect 309424 234335 309430 234347
rect 271658 234307 309430 234335
rect 271658 234295 271664 234307
rect 309424 234295 309430 234307
rect 309482 234295 309488 234347
rect 284656 234221 284662 234273
rect 284714 234261 284720 234273
rect 317488 234261 317494 234273
rect 284714 234233 317494 234261
rect 284714 234221 284720 234233
rect 317488 234221 317494 234233
rect 317546 234221 317552 234273
rect 284272 234147 284278 234199
rect 284330 234187 284336 234199
rect 319120 234187 319126 234199
rect 284330 234159 319126 234187
rect 284330 234147 284336 234159
rect 319120 234147 319126 234159
rect 319178 234147 319184 234199
rect 268816 234073 268822 234125
rect 268874 234113 268880 234125
rect 301936 234113 301942 234125
rect 268874 234085 301942 234113
rect 268874 234073 268880 234085
rect 301936 234073 301942 234085
rect 301994 234073 302000 234125
rect 269584 233999 269590 234051
rect 269642 234039 269648 234051
rect 300304 234039 300310 234051
rect 269642 234011 300310 234039
rect 269642 233999 269648 234011
rect 300304 233999 300310 234011
rect 300362 233999 300368 234051
rect 285136 233925 285142 233977
rect 285194 233965 285200 233977
rect 316144 233965 316150 233977
rect 285194 233937 316150 233965
rect 285194 233925 285200 233937
rect 316144 233925 316150 233937
rect 316202 233925 316208 233977
rect 274864 233851 274870 233903
rect 274922 233891 274928 233903
rect 288592 233891 288598 233903
rect 274922 233863 288598 233891
rect 274922 233851 274928 233863
rect 288592 233851 288598 233863
rect 288650 233851 288656 233903
rect 292528 233851 292534 233903
rect 292586 233891 292592 233903
rect 320560 233891 320566 233903
rect 292586 233863 320566 233891
rect 292586 233851 292592 233863
rect 320560 233851 320566 233863
rect 320618 233851 320624 233903
rect 293104 233777 293110 233829
rect 293162 233817 293168 233829
rect 321424 233817 321430 233829
rect 293162 233789 321430 233817
rect 293162 233777 293168 233789
rect 321424 233777 321430 233789
rect 321482 233777 321488 233829
rect 209776 233703 209782 233755
rect 209834 233743 209840 233755
rect 212176 233743 212182 233755
rect 209834 233715 212182 233743
rect 209834 233703 209840 233715
rect 212176 233703 212182 233715
rect 212234 233703 212240 233755
rect 238048 233703 238054 233755
rect 238106 233743 238112 233755
rect 239056 233743 239062 233755
rect 238106 233715 239062 233743
rect 238106 233703 238112 233715
rect 239056 233703 239062 233715
rect 239114 233703 239120 233755
rect 270064 233703 270070 233755
rect 270122 233743 270128 233755
rect 298576 233743 298582 233755
rect 270122 233715 298582 233743
rect 270122 233703 270128 233715
rect 298576 233703 298582 233715
rect 298634 233703 298640 233755
rect 305584 233703 305590 233755
rect 305642 233743 305648 233755
rect 308704 233743 308710 233755
rect 305642 233715 308710 233743
rect 305642 233703 305648 233715
rect 308704 233703 308710 233715
rect 308762 233703 308768 233755
rect 208144 233629 208150 233681
rect 208202 233669 208208 233681
rect 213520 233669 213526 233681
rect 208202 233641 213526 233669
rect 208202 233629 208208 233641
rect 213520 233629 213526 233641
rect 213578 233629 213584 233681
rect 270640 233629 270646 233681
rect 270698 233669 270704 233681
rect 298480 233669 298486 233681
rect 270698 233641 298486 233669
rect 270698 233629 270704 233641
rect 298480 233629 298486 233641
rect 298538 233629 298544 233681
rect 316912 233669 316918 233681
rect 307906 233641 316918 233669
rect 209968 233555 209974 233607
rect 210026 233595 210032 233607
rect 213136 233595 213142 233607
rect 210026 233567 213142 233595
rect 210026 233555 210032 233567
rect 213136 233555 213142 233567
rect 213194 233555 213200 233607
rect 269104 233555 269110 233607
rect 269162 233595 269168 233607
rect 297040 233595 297046 233607
rect 269162 233567 297046 233595
rect 269162 233555 269168 233567
rect 297040 233555 297046 233567
rect 297098 233555 297104 233607
rect 298192 233555 298198 233607
rect 298250 233595 298256 233607
rect 298250 233567 299486 233595
rect 298250 233555 298256 233567
rect 210256 233481 210262 233533
rect 210314 233521 210320 233533
rect 210928 233521 210934 233533
rect 210314 233493 210934 233521
rect 210314 233481 210320 233493
rect 210928 233481 210934 233493
rect 210986 233481 210992 233533
rect 211299 233526 211374 233532
rect 211299 233514 211307 233526
rect 211298 233486 211307 233514
rect 211299 233474 211307 233486
rect 211359 233514 211374 233526
rect 213904 233514 213910 233533
rect 211359 233486 213910 233514
rect 211359 233474 211374 233486
rect 213904 233481 213910 233486
rect 213962 233481 213968 233533
rect 299458 233521 299486 233567
rect 307906 233521 307934 233641
rect 316912 233629 316918 233641
rect 316970 233629 316976 233681
rect 299458 233493 307934 233521
rect 211299 233465 211374 233474
rect 144016 233259 144022 233311
rect 144074 233299 144080 233311
rect 165520 233299 165526 233311
rect 144074 233271 165526 233299
rect 144074 233259 144080 233271
rect 165520 233259 165526 233271
rect 165578 233259 165584 233311
rect 206512 233185 206518 233237
rect 206570 233225 206576 233237
rect 206608 233225 206614 233237
rect 206570 233197 206614 233225
rect 206570 233185 206576 233197
rect 206608 233185 206614 233197
rect 206666 233185 206672 233237
rect 645712 233185 645718 233237
rect 645770 233225 645776 233237
rect 649744 233225 649750 233237
rect 645770 233197 649750 233225
rect 645770 233185 645776 233197
rect 649744 233185 649750 233197
rect 649802 233185 649808 233237
rect 645808 233111 645814 233163
rect 645866 233151 645872 233163
rect 649936 233151 649942 233163
rect 645866 233123 649942 233151
rect 645866 233111 645872 233123
rect 649936 233111 649942 233123
rect 649994 233111 650000 233163
rect 645136 233037 645142 233089
rect 645194 233077 645200 233089
rect 650416 233077 650422 233089
rect 645194 233049 650422 233077
rect 645194 233037 645200 233049
rect 650416 233037 650422 233049
rect 650474 233037 650480 233089
rect 645328 232963 645334 233015
rect 645386 233003 645392 233015
rect 650128 233003 650134 233015
rect 645386 232975 650134 233003
rect 645386 232963 645392 232975
rect 650128 232963 650134 232975
rect 650186 232963 650192 233015
rect 645232 232889 645238 232941
rect 645290 232929 645296 232941
rect 650608 232929 650614 232941
rect 645290 232901 650614 232929
rect 645290 232889 645296 232901
rect 650608 232889 650614 232901
rect 650666 232889 650672 232941
rect 205072 232593 205078 232645
rect 205130 232593 205136 232645
rect 205090 232497 205118 232593
rect 205072 232445 205078 232497
rect 205130 232445 205136 232497
rect 42064 231039 42070 231091
rect 42122 231079 42128 231091
rect 42928 231079 42934 231091
rect 42122 231051 42934 231079
rect 42122 231039 42128 231051
rect 42928 231039 42934 231051
rect 42986 231039 42992 231091
rect 206896 230669 206902 230721
rect 206954 230709 206960 230721
rect 207088 230709 207094 230721
rect 206954 230681 207094 230709
rect 206954 230669 206960 230681
rect 207088 230669 207094 230681
rect 207146 230669 207152 230721
rect 144016 230521 144022 230573
rect 144074 230561 144080 230573
rect 151120 230561 151126 230573
rect 144074 230533 151126 230561
rect 144074 230521 144080 230533
rect 151120 230521 151126 230533
rect 151178 230521 151184 230573
rect 206320 230521 206326 230573
rect 206378 230561 206384 230573
rect 206896 230561 206902 230573
rect 206378 230533 206902 230561
rect 206378 230521 206384 230533
rect 206896 230521 206902 230533
rect 206954 230521 206960 230573
rect 144112 230447 144118 230499
rect 144170 230487 144176 230499
rect 202960 230487 202966 230499
rect 144170 230459 202966 230487
rect 144170 230447 144176 230459
rect 202960 230447 202966 230459
rect 203018 230447 203024 230499
rect 144016 227709 144022 227761
rect 144074 227749 144080 227761
rect 188560 227749 188566 227761
rect 144074 227721 188566 227749
rect 144074 227709 144080 227721
rect 188560 227709 188566 227721
rect 188618 227709 188624 227761
rect 144112 227635 144118 227687
rect 144170 227675 144176 227687
rect 194320 227675 194326 227687
rect 144170 227647 194326 227675
rect 144170 227635 144176 227647
rect 194320 227635 194326 227647
rect 194378 227635 194384 227687
rect 144208 227561 144214 227613
rect 144266 227601 144272 227613
rect 197200 227601 197206 227613
rect 144266 227573 197206 227601
rect 144266 227561 144272 227573
rect 197200 227561 197206 227573
rect 197258 227561 197264 227613
rect 204880 227117 204886 227169
rect 204938 227157 204944 227169
rect 205648 227157 205654 227169
rect 204938 227129 205654 227157
rect 204938 227117 204944 227129
rect 205648 227117 205654 227129
rect 205706 227117 205712 227169
rect 146800 225637 146806 225689
rect 146858 225677 146864 225689
rect 156880 225677 156886 225689
rect 146858 225649 156886 225677
rect 146858 225637 146864 225649
rect 156880 225637 156886 225649
rect 156938 225637 156944 225689
rect 666832 225045 666838 225097
rect 666890 225085 666896 225097
rect 674704 225085 674710 225097
rect 666890 225057 674710 225085
rect 666890 225045 666896 225057
rect 674704 225045 674710 225057
rect 674762 225045 674768 225097
rect 146800 224675 146806 224727
rect 146858 224715 146864 224727
rect 200080 224715 200086 224727
rect 146858 224687 200086 224715
rect 146858 224675 146864 224687
rect 200080 224675 200086 224687
rect 200138 224675 200144 224727
rect 141040 224601 141046 224653
rect 141098 224641 141104 224653
rect 199696 224641 199702 224653
rect 141098 224613 199702 224641
rect 141098 224601 141104 224613
rect 199696 224601 199702 224613
rect 199754 224601 199760 224653
rect 146416 224527 146422 224579
rect 146474 224567 146480 224579
rect 201712 224567 201718 224579
rect 146474 224539 201718 224567
rect 146474 224527 146480 224539
rect 201712 224527 201718 224539
rect 201770 224527 201776 224579
rect 149680 224453 149686 224505
rect 149738 224493 149744 224505
rect 201616 224493 201622 224505
rect 149738 224465 201622 224493
rect 149738 224453 149744 224465
rect 201616 224453 201622 224465
rect 201674 224453 201680 224505
rect 152560 224379 152566 224431
rect 152618 224419 152624 224431
rect 201808 224419 201814 224431
rect 152618 224391 201814 224419
rect 152618 224379 152624 224391
rect 201808 224379 201814 224391
rect 201866 224379 201872 224431
rect 669616 224305 669622 224357
rect 669674 224345 669680 224357
rect 674416 224345 674422 224357
rect 669674 224317 674422 224345
rect 669674 224305 669680 224317
rect 674416 224305 674422 224317
rect 674474 224305 674480 224357
rect 669520 224009 669526 224061
rect 669578 224049 669584 224061
rect 674704 224049 674710 224061
rect 669578 224021 674710 224049
rect 669578 224009 669584 224021
rect 674704 224009 674710 224021
rect 674762 224009 674768 224061
rect 205744 223121 205750 223173
rect 205802 223161 205808 223173
rect 206128 223161 206134 223173
rect 205802 223133 206134 223161
rect 205802 223121 205808 223133
rect 206128 223121 206134 223133
rect 206186 223121 206192 223173
rect 146704 221937 146710 221989
rect 146762 221977 146768 221989
rect 177040 221977 177046 221989
rect 146762 221949 177046 221977
rect 146762 221937 146768 221949
rect 177040 221937 177046 221949
rect 177098 221937 177104 221989
rect 146800 221863 146806 221915
rect 146858 221903 146864 221915
rect 179920 221903 179926 221915
rect 146858 221875 179926 221903
rect 146858 221863 146864 221875
rect 179920 221863 179926 221875
rect 179978 221863 179984 221915
rect 144400 221789 144406 221841
rect 144458 221829 144464 221841
rect 182800 221829 182806 221841
rect 144458 221801 182806 221829
rect 144458 221789 144464 221801
rect 182800 221789 182806 221801
rect 182858 221789 182864 221841
rect 155440 221715 155446 221767
rect 155498 221755 155504 221767
rect 198832 221755 198838 221767
rect 155498 221727 198838 221755
rect 155498 221715 155504 221727
rect 198832 221715 198838 221727
rect 198890 221715 198896 221767
rect 161200 221641 161206 221693
rect 161258 221681 161264 221693
rect 210160 221681 210166 221693
rect 161258 221653 210166 221681
rect 161258 221641 161264 221653
rect 210160 221641 210166 221653
rect 210218 221641 210224 221693
rect 164080 221567 164086 221619
rect 164138 221607 164144 221619
rect 201712 221607 201718 221619
rect 164138 221579 201718 221607
rect 164138 221567 164144 221579
rect 201712 221567 201718 221579
rect 201770 221567 201776 221619
rect 166960 221493 166966 221545
rect 167018 221533 167024 221545
rect 201616 221533 201622 221545
rect 167018 221505 201622 221533
rect 167018 221493 167024 221505
rect 201616 221493 201622 221505
rect 201674 221493 201680 221545
rect 169840 221419 169846 221471
rect 169898 221459 169904 221471
rect 196048 221459 196054 221471
rect 169898 221431 196054 221459
rect 169898 221419 169904 221431
rect 196048 221419 196054 221431
rect 196106 221419 196112 221471
rect 144400 218903 144406 218955
rect 144458 218943 144464 218955
rect 174256 218943 174262 218955
rect 144458 218915 174262 218943
rect 144458 218903 144464 218915
rect 174256 218903 174262 218915
rect 174314 218903 174320 218955
rect 175600 218829 175606 218881
rect 175658 218869 175664 218881
rect 200656 218869 200662 218881
rect 175658 218841 200662 218869
rect 175658 218829 175664 218841
rect 200656 218829 200662 218841
rect 200714 218829 200720 218881
rect 178480 218755 178486 218807
rect 178538 218795 178544 218807
rect 201712 218795 201718 218807
rect 178538 218767 201718 218795
rect 178538 218755 178544 218767
rect 201712 218755 201718 218767
rect 201770 218755 201776 218807
rect 181360 218681 181366 218733
rect 181418 218721 181424 218733
rect 210160 218721 210166 218733
rect 181418 218693 210166 218721
rect 181418 218681 181424 218693
rect 210160 218681 210166 218693
rect 210218 218681 210224 218733
rect 184240 218607 184246 218659
rect 184298 218647 184304 218659
rect 201616 218647 201622 218659
rect 184298 218619 201622 218647
rect 184298 218607 184304 218619
rect 201616 218607 201622 218619
rect 201674 218607 201680 218659
rect 42448 216461 42454 216513
rect 42506 216501 42512 216513
rect 45136 216501 45142 216513
rect 42506 216473 45142 216501
rect 42506 216461 42512 216473
rect 45136 216461 45142 216473
rect 45194 216461 45200 216513
rect 146800 216313 146806 216365
rect 146858 216353 146864 216365
rect 154000 216353 154006 216365
rect 146858 216325 154006 216353
rect 146858 216313 146864 216325
rect 154000 216313 154006 216325
rect 154058 216313 154064 216365
rect 645424 216017 645430 216069
rect 645482 216057 645488 216069
rect 645808 216057 645814 216069
rect 645482 216029 645814 216057
rect 645482 216017 645488 216029
rect 645808 216017 645814 216029
rect 645866 216017 645872 216069
rect 187120 215943 187126 215995
rect 187178 215983 187184 215995
rect 210160 215983 210166 215995
rect 187178 215955 210166 215983
rect 187178 215943 187184 215955
rect 210160 215943 210166 215955
rect 210218 215943 210224 215995
rect 674128 215943 674134 215995
rect 674186 215983 674192 215995
rect 674512 215983 674518 215995
rect 674186 215955 674518 215983
rect 674186 215943 674192 215955
rect 674512 215943 674518 215955
rect 674570 215943 674576 215995
rect 192880 215869 192886 215921
rect 192938 215909 192944 215921
rect 201712 215909 201718 215921
rect 192938 215881 201718 215909
rect 192938 215869 192944 215881
rect 201712 215869 201718 215881
rect 201770 215869 201776 215921
rect 42832 215721 42838 215773
rect 42890 215761 42896 215773
rect 45040 215761 45046 215773
rect 42890 215733 45046 215761
rect 42890 215721 42896 215733
rect 45040 215721 45046 215733
rect 45098 215721 45104 215773
rect 42832 215203 42838 215255
rect 42890 215243 42896 215255
rect 44656 215243 44662 215255
rect 42890 215215 44662 215243
rect 42890 215203 42896 215215
rect 44656 215203 44662 215215
rect 44714 215203 44720 215255
rect 206032 213501 206038 213553
rect 206090 213541 206096 213553
rect 206320 213541 206326 213553
rect 206090 213513 206326 213541
rect 206090 213501 206096 213513
rect 206320 213501 206326 213513
rect 206378 213501 206384 213553
rect 146800 213205 146806 213257
rect 146858 213245 146864 213257
rect 168496 213245 168502 213257
rect 146858 213217 168502 213245
rect 146858 213205 146864 213217
rect 168496 213205 168502 213217
rect 168554 213205 168560 213257
rect 144208 213131 144214 213183
rect 144266 213171 144272 213183
rect 171376 213171 171382 213183
rect 144266 213143 171382 213171
rect 144266 213131 144272 213143
rect 171376 213131 171382 213143
rect 171434 213131 171440 213183
rect 146800 210245 146806 210297
rect 146858 210285 146864 210297
rect 148240 210285 148246 210297
rect 146858 210257 148246 210285
rect 146858 210245 146864 210257
rect 148240 210245 148246 210257
rect 148298 210245 148304 210297
rect 647920 210245 647926 210297
rect 647978 210285 647984 210297
rect 677008 210285 677014 210297
rect 647978 210257 677014 210285
rect 647978 210245 647984 210257
rect 677008 210245 677014 210257
rect 677066 210245 677072 210297
rect 146704 207433 146710 207485
rect 146762 207473 146768 207485
rect 165616 207473 165622 207485
rect 146762 207445 165622 207473
rect 146762 207433 146768 207445
rect 165616 207433 165622 207445
rect 165674 207433 165680 207485
rect 146800 207359 146806 207411
rect 146858 207399 146864 207411
rect 203056 207399 203062 207411
rect 146858 207371 203062 207399
rect 146858 207359 146864 207371
rect 203056 207359 203062 207371
rect 203114 207359 203120 207411
rect 645424 207285 645430 207337
rect 645482 207325 645488 207337
rect 645808 207325 645814 207337
rect 645482 207297 645814 207325
rect 645482 207285 645488 207297
rect 645808 207285 645814 207297
rect 645866 207285 645872 207337
rect 42448 204399 42454 204451
rect 42506 204439 42512 204451
rect 50320 204439 50326 204451
rect 42506 204411 50326 204439
rect 42506 204399 42512 204411
rect 50320 204399 50326 204411
rect 50378 204399 50384 204451
rect 674992 204399 674998 204451
rect 675050 204439 675056 204451
rect 675376 204439 675382 204451
rect 675050 204411 675382 204439
rect 675050 204399 675056 204411
rect 675376 204399 675382 204411
rect 675434 204399 675440 204451
rect 146800 201661 146806 201713
rect 146858 201701 146864 201713
rect 159760 201701 159766 201713
rect 146858 201673 159766 201701
rect 146858 201661 146864 201673
rect 159760 201661 159766 201673
rect 159818 201661 159824 201713
rect 144976 201587 144982 201639
rect 145034 201627 145040 201639
rect 162640 201627 162646 201639
rect 145034 201599 162646 201627
rect 145034 201587 145040 201599
rect 162640 201587 162646 201599
rect 162698 201587 162704 201639
rect 674128 201291 674134 201343
rect 674186 201331 674192 201343
rect 675376 201331 675382 201343
rect 674186 201303 675382 201331
rect 674186 201291 674192 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 40048 200107 40054 200159
rect 40106 200147 40112 200159
rect 43120 200147 43126 200159
rect 40106 200119 43126 200147
rect 40106 200107 40112 200119
rect 43120 200107 43126 200119
rect 43178 200107 43184 200159
rect 40144 198997 40150 199049
rect 40202 199037 40208 199049
rect 42352 199037 42358 199049
rect 40202 199009 42358 199037
rect 40202 198997 40208 199009
rect 42352 198997 42358 199009
rect 42410 198997 42416 199049
rect 39952 198775 39958 198827
rect 40010 198815 40016 198827
rect 43312 198815 43318 198827
rect 40010 198787 43318 198815
rect 40010 198775 40016 198787
rect 43312 198775 43318 198787
rect 43370 198775 43376 198827
rect 40240 198701 40246 198753
rect 40298 198741 40304 198753
rect 41008 198741 41014 198753
rect 40298 198713 41014 198741
rect 40298 198701 40304 198713
rect 41008 198701 41014 198713
rect 41066 198701 41072 198753
rect 146800 198701 146806 198753
rect 146858 198741 146864 198753
rect 191440 198741 191446 198753
rect 146858 198713 191446 198741
rect 146858 198701 146864 198713
rect 191440 198701 191446 198713
rect 191498 198701 191504 198753
rect 674704 197591 674710 197643
rect 674762 197631 674768 197643
rect 675376 197631 675382 197643
rect 674762 197603 675382 197631
rect 674762 197591 674768 197603
rect 675376 197591 675382 197603
rect 675434 197591 675440 197643
rect 42064 197369 42070 197421
rect 42122 197369 42128 197421
rect 42082 197199 42110 197369
rect 42064 197147 42070 197199
rect 42122 197147 42128 197199
rect 674512 196999 674518 197051
rect 674570 197039 674576 197051
rect 675472 197039 675478 197051
rect 674570 197011 675478 197039
rect 674570 196999 674576 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 42352 196851 42358 196903
rect 42410 196891 42416 196903
rect 43216 196891 43222 196903
rect 42410 196863 43222 196891
rect 42410 196851 42416 196863
rect 43216 196851 43222 196863
rect 43274 196851 43280 196903
rect 674608 196555 674614 196607
rect 674666 196595 674672 196607
rect 675376 196595 675382 196607
rect 674666 196567 675382 196595
rect 674666 196555 674672 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 146800 195815 146806 195867
rect 146858 195855 146864 195867
rect 185680 195855 185686 195867
rect 146858 195827 185686 195855
rect 146858 195815 146864 195827
rect 185680 195815 185686 195827
rect 185738 195815 185744 195867
rect 42448 195593 42454 195645
rect 42506 195593 42512 195645
rect 42160 195297 42166 195349
rect 42218 195337 42224 195349
rect 42466 195337 42494 195593
rect 42218 195309 42494 195337
rect 42218 195297 42224 195309
rect 42928 194779 42934 194831
rect 42986 194819 42992 194831
rect 43216 194819 43222 194831
rect 42986 194791 43222 194819
rect 42986 194779 42992 194791
rect 43216 194779 43222 194791
rect 43274 194779 43280 194831
rect 42832 194705 42838 194757
rect 42890 194745 42896 194757
rect 43312 194745 43318 194757
rect 42890 194717 43318 194745
rect 42890 194705 42896 194717
rect 43312 194705 43318 194717
rect 43370 194705 43376 194757
rect 42064 194483 42070 194535
rect 42122 194523 42128 194535
rect 44752 194523 44758 194535
rect 42122 194495 44758 194523
rect 42122 194483 42128 194495
rect 44752 194483 44758 194495
rect 44810 194483 44816 194535
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 43120 193487 43126 193499
rect 42122 193459 43126 193487
rect 42122 193447 42128 193459
rect 43120 193447 43126 193459
rect 43178 193447 43184 193499
rect 206896 192929 206902 192981
rect 206954 192969 206960 192981
rect 206992 192969 206998 192981
rect 206954 192941 206998 192969
rect 206954 192929 206960 192941
rect 206992 192929 206998 192941
rect 207050 192929 207056 192981
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 43024 192229 43030 192241
rect 42218 192201 43030 192229
rect 42218 192189 42224 192201
rect 43024 192189 43030 192201
rect 43082 192189 43088 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 42928 191489 42934 191501
rect 42122 191461 42934 191489
rect 42122 191449 42128 191461
rect 42928 191449 42934 191461
rect 42986 191449 42992 191501
rect 146704 190191 146710 190243
rect 146762 190231 146768 190243
rect 151216 190231 151222 190243
rect 146762 190203 151222 190231
rect 146762 190191 146768 190203
rect 151216 190191 151222 190203
rect 151274 190191 151280 190243
rect 146800 190117 146806 190169
rect 146858 190157 146864 190169
rect 148432 190157 148438 190169
rect 146858 190129 148438 190157
rect 146858 190117 146864 190129
rect 148432 190117 148438 190129
rect 148490 190117 148496 190169
rect 42160 187675 42166 187727
rect 42218 187715 42224 187727
rect 42832 187715 42838 187727
rect 42218 187687 42838 187715
rect 42218 187675 42224 187687
rect 42832 187675 42838 187687
rect 42890 187675 42896 187727
rect 146800 187231 146806 187283
rect 146858 187271 146864 187283
rect 197296 187271 197302 187283
rect 146858 187243 197302 187271
rect 146858 187231 146864 187243
rect 197296 187231 197302 187243
rect 197354 187231 197360 187283
rect 146800 184345 146806 184397
rect 146858 184385 146864 184397
rect 194416 184385 194422 184397
rect 146858 184357 194422 184385
rect 146858 184345 146864 184357
rect 194416 184345 194422 184357
rect 194474 184345 194480 184397
rect 144496 181533 144502 181585
rect 144554 181573 144560 181585
rect 148528 181573 148534 181585
rect 144554 181545 148534 181573
rect 144554 181533 144560 181545
rect 148528 181533 148534 181545
rect 148586 181533 148592 181585
rect 144016 181459 144022 181511
rect 144074 181499 144080 181511
rect 188656 181499 188662 181511
rect 144074 181471 188662 181499
rect 144074 181459 144080 181471
rect 188656 181459 188662 181471
rect 188714 181459 188720 181511
rect 661072 179313 661078 179365
rect 661130 179353 661136 179365
rect 674416 179353 674422 179365
rect 661130 179325 674422 179353
rect 661130 179313 661136 179325
rect 674416 179313 674422 179325
rect 674474 179313 674480 179365
rect 666640 178795 666646 178847
rect 666698 178835 666704 178847
rect 674416 178835 674422 178847
rect 666698 178807 674422 178835
rect 666698 178795 666704 178807
rect 674416 178795 674422 178807
rect 674474 178795 674480 178847
rect 145264 178647 145270 178699
rect 145322 178687 145328 178699
rect 148624 178687 148630 178699
rect 145322 178659 148630 178687
rect 145322 178647 145328 178659
rect 148624 178647 148630 178659
rect 148682 178647 148688 178699
rect 655216 178647 655222 178699
rect 655274 178687 655280 178699
rect 674608 178687 674614 178699
rect 655274 178659 674614 178687
rect 655274 178647 655280 178659
rect 674608 178647 674614 178659
rect 674666 178647 674672 178699
rect 146800 178573 146806 178625
rect 146858 178613 146864 178625
rect 191536 178613 191542 178625
rect 146858 178585 191542 178613
rect 146858 178573 146864 178585
rect 191536 178573 191542 178585
rect 191594 178573 191600 178625
rect 146800 175835 146806 175887
rect 146858 175875 146864 175887
rect 148720 175875 148726 175887
rect 146858 175847 148726 175875
rect 146858 175835 146864 175847
rect 148720 175835 148726 175847
rect 148778 175835 148784 175887
rect 144112 175687 144118 175739
rect 144170 175727 144176 175739
rect 185776 175727 185782 175739
rect 144170 175699 185782 175727
rect 144170 175687 144176 175699
rect 185776 175687 185782 175699
rect 185834 175687 185840 175739
rect 144784 172801 144790 172853
rect 144842 172841 144848 172853
rect 162736 172841 162742 172853
rect 144842 172813 162742 172841
rect 144842 172801 144848 172813
rect 162736 172801 162742 172813
rect 162794 172801 162800 172853
rect 146800 169915 146806 169967
rect 146858 169955 146864 169967
rect 159856 169955 159862 169967
rect 146858 169927 159862 169955
rect 146858 169915 146864 169927
rect 159856 169915 159862 169927
rect 159914 169915 159920 169967
rect 206704 169841 206710 169893
rect 206762 169881 206768 169893
rect 206992 169881 206998 169893
rect 206762 169853 206998 169881
rect 206762 169841 206768 169853
rect 206992 169841 206998 169853
rect 207050 169841 207056 169893
rect 646864 167399 646870 167451
rect 646922 167439 646928 167451
rect 674704 167439 674710 167451
rect 646922 167411 674710 167439
rect 646922 167399 646928 167411
rect 674704 167399 674710 167411
rect 674762 167399 674768 167451
rect 646288 167177 646294 167229
rect 646346 167217 646352 167229
rect 674704 167217 674710 167229
rect 646346 167189 674710 167217
rect 646346 167177 646352 167189
rect 674704 167177 674710 167189
rect 674762 167177 674768 167229
rect 146800 167103 146806 167155
rect 146858 167143 146864 167155
rect 156976 167143 156982 167155
rect 146858 167115 156982 167143
rect 146858 167103 146864 167115
rect 156976 167103 156982 167115
rect 157034 167103 157040 167155
rect 647920 167103 647926 167155
rect 647978 167143 647984 167155
rect 674608 167143 674614 167155
rect 647978 167115 674614 167143
rect 647978 167103 647984 167115
rect 674608 167103 674614 167115
rect 674666 167103 674672 167155
rect 144784 167029 144790 167081
rect 144842 167069 144848 167081
rect 148816 167069 148822 167081
rect 144842 167041 148822 167069
rect 144842 167029 144848 167041
rect 148816 167029 148822 167041
rect 148874 167029 148880 167081
rect 144784 164143 144790 164195
rect 144842 164183 144848 164195
rect 148912 164183 148918 164195
rect 144842 164155 148918 164183
rect 144842 164143 144848 164155
rect 148912 164143 148918 164155
rect 148970 164143 148976 164195
rect 144976 162737 144982 162789
rect 145034 162777 145040 162789
rect 146704 162777 146710 162789
rect 145034 162749 146710 162777
rect 145034 162737 145040 162749
rect 146704 162737 146710 162749
rect 146762 162737 146768 162789
rect 144880 161257 144886 161309
rect 144938 161297 144944 161309
rect 149008 161297 149014 161309
rect 144938 161269 149014 161297
rect 144938 161257 144944 161269
rect 149008 161257 149014 161269
rect 149066 161257 149072 161309
rect 675472 160961 675478 161013
rect 675530 160961 675536 161013
rect 675490 160791 675518 160961
rect 675472 160739 675478 160791
rect 675530 160739 675536 160791
rect 675088 159555 675094 159607
rect 675146 159595 675152 159607
rect 675280 159595 675286 159607
rect 675146 159567 675286 159595
rect 675146 159555 675152 159567
rect 675280 159555 675286 159567
rect 675338 159555 675344 159607
rect 144880 158445 144886 158497
rect 144938 158485 144944 158497
rect 149104 158485 149110 158497
rect 144938 158457 149110 158485
rect 144938 158445 144944 158457
rect 149104 158445 149110 158457
rect 149162 158445 149168 158497
rect 144880 155559 144886 155611
rect 144938 155599 144944 155611
rect 200176 155599 200182 155611
rect 144938 155571 200182 155599
rect 144938 155559 144944 155571
rect 200176 155559 200182 155571
rect 200234 155559 200240 155611
rect 674032 153339 674038 153391
rect 674090 153379 674096 153391
rect 675472 153379 675478 153391
rect 674090 153351 675478 153379
rect 674090 153339 674096 153351
rect 675472 153339 675478 153351
rect 675530 153339 675536 153391
rect 144880 152747 144886 152799
rect 144938 152787 144944 152799
rect 180016 152787 180022 152799
rect 144938 152759 180022 152787
rect 144938 152747 144944 152759
rect 180016 152747 180022 152759
rect 180074 152747 180080 152799
rect 674224 152747 674230 152799
rect 674282 152787 674288 152799
rect 675376 152787 675382 152799
rect 674282 152759 675382 152787
rect 674282 152747 674288 152759
rect 675376 152747 675382 152759
rect 675434 152747 675440 152799
rect 144784 152673 144790 152725
rect 144842 152713 144848 152725
rect 182896 152713 182902 152725
rect 144842 152685 182902 152713
rect 144842 152673 144848 152685
rect 182896 152673 182902 152685
rect 182954 152673 182960 152725
rect 673936 152007 673942 152059
rect 673994 152047 674000 152059
rect 675472 152047 675478 152059
rect 673994 152019 675478 152047
rect 673994 152007 674000 152019
rect 675472 152007 675478 152019
rect 675530 152007 675536 152059
rect 674128 151489 674134 151541
rect 674186 151529 674192 151541
rect 675376 151529 675382 151541
rect 674186 151501 675382 151529
rect 674186 151489 674192 151501
rect 675376 151489 675382 151501
rect 675434 151489 675440 151541
rect 144880 149787 144886 149839
rect 144938 149827 144944 149839
rect 177136 149827 177142 149839
rect 144938 149799 177142 149827
rect 144938 149787 144944 149799
rect 177136 149787 177142 149799
rect 177194 149787 177200 149839
rect 144880 146901 144886 146953
rect 144938 146941 144944 146953
rect 174352 146941 174358 146953
rect 144938 146913 174358 146941
rect 144938 146901 144944 146913
rect 174352 146901 174358 146913
rect 174410 146901 174416 146953
rect 144496 146087 144502 146139
rect 144554 146127 144560 146139
rect 144880 146127 144886 146139
rect 144554 146099 144886 146127
rect 144554 146087 144560 146099
rect 144880 146087 144886 146099
rect 144938 146087 144944 146139
rect 146128 144607 146134 144659
rect 146186 144647 146192 144659
rect 146320 144647 146326 144659
rect 146186 144619 146326 144647
rect 146186 144607 146192 144619
rect 146320 144607 146326 144619
rect 146378 144607 146384 144659
rect 144304 144459 144310 144511
rect 144362 144499 144368 144511
rect 146128 144499 146134 144511
rect 144362 144471 146134 144499
rect 144362 144459 144368 144471
rect 146128 144459 146134 144471
rect 146186 144459 146192 144511
rect 144496 144311 144502 144363
rect 144554 144351 144560 144363
rect 154096 144351 154102 144363
rect 144554 144323 154102 144351
rect 144554 144311 144560 144323
rect 154096 144311 154102 144323
rect 154154 144311 154160 144363
rect 144304 144015 144310 144067
rect 144362 144055 144368 144067
rect 208720 144055 208726 144067
rect 144362 144027 208726 144055
rect 144362 144015 144368 144027
rect 208720 144015 208726 144027
rect 208778 144015 208784 144067
rect 144304 141647 144310 141699
rect 144362 141687 144368 141699
rect 171568 141687 171574 141699
rect 144362 141659 171574 141687
rect 144362 141647 144368 141659
rect 171568 141647 171574 141659
rect 171626 141647 171632 141699
rect 144304 141203 144310 141255
rect 144362 141243 144368 141255
rect 149200 141243 149206 141255
rect 144362 141215 149206 141243
rect 144362 141203 144368 141215
rect 149200 141203 149206 141215
rect 149258 141203 149264 141255
rect 645424 141203 645430 141255
rect 645482 141243 645488 141255
rect 645808 141243 645814 141255
rect 645482 141215 645814 141243
rect 645482 141203 645488 141215
rect 645808 141203 645814 141215
rect 645866 141203 645872 141255
rect 144496 141129 144502 141181
rect 144554 141169 144560 141181
rect 208816 141169 208822 141181
rect 144554 141141 208822 141169
rect 144554 141129 144560 141141
rect 208816 141129 208822 141141
rect 208874 141129 208880 141181
rect 645136 141055 645142 141107
rect 645194 141055 645200 141107
rect 645232 141055 645238 141107
rect 645290 141055 645296 141107
rect 645424 141055 645430 141107
rect 645482 141095 645488 141107
rect 645808 141095 645814 141107
rect 645482 141067 645814 141095
rect 645482 141055 645488 141067
rect 645808 141055 645814 141067
rect 645866 141055 645872 141107
rect 144496 140907 144502 140959
rect 144554 140947 144560 140959
rect 146320 140947 146326 140959
rect 144554 140919 146326 140947
rect 144554 140907 144560 140919
rect 146320 140907 146326 140919
rect 146378 140907 146384 140959
rect 645154 140589 645182 141055
rect 645250 140811 645278 141055
rect 645232 140759 645238 140811
rect 645290 140759 645296 140811
rect 645136 140537 645142 140589
rect 645194 140537 645200 140589
rect 144304 138243 144310 138295
rect 144362 138283 144368 138295
rect 168592 138283 168598 138295
rect 144362 138255 168598 138283
rect 144362 138243 144368 138255
rect 168592 138243 168598 138255
rect 168650 138243 168656 138295
rect 144880 137059 144886 137111
rect 144938 137099 144944 137111
rect 144938 137071 145022 137099
rect 144938 137059 144944 137071
rect 144688 136911 144694 136963
rect 144746 136951 144752 136963
rect 144880 136951 144886 136963
rect 144746 136923 144886 136951
rect 144746 136911 144752 136923
rect 144880 136911 144886 136923
rect 144938 136911 144944 136963
rect 144994 136877 145022 137071
rect 144802 136849 145022 136877
rect 144802 136741 144830 136849
rect 144784 136689 144790 136741
rect 144842 136689 144848 136741
rect 146896 135949 146902 136001
rect 146954 135989 146960 136001
rect 149296 135989 149302 136001
rect 146954 135961 149302 135989
rect 146954 135949 146960 135961
rect 149296 135949 149302 135961
rect 149354 135949 149360 136001
rect 144304 135431 144310 135483
rect 144362 135471 144368 135483
rect 144362 135443 148094 135471
rect 144362 135431 144368 135443
rect 148066 135397 148094 135443
rect 208912 135397 208918 135409
rect 148066 135369 208918 135397
rect 208912 135357 208918 135369
rect 208970 135357 208976 135409
rect 144496 134987 144502 135039
rect 144554 135027 144560 135039
rect 146896 135027 146902 135039
rect 144554 134999 146902 135027
rect 144554 134987 144560 134999
rect 146896 134987 146902 134999
rect 146954 134987 146960 135039
rect 663760 133581 663766 133633
rect 663818 133621 663824 133633
rect 674416 133621 674422 133633
rect 663818 133593 674422 133621
rect 663818 133581 663824 133593
rect 674416 133581 674422 133593
rect 674474 133581 674480 133633
rect 144304 132915 144310 132967
rect 144362 132955 144368 132967
rect 165712 132955 165718 132967
rect 144362 132927 165718 132955
rect 144362 132915 144368 132927
rect 165712 132915 165718 132927
rect 165770 132915 165776 132967
rect 655312 132767 655318 132819
rect 655370 132807 655376 132819
rect 676912 132807 676918 132819
rect 655370 132779 676918 132807
rect 655370 132767 655376 132779
rect 676912 132767 676918 132779
rect 676970 132767 676976 132819
rect 655120 132619 655126 132671
rect 655178 132659 655184 132671
rect 676816 132659 676822 132671
rect 655178 132631 676822 132659
rect 655178 132619 655184 132631
rect 676816 132619 676822 132631
rect 676874 132619 676880 132671
rect 144304 132545 144310 132597
rect 144362 132585 144368 132597
rect 209008 132585 209014 132597
rect 144362 132557 209014 132585
rect 144362 132545 144368 132557
rect 209008 132545 209014 132557
rect 209066 132545 209072 132597
rect 144496 132471 144502 132523
rect 144554 132511 144560 132523
rect 209104 132511 209110 132523
rect 144554 132483 209110 132511
rect 144554 132471 144560 132483
rect 209104 132471 209110 132483
rect 209162 132471 209168 132523
rect 647632 132471 647638 132523
rect 647690 132511 647696 132523
rect 674416 132511 674422 132523
rect 647690 132483 674422 132511
rect 647690 132471 647696 132483
rect 674416 132471 674422 132483
rect 674474 132471 674480 132523
rect 144496 129659 144502 129711
rect 144554 129699 144560 129711
rect 151408 129699 151414 129711
rect 144554 129671 151414 129699
rect 144554 129659 144560 129671
rect 151408 129659 151414 129671
rect 151466 129659 151472 129711
rect 144304 129585 144310 129637
rect 144362 129625 144368 129637
rect 208624 129625 208630 129637
rect 144362 129597 208630 129625
rect 144362 129585 144368 129597
rect 208624 129585 208630 129597
rect 208682 129585 208688 129637
rect 144496 129511 144502 129563
rect 144554 129551 144560 129563
rect 144880 129551 144886 129563
rect 144554 129523 144886 129551
rect 144554 129511 144560 129523
rect 144880 129511 144886 129523
rect 144938 129511 144944 129563
rect 144880 129363 144886 129415
rect 144938 129403 144944 129415
rect 146128 129403 146134 129415
rect 144938 129375 146134 129403
rect 144938 129363 144944 129375
rect 146128 129363 146134 129375
rect 146186 129363 146192 129415
rect 146128 128475 146134 128527
rect 146186 128515 146192 128527
rect 146512 128515 146518 128527
rect 146186 128487 146518 128515
rect 146186 128475 146192 128487
rect 146512 128475 146518 128487
rect 146570 128475 146576 128527
rect 144016 126995 144022 127047
rect 144074 126995 144080 127047
rect 144112 126995 144118 127047
rect 144170 126995 144176 127047
rect 144208 126995 144214 127047
rect 144266 126995 144272 127047
rect 144034 126825 144062 126995
rect 144130 126825 144158 126995
rect 144226 126825 144254 126995
rect 144304 126921 144310 126973
rect 144362 126961 144368 126973
rect 144362 126933 146846 126961
rect 144362 126921 144368 126933
rect 144016 126773 144022 126825
rect 144074 126773 144080 126825
rect 144112 126773 144118 126825
rect 144170 126773 144176 126825
rect 144208 126773 144214 126825
rect 144266 126773 144272 126825
rect 146320 126773 146326 126825
rect 146378 126773 146384 126825
rect 146818 126813 146846 126933
rect 146992 126847 146998 126899
rect 147050 126887 147056 126899
rect 149392 126887 149398 126899
rect 147050 126859 149398 126887
rect 147050 126847 147056 126859
rect 149392 126847 149398 126859
rect 149450 126847 149456 126899
rect 203152 126813 203158 126825
rect 146818 126785 203158 126813
rect 203152 126773 203158 126785
rect 203210 126773 203216 126825
rect 143920 126699 143926 126751
rect 143978 126739 143984 126751
rect 146338 126739 146366 126773
rect 143978 126711 146366 126739
rect 143978 126699 143984 126711
rect 146512 126699 146518 126751
rect 146570 126739 146576 126751
rect 208528 126739 208534 126751
rect 146570 126711 208534 126739
rect 146570 126699 146576 126711
rect 208528 126699 208534 126711
rect 208586 126699 208592 126751
rect 145072 126625 145078 126677
rect 145130 126665 145136 126677
rect 146320 126665 146326 126677
rect 145130 126637 146326 126665
rect 145130 126625 145136 126637
rect 146320 126625 146326 126637
rect 146378 126625 146384 126677
rect 645520 126625 645526 126677
rect 645578 126665 645584 126677
rect 645808 126665 645814 126677
rect 645578 126637 645814 126665
rect 645578 126625 645584 126637
rect 645808 126625 645814 126637
rect 645866 126625 645872 126677
rect 143920 126477 143926 126529
rect 143978 126517 143984 126529
rect 145072 126517 145078 126529
rect 143978 126489 145078 126517
rect 143978 126477 143984 126489
rect 145072 126477 145078 126489
rect 145130 126477 145136 126529
rect 144592 125367 144598 125419
rect 144650 125407 144656 125419
rect 146512 125407 146518 125419
rect 144650 125379 146518 125407
rect 144650 125367 144656 125379
rect 146512 125367 146518 125379
rect 146570 125367 146576 125419
rect 39856 125293 39862 125345
rect 39914 125333 39920 125345
rect 42928 125333 42934 125345
rect 39914 125305 42934 125333
rect 39914 125293 39920 125305
rect 42928 125293 42934 125305
rect 42986 125293 42992 125345
rect 144400 125219 144406 125271
rect 144458 125259 144464 125271
rect 144592 125259 144598 125271
rect 144458 125231 144598 125259
rect 144458 125219 144464 125231
rect 144592 125219 144598 125231
rect 144650 125219 144656 125271
rect 146320 124997 146326 125049
rect 146378 125037 146384 125049
rect 146378 125009 146462 125037
rect 146378 124997 146384 125009
rect 146128 124849 146134 124901
rect 146186 124889 146192 124901
rect 146320 124889 146326 124901
rect 146186 124861 146326 124889
rect 146186 124849 146192 124861
rect 146320 124849 146326 124861
rect 146378 124849 146384 124901
rect 146128 124701 146134 124753
rect 146186 124741 146192 124753
rect 146434 124741 146462 125009
rect 146186 124713 146462 124741
rect 146186 124701 146192 124713
rect 144304 123961 144310 124013
rect 144362 124001 144368 124013
rect 197392 124001 197398 124013
rect 144362 123973 197398 124001
rect 144362 123961 144368 123973
rect 197392 123961 197398 123973
rect 197450 123961 197456 124013
rect 144400 123887 144406 123939
rect 144458 123927 144464 123939
rect 200272 123927 200278 123939
rect 144458 123899 200278 123927
rect 144458 123887 144464 123899
rect 200272 123887 200278 123899
rect 200330 123887 200336 123939
rect 645808 121223 645814 121275
rect 645866 121263 645872 121275
rect 676816 121263 676822 121275
rect 645866 121235 676822 121263
rect 645866 121223 645872 121235
rect 676816 121223 676822 121235
rect 676874 121223 676880 121275
rect 645904 121149 645910 121201
rect 645962 121189 645968 121201
rect 674704 121189 674710 121201
rect 645962 121161 674710 121189
rect 645962 121149 645968 121161
rect 674704 121149 674710 121161
rect 674762 121149 674768 121201
rect 144400 121075 144406 121127
rect 144458 121115 144464 121127
rect 149488 121115 149494 121127
rect 144458 121087 149494 121115
rect 144458 121075 144464 121087
rect 149488 121075 149494 121087
rect 149546 121075 149552 121127
rect 646000 121075 646006 121127
rect 646058 121115 646064 121127
rect 676912 121115 676918 121127
rect 646058 121087 676918 121115
rect 646058 121075 646064 121087
rect 676912 121075 676918 121087
rect 676970 121075 676976 121127
rect 144304 121001 144310 121053
rect 144362 121041 144368 121053
rect 149584 121041 149590 121053
rect 144362 121013 149590 121041
rect 144362 121001 144368 121013
rect 149584 121001 149590 121013
rect 149642 121001 149648 121053
rect 144400 120927 144406 120979
rect 144458 120967 144464 120979
rect 144592 120967 144598 120979
rect 144458 120939 144598 120967
rect 144458 120927 144464 120939
rect 144592 120927 144598 120939
rect 144650 120927 144656 120979
rect 207088 120927 207094 120979
rect 207146 120967 207152 120979
rect 207184 120967 207190 120979
rect 207146 120939 207190 120967
rect 207146 120927 207152 120939
rect 207184 120927 207190 120939
rect 207242 120927 207248 120979
rect 144304 118411 144310 118463
rect 144362 118411 144368 118463
rect 144322 118303 144350 118411
rect 144226 118275 144350 118303
rect 144226 118155 144254 118275
rect 144400 118263 144406 118315
rect 144458 118303 144464 118315
rect 171472 118303 171478 118315
rect 144458 118275 171478 118303
rect 144458 118263 144464 118275
rect 171472 118263 171478 118275
rect 171530 118263 171536 118315
rect 144304 118189 144310 118241
rect 144362 118229 144368 118241
rect 188752 118229 188758 118241
rect 144362 118201 188758 118229
rect 144362 118189 144368 118201
rect 188752 118189 188758 118201
rect 188810 118189 188816 118241
rect 144226 118127 144542 118155
rect 144514 118007 144542 118127
rect 144592 118115 144598 118167
rect 144650 118155 144656 118167
rect 194512 118155 194518 118167
rect 144650 118127 194518 118155
rect 144650 118115 144656 118127
rect 194512 118115 194518 118127
rect 194570 118115 194576 118167
rect 144592 118007 144598 118019
rect 144514 117979 144598 118007
rect 144592 117967 144598 117979
rect 144650 117967 144656 118019
rect 144304 116191 144310 116243
rect 144362 116231 144368 116243
rect 149680 116231 149686 116243
rect 144362 116203 149686 116231
rect 144362 116191 144368 116203
rect 149680 116191 149686 116203
rect 149738 116191 149744 116243
rect 144304 115525 144310 115577
rect 144362 115565 144368 115577
rect 148144 115565 148150 115577
rect 144362 115537 148150 115565
rect 144362 115525 144368 115537
rect 148144 115525 148150 115537
rect 148202 115525 148208 115577
rect 144304 115377 144310 115429
rect 144362 115417 144368 115429
rect 146128 115417 146134 115429
rect 144362 115389 146134 115417
rect 144362 115377 144368 115389
rect 146128 115377 146134 115389
rect 146186 115377 146192 115429
rect 146128 115007 146134 115059
rect 146186 115047 146192 115059
rect 146896 115047 146902 115059
rect 146186 115019 146902 115047
rect 146186 115007 146192 115019
rect 146896 115007 146902 115019
rect 146954 115007 146960 115059
rect 674512 114119 674518 114171
rect 674570 114159 674576 114171
rect 675376 114159 675382 114171
rect 674570 114131 675382 114159
rect 674570 114119 674576 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 674320 113601 674326 113653
rect 674378 113641 674384 113653
rect 675088 113641 675094 113653
rect 674378 113613 675094 113641
rect 674378 113601 674384 113613
rect 675088 113601 675094 113613
rect 675146 113601 675152 113653
rect 144304 112639 144310 112691
rect 144362 112679 144368 112691
rect 147952 112679 147958 112691
rect 144362 112651 147958 112679
rect 144362 112639 144368 112651
rect 147952 112639 147958 112651
rect 148010 112639 148016 112691
rect 144304 112417 144310 112469
rect 144362 112457 144368 112469
rect 148048 112457 148054 112469
rect 144362 112429 148054 112457
rect 144362 112417 144368 112429
rect 148048 112417 148054 112429
rect 148106 112417 148112 112469
rect 144400 112343 144406 112395
rect 144458 112383 144464 112395
rect 191632 112383 191638 112395
rect 144458 112355 191638 112383
rect 144458 112343 144464 112355
rect 191632 112343 191638 112355
rect 191690 112343 191696 112395
rect 674224 111825 674230 111877
rect 674282 111865 674288 111877
rect 675088 111865 675094 111877
rect 674282 111837 675094 111865
rect 674282 111825 674288 111837
rect 675088 111825 675094 111837
rect 675146 111825 675152 111877
rect 674704 111307 674710 111359
rect 674762 111347 674768 111359
rect 675376 111347 675382 111359
rect 674762 111319 675382 111347
rect 674762 111307 674768 111319
rect 675376 111307 675382 111319
rect 675434 111307 675440 111359
rect 674800 111233 674806 111285
rect 674858 111273 674864 111285
rect 675088 111273 675094 111285
rect 674858 111245 675094 111273
rect 674858 111233 674864 111245
rect 675088 111233 675094 111245
rect 675146 111233 675152 111285
rect 144400 109531 144406 109583
rect 144458 109571 144464 109583
rect 147856 109571 147862 109583
rect 144458 109543 147862 109571
rect 144458 109531 144464 109543
rect 147856 109531 147862 109543
rect 147914 109531 147920 109583
rect 144304 109457 144310 109509
rect 144362 109497 144368 109509
rect 185872 109497 185878 109509
rect 144362 109469 185878 109497
rect 144362 109457 144368 109469
rect 185872 109457 185878 109469
rect 185930 109457 185936 109509
rect 144400 109383 144406 109435
rect 144458 109423 144464 109435
rect 144592 109423 144598 109435
rect 144458 109395 144598 109423
rect 144458 109383 144464 109395
rect 144592 109383 144598 109395
rect 144650 109383 144656 109435
rect 674896 107533 674902 107585
rect 674954 107573 674960 107585
rect 675376 107573 675382 107585
rect 674954 107545 675382 107573
rect 674954 107533 674960 107545
rect 675376 107533 675382 107545
rect 675434 107533 675440 107585
rect 143824 106941 143830 106993
rect 143882 106981 143888 106993
rect 144400 106981 144406 106993
rect 143882 106953 144406 106981
rect 143882 106941 143888 106953
rect 144400 106941 144406 106953
rect 144458 106941 144464 106993
rect 144304 106867 144310 106919
rect 144362 106907 144368 106919
rect 162832 106907 162838 106919
rect 144362 106879 162838 106907
rect 144362 106867 144368 106879
rect 162832 106867 162838 106879
rect 162890 106867 162896 106919
rect 673936 106867 673942 106919
rect 673994 106907 674000 106919
rect 675472 106907 675478 106919
rect 673994 106879 675478 106907
rect 673994 106867 674000 106879
rect 675472 106867 675478 106879
rect 675530 106867 675536 106919
rect 143920 106793 143926 106845
rect 143978 106833 143984 106845
rect 146512 106833 146518 106845
rect 143978 106805 146518 106833
rect 143978 106793 143984 106805
rect 146512 106793 146518 106805
rect 146570 106793 146576 106845
rect 144304 106719 144310 106771
rect 144362 106759 144368 106771
rect 145072 106759 145078 106771
rect 144362 106731 145078 106759
rect 144362 106719 144368 106731
rect 145072 106719 145078 106731
rect 145130 106719 145136 106771
rect 144592 106571 144598 106623
rect 144650 106611 144656 106623
rect 147760 106611 147766 106623
rect 144650 106583 147766 106611
rect 144650 106571 144656 106583
rect 147760 106571 147766 106583
rect 147818 106571 147824 106623
rect 645520 106497 645526 106549
rect 645578 106537 645584 106549
rect 645904 106537 645910 106549
rect 645578 106509 645910 106537
rect 645578 106497 645584 106509
rect 645904 106497 645910 106509
rect 645962 106497 645968 106549
rect 668176 106497 668182 106549
rect 668234 106537 668240 106549
rect 675088 106537 675094 106549
rect 668234 106509 675094 106537
rect 668234 106497 668240 106509
rect 675088 106497 675094 106509
rect 675146 106497 675152 106549
rect 143920 106423 143926 106475
rect 143978 106463 143984 106475
rect 144592 106463 144598 106475
rect 143978 106435 144598 106463
rect 143978 106423 143984 106435
rect 144592 106423 144598 106435
rect 144650 106423 144656 106475
rect 146512 106423 146518 106475
rect 146570 106463 146576 106475
rect 159952 106463 159958 106475
rect 146570 106435 159958 106463
rect 146570 106423 146576 106435
rect 159952 106423 159958 106435
rect 160010 106423 160016 106475
rect 674416 106349 674422 106401
rect 674474 106389 674480 106401
rect 675376 106389 675382 106401
rect 674474 106361 675382 106389
rect 674474 106349 674480 106361
rect 675376 106349 675382 106361
rect 675434 106349 675440 106401
rect 146320 104795 146326 104847
rect 146378 104835 146384 104847
rect 146896 104835 146902 104847
rect 146378 104807 146902 104835
rect 146378 104795 146384 104807
rect 146896 104795 146902 104807
rect 146954 104795 146960 104847
rect 645424 104499 645430 104551
rect 645482 104539 645488 104551
rect 665200 104539 665206 104551
rect 645482 104511 665206 104539
rect 645482 104499 645488 104511
rect 665200 104499 665206 104511
rect 665258 104499 665264 104551
rect 659536 104425 659542 104477
rect 659594 104465 659600 104477
rect 665296 104465 665302 104477
rect 659594 104437 665302 104465
rect 659594 104425 659600 104437
rect 665296 104425 665302 104437
rect 665354 104425 665360 104477
rect 146512 104351 146518 104403
rect 146570 104391 146576 104403
rect 160048 104391 160054 104403
rect 146570 104363 160054 104391
rect 146570 104351 146576 104363
rect 160048 104351 160054 104363
rect 160106 104351 160112 104403
rect 146320 103685 146326 103737
rect 146378 103725 146384 103737
rect 208432 103725 208438 103737
rect 146378 103697 208438 103725
rect 146378 103685 146384 103697
rect 208432 103685 208438 103697
rect 208490 103685 208496 103737
rect 146128 103611 146134 103663
rect 146186 103651 146192 103663
rect 204592 103651 204598 103663
rect 146186 103623 204598 103651
rect 146186 103611 146192 103623
rect 204592 103611 204598 103623
rect 204650 103611 204656 103663
rect 145072 103537 145078 103589
rect 145130 103577 145136 103589
rect 204688 103577 204694 103589
rect 145130 103549 204694 103577
rect 145130 103537 145136 103549
rect 204688 103537 204694 103549
rect 204746 103537 204752 103589
rect 146896 103463 146902 103515
rect 146954 103503 146960 103515
rect 204496 103503 204502 103515
rect 146954 103475 204502 103503
rect 146954 103463 146960 103475
rect 204496 103463 204502 103475
rect 204554 103463 204560 103515
rect 143824 103389 143830 103441
rect 143882 103429 143888 103441
rect 145072 103429 145078 103441
rect 143882 103401 145078 103429
rect 143882 103389 143888 103401
rect 145072 103389 145078 103401
rect 145130 103389 145136 103441
rect 146512 101539 146518 101591
rect 146570 101579 146576 101591
rect 157072 101579 157078 101591
rect 146570 101551 157078 101579
rect 146570 101539 146576 101551
rect 157072 101539 157078 101551
rect 157130 101539 157136 101591
rect 146320 100799 146326 100851
rect 146378 100839 146384 100851
rect 151312 100839 151318 100851
rect 146378 100811 151318 100839
rect 146378 100799 146384 100811
rect 151312 100799 151318 100811
rect 151370 100799 151376 100851
rect 145072 100725 145078 100777
rect 145130 100765 145136 100777
rect 194704 100765 194710 100777
rect 145130 100737 194710 100765
rect 145130 100725 145136 100737
rect 194704 100725 194710 100737
rect 194762 100725 194768 100777
rect 144400 100651 144406 100703
rect 144458 100691 144464 100703
rect 201712 100691 201718 100703
rect 144458 100663 201718 100691
rect 144458 100651 144464 100663
rect 201712 100651 201718 100663
rect 201770 100651 201776 100703
rect 144592 100577 144598 100629
rect 144650 100617 144656 100629
rect 204592 100617 204598 100629
rect 144650 100589 204598 100617
rect 144650 100577 144656 100589
rect 204592 100577 204598 100589
rect 204650 100577 204656 100629
rect 151120 100503 151126 100555
rect 151178 100543 151184 100555
rect 198352 100543 198358 100555
rect 151178 100515 198358 100543
rect 151178 100503 151184 100515
rect 198352 100503 198358 100515
rect 198410 100503 198416 100555
rect 159760 100429 159766 100481
rect 159818 100469 159824 100481
rect 210160 100469 210166 100481
rect 159818 100441 210166 100469
rect 159818 100429 159824 100441
rect 210160 100429 210166 100441
rect 210218 100429 210224 100481
rect 146512 98061 146518 98113
rect 146570 98101 146576 98113
rect 180112 98101 180118 98113
rect 146570 98073 180118 98101
rect 146570 98061 146576 98073
rect 180112 98061 180118 98073
rect 180170 98061 180176 98113
rect 146320 97987 146326 98039
rect 146378 98027 146384 98039
rect 182992 98027 182998 98039
rect 146378 97999 182998 98027
rect 146378 97987 146384 97999
rect 182992 97987 182998 97999
rect 183050 97987 183056 98039
rect 146128 97913 146134 97965
rect 146186 97953 146192 97965
rect 208336 97953 208342 97965
rect 146186 97925 208342 97953
rect 146186 97913 146192 97925
rect 208336 97913 208342 97925
rect 208394 97913 208400 97965
rect 154000 97839 154006 97891
rect 154058 97879 154064 97891
rect 200752 97879 200758 97891
rect 154058 97851 200758 97879
rect 154058 97839 154064 97851
rect 200752 97839 200758 97851
rect 200810 97839 200816 97891
rect 156880 97765 156886 97817
rect 156938 97805 156944 97817
rect 200560 97805 200566 97817
rect 156938 97777 200566 97805
rect 156938 97765 156944 97777
rect 200560 97765 200566 97777
rect 200618 97765 200624 97817
rect 171376 97691 171382 97743
rect 171434 97731 171440 97743
rect 201712 97731 201718 97743
rect 171434 97703 201718 97731
rect 171434 97691 171440 97703
rect 201712 97691 201718 97703
rect 201770 97691 201776 97743
rect 174256 97617 174262 97669
rect 174314 97657 174320 97669
rect 210160 97657 210166 97669
rect 174314 97629 210166 97657
rect 174314 97617 174320 97629
rect 210160 97617 210166 97629
rect 210218 97617 210224 97669
rect 182800 97543 182806 97595
rect 182858 97583 182864 97595
rect 201040 97583 201046 97595
rect 182858 97555 201046 97583
rect 182858 97543 182864 97555
rect 201040 97543 201046 97555
rect 201098 97543 201104 97595
rect 146512 95101 146518 95153
rect 146570 95141 146576 95153
rect 174448 95141 174454 95153
rect 146570 95113 174454 95141
rect 146570 95101 146576 95113
rect 174448 95101 174454 95113
rect 174506 95101 174512 95153
rect 146320 95027 146326 95079
rect 146378 95067 146384 95079
rect 177232 95067 177238 95079
rect 146378 95039 177238 95067
rect 146378 95027 146384 95039
rect 177232 95027 177238 95039
rect 177290 95027 177296 95079
rect 144208 94879 144214 94931
rect 144266 94919 144272 94931
rect 201616 94919 201622 94931
rect 144266 94891 201622 94919
rect 144266 94879 144272 94891
rect 201616 94879 201622 94891
rect 201674 94879 201680 94931
rect 151216 94805 151222 94857
rect 151274 94845 151280 94857
rect 195472 94845 195478 94857
rect 151274 94817 195478 94845
rect 151274 94805 151280 94817
rect 195472 94805 195478 94817
rect 195530 94805 195536 94857
rect 165616 94731 165622 94783
rect 165674 94771 165680 94783
rect 201712 94771 201718 94783
rect 165674 94743 201718 94771
rect 165674 94731 165680 94743
rect 201712 94731 201718 94743
rect 201770 94731 201776 94783
rect 168496 94657 168502 94709
rect 168554 94697 168560 94709
rect 210160 94697 210166 94709
rect 168554 94669 210166 94697
rect 168554 94657 168560 94669
rect 210160 94657 210166 94669
rect 210218 94657 210224 94709
rect 144016 94583 144022 94635
rect 144074 94623 144080 94635
rect 194800 94623 194806 94635
rect 144074 94595 194806 94623
rect 144074 94583 144080 94595
rect 194800 94583 194806 94595
rect 194858 94583 194864 94635
rect 651280 93695 651286 93747
rect 651338 93735 651344 93747
rect 659536 93735 659542 93747
rect 651338 93707 659542 93735
rect 651338 93695 651344 93707
rect 659536 93695 659542 93707
rect 659594 93695 659600 93747
rect 646384 92659 646390 92711
rect 646442 92699 646448 92711
rect 659824 92699 659830 92711
rect 646442 92671 659830 92699
rect 646442 92659 646448 92671
rect 659824 92659 659830 92671
rect 659882 92659 659888 92711
rect 647440 92585 647446 92637
rect 647498 92625 647504 92637
rect 661744 92625 661750 92637
rect 647498 92597 661750 92625
rect 647498 92585 647504 92597
rect 661744 92585 661750 92597
rect 661802 92585 661808 92637
rect 646192 92511 646198 92563
rect 646250 92551 646256 92563
rect 660688 92551 660694 92563
rect 646250 92523 660694 92551
rect 646250 92511 646256 92523
rect 660688 92511 660694 92523
rect 660746 92511 660752 92563
rect 647824 92363 647830 92415
rect 647882 92403 647888 92415
rect 663088 92403 663094 92415
rect 647882 92375 663094 92403
rect 647882 92363 647888 92375
rect 663088 92363 663094 92375
rect 663146 92363 663152 92415
rect 647248 92289 647254 92341
rect 647306 92329 647312 92341
rect 661168 92329 661174 92341
rect 647306 92301 661174 92329
rect 647306 92289 647312 92301
rect 661168 92289 661174 92301
rect 661226 92289 661232 92341
rect 146320 92215 146326 92267
rect 146378 92255 146384 92267
rect 154000 92255 154006 92267
rect 146378 92227 154006 92255
rect 146378 92215 146384 92227
rect 154000 92215 154006 92227
rect 154058 92215 154064 92267
rect 647728 92215 647734 92267
rect 647786 92255 647792 92267
rect 662512 92255 662518 92267
rect 647786 92227 662518 92255
rect 647786 92215 647792 92227
rect 662512 92215 662518 92227
rect 662570 92215 662576 92267
rect 146512 92141 146518 92193
rect 146570 92181 146576 92193
rect 171376 92181 171382 92193
rect 146570 92153 171382 92181
rect 146570 92141 146576 92153
rect 171376 92141 171382 92153
rect 171434 92141 171440 92193
rect 646672 92141 646678 92193
rect 646730 92181 646736 92193
rect 658864 92181 658870 92193
rect 646730 92153 658870 92181
rect 646730 92141 646736 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 144112 92067 144118 92119
rect 144170 92107 144176 92119
rect 210160 92107 210166 92119
rect 144170 92079 210166 92107
rect 144170 92067 144176 92079
rect 210160 92067 210166 92079
rect 210218 92067 210224 92119
rect 188656 91771 188662 91823
rect 188714 91811 188720 91823
rect 201712 91811 201718 91823
rect 188714 91783 201718 91811
rect 188714 91771 188720 91783
rect 201712 91771 201718 91783
rect 201770 91771 201776 91823
rect 146128 89403 146134 89455
rect 146186 89443 146192 89455
rect 151120 89443 151126 89455
rect 146186 89415 151126 89443
rect 146186 89403 146192 89415
rect 151120 89403 151126 89415
rect 151178 89403 151184 89455
rect 146512 89329 146518 89381
rect 146570 89369 146576 89381
rect 165616 89369 165622 89381
rect 146570 89341 165622 89369
rect 146570 89329 146576 89341
rect 165616 89329 165622 89341
rect 165674 89329 165680 89381
rect 146320 89255 146326 89307
rect 146378 89295 146384 89307
rect 168496 89295 168502 89307
rect 146378 89267 168502 89295
rect 146378 89255 146384 89267
rect 168496 89255 168502 89267
rect 168554 89255 168560 89307
rect 156976 89181 156982 89233
rect 157034 89221 157040 89233
rect 197872 89221 197878 89233
rect 157034 89193 197878 89221
rect 157034 89181 157040 89193
rect 197872 89181 197878 89193
rect 197930 89181 197936 89233
rect 159856 89107 159862 89159
rect 159914 89147 159920 89159
rect 201808 89147 201814 89159
rect 159914 89119 201814 89147
rect 159914 89107 159920 89119
rect 201808 89107 201814 89119
rect 201866 89107 201872 89159
rect 162736 89033 162742 89085
rect 162794 89073 162800 89085
rect 201616 89073 201622 89085
rect 162794 89045 201622 89073
rect 162794 89033 162800 89045
rect 201616 89033 201622 89045
rect 201674 89033 201680 89085
rect 185776 88959 185782 89011
rect 185834 88999 185840 89011
rect 201328 88999 201334 89011
rect 185834 88971 201334 88999
rect 185834 88959 185840 88971
rect 201328 88959 201334 88971
rect 201386 88959 201392 89011
rect 191536 88885 191542 88937
rect 191594 88925 191600 88937
rect 201712 88925 201718 88937
rect 191594 88897 201718 88925
rect 191594 88885 191600 88897
rect 201712 88885 201718 88897
rect 201770 88885 201776 88937
rect 650608 87331 650614 87383
rect 650666 87371 650672 87383
rect 659344 87371 659350 87383
rect 650666 87343 659350 87371
rect 650666 87331 650672 87343
rect 659344 87331 659350 87343
rect 659402 87331 659408 87383
rect 658000 87297 658006 87309
rect 657058 87269 658006 87297
rect 657058 87161 657086 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 657040 87109 657046 87161
rect 657098 87109 657104 87161
rect 645424 87035 645430 87087
rect 645482 87075 645488 87087
rect 663280 87075 663286 87087
rect 645482 87047 663286 87075
rect 645482 87035 645488 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 645808 86961 645814 87013
rect 645866 87001 645872 87013
rect 650992 87001 650998 87013
rect 645866 86973 650998 87001
rect 645866 86961 645872 86973
rect 650992 86961 650998 86973
rect 651050 86961 651056 87013
rect 645424 86887 645430 86939
rect 645482 86927 645488 86939
rect 645904 86927 645910 86939
rect 645482 86899 645910 86927
rect 645482 86887 645488 86899
rect 645904 86887 645910 86899
rect 645962 86887 645968 86939
rect 645808 86443 645814 86495
rect 645866 86483 645872 86495
rect 651088 86483 651094 86495
rect 645866 86455 651094 86483
rect 645866 86443 645872 86455
rect 651088 86443 651094 86455
rect 651146 86443 651152 86495
rect 154096 86369 154102 86421
rect 154154 86409 154160 86421
rect 196048 86409 196054 86421
rect 154154 86381 196054 86409
rect 154154 86369 154160 86381
rect 196048 86369 196054 86381
rect 196106 86369 196112 86421
rect 645424 86369 645430 86421
rect 645482 86409 645488 86421
rect 646096 86409 646102 86421
rect 645482 86381 646102 86409
rect 645482 86369 645488 86381
rect 646096 86369 646102 86381
rect 646154 86369 646160 86421
rect 174352 86295 174358 86347
rect 174410 86335 174416 86347
rect 201808 86335 201814 86347
rect 174410 86307 201814 86335
rect 174410 86295 174416 86307
rect 201808 86295 201814 86307
rect 201866 86295 201872 86347
rect 177136 86221 177142 86273
rect 177194 86261 177200 86273
rect 198736 86261 198742 86273
rect 177194 86233 198742 86261
rect 177194 86221 177200 86233
rect 198736 86221 198742 86233
rect 198794 86221 198800 86273
rect 180016 86147 180022 86199
rect 180074 86187 180080 86199
rect 201712 86187 201718 86199
rect 180074 86159 201718 86187
rect 180074 86147 180080 86159
rect 201712 86147 201718 86159
rect 201770 86147 201776 86199
rect 182896 86073 182902 86125
rect 182954 86113 182960 86125
rect 201616 86113 201622 86125
rect 182954 86085 201622 86113
rect 182954 86073 182960 86085
rect 201616 86073 201622 86085
rect 201674 86073 201680 86125
rect 645424 85185 645430 85237
rect 645482 85225 645488 85237
rect 650896 85225 650902 85237
rect 645482 85197 650902 85225
rect 645482 85185 645488 85197
rect 650896 85185 650902 85197
rect 650954 85185 650960 85237
rect 146512 84963 146518 85015
rect 146570 85003 146576 85015
rect 197776 85003 197782 85015
rect 146570 84975 197782 85003
rect 146570 84963 146576 84975
rect 197776 84963 197782 84975
rect 197834 84963 197840 85015
rect 151408 83483 151414 83535
rect 151466 83523 151472 83535
rect 201520 83523 201526 83535
rect 151466 83495 201526 83523
rect 151466 83483 151472 83495
rect 201520 83483 201526 83495
rect 201578 83483 201584 83535
rect 165712 83409 165718 83461
rect 165770 83449 165776 83461
rect 201808 83449 201814 83461
rect 165770 83421 201814 83449
rect 165770 83409 165776 83421
rect 201808 83409 201814 83421
rect 201866 83409 201872 83461
rect 645424 83409 645430 83461
rect 645482 83449 645488 83461
rect 657040 83449 657046 83461
rect 645482 83421 657046 83449
rect 645482 83409 645488 83421
rect 657040 83409 657046 83421
rect 657098 83409 657104 83461
rect 168592 83335 168598 83387
rect 168650 83375 168656 83387
rect 201616 83375 201622 83387
rect 168650 83347 201622 83375
rect 168650 83335 168656 83347
rect 201616 83335 201622 83347
rect 201674 83335 201680 83387
rect 171568 83261 171574 83313
rect 171626 83301 171632 83313
rect 201712 83301 201718 83313
rect 171626 83273 201718 83301
rect 171626 83261 171632 83273
rect 201712 83261 201718 83273
rect 201770 83261 201776 83313
rect 146512 82077 146518 82129
rect 146570 82117 146576 82129
rect 201712 82117 201718 82129
rect 146570 82089 201718 82117
rect 146570 82077 146576 82089
rect 201712 82077 201718 82089
rect 201770 82077 201776 82129
rect 645424 81855 645430 81907
rect 645482 81895 645488 81907
rect 663280 81895 663286 81907
rect 645482 81867 663286 81895
rect 645482 81855 645488 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 645808 81781 645814 81833
rect 645866 81821 645872 81833
rect 663376 81821 663382 81833
rect 645866 81793 663382 81821
rect 645866 81781 645872 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 647536 81633 647542 81685
rect 647594 81673 647600 81685
rect 661072 81673 661078 81685
rect 647594 81645 661078 81673
rect 647594 81633 647600 81645
rect 661072 81633 661078 81645
rect 661130 81633 661136 81685
rect 645424 81263 645430 81315
rect 645482 81303 645488 81315
rect 657520 81303 657526 81315
rect 645482 81275 657526 81303
rect 645482 81263 645488 81275
rect 657520 81263 657526 81275
rect 657578 81263 657584 81315
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 188752 80301 188758 80353
rect 188810 80341 188816 80353
rect 210160 80341 210166 80353
rect 188810 80313 210166 80341
rect 188810 80301 188816 80313
rect 210160 80301 210166 80313
rect 210218 80301 210224 80353
rect 645424 80153 645430 80205
rect 645482 80193 645488 80205
rect 656944 80193 656950 80205
rect 645482 80165 656950 80193
rect 645482 80153 645488 80165
rect 656944 80153 656950 80165
rect 657002 80153 657008 80205
rect 645904 79043 645910 79095
rect 645962 79083 645968 79095
rect 651184 79083 651190 79095
rect 645962 79055 651190 79083
rect 645962 79043 645968 79055
rect 651184 79043 651190 79055
rect 651242 79043 651248 79095
rect 645424 78895 645430 78947
rect 645482 78935 645488 78947
rect 658864 78935 658870 78947
rect 645482 78907 658870 78935
rect 645482 78895 645488 78907
rect 658864 78895 658870 78907
rect 658922 78895 658928 78947
rect 645808 78377 645814 78429
rect 645866 78417 645872 78429
rect 662512 78417 662518 78429
rect 645866 78389 662518 78417
rect 645866 78377 645872 78389
rect 662512 78377 662518 78389
rect 662570 78377 662576 78429
rect 646000 78007 646006 78059
rect 646058 78047 646064 78059
rect 660688 78047 660694 78059
rect 646058 78019 660694 78047
rect 646058 78007 646064 78019
rect 660688 78007 660694 78019
rect 660746 78007 660752 78059
rect 146320 77859 146326 77911
rect 146378 77899 146384 77911
rect 190000 77899 190006 77911
rect 146378 77871 190006 77899
rect 146378 77859 146384 77871
rect 190000 77859 190006 77871
rect 190058 77859 190064 77911
rect 146512 77785 146518 77837
rect 146570 77825 146576 77837
rect 208240 77825 208246 77837
rect 146570 77797 208246 77825
rect 146570 77785 146576 77797
rect 208240 77785 208246 77797
rect 208298 77785 208304 77837
rect 157072 77711 157078 77763
rect 157130 77751 157136 77763
rect 196912 77751 196918 77763
rect 157130 77723 196918 77751
rect 157130 77711 157136 77723
rect 196912 77711 196918 77723
rect 196970 77711 196976 77763
rect 647632 77711 647638 77763
rect 647690 77751 647696 77763
rect 659440 77751 659446 77763
rect 647690 77723 659446 77751
rect 647690 77711 647696 77723
rect 659440 77711 659446 77723
rect 659498 77711 659504 77763
rect 160048 77637 160054 77689
rect 160106 77677 160112 77689
rect 201616 77677 201622 77689
rect 160106 77649 201622 77677
rect 160106 77637 160112 77649
rect 201616 77637 201622 77649
rect 201674 77637 201680 77689
rect 645424 77637 645430 77689
rect 645482 77677 645488 77689
rect 650992 77677 650998 77689
rect 645482 77649 650998 77677
rect 645482 77637 645488 77649
rect 650992 77637 650998 77649
rect 651050 77637 651056 77689
rect 162832 77563 162838 77615
rect 162890 77603 162896 77615
rect 200272 77603 200278 77615
rect 162890 77575 200278 77603
rect 162890 77563 162896 77575
rect 200272 77563 200278 77575
rect 200330 77563 200336 77615
rect 185872 77489 185878 77541
rect 185930 77529 185936 77541
rect 210160 77529 210166 77541
rect 185930 77501 210166 77529
rect 185930 77489 185936 77501
rect 210160 77489 210166 77501
rect 210218 77489 210224 77541
rect 191632 77415 191638 77467
rect 191690 77455 191696 77467
rect 201712 77455 201718 77467
rect 191690 77427 201718 77455
rect 191690 77415 191696 77427
rect 201712 77415 201718 77427
rect 201770 77415 201776 77467
rect 645424 77267 645430 77319
rect 645482 77307 645488 77319
rect 662896 77307 662902 77319
rect 645482 77279 662902 77307
rect 645482 77267 645488 77279
rect 662896 77267 662902 77279
rect 662954 77267 662960 77319
rect 190000 77193 190006 77245
rect 190058 77233 190064 77245
rect 201712 77233 201718 77245
rect 190058 77205 201718 77233
rect 190058 77193 190064 77205
rect 201712 77193 201718 77205
rect 201770 77193 201776 77245
rect 645904 76971 645910 77023
rect 645962 77011 645968 77023
rect 661744 77011 661750 77023
rect 645962 76983 661750 77011
rect 645962 76971 645968 76983
rect 661744 76971 661750 76983
rect 661802 76971 661808 77023
rect 645424 76897 645430 76949
rect 645482 76937 645488 76949
rect 658288 76937 658294 76949
rect 645482 76909 658294 76937
rect 645482 76897 645488 76909
rect 658288 76897 658294 76909
rect 658346 76897 658352 76949
rect 645808 76675 645814 76727
rect 645866 76715 645872 76727
rect 650896 76715 650902 76727
rect 645866 76687 650902 76715
rect 645866 76675 645872 76687
rect 650896 76675 650902 76687
rect 650954 76675 650960 76727
rect 640720 76231 640726 76283
rect 640778 76271 640784 76283
rect 651280 76271 651286 76283
rect 640778 76243 651286 76271
rect 640778 76231 640784 76243
rect 651280 76231 651286 76243
rect 651338 76231 651344 76283
rect 645424 75491 645430 75543
rect 645482 75531 645488 75543
rect 656848 75531 656854 75543
rect 645482 75503 656854 75531
rect 645482 75491 645488 75503
rect 656848 75491 656854 75503
rect 656906 75491 656912 75543
rect 146320 75269 146326 75321
rect 146378 75309 146384 75321
rect 146378 75281 148190 75309
rect 146378 75269 146384 75281
rect 146128 75195 146134 75247
rect 146186 75235 146192 75247
rect 146512 75235 146518 75247
rect 146186 75207 146518 75235
rect 146186 75195 146192 75207
rect 146512 75195 146518 75207
rect 146570 75195 146576 75247
rect 144016 75121 144022 75173
rect 144074 75161 144080 75173
rect 144074 75133 146270 75161
rect 144074 75121 144080 75133
rect 144208 75047 144214 75099
rect 144266 75087 144272 75099
rect 146128 75087 146134 75099
rect 144266 75059 146134 75087
rect 144266 75047 144272 75059
rect 146128 75047 146134 75059
rect 146186 75047 146192 75099
rect 146242 75087 146270 75133
rect 148162 75087 148190 75281
rect 160048 75087 160054 75099
rect 146242 75059 148094 75087
rect 148162 75059 160054 75087
rect 144112 74973 144118 75025
rect 144170 75013 144176 75025
rect 146320 75013 146326 75025
rect 144170 74985 146326 75013
rect 144170 74973 144176 74985
rect 146320 74973 146326 74985
rect 146378 74973 146384 75025
rect 148066 75013 148094 75059
rect 160048 75047 160054 75059
rect 160106 75047 160112 75099
rect 156400 75013 156406 75025
rect 148066 74985 156406 75013
rect 156400 74973 156406 74985
rect 156458 74973 156464 75025
rect 144400 74899 144406 74951
rect 144458 74939 144464 74951
rect 161488 74939 161494 74951
rect 144458 74911 161494 74939
rect 144458 74899 144464 74911
rect 161488 74899 161494 74911
rect 161546 74899 161552 74951
rect 154000 74825 154006 74877
rect 154058 74865 154064 74877
rect 201520 74865 201526 74877
rect 154058 74837 201526 74865
rect 154058 74825 154064 74837
rect 201520 74825 201526 74837
rect 201578 74825 201584 74877
rect 174448 74751 174454 74803
rect 174506 74791 174512 74803
rect 201808 74791 201814 74803
rect 174506 74763 201814 74791
rect 174506 74751 174512 74763
rect 201808 74751 201814 74763
rect 201866 74751 201872 74803
rect 177232 74677 177238 74729
rect 177290 74717 177296 74729
rect 210160 74717 210166 74729
rect 177290 74689 210166 74717
rect 177290 74677 177296 74689
rect 210160 74677 210166 74689
rect 210218 74677 210224 74729
rect 180112 74603 180118 74655
rect 180170 74643 180176 74655
rect 201616 74643 201622 74655
rect 180170 74615 201622 74643
rect 180170 74603 180176 74615
rect 201616 74603 201622 74615
rect 201674 74603 201680 74655
rect 182992 74529 182998 74581
rect 183050 74569 183056 74581
rect 201712 74569 201718 74581
rect 183050 74541 201718 74569
rect 183050 74529 183056 74541
rect 201712 74529 201718 74541
rect 201770 74529 201776 74581
rect 144400 74455 144406 74507
rect 144458 74495 144464 74507
rect 148336 74495 148342 74507
rect 144458 74467 148342 74495
rect 144458 74455 144464 74467
rect 148336 74455 148342 74467
rect 148394 74455 148400 74507
rect 144208 74011 144214 74063
rect 144266 74051 144272 74063
rect 146704 74051 146710 74063
rect 144266 74023 146710 74051
rect 144266 74011 144272 74023
rect 146704 74011 146710 74023
rect 146762 74011 146768 74063
rect 645424 72975 645430 73027
rect 645482 73015 645488 73027
rect 663376 73015 663382 73027
rect 645482 72987 663382 73015
rect 645482 72975 645488 72987
rect 663376 72975 663382 72987
rect 663434 72975 663440 73027
rect 645808 72309 645814 72361
rect 645866 72349 645872 72361
rect 660112 72349 660118 72361
rect 645866 72321 660118 72349
rect 645866 72309 645872 72321
rect 660112 72309 660118 72321
rect 660170 72309 660176 72361
rect 645424 72087 645430 72139
rect 645482 72127 645488 72139
rect 663184 72127 663190 72139
rect 645482 72099 663190 72127
rect 645482 72087 645488 72099
rect 663184 72087 663190 72099
rect 663242 72087 663248 72139
rect 146704 72013 146710 72065
rect 146762 72053 146768 72065
rect 153904 72053 153910 72065
rect 146762 72025 153910 72053
rect 146762 72013 146768 72025
rect 153904 72013 153910 72025
rect 153962 72013 153968 72065
rect 151120 71939 151126 71991
rect 151178 71979 151184 71991
rect 200368 71979 200374 71991
rect 151178 71951 200374 71979
rect 151178 71939 151184 71951
rect 200368 71939 200374 71951
rect 200426 71939 200432 71991
rect 209776 71939 209782 71991
rect 209834 71979 209840 71991
rect 210160 71979 210166 71991
rect 209834 71951 210166 71979
rect 209834 71939 209840 71951
rect 210160 71939 210166 71951
rect 210218 71939 210224 71991
rect 161488 71865 161494 71917
rect 161546 71905 161552 71917
rect 201808 71905 201814 71917
rect 161546 71877 201814 71905
rect 161546 71865 161552 71877
rect 201808 71865 201814 71877
rect 201866 71865 201872 71917
rect 165616 71791 165622 71843
rect 165674 71831 165680 71843
rect 201616 71831 201622 71843
rect 165674 71803 201622 71831
rect 165674 71791 165680 71803
rect 201616 71791 201622 71803
rect 201674 71791 201680 71843
rect 209776 71791 209782 71843
rect 209834 71831 209840 71843
rect 209968 71831 209974 71843
rect 209834 71803 209974 71831
rect 209834 71791 209840 71803
rect 209968 71791 209974 71803
rect 210026 71791 210032 71843
rect 168496 71717 168502 71769
rect 168554 71757 168560 71769
rect 201712 71757 201718 71769
rect 168554 71729 201718 71757
rect 168554 71717 168560 71729
rect 201712 71717 201718 71729
rect 201770 71717 201776 71769
rect 171376 71643 171382 71695
rect 171434 71683 171440 71695
rect 209968 71683 209974 71695
rect 171434 71655 209974 71683
rect 171434 71643 171440 71655
rect 209968 71643 209974 71655
rect 210026 71643 210032 71695
rect 146704 70903 146710 70955
rect 146762 70943 146768 70955
rect 149776 70943 149782 70955
rect 146762 70915 149782 70943
rect 146762 70903 146768 70915
rect 149776 70903 149782 70915
rect 149834 70903 149840 70955
rect 144112 69497 144118 69549
rect 144170 69537 144176 69549
rect 145648 69537 145654 69549
rect 144170 69509 145654 69537
rect 144170 69497 144176 69509
rect 145648 69497 145654 69509
rect 145706 69497 145712 69549
rect 145456 69349 145462 69401
rect 145514 69389 145520 69401
rect 145648 69389 145654 69401
rect 145514 69361 145654 69389
rect 145514 69349 145520 69361
rect 145648 69349 145654 69361
rect 145706 69349 145712 69401
rect 145456 69201 145462 69253
rect 145514 69241 145520 69253
rect 145840 69241 145846 69253
rect 145514 69213 145846 69241
rect 145514 69201 145520 69213
rect 145840 69201 145846 69213
rect 145898 69201 145904 69253
rect 144016 69127 144022 69179
rect 144074 69167 144080 69179
rect 144074 69139 146942 69167
rect 144074 69127 144080 69139
rect 146914 69093 146942 69139
rect 201808 69093 201814 69105
rect 146914 69065 201814 69093
rect 201808 69053 201814 69065
rect 201866 69053 201872 69105
rect 149776 68979 149782 69031
rect 149834 69019 149840 69031
rect 201616 69019 201622 69031
rect 149834 68991 201622 69019
rect 149834 68979 149840 68991
rect 201616 68979 201622 68991
rect 201674 68979 201680 69031
rect 153904 68905 153910 68957
rect 153962 68945 153968 68957
rect 201712 68945 201718 68957
rect 153962 68917 201718 68945
rect 153962 68905 153968 68917
rect 201712 68905 201718 68917
rect 201770 68905 201776 68957
rect 156400 68831 156406 68883
rect 156458 68871 156464 68883
rect 196240 68871 196246 68883
rect 156458 68843 196246 68871
rect 156458 68831 156464 68843
rect 196240 68831 196246 68843
rect 196298 68831 196304 68883
rect 160048 68757 160054 68809
rect 160106 68797 160112 68809
rect 195472 68797 195478 68809
rect 160106 68769 195478 68797
rect 160106 68757 160112 68769
rect 195472 68757 195478 68769
rect 195530 68757 195536 68809
rect 146704 67351 146710 67403
rect 146762 67391 146768 67403
rect 152656 67391 152662 67403
rect 146762 67363 152662 67391
rect 146762 67351 146768 67363
rect 152656 67351 152662 67363
rect 152714 67351 152720 67403
rect 145840 66389 145846 66441
rect 145898 66429 145904 66441
rect 158320 66429 158326 66441
rect 145898 66401 158326 66429
rect 145898 66389 145904 66401
rect 158320 66389 158326 66401
rect 158378 66389 158384 66441
rect 146800 66241 146806 66293
rect 146858 66281 146864 66293
rect 146858 66253 149822 66281
rect 146858 66241 146864 66253
rect 149794 66207 149822 66253
rect 645520 66241 645526 66293
rect 645578 66281 645584 66293
rect 646096 66281 646102 66293
rect 645578 66253 646102 66281
rect 645578 66241 645584 66253
rect 646096 66241 646102 66253
rect 646154 66241 646160 66293
rect 201712 66207 201718 66219
rect 149794 66179 201718 66207
rect 201712 66167 201718 66179
rect 201770 66167 201776 66219
rect 152656 66093 152662 66145
rect 152714 66133 152720 66145
rect 198544 66133 198550 66145
rect 152714 66105 198550 66133
rect 152714 66093 152720 66105
rect 198544 66093 198550 66105
rect 198602 66093 198608 66145
rect 158320 66019 158326 66071
rect 158378 66059 158384 66071
rect 193648 66059 193654 66071
rect 158378 66031 193654 66059
rect 158378 66019 158384 66031
rect 193648 66019 193654 66031
rect 193706 66019 193712 66071
rect 145648 64835 145654 64887
rect 145706 64835 145712 64887
rect 146704 64835 146710 64887
rect 146762 64875 146768 64887
rect 201712 64875 201718 64887
rect 146762 64847 201718 64875
rect 146762 64835 146768 64847
rect 201712 64835 201718 64847
rect 201770 64835 201776 64887
rect 144496 64613 144502 64665
rect 144554 64653 144560 64665
rect 144688 64653 144694 64665
rect 144554 64625 144694 64653
rect 144554 64613 144560 64625
rect 144688 64613 144694 64625
rect 144746 64613 144752 64665
rect 144784 64613 144790 64665
rect 144842 64653 144848 64665
rect 145552 64653 145558 64665
rect 144842 64625 145558 64653
rect 144842 64613 144848 64625
rect 145552 64613 145558 64625
rect 145610 64613 145616 64665
rect 144688 64465 144694 64517
rect 144746 64505 144752 64517
rect 145666 64505 145694 64835
rect 146800 64761 146806 64813
rect 146858 64801 146864 64813
rect 201808 64801 201814 64813
rect 146858 64773 201814 64801
rect 146858 64761 146864 64773
rect 201808 64761 201814 64773
rect 201866 64761 201872 64813
rect 144746 64477 145694 64505
rect 144746 64465 144752 64477
rect 144208 64391 144214 64443
rect 144266 64431 144272 64443
rect 145936 64431 145942 64443
rect 144266 64403 145942 64431
rect 144266 64391 144272 64403
rect 145936 64391 145942 64403
rect 145994 64391 146000 64443
rect 146896 63355 146902 63407
rect 146954 63395 146960 63407
rect 195472 63395 195478 63407
rect 146954 63367 195478 63395
rect 146954 63355 146960 63367
rect 195472 63355 195478 63367
rect 195530 63355 195536 63407
rect 209392 62763 209398 62815
rect 209450 62803 209456 62815
rect 210256 62803 210262 62815
rect 209450 62775 210262 62803
rect 209450 62763 209456 62775
rect 210256 62763 210262 62775
rect 210314 62763 210320 62815
rect 209488 62615 209494 62667
rect 209546 62655 209552 62667
rect 210256 62655 210262 62667
rect 209546 62627 210262 62655
rect 209546 62615 209552 62627
rect 210256 62615 210262 62627
rect 210314 62615 210320 62667
rect 146800 62467 146806 62519
rect 146858 62507 146864 62519
rect 149776 62507 149782 62519
rect 146858 62479 149782 62507
rect 146858 62467 146864 62479
rect 149776 62467 149782 62479
rect 149834 62467 149840 62519
rect 160528 60765 160534 60817
rect 160586 60805 160592 60817
rect 201712 60805 201718 60817
rect 160586 60777 201718 60805
rect 160586 60765 160592 60777
rect 201712 60765 201718 60777
rect 201770 60765 201776 60817
rect 156304 60691 156310 60743
rect 156362 60731 156368 60743
rect 201616 60731 201622 60743
rect 156362 60703 201622 60731
rect 156362 60691 156368 60703
rect 201616 60691 201622 60703
rect 201674 60691 201680 60743
rect 152656 60617 152662 60669
rect 152714 60657 152720 60669
rect 195472 60657 195478 60669
rect 152714 60629 195478 60657
rect 152714 60617 152720 60629
rect 195472 60617 195478 60629
rect 195530 60617 195536 60669
rect 151120 60543 151126 60595
rect 151178 60583 151184 60595
rect 201520 60583 201526 60595
rect 151178 60555 201526 60583
rect 151178 60543 151184 60555
rect 201520 60543 201526 60555
rect 201578 60543 201584 60595
rect 148336 60469 148342 60521
rect 148394 60509 148400 60521
rect 201808 60509 201814 60521
rect 148394 60481 201814 60509
rect 148394 60469 148400 60481
rect 201808 60469 201814 60481
rect 201866 60469 201872 60521
rect 146896 60395 146902 60447
rect 146954 60435 146960 60447
rect 209968 60435 209974 60447
rect 146954 60407 209974 60435
rect 146954 60395 146960 60407
rect 209968 60395 209974 60407
rect 210026 60395 210032 60447
rect 149776 60321 149782 60373
rect 149834 60361 149840 60373
rect 198352 60361 198358 60373
rect 149834 60333 198358 60361
rect 149834 60321 149840 60333
rect 198352 60321 198358 60333
rect 198410 60321 198416 60373
rect 146800 59581 146806 59633
rect 146858 59621 146864 59633
rect 160528 59621 160534 59633
rect 146858 59593 160534 59621
rect 146858 59581 146864 59593
rect 160528 59581 160534 59593
rect 160586 59581 160592 59633
rect 146800 58989 146806 59041
rect 146858 59029 146864 59041
rect 201712 59029 201718 59041
rect 146858 59001 201718 59029
rect 146858 58989 146864 59001
rect 201712 58989 201718 59001
rect 201770 58989 201776 59041
rect 146800 57065 146806 57117
rect 146858 57105 146864 57117
rect 156304 57105 156310 57117
rect 146858 57077 156310 57105
rect 146858 57065 146864 57077
rect 156304 57065 156310 57077
rect 156362 57065 156368 57117
rect 144112 56917 144118 56969
rect 144170 56957 144176 56969
rect 146800 56957 146806 56969
rect 144170 56929 146806 56957
rect 144170 56917 144176 56929
rect 146800 56917 146806 56929
rect 146858 56917 146864 56969
rect 144016 56473 144022 56525
rect 144074 56513 144080 56525
rect 152656 56513 152662 56525
rect 144074 56485 152662 56513
rect 144074 56473 144080 56485
rect 152656 56473 152662 56485
rect 152714 56473 152720 56525
rect 144784 54623 144790 54675
rect 144842 54663 144848 54675
rect 151120 54663 151126 54675
rect 144842 54635 151126 54663
rect 144842 54623 144848 54635
rect 151120 54623 151126 54635
rect 151178 54623 151184 54675
rect 144208 54327 144214 54379
rect 144266 54367 144272 54379
rect 144592 54367 144598 54379
rect 144266 54339 144598 54367
rect 144266 54327 144272 54339
rect 144592 54327 144598 54339
rect 144650 54327 144656 54379
rect 210256 54327 210262 54379
rect 210314 54367 210320 54379
rect 210314 54339 219422 54367
rect 210314 54327 210320 54339
rect 219394 54305 219422 54339
rect 209296 54253 209302 54305
rect 209354 54293 209360 54305
rect 217456 54293 217462 54305
rect 209354 54265 217462 54293
rect 209354 54253 209360 54265
rect 217456 54253 217462 54265
rect 217514 54253 217520 54305
rect 219376 54253 219382 54305
rect 219434 54253 219440 54305
rect 209776 54179 209782 54231
rect 209834 54219 209840 54231
rect 219184 54219 219190 54231
rect 209834 54191 219190 54219
rect 209834 54179 209840 54191
rect 219184 54179 219190 54191
rect 219242 54179 219248 54231
rect 144496 54105 144502 54157
rect 144554 54145 144560 54157
rect 148336 54145 148342 54157
rect 144554 54117 148342 54145
rect 144554 54105 144560 54117
rect 148336 54105 148342 54117
rect 148394 54105 148400 54157
rect 209680 54105 209686 54157
rect 209738 54145 209744 54157
rect 213760 54145 213766 54157
rect 209738 54117 213766 54145
rect 209738 54105 209744 54117
rect 213760 54105 213766 54117
rect 213818 54105 213824 54157
rect 205648 53957 205654 54009
rect 205706 53997 205712 54009
rect 218176 53997 218182 54009
rect 205706 53969 218182 53997
rect 205706 53957 205712 53969
rect 218176 53957 218182 53969
rect 218234 53957 218240 54009
rect 208336 53883 208342 53935
rect 208394 53923 208400 53935
rect 214960 53923 214966 53935
rect 208394 53895 214966 53923
rect 208394 53883 208400 53895
rect 214960 53883 214966 53895
rect 215018 53883 215024 53935
rect 261904 53923 261910 53935
rect 241858 53895 261910 53923
rect 210352 53809 210358 53861
rect 210410 53849 210416 53861
rect 221392 53849 221398 53861
rect 210410 53821 221398 53849
rect 210410 53809 210416 53821
rect 221392 53809 221398 53821
rect 221450 53809 221456 53861
rect 231760 53809 231766 53861
rect 231818 53849 231824 53861
rect 241858 53849 241886 53895
rect 261904 53883 261910 53895
rect 261962 53883 261968 53935
rect 282160 53923 282166 53935
rect 262210 53895 282166 53923
rect 231818 53821 241886 53849
rect 231818 53809 231824 53821
rect 262000 53809 262006 53861
rect 262058 53849 262064 53861
rect 262058 53821 262142 53849
rect 262058 53809 262064 53821
rect 209968 53735 209974 53787
rect 210026 53775 210032 53787
rect 219184 53775 219190 53787
rect 210026 53747 219190 53775
rect 210026 53735 210032 53747
rect 219184 53735 219190 53747
rect 219242 53735 219248 53787
rect 262114 53775 262142 53821
rect 262210 53775 262238 53895
rect 282160 53883 282166 53895
rect 282218 53883 282224 53935
rect 262114 53747 262238 53775
rect 210160 53661 210166 53713
rect 210218 53701 210224 53713
rect 210218 53673 221822 53701
rect 210218 53661 210224 53673
rect 207952 53587 207958 53639
rect 208010 53627 208016 53639
rect 221794 53627 221822 53673
rect 231760 53627 231766 53639
rect 208010 53599 216398 53627
rect 221794 53599 231766 53627
rect 208010 53587 208016 53599
rect 216370 53565 216398 53599
rect 231760 53587 231766 53599
rect 231818 53587 231824 53639
rect 209392 53513 209398 53565
rect 209450 53553 209456 53565
rect 215248 53553 215254 53565
rect 209450 53525 215254 53553
rect 209450 53513 209456 53525
rect 215248 53513 215254 53525
rect 215306 53513 215312 53565
rect 216352 53513 216358 53565
rect 216410 53513 216416 53565
rect 351280 53553 351286 53565
rect 219010 53525 351286 53553
rect 209488 53439 209494 53491
rect 209546 53479 209552 53491
rect 218896 53479 218902 53491
rect 209546 53451 218902 53479
rect 209546 53439 209552 53451
rect 218896 53439 218902 53451
rect 218954 53439 218960 53491
rect 210640 53365 210646 53417
rect 210698 53405 210704 53417
rect 219010 53405 219038 53525
rect 351280 53513 351286 53525
rect 351338 53513 351344 53565
rect 219184 53439 219190 53491
rect 219242 53479 219248 53491
rect 384400 53479 384406 53491
rect 219242 53451 384406 53479
rect 219242 53439 219248 53451
rect 384400 53439 384406 53451
rect 384458 53439 384464 53491
rect 210698 53377 219038 53405
rect 210698 53365 210704 53377
rect 219376 53365 219382 53417
rect 219434 53405 219440 53417
rect 467440 53405 467446 53417
rect 219434 53377 467446 53405
rect 219434 53365 219440 53377
rect 467440 53365 467446 53377
rect 467498 53365 467504 53417
rect 469360 53365 469366 53417
rect 469418 53405 469424 53417
rect 501040 53405 501046 53417
rect 469418 53377 501046 53405
rect 469418 53365 469424 53377
rect 501040 53365 501046 53377
rect 501098 53365 501104 53417
rect 210256 53291 210262 53343
rect 210314 53331 210320 53343
rect 219664 53331 219670 53343
rect 210314 53303 219670 53331
rect 210314 53291 210320 53303
rect 219664 53291 219670 53303
rect 219722 53291 219728 53343
rect 221392 53291 221398 53343
rect 221450 53331 221456 53343
rect 501136 53331 501142 53343
rect 221450 53303 501142 53331
rect 221450 53291 221456 53303
rect 501136 53291 501142 53303
rect 501194 53291 501200 53343
rect 204880 53217 204886 53269
rect 204938 53257 204944 53269
rect 215632 53257 215638 53269
rect 204938 53229 215638 53257
rect 204938 53217 204944 53229
rect 215632 53217 215638 53229
rect 215690 53217 215696 53269
rect 292258 53229 292478 53257
rect 210448 53143 210454 53195
rect 210506 53183 210512 53195
rect 213424 53183 213430 53195
rect 210506 53155 213430 53183
rect 210506 53143 210512 53155
rect 213424 53143 213430 53155
rect 213482 53143 213488 53195
rect 251920 53143 251926 53195
rect 251978 53183 251984 53195
rect 292258 53183 292286 53229
rect 251978 53155 262046 53183
rect 251978 53143 251984 53155
rect 208048 53069 208054 53121
rect 208106 53109 208112 53121
rect 220336 53109 220342 53121
rect 208106 53081 220342 53109
rect 208106 53069 208112 53081
rect 220336 53069 220342 53081
rect 220394 53069 220400 53121
rect 262018 53109 262046 53155
rect 267778 53155 292286 53183
rect 292450 53183 292478 53229
rect 315664 53217 315670 53269
rect 315722 53257 315728 53269
rect 368560 53257 368566 53269
rect 315722 53229 368566 53257
rect 315722 53217 315728 53229
rect 368560 53217 368566 53229
rect 368618 53217 368624 53269
rect 388816 53217 388822 53269
rect 388874 53257 388880 53269
rect 408976 53257 408982 53269
rect 388874 53229 408982 53257
rect 388874 53217 388880 53229
rect 408976 53217 408982 53229
rect 409034 53217 409040 53269
rect 429154 53229 449246 53257
rect 292450 53155 302366 53183
rect 267778 53109 267806 53155
rect 262018 53081 267806 53109
rect 302338 53109 302366 53155
rect 368656 53143 368662 53195
rect 368714 53183 368720 53195
rect 388720 53183 388726 53195
rect 368714 53155 388726 53183
rect 368714 53143 368720 53155
rect 388720 53143 388726 53155
rect 388778 53143 388784 53195
rect 302338 53081 302462 53109
rect 216976 52995 216982 53047
rect 217034 53035 217040 53047
rect 302434 53035 302462 53081
rect 315664 53035 315670 53047
rect 217034 53007 241886 53035
rect 302434 53007 315670 53035
rect 217034 52995 217040 53007
rect 241858 52961 241886 53007
rect 315664 52995 315670 53007
rect 315722 52995 315728 53047
rect 409072 52995 409078 53047
rect 409130 53035 409136 53047
rect 429154 53035 429182 53229
rect 449218 53183 449246 53229
rect 449314 53229 463646 53257
rect 449314 53183 449342 53229
rect 449218 53155 449342 53183
rect 463618 53183 463646 53229
rect 469360 53183 469366 53195
rect 463618 53155 469366 53183
rect 469360 53143 469366 53155
rect 469418 53143 469424 53195
rect 501040 53143 501046 53195
rect 501098 53183 501104 53195
rect 509680 53183 509686 53195
rect 501098 53155 509686 53183
rect 501098 53143 501104 53155
rect 509680 53143 509686 53155
rect 509738 53143 509744 53195
rect 409130 53007 429182 53035
rect 409130 52995 409136 53007
rect 251920 52961 251926 52973
rect 241858 52933 251926 52961
rect 251920 52921 251926 52933
rect 251978 52921 251984 52973
rect 159952 52847 159958 52899
rect 160010 52887 160016 52899
rect 217264 52887 217270 52899
rect 160010 52859 217270 52887
rect 160010 52847 160016 52859
rect 217264 52847 217270 52859
rect 217322 52847 217328 52899
rect 211600 52773 211606 52825
rect 211658 52813 211664 52825
rect 219952 52813 219958 52825
rect 211658 52785 219958 52813
rect 211658 52773 211664 52785
rect 219952 52773 219958 52785
rect 220010 52773 220016 52825
rect 151312 52699 151318 52751
rect 151370 52739 151376 52751
rect 216496 52739 216502 52751
rect 151370 52711 216502 52739
rect 151370 52699 151376 52711
rect 216496 52699 216502 52711
rect 216554 52699 216560 52751
rect 212272 52477 212278 52529
rect 212330 52517 212336 52529
rect 213424 52517 213430 52529
rect 212330 52489 213430 52517
rect 212330 52477 212336 52489
rect 213424 52477 213430 52489
rect 213482 52477 213488 52529
rect 211216 52403 211222 52455
rect 211274 52443 211280 52455
rect 213808 52443 213814 52455
rect 211274 52415 213814 52443
rect 211274 52403 211280 52415
rect 213808 52403 213814 52415
rect 213866 52403 213872 52455
rect 203056 52329 203062 52381
rect 203114 52369 203120 52381
rect 226576 52369 226582 52381
rect 203114 52341 226582 52369
rect 203114 52329 203120 52341
rect 226576 52329 226582 52341
rect 226634 52329 226640 52381
rect 146512 52255 146518 52307
rect 146570 52295 146576 52307
rect 225712 52295 225718 52307
rect 146570 52267 225718 52295
rect 146570 52255 146576 52267
rect 225712 52255 225718 52267
rect 225770 52255 225776 52307
rect 171472 52181 171478 52233
rect 171530 52221 171536 52233
rect 219856 52221 219862 52233
rect 171530 52193 219862 52221
rect 171530 52181 171536 52193
rect 219856 52181 219862 52193
rect 219914 52181 219920 52233
rect 146320 52107 146326 52159
rect 146378 52147 146384 52159
rect 226960 52147 226966 52159
rect 146378 52119 226966 52147
rect 146378 52107 146384 52119
rect 226960 52107 226966 52119
rect 227018 52107 227024 52159
rect 144208 52033 144214 52085
rect 144266 52073 144272 52085
rect 220912 52073 220918 52085
rect 144266 52045 220918 52073
rect 144266 52033 144272 52045
rect 220912 52033 220918 52045
rect 220970 52033 220976 52085
rect 145072 51959 145078 52011
rect 145130 51999 145136 52011
rect 203056 51999 203062 52011
rect 145130 51971 203062 51999
rect 145130 51959 145136 51971
rect 203056 51959 203062 51971
rect 203114 51959 203120 52011
rect 213346 51971 213566 51999
rect 146128 51885 146134 51937
rect 146186 51925 146192 51937
rect 213346 51925 213374 51971
rect 146186 51897 213374 51925
rect 213538 51925 213566 51971
rect 227536 51925 227542 51937
rect 213538 51897 227542 51925
rect 146186 51885 146192 51897
rect 227536 51885 227542 51897
rect 227594 51885 227600 51937
rect 213424 51811 213430 51863
rect 213482 51851 213488 51863
rect 213482 51823 219902 51851
rect 213482 51811 213488 51823
rect 213808 51737 213814 51789
rect 213866 51777 213872 51789
rect 219874 51777 219902 51823
rect 219952 51811 219958 51863
rect 220010 51851 220016 51863
rect 645520 51851 645526 51863
rect 220010 51823 645526 51851
rect 220010 51811 220016 51823
rect 645520 51811 645526 51823
rect 645578 51811 645584 51863
rect 645712 51777 645718 51789
rect 213866 51749 219326 51777
rect 219874 51749 645718 51777
rect 213866 51737 213872 51749
rect 209872 51663 209878 51715
rect 209930 51703 209936 51715
rect 214096 51703 214102 51715
rect 209930 51675 214102 51703
rect 209930 51663 209936 51675
rect 214096 51663 214102 51675
rect 214154 51663 214160 51715
rect 219298 51703 219326 51749
rect 645712 51737 645718 51749
rect 645770 51737 645776 51789
rect 639664 51703 639670 51715
rect 219298 51675 639670 51703
rect 639664 51663 639670 51675
rect 639722 51663 639728 51715
rect 209584 51589 209590 51641
rect 209642 51629 209648 51641
rect 214480 51629 214486 51641
rect 209642 51601 214486 51629
rect 209642 51589 209648 51601
rect 214480 51589 214486 51601
rect 214538 51589 214544 51641
rect 144976 51441 144982 51493
rect 145034 51481 145040 51493
rect 233584 51481 233590 51493
rect 145034 51453 233590 51481
rect 145034 51441 145040 51453
rect 233584 51441 233590 51453
rect 233642 51441 233648 51493
rect 145168 51367 145174 51419
rect 145226 51407 145232 51419
rect 234544 51407 234550 51419
rect 145226 51379 234550 51407
rect 145226 51367 145232 51379
rect 234544 51367 234550 51379
rect 234602 51367 234608 51419
rect 145360 51293 145366 51345
rect 145418 51333 145424 51345
rect 235792 51333 235798 51345
rect 145418 51305 235798 51333
rect 145418 51293 145424 51305
rect 235792 51293 235798 51305
rect 235850 51293 235856 51345
rect 145648 51219 145654 51271
rect 145706 51259 145712 51271
rect 235312 51259 235318 51271
rect 145706 51231 235318 51259
rect 145706 51219 145712 51231
rect 235312 51219 235318 51231
rect 235370 51219 235376 51271
rect 146032 51145 146038 51197
rect 146090 51185 146096 51197
rect 232336 51185 232342 51197
rect 146090 51157 232342 51185
rect 146090 51145 146096 51157
rect 232336 51145 232342 51157
rect 232394 51145 232400 51197
rect 146224 51071 146230 51123
rect 146282 51111 146288 51123
rect 231376 51111 231382 51123
rect 146282 51083 231382 51111
rect 146282 51071 146288 51083
rect 231376 51071 231382 51083
rect 231434 51071 231440 51123
rect 146416 50997 146422 51049
rect 146474 51037 146480 51049
rect 231952 51037 231958 51049
rect 146474 51009 231958 51037
rect 146474 50997 146480 51009
rect 231952 50997 231958 51009
rect 232010 50997 232016 51049
rect 146608 50923 146614 50975
rect 146666 50963 146672 50975
rect 230896 50963 230902 50975
rect 146666 50935 230902 50963
rect 146666 50923 146672 50935
rect 230896 50923 230902 50935
rect 230954 50923 230960 50975
rect 144880 50849 144886 50901
rect 144938 50889 144944 50901
rect 230128 50889 230134 50901
rect 144938 50861 230134 50889
rect 144938 50849 144944 50861
rect 230128 50849 230134 50861
rect 230186 50849 230192 50901
rect 145264 50775 145270 50827
rect 145322 50815 145328 50827
rect 228784 50815 228790 50827
rect 145322 50787 228790 50815
rect 145322 50775 145328 50787
rect 228784 50775 228790 50787
rect 228842 50775 228848 50827
rect 146704 50701 146710 50753
rect 146762 50741 146768 50753
rect 228688 50741 228694 50753
rect 146762 50713 228694 50741
rect 146762 50701 146768 50713
rect 228688 50701 228694 50713
rect 228746 50701 228752 50753
rect 145936 50627 145942 50679
rect 145994 50667 146000 50679
rect 229168 50667 229174 50679
rect 145994 50639 229174 50667
rect 145994 50627 146000 50639
rect 229168 50627 229174 50639
rect 229226 50627 229232 50679
rect 144400 50553 144406 50605
rect 144458 50593 144464 50605
rect 208048 50593 208054 50605
rect 144458 50565 208054 50593
rect 144458 50553 144464 50565
rect 208048 50553 208054 50565
rect 208106 50553 208112 50605
rect 208240 50553 208246 50605
rect 208298 50593 208304 50605
rect 216112 50593 216118 50605
rect 208298 50565 216118 50593
rect 208298 50553 208304 50565
rect 216112 50553 216118 50565
rect 216170 50553 216176 50605
rect 144688 50479 144694 50531
rect 144746 50519 144752 50531
rect 208336 50519 208342 50531
rect 144746 50491 208342 50519
rect 144746 50479 144752 50491
rect 208336 50479 208342 50491
rect 208394 50479 208400 50531
rect 208432 50479 208438 50531
rect 208490 50519 208496 50531
rect 216880 50519 216886 50531
rect 208490 50491 216886 50519
rect 208490 50479 208496 50491
rect 216880 50479 216886 50491
rect 216938 50479 216944 50531
rect 145552 50405 145558 50457
rect 145610 50445 145616 50457
rect 211504 50445 211510 50457
rect 145610 50417 211510 50445
rect 145610 50405 145616 50417
rect 211504 50405 211510 50417
rect 211562 50405 211568 50457
rect 144304 50331 144310 50383
rect 144362 50371 144368 50383
rect 209104 50371 209110 50383
rect 144362 50343 209110 50371
rect 144362 50331 144368 50343
rect 209104 50331 209110 50343
rect 209162 50331 209168 50383
rect 209392 50331 209398 50383
rect 209450 50371 209456 50383
rect 221488 50371 221494 50383
rect 209450 50343 221494 50371
rect 209450 50331 209456 50343
rect 221488 50331 221494 50343
rect 221546 50331 221552 50383
rect 144784 50257 144790 50309
rect 144842 50297 144848 50309
rect 235408 50297 235414 50309
rect 144842 50269 235414 50297
rect 144842 50257 144848 50269
rect 235408 50257 235414 50269
rect 235466 50257 235472 50309
rect 145744 50183 145750 50235
rect 145802 50223 145808 50235
rect 234928 50223 234934 50235
rect 145802 50195 234934 50223
rect 145802 50183 145808 50195
rect 234928 50183 234934 50195
rect 234986 50183 234992 50235
rect 145840 50109 145846 50161
rect 145898 50149 145904 50161
rect 232720 50149 232726 50161
rect 145898 50121 232726 50149
rect 145898 50109 145904 50121
rect 232720 50109 232726 50121
rect 232778 50109 232784 50161
rect 209104 50035 209110 50087
rect 209162 50075 209168 50087
rect 223888 50075 223894 50087
rect 209162 50047 223894 50075
rect 209162 50035 209168 50047
rect 223888 50035 223894 50047
rect 223946 50035 223952 50087
rect 208048 49961 208054 50013
rect 208106 50001 208112 50013
rect 225328 50001 225334 50013
rect 208106 49973 225334 50001
rect 208106 49961 208112 49973
rect 225328 49961 225334 49973
rect 225386 49961 225392 50013
rect 146800 49887 146806 49939
rect 146858 49927 146864 49939
rect 241168 49927 241174 49939
rect 146858 49899 241174 49927
rect 146858 49887 146864 49899
rect 241168 49887 241174 49899
rect 241226 49887 241232 49939
rect 145360 49813 145366 49865
rect 145418 49853 145424 49865
rect 244144 49853 244150 49865
rect 145418 49825 244150 49853
rect 145418 49813 145424 49825
rect 244144 49813 244150 49825
rect 244202 49813 244208 49865
rect 208336 49739 208342 49791
rect 208394 49779 208400 49791
rect 226096 49779 226102 49791
rect 208394 49751 226102 49779
rect 208394 49739 208400 49751
rect 226096 49739 226102 49751
rect 226154 49739 226160 49791
rect 145456 49665 145462 49717
rect 145514 49705 145520 49717
rect 237136 49705 237142 49717
rect 145514 49677 237142 49705
rect 145514 49665 145520 49677
rect 237136 49665 237142 49677
rect 237194 49665 237200 49717
rect 211504 49591 211510 49643
rect 211562 49631 211568 49643
rect 226480 49631 226486 49643
rect 211562 49603 226486 49631
rect 211562 49591 211568 49603
rect 226480 49591 226486 49603
rect 226538 49591 226544 49643
rect 220240 49039 220246 49051
rect 218530 49011 220246 49039
rect 208912 48925 208918 48977
rect 208970 48965 208976 48977
rect 218530 48965 218558 49011
rect 220240 48999 220246 49011
rect 220298 48999 220304 49051
rect 509680 48999 509686 49051
rect 509738 49039 509744 49051
rect 525904 49039 525910 49051
rect 509738 49011 525910 49039
rect 509738 48999 509744 49011
rect 525904 48999 525910 49011
rect 525962 48999 525968 49051
rect 208970 48937 218558 48965
rect 208970 48925 208976 48937
rect 218608 48925 218614 48977
rect 218666 48965 218672 48977
rect 645616 48965 645622 48977
rect 218666 48937 645622 48965
rect 218666 48925 218672 48937
rect 645616 48925 645622 48937
rect 645674 48925 645680 48977
rect 210064 48851 210070 48903
rect 210122 48891 210128 48903
rect 220720 48891 220726 48903
rect 210122 48863 220726 48891
rect 210122 48851 210128 48863
rect 220720 48851 220726 48863
rect 220778 48851 220784 48903
rect 501136 48851 501142 48903
rect 501194 48891 501200 48903
rect 507088 48891 507094 48903
rect 501194 48863 507094 48891
rect 501194 48851 501200 48863
rect 507088 48851 507094 48863
rect 507146 48851 507152 48903
rect 208144 48777 208150 48829
rect 208202 48817 208208 48829
rect 220048 48817 220054 48829
rect 208202 48789 220054 48817
rect 208202 48777 208208 48789
rect 220048 48777 220054 48789
rect 220106 48777 220112 48829
rect 220240 48777 220246 48829
rect 220298 48817 220304 48829
rect 223504 48817 223510 48829
rect 220298 48789 223510 48817
rect 220298 48777 220304 48789
rect 223504 48777 223510 48789
rect 223562 48777 223568 48829
rect 208528 48703 208534 48755
rect 208586 48743 208592 48755
rect 221680 48743 221686 48755
rect 208586 48715 221686 48743
rect 208586 48703 208592 48715
rect 221680 48703 221686 48715
rect 221738 48703 221744 48755
rect 222256 48703 222262 48755
rect 222314 48743 222320 48755
rect 645232 48743 645238 48755
rect 222314 48715 645238 48743
rect 222314 48703 222320 48715
rect 645232 48703 645238 48715
rect 645290 48703 645296 48755
rect 209008 48629 209014 48681
rect 209066 48669 209072 48681
rect 222448 48669 222454 48681
rect 209066 48641 222454 48669
rect 209066 48629 209072 48641
rect 222448 48629 222454 48641
rect 222506 48629 222512 48681
rect 222928 48629 222934 48681
rect 222986 48669 222992 48681
rect 645136 48669 645142 48681
rect 222986 48641 645142 48669
rect 222986 48629 222992 48641
rect 645136 48629 645142 48641
rect 645194 48629 645200 48681
rect 188560 48555 188566 48607
rect 188618 48595 188624 48607
rect 239344 48595 239350 48607
rect 188618 48567 239350 48595
rect 188618 48555 188624 48567
rect 239344 48555 239350 48567
rect 239402 48555 239408 48607
rect 185680 48481 185686 48533
rect 185738 48521 185744 48533
rect 240208 48521 240214 48533
rect 185738 48493 240214 48521
rect 185738 48481 185744 48493
rect 240208 48481 240214 48493
rect 240266 48481 240272 48533
rect 194320 48407 194326 48459
rect 194378 48447 194384 48459
rect 239728 48447 239734 48459
rect 194378 48419 239734 48447
rect 194378 48407 194384 48419
rect 239728 48407 239734 48419
rect 239786 48407 239792 48459
rect 197200 48333 197206 48385
rect 197258 48373 197264 48385
rect 239824 48373 239830 48385
rect 197258 48345 239830 48373
rect 197258 48333 197264 48345
rect 239824 48333 239830 48345
rect 239882 48333 239888 48385
rect 162640 48259 162646 48311
rect 162698 48299 162704 48311
rect 241552 48299 241558 48311
rect 162698 48271 241558 48299
rect 162698 48259 162704 48271
rect 241552 48259 241558 48271
rect 241610 48259 241616 48311
rect 149296 48185 149302 48237
rect 149354 48225 149360 48237
rect 209200 48225 209206 48237
rect 149354 48197 209206 48225
rect 149354 48185 149360 48197
rect 209200 48185 209206 48197
rect 209258 48185 209264 48237
rect 209296 48185 209302 48237
rect 209354 48225 209360 48237
rect 222736 48225 222742 48237
rect 209354 48197 222742 48225
rect 209354 48185 209360 48197
rect 222736 48185 222742 48197
rect 222794 48185 222800 48237
rect 224080 48185 224086 48237
rect 224138 48225 224144 48237
rect 645328 48225 645334 48237
rect 224138 48197 645334 48225
rect 224138 48185 224144 48197
rect 645328 48185 645334 48197
rect 645386 48185 645392 48237
rect 149200 48111 149206 48163
rect 149258 48151 149264 48163
rect 208528 48151 208534 48163
rect 149258 48123 208534 48151
rect 149258 48111 149264 48123
rect 208528 48111 208534 48123
rect 208586 48111 208592 48163
rect 208624 48111 208630 48163
rect 208682 48151 208688 48163
rect 222064 48151 222070 48163
rect 208682 48123 222070 48151
rect 208682 48111 208688 48123
rect 222064 48111 222070 48123
rect 222122 48111 222128 48163
rect 148144 48037 148150 48089
rect 148202 48077 148208 48089
rect 219088 48077 219094 48089
rect 148202 48049 219094 48077
rect 148202 48037 148208 48049
rect 219088 48037 219094 48049
rect 219146 48037 219152 48089
rect 149392 47963 149398 48015
rect 149450 48003 149456 48015
rect 221296 48003 221302 48015
rect 149450 47975 221302 48003
rect 149450 47963 149456 47975
rect 221296 47963 221302 47975
rect 221354 47963 221360 48015
rect 149488 47889 149494 47941
rect 149546 47929 149552 47941
rect 220528 47929 220534 47941
rect 149546 47901 220534 47929
rect 149546 47889 149552 47901
rect 220528 47889 220534 47901
rect 220586 47889 220592 47941
rect 149680 47815 149686 47867
rect 149738 47855 149744 47867
rect 219472 47855 219478 47867
rect 149738 47827 219478 47855
rect 149738 47815 149744 47827
rect 219472 47815 219478 47827
rect 219530 47815 219536 47867
rect 149584 47741 149590 47793
rect 149642 47781 149648 47793
rect 220144 47781 220150 47793
rect 149642 47753 220150 47781
rect 149642 47741 149648 47753
rect 220144 47741 220150 47753
rect 220202 47741 220208 47793
rect 147856 47667 147862 47719
rect 147914 47707 147920 47719
rect 218032 47707 218038 47719
rect 147914 47679 218038 47707
rect 147914 47667 147920 47679
rect 218032 47667 218038 47679
rect 218090 47667 218096 47719
rect 147760 47593 147766 47645
rect 147818 47633 147824 47645
rect 217648 47633 217654 47645
rect 147818 47605 217654 47633
rect 147818 47593 147824 47605
rect 217648 47593 217654 47605
rect 217706 47593 217712 47645
rect 148048 47519 148054 47571
rect 148106 47559 148112 47571
rect 218320 47559 218326 47571
rect 148106 47531 218326 47559
rect 148106 47519 148112 47531
rect 218320 47519 218326 47531
rect 218378 47519 218384 47571
rect 623440 47519 623446 47571
rect 623498 47559 623504 47571
rect 640720 47559 640726 47571
rect 623498 47531 640726 47559
rect 623498 47519 623504 47531
rect 640720 47519 640726 47531
rect 640778 47519 640784 47571
rect 147952 47445 147958 47497
rect 148010 47485 148016 47497
rect 218704 47485 218710 47497
rect 148010 47457 218710 47485
rect 148010 47445 148016 47457
rect 218704 47445 218710 47457
rect 218762 47445 218768 47497
rect 177040 47371 177046 47423
rect 177098 47411 177104 47423
rect 238000 47411 238006 47423
rect 177098 47383 238006 47411
rect 177098 47371 177104 47383
rect 238000 47371 238006 47383
rect 238058 47371 238064 47423
rect 179920 47297 179926 47349
rect 179978 47337 179984 47349
rect 238576 47337 238582 47349
rect 179978 47309 238582 47337
rect 179978 47297 179984 47309
rect 238576 47297 238582 47309
rect 238634 47297 238640 47349
rect 200080 47223 200086 47275
rect 200138 47263 200144 47275
rect 238960 47263 238966 47275
rect 200138 47235 238966 47263
rect 200138 47223 200144 47235
rect 238960 47223 238966 47235
rect 239018 47223 239024 47275
rect 148528 47149 148534 47201
rect 148586 47189 148592 47201
rect 230992 47189 230998 47201
rect 148586 47161 230998 47189
rect 148586 47149 148592 47161
rect 230992 47149 230998 47161
rect 231050 47149 231056 47201
rect 148240 47075 148246 47127
rect 148298 47115 148304 47127
rect 236368 47115 236374 47127
rect 148298 47087 236374 47115
rect 148298 47075 148304 47087
rect 236368 47075 236374 47087
rect 236426 47075 236432 47127
rect 149104 47001 149110 47053
rect 149162 47041 149168 47053
rect 233296 47041 233302 47053
rect 149162 47013 233302 47041
rect 149162 47001 149168 47013
rect 233296 47001 233302 47013
rect 233354 47001 233360 47053
rect 149008 46927 149014 46979
rect 149066 46967 149072 46979
rect 234160 46967 234166 46979
rect 149066 46939 234166 46967
rect 149066 46927 149072 46939
rect 234160 46927 234166 46939
rect 234218 46927 234224 46979
rect 148720 46853 148726 46905
rect 148778 46893 148784 46905
rect 229744 46893 229750 46905
rect 148778 46865 229750 46893
rect 148778 46853 148784 46865
rect 229744 46853 229750 46865
rect 229802 46853 229808 46905
rect 148624 46779 148630 46831
rect 148682 46819 148688 46831
rect 230512 46819 230518 46831
rect 148682 46791 230518 46819
rect 148682 46779 148688 46791
rect 230512 46779 230518 46791
rect 230570 46779 230576 46831
rect 148816 46705 148822 46757
rect 148874 46745 148880 46757
rect 228304 46745 228310 46757
rect 148874 46717 228310 46745
rect 148874 46705 148880 46717
rect 228304 46705 228310 46717
rect 228362 46705 228368 46757
rect 209200 46631 209206 46683
rect 209258 46671 209264 46683
rect 223120 46671 223126 46683
rect 209258 46643 223126 46671
rect 209258 46631 209264 46643
rect 223120 46631 223126 46643
rect 223178 46631 223184 46683
rect 148912 46557 148918 46609
rect 148970 46597 148976 46609
rect 227920 46597 227926 46609
rect 148970 46569 227926 46597
rect 148970 46557 148976 46569
rect 227920 46557 227926 46569
rect 227978 46557 227984 46609
rect 148432 46483 148438 46535
rect 148490 46523 148496 46535
rect 233104 46523 233110 46535
rect 148490 46495 233110 46523
rect 148490 46483 148496 46495
rect 233104 46483 233110 46495
rect 233162 46483 233168 46535
rect 208816 46409 208822 46461
rect 208874 46449 208880 46461
rect 224656 46449 224662 46461
rect 208874 46421 224662 46449
rect 208874 46409 208880 46421
rect 224656 46409 224662 46421
rect 224714 46409 224720 46461
rect 208720 46335 208726 46387
rect 208778 46375 208784 46387
rect 224944 46375 224950 46387
rect 208778 46347 224950 46375
rect 208778 46335 208784 46347
rect 224944 46335 224950 46347
rect 225002 46335 225008 46387
rect 208528 46261 208534 46313
rect 208586 46301 208592 46313
rect 224272 46301 224278 46313
rect 208586 46273 224278 46301
rect 208586 46261 208592 46273
rect 224272 46261 224278 46273
rect 224330 46261 224336 46313
rect 191440 46187 191446 46239
rect 191498 46227 191504 46239
rect 240784 46227 240790 46239
rect 191498 46199 240790 46227
rect 191498 46187 191504 46199
rect 240784 46187 240790 46199
rect 240842 46187 240848 46239
rect 206992 46039 206998 46091
rect 207050 46079 207056 46091
rect 465808 46079 465814 46091
rect 207050 46051 465814 46079
rect 207050 46039 207056 46051
rect 465808 46039 465814 46051
rect 465866 46039 465872 46091
rect 384400 45373 384406 45425
rect 384458 45413 384464 45425
rect 388816 45413 388822 45425
rect 384458 45385 388822 45413
rect 384458 45373 384464 45385
rect 388816 45373 388822 45385
rect 388874 45373 388880 45425
rect 212080 45003 212086 45055
rect 212138 45043 212144 45055
rect 297232 45043 297238 45055
rect 212138 45015 297238 45043
rect 212138 45003 212144 45015
rect 297232 45003 297238 45015
rect 297290 45003 297296 45055
rect 211408 44929 211414 44981
rect 211466 44969 211472 44981
rect 361744 44969 361750 44981
rect 211466 44941 361750 44969
rect 211466 44929 211472 44941
rect 361744 44929 361750 44941
rect 361802 44929 361808 44981
rect 213904 44855 213910 44907
rect 213962 44895 213968 44907
rect 455728 44895 455734 44907
rect 213962 44867 455734 44895
rect 213962 44855 213968 44867
rect 455728 44855 455734 44867
rect 455786 44855 455792 44907
rect 211696 44781 211702 44833
rect 211754 44821 211760 44833
rect 362800 44821 362806 44833
rect 211754 44793 362806 44821
rect 211754 44781 211760 44793
rect 362800 44781 362806 44793
rect 362858 44781 362864 44833
rect 212464 44633 212470 44685
rect 212522 44673 212528 44685
rect 310096 44673 310102 44685
rect 212522 44645 310102 44673
rect 212522 44633 212528 44645
rect 310096 44633 310102 44645
rect 310154 44633 310160 44685
rect 507088 43301 507094 43353
rect 507146 43341 507152 43353
rect 507146 43313 520382 43341
rect 507146 43301 507152 43313
rect 215056 43227 215062 43279
rect 215114 43267 215120 43279
rect 518704 43267 518710 43279
rect 215114 43239 518710 43267
rect 215114 43227 215120 43239
rect 518704 43227 518710 43239
rect 518762 43227 518768 43279
rect 520354 43205 520382 43313
rect 520336 43153 520342 43205
rect 520394 43153 520400 43205
rect 206896 42265 206902 42317
rect 206954 42305 206960 42317
rect 405520 42305 405526 42317
rect 206954 42277 405526 42305
rect 206954 42265 206960 42277
rect 405520 42265 405526 42277
rect 405578 42265 405584 42317
rect 213616 42191 213622 42243
rect 213674 42231 213680 42243
rect 460048 42231 460054 42243
rect 213674 42203 460054 42231
rect 213674 42191 213680 42203
rect 460048 42191 460054 42203
rect 460106 42191 460112 42243
rect 214288 42117 214294 42169
rect 214346 42157 214352 42169
rect 514864 42157 514870 42169
rect 214346 42129 514870 42157
rect 214346 42117 214352 42129
rect 514864 42117 514870 42129
rect 514922 42117 514928 42169
rect 404368 41525 404374 41577
rect 404426 41565 404432 41577
rect 409378 41565 409406 41786
rect 404426 41537 409406 41565
rect 404426 41525 404432 41537
rect 334096 40859 334102 40911
rect 334154 40899 334160 40911
rect 344176 40899 344182 40911
rect 334154 40871 344182 40899
rect 334154 40859 334160 40871
rect 344176 40859 344182 40871
rect 344234 40859 344240 40911
rect 388816 40267 388822 40319
rect 388874 40307 388880 40319
rect 394576 40307 394582 40319
rect 388874 40279 394582 40307
rect 388874 40267 388880 40279
rect 394576 40267 394582 40279
rect 394634 40267 394640 40319
rect 394576 37381 394582 37433
rect 394634 37421 394640 37433
rect 404368 37421 404374 37433
rect 394634 37393 404374 37421
rect 394634 37381 394640 37393
rect 404368 37381 404374 37393
rect 404426 37381 404432 37433
<< via1 >>
rect 434998 1008039 435050 1008091
rect 470806 1008039 470858 1008091
rect 434710 1005523 434762 1005575
rect 472150 1005523 472202 1005575
rect 367222 1005375 367274 1005427
rect 383638 1005375 383690 1005427
rect 434902 1005375 434954 1005427
rect 459286 1005375 459338 1005427
rect 436918 1005301 436970 1005353
rect 471382 1005301 471434 1005353
rect 164278 1005227 164330 1005279
rect 172822 1005227 172874 1005279
rect 316822 1005227 316874 1005279
rect 331222 1005227 331274 1005279
rect 434614 1005227 434666 1005279
rect 472246 1005227 472298 1005279
rect 218806 1005153 218858 1005205
rect 222742 1005153 222794 1005205
rect 434806 1005153 434858 1005205
rect 443734 1005153 443786 1005205
rect 443542 1003673 443594 1003725
rect 463798 1003673 463850 1003725
rect 377686 1003229 377738 1003281
rect 467062 1003229 467114 1003281
rect 160438 1003155 160490 1003207
rect 164278 1003155 164330 1003207
rect 211798 1003155 211850 1003207
rect 213814 1003155 213866 1003207
rect 359062 1003155 359114 1003207
rect 362518 1003155 362570 1003207
rect 367222 1003155 367274 1003207
rect 426070 1003155 426122 1003207
rect 429238 1003155 429290 1003207
rect 434614 1003155 434666 1003207
rect 439222 1003155 439274 1003207
rect 466582 1003155 466634 1003207
rect 518614 1003229 518666 1003281
rect 449206 1003081 449258 1003133
rect 467830 1003081 467882 1003133
rect 502390 1003081 502442 1003133
rect 425398 1003007 425450 1003059
rect 430198 1003007 430250 1003059
rect 430294 1003007 430346 1003059
rect 434902 1003007 434954 1003059
rect 439126 1003007 439178 1003059
rect 463510 1003007 463562 1003059
rect 501334 1003007 501386 1003059
rect 518806 1003155 518858 1003207
rect 502966 1003081 503018 1003133
rect 518710 1003081 518762 1003133
rect 504022 1003007 504074 1003059
rect 518422 1003007 518474 1003059
rect 424342 1002933 424394 1002985
rect 463606 1002933 463658 1002985
rect 554902 1002933 554954 1002985
rect 573046 1002933 573098 1002985
rect 299350 1002859 299402 1002911
rect 308854 1002859 308906 1002911
rect 428758 1002859 428810 1002911
rect 434710 1002859 434762 1002911
rect 161494 1002785 161546 1002837
rect 169942 1002785 169994 1002837
rect 299446 1002785 299498 1002837
rect 309334 1002785 309386 1002837
rect 428278 1002785 428330 1002837
rect 434806 1002785 434858 1002837
rect 554326 1002785 554378 1002837
rect 572854 1002785 572906 1002837
rect 299254 1002711 299306 1002763
rect 308278 1002711 308330 1002763
rect 423766 1002711 423818 1002763
rect 439126 1002711 439178 1002763
rect 424822 1002637 424874 1002689
rect 439222 1002637 439274 1002689
rect 361270 1002563 361322 1002615
rect 368854 1002563 368906 1002615
rect 427702 1002563 427754 1002615
rect 435190 1002563 435242 1002615
rect 553750 1002563 553802 1002615
rect 572950 1002563 573002 1002615
rect 361846 1002489 361898 1002541
rect 368662 1002489 368714 1002541
rect 426646 1002489 426698 1002541
rect 435094 1002489 435146 1002541
rect 143734 1002341 143786 1002393
rect 151126 1002415 151178 1002467
rect 427126 1002415 427178 1002467
rect 443638 1002415 443690 1002467
rect 146806 1002341 146858 1002393
rect 152758 1002341 152810 1002393
rect 143926 1002267 143978 1002319
rect 175702 1002267 175754 1002319
rect 255478 1002341 255530 1002393
rect 363478 1002341 363530 1002393
rect 377110 1002341 377162 1002393
rect 431926 1002341 431978 1002393
rect 434998 1002341 435050 1002393
rect 503446 1002341 503498 1002393
rect 514006 1002341 514058 1002393
rect 553270 1002341 553322 1002393
rect 567478 1002341 567530 1002393
rect 246646 1002267 246698 1002319
rect 253846 1002267 253898 1002319
rect 362902 1002267 362954 1002319
rect 368758 1002267 368810 1002319
rect 377686 1002267 377738 1002319
rect 383446 1002267 383498 1002319
rect 430198 1002267 430250 1002319
rect 449206 1002267 449258 1002319
rect 489526 1002267 489578 1002319
rect 519862 1002267 519914 1002319
rect 555382 1002267 555434 1002319
rect 567382 1002267 567434 1002319
rect 246550 1002193 246602 1002245
rect 506230 1001453 506282 1001505
rect 518518 1001453 518570 1001505
rect 557782 1001305 557834 1001357
rect 571030 1001305 571082 1001357
rect 465718 1001009 465770 1001061
rect 472630 1001009 472682 1001061
rect 443638 1000935 443690 1000987
rect 472438 1000935 472490 1000987
rect 507862 1000935 507914 1000987
rect 512662 1000935 512714 1000987
rect 356374 1000861 356426 1000913
rect 377206 1000861 377258 1000913
rect 429910 1000861 429962 1000913
rect 472630 1000861 472682 1000913
rect 552310 1000861 552362 1000913
rect 573238 1000861 573290 1000913
rect 143830 1000787 143882 1000839
rect 157654 1000787 157706 1000839
rect 195190 1000787 195242 1000839
rect 209110 1000787 209162 1000839
rect 360214 1000787 360266 1000839
rect 383638 1000787 383690 1000839
rect 430966 1000787 431018 1000839
rect 472534 1000787 472586 1000839
rect 500758 1000787 500810 1000839
rect 523318 1000787 523370 1000839
rect 552982 1000787 553034 1000839
rect 575158 1000787 575210 1000839
rect 506902 1000639 506954 1000691
rect 512086 1000639 512138 1000691
rect 610678 999751 610730 999803
rect 625846 999751 625898 999803
rect 502006 999677 502058 999729
rect 512086 999677 512138 999729
rect 609046 999677 609098 999729
rect 625750 999677 625802 999729
rect 247030 999603 247082 999655
rect 258838 999603 258890 999655
rect 610582 999603 610634 999655
rect 625654 999603 625706 999655
rect 246742 999529 246794 999581
rect 258358 999529 258410 999581
rect 298294 999529 298346 999581
rect 312118 999529 312170 999581
rect 504694 999529 504746 999581
rect 512086 999529 512138 999581
rect 596278 999529 596330 999581
rect 625558 999529 625610 999581
rect 92566 999455 92618 999507
rect 92374 999381 92426 999433
rect 106294 999381 106346 999433
rect 143734 999455 143786 999507
rect 155542 999455 155594 999507
rect 246838 999455 246890 999507
rect 260470 999455 260522 999507
rect 298390 999455 298442 999507
rect 310486 999455 310538 999507
rect 593302 999455 593354 999507
rect 625846 999455 625898 999507
rect 126646 999381 126698 999433
rect 144022 999381 144074 999433
rect 146806 999381 146858 999433
rect 195094 999381 195146 999433
rect 206902 999381 206954 999433
rect 246934 999381 246986 999433
rect 279286 999381 279338 999433
rect 298102 999381 298154 999433
rect 309910 999381 309962 999433
rect 357142 999381 357194 999433
rect 313750 999307 313802 999359
rect 331126 999307 331178 999359
rect 377110 999381 377162 999433
rect 383542 999381 383594 999433
rect 459286 999381 459338 999433
rect 383158 999307 383210 999359
rect 500182 999381 500234 999433
rect 515830 999381 515882 999433
rect 596182 999381 596234 999433
rect 625462 999381 625514 999433
rect 464758 999307 464810 999359
rect 302998 999233 303050 999285
rect 304342 999233 304394 999285
rect 304918 999233 304970 999285
rect 364534 999159 364586 999211
rect 380182 999159 380234 999211
rect 557206 999085 557258 999137
rect 573814 999085 573866 999137
rect 558838 998937 558890 998989
rect 573526 998937 573578 998989
rect 368854 998641 368906 998693
rect 374518 998641 374570 998693
rect 377206 997827 377258 997879
rect 383062 997827 383114 997879
rect 314806 997679 314858 997731
rect 365206 997679 365258 997731
rect 555958 997679 556010 997731
rect 593302 997679 593354 997731
rect 331126 997605 331178 997657
rect 364534 997605 364586 997657
rect 567478 997605 567530 997657
rect 596182 997605 596234 997657
rect 567382 997531 567434 997583
rect 596278 997531 596330 997583
rect 571030 997457 571082 997509
rect 610582 997457 610634 997509
rect 558166 997383 558218 997435
rect 609046 997383 609098 997435
rect 559414 997309 559466 997361
rect 610678 997309 610730 997361
rect 463510 997161 463562 997213
rect 465334 997161 465386 997213
rect 298102 997087 298154 997139
rect 313750 997087 313802 997139
rect 368758 997087 368810 997139
rect 377110 997087 377162 997139
rect 507286 996569 507338 996621
rect 523414 996569 523466 996621
rect 144118 996495 144170 996547
rect 156022 996495 156074 996547
rect 195766 996495 195818 996547
rect 205270 996495 205322 996547
rect 247126 996495 247178 996547
rect 259990 996495 260042 996547
rect 368662 996495 368714 996547
rect 377206 996495 377258 996547
rect 505654 996495 505706 996547
rect 521206 996495 521258 996547
rect 210166 996421 210218 996473
rect 225430 996421 225482 996473
rect 313174 996421 313226 996473
rect 363958 996421 364010 996473
rect 280246 996199 280298 996251
rect 107926 996125 107978 996177
rect 159766 996125 159818 996177
rect 178486 996125 178538 996177
rect 198646 996125 198698 996177
rect 204022 996125 204074 996177
rect 107542 996051 107594 996103
rect 159190 996051 159242 996103
rect 210166 996051 210218 996103
rect 262102 996125 262154 996177
rect 263062 996125 263114 996177
rect 314806 996125 314858 996177
rect 368662 996125 368714 996177
rect 432598 996199 432650 996251
rect 508342 996199 508394 996251
rect 432502 996125 432554 996177
rect 509590 996125 509642 996177
rect 225430 996051 225482 996103
rect 262006 996051 262058 996103
rect 313174 996051 313226 996103
rect 380182 996051 380234 996103
rect 434998 996051 435050 996103
rect 470806 996051 470858 996103
rect 508534 996051 508586 996103
rect 518422 996125 518474 996177
rect 561046 996125 561098 996177
rect 559798 996051 559850 996103
rect 108982 995977 109034 996029
rect 160438 995977 160490 996029
rect 178486 995977 178538 996029
rect 210646 995977 210698 996029
rect 222742 995977 222794 996029
rect 263254 995977 263306 996029
rect 94966 995903 95018 995955
rect 102934 995903 102986 995955
rect 146806 995903 146858 995955
rect 152086 995903 152138 995955
rect 172822 995903 172874 995955
rect 211798 995903 211850 995955
rect 97846 995829 97898 995881
rect 144022 995829 144074 995881
rect 82294 995755 82346 995807
rect 91510 995755 91562 995807
rect 92278 995755 92330 995807
rect 93526 995755 93578 995807
rect 97942 995755 97994 995807
rect 137398 995755 137450 995807
rect 137974 995755 138026 995807
rect 143638 995755 143690 995807
rect 149590 995755 149642 995807
rect 154870 995755 154922 995807
rect 183766 995755 183818 995807
rect 198646 995829 198698 995881
rect 202486 995829 202538 995881
rect 254518 995829 254570 995881
rect 299446 995977 299498 996029
rect 363958 995977 364010 996029
rect 430966 995977 431018 996029
rect 436918 995977 436970 996029
rect 560182 995977 560234 996029
rect 471382 995903 471434 995955
rect 508342 995903 508394 995955
rect 510550 995903 510602 995955
rect 515734 995903 515786 995955
rect 523702 995903 523754 995955
rect 299254 995829 299306 995881
rect 383446 995829 383498 995881
rect 472438 995829 472490 995881
rect 523894 995829 523946 995881
rect 561910 995903 561962 995955
rect 569782 995903 569834 995955
rect 625462 995903 625514 995955
rect 625654 995829 625706 995881
rect 205654 995755 205706 995807
rect 239542 995755 239594 995807
rect 240886 995755 240938 995807
rect 246646 995755 246698 995807
rect 246934 995755 246986 995807
rect 257686 995755 257738 995807
rect 283798 995755 283850 995807
rect 290710 995755 290762 995807
rect 291190 995755 291242 995807
rect 306070 995755 306122 995807
rect 366742 995755 366794 995807
rect 371638 995755 371690 995807
rect 383638 995755 383690 995807
rect 384982 995755 385034 995807
rect 388822 995755 388874 995807
rect 472630 995755 472682 995807
rect 473302 995755 473354 995807
rect 476950 995755 477002 995807
rect 511126 995755 511178 995807
rect 515638 995755 515690 995807
rect 524182 995755 524234 995807
rect 525334 995755 525386 995807
rect 528406 995755 528458 995807
rect 529846 995755 529898 995807
rect 559798 995755 559850 995807
rect 564598 995755 564650 995807
rect 625846 995755 625898 995807
rect 627094 995755 627146 995807
rect 629590 995755 629642 995807
rect 631510 995755 631562 995807
rect 89782 995681 89834 995733
rect 92374 995681 92426 995733
rect 136726 995681 136778 995733
rect 151702 995681 151754 995733
rect 175702 995681 175754 995733
rect 185206 995681 185258 995733
rect 194422 995681 194474 995733
rect 195094 995681 195146 995733
rect 198454 995681 198506 995733
rect 202966 995681 203018 995733
rect 240310 995681 240362 995733
rect 246550 995681 246602 995733
rect 247606 995681 247658 995733
rect 256150 995681 256202 995733
rect 291766 995681 291818 995733
rect 306454 995681 306506 995733
rect 366166 995681 366218 995733
rect 371734 995681 371786 995733
rect 383542 995681 383594 995733
rect 386038 995681 386090 995733
rect 472534 995681 472586 995733
rect 474646 995681 474698 995733
rect 523990 995681 524042 995733
rect 524758 995681 524810 995733
rect 625750 995681 625802 995733
rect 626518 995681 626570 995733
rect 93814 995607 93866 995659
rect 98998 995607 99050 995659
rect 142966 995607 143018 995659
rect 143734 995607 143786 995659
rect 192502 995607 192554 995659
rect 195190 995607 195242 995659
rect 297334 995607 297386 995659
rect 298006 995607 298058 995659
rect 383734 995607 383786 995659
rect 384406 995607 384458 995659
rect 472726 995607 472778 995659
rect 474070 995607 474122 995659
rect 141046 995533 141098 995585
rect 143830 995533 143882 995585
rect 185110 995533 185162 995585
rect 198646 995533 198698 995585
rect 286774 995533 286826 995585
rect 81622 995459 81674 995511
rect 102454 995459 102506 995511
rect 184054 995459 184106 995511
rect 195766 995459 195818 995511
rect 245686 995459 245738 995511
rect 246742 995459 246794 995511
rect 287446 995459 287498 995511
rect 290710 995459 290762 995511
rect 295414 995533 295466 995585
rect 298294 995533 298346 995585
rect 383158 995533 383210 995585
rect 392374 995533 392426 995585
rect 466582 995533 466634 995585
rect 478390 995607 478442 995659
rect 523798 995607 523850 995659
rect 526102 995607 526154 995659
rect 560182 995607 560234 995659
rect 564502 995607 564554 995659
rect 625558 995607 625610 995659
rect 630166 995607 630218 995659
rect 523606 995533 523658 995585
rect 527830 995533 527882 995585
rect 625942 995533 625994 995585
rect 627862 995533 627914 995585
rect 299350 995459 299402 995511
rect 518806 995459 518858 995511
rect 532822 995459 532874 995511
rect 287926 995385 287978 995437
rect 306550 995385 306602 995437
rect 383158 995385 383210 995437
rect 390454 995385 390506 995437
rect 403126 995385 403178 995437
rect 518614 995385 518666 995437
rect 533398 995385 533450 995437
rect 518710 995311 518762 995363
rect 535558 995311 535610 995363
rect 523414 995237 523466 995289
rect 537382 995237 537434 995289
rect 523318 995163 523370 995215
rect 534358 995163 534410 995215
rect 66838 995089 66890 995141
rect 349654 995089 349706 995141
rect 519862 995089 519914 995141
rect 530710 995089 530762 995141
rect 532726 995089 532778 995141
rect 555382 995089 555434 995141
rect 649366 995089 649418 995141
rect 233302 995015 233354 995067
rect 247798 995015 247850 995067
rect 279286 995015 279338 995067
rect 609046 995015 609098 995067
rect 524086 994645 524138 994697
rect 531190 994645 531242 994697
rect 290902 994275 290954 994327
rect 299158 994275 299210 994327
rect 463702 994127 463754 994179
rect 479158 994127 479210 994179
rect 235798 993979 235850 994031
rect 247606 993979 247658 994031
rect 180502 993905 180554 993957
rect 198646 993905 198698 993957
rect 234934 993905 234986 993957
rect 250486 993905 250538 993957
rect 77686 993831 77738 993883
rect 97846 993831 97898 993883
rect 132118 993831 132170 993883
rect 149686 993831 149738 993883
rect 182998 993831 183050 993883
rect 208150 993831 208202 993883
rect 232150 993831 232202 993883
rect 246934 993831 246986 993883
rect 561622 993831 561674 993883
rect 641014 993831 641066 993883
rect 80182 993757 80234 993809
rect 105334 993757 105386 993809
rect 129334 993757 129386 993809
rect 149590 993757 149642 993809
rect 181366 993757 181418 993809
rect 209782 993757 209834 993809
rect 231478 993757 231530 993809
rect 247126 993757 247178 993809
rect 521302 993757 521354 993809
rect 538966 993757 539018 993809
rect 78358 993683 78410 993735
rect 106966 993683 107018 993735
rect 128470 993683 128522 993735
rect 157270 993683 157322 993735
rect 179830 993683 179882 993735
rect 208726 993683 208778 993735
rect 234358 993683 234410 993735
rect 259414 993683 259466 993735
rect 282838 993683 282890 993735
rect 311542 993683 311594 993735
rect 374518 993683 374570 993735
rect 392086 993683 392138 993735
rect 532726 993683 532778 993735
rect 632374 993683 632426 993735
rect 77302 993609 77354 993661
rect 105910 993609 105962 993661
rect 129718 993609 129770 993661
rect 158230 993609 158282 993661
rect 185398 993609 185450 993661
rect 236758 993609 236810 993661
rect 61846 993535 61898 993587
rect 82582 993535 82634 993587
rect 133942 993535 133994 993587
rect 143926 993535 143978 993587
rect 62038 993461 62090 993513
rect 83446 993461 83498 993513
rect 92566 993461 92618 993513
rect 284374 993609 284426 993661
rect 312790 993609 312842 993661
rect 365782 993609 365834 993661
rect 398806 993609 398858 993661
rect 443734 993609 443786 993661
rect 487798 993609 487850 993661
rect 531190 993609 531242 993661
rect 633046 993609 633098 993661
rect 328246 993535 328298 993587
rect 288118 993387 288170 993439
rect 328438 993387 328490 993439
rect 348406 993461 348458 993513
rect 348502 993387 348554 993439
rect 408982 993461 409034 993513
rect 423382 993535 423434 993587
rect 443446 993461 443498 993513
rect 449206 993461 449258 993513
rect 642262 993461 642314 993513
rect 650326 993461 650378 993513
rect 403126 993387 403178 993439
rect 408886 993387 408938 993439
rect 449398 993387 449450 993439
rect 463702 993387 463754 993439
rect 479158 993387 479210 993439
rect 489526 993387 489578 993439
rect 362902 993313 362954 993365
rect 382966 993313 383018 993365
rect 383062 993239 383114 993291
rect 422134 992721 422186 992773
rect 426262 992721 426314 992773
rect 73462 992129 73514 992181
rect 110230 992129 110282 992181
rect 604726 991907 604778 991959
rect 605782 991907 605834 991959
rect 605782 991611 605834 991663
rect 619798 991611 619850 991663
rect 105814 990427 105866 990479
rect 109558 990427 109610 990479
rect 371638 989391 371690 989443
rect 397846 989391 397898 989443
rect 437782 989391 437834 989443
rect 462742 989391 462794 989443
rect 515638 989391 515690 989443
rect 527638 989391 527690 989443
rect 569686 989391 569738 989443
rect 592438 989391 592490 989443
rect 154486 989317 154538 989369
rect 161686 989317 161738 989369
rect 203158 989317 203210 989369
rect 213334 989317 213386 989369
rect 270742 989317 270794 989369
rect 284278 989317 284330 989369
rect 319606 989317 319658 989369
rect 349174 989317 349226 989369
rect 371542 989317 371594 989369
rect 414070 989317 414122 989369
rect 437878 989317 437930 989369
rect 478966 989317 479018 989369
rect 515542 989317 515594 989369
rect 543766 989317 543818 989369
rect 569878 989317 569930 989369
rect 608758 989317 608810 989369
rect 89590 989243 89642 989295
rect 109366 989243 109418 989295
rect 138262 989243 138314 989295
rect 161494 989243 161546 989295
rect 216022 989243 216074 989295
rect 235606 989243 235658 989295
rect 267862 989243 267914 989295
rect 300502 989243 300554 989295
rect 319702 989243 319754 989295
rect 365398 989243 365450 989295
rect 371734 989243 371786 989295
rect 430294 989243 430346 989295
rect 437974 989243 438026 989295
rect 495190 989243 495242 989295
rect 515734 989243 515786 989295
rect 560086 989243 560138 989295
rect 569782 989243 569834 989295
rect 624982 989243 625034 989295
rect 634294 989243 634346 989295
rect 649846 989243 649898 989295
rect 64822 988503 64874 988555
rect 66838 988503 66890 988555
rect 50422 988281 50474 988333
rect 122038 988281 122090 988333
rect 331222 988281 331274 988333
rect 332566 988281 332618 988333
rect 47638 988207 47690 988259
rect 186934 988207 186986 988259
rect 44758 988133 44810 988185
rect 251830 988133 251882 988185
rect 44854 988059 44906 988111
rect 316726 988059 316778 988111
rect 44950 987985 45002 988037
rect 381622 987985 381674 988037
rect 45046 987911 45098 987963
rect 446518 987911 446570 987963
rect 43126 987837 43178 987889
rect 511414 987837 511466 987889
rect 65110 986727 65162 986779
rect 93526 986727 93578 986779
rect 47542 986653 47594 986705
rect 109174 986653 109226 986705
rect 619798 986653 619850 986705
rect 650230 986653 650282 986705
rect 47446 986579 47498 986631
rect 107542 986579 107594 986631
rect 609046 986579 609098 986631
rect 650134 986579 650186 986631
rect 44566 986505 44618 986557
rect 107926 986505 107978 986557
rect 564502 986505 564554 986557
rect 658006 986505 658058 986557
rect 65206 986431 65258 986483
rect 145366 986431 145418 986483
rect 565846 986431 565898 986483
rect 658102 986431 658154 986483
rect 65014 986357 65066 986409
rect 197206 986357 197258 986409
rect 267862 986357 267914 986409
rect 290902 986357 290954 986409
rect 564598 986357 564650 986409
rect 660886 986357 660938 986409
rect 225526 984951 225578 985003
rect 233206 984951 233258 985003
rect 632374 983693 632426 983745
rect 674518 983693 674570 983745
rect 633046 983619 633098 983671
rect 674326 983619 674378 983671
rect 64726 983545 64778 983597
rect 225526 983545 225578 983597
rect 515830 983545 515882 983597
rect 649558 983545 649610 983597
rect 64918 983471 64970 983523
rect 267862 983471 267914 983523
rect 426262 983471 426314 983523
rect 649462 983471 649514 983523
rect 53686 973481 53738 973533
rect 59446 973481 59498 973533
rect 42166 967265 42218 967317
rect 43126 967265 43178 967317
rect 42166 960901 42218 960953
rect 42838 960901 42890 960953
rect 42742 959051 42794 959103
rect 59542 959051 59594 959103
rect 675094 958385 675146 958437
rect 675382 958385 675434 958437
rect 675190 956979 675242 957031
rect 675478 956979 675530 957031
rect 669526 954685 669578 954737
rect 675382 954685 675434 954737
rect 674134 953871 674186 953923
rect 675478 953871 675530 953923
rect 42166 953205 42218 953257
rect 42454 953205 42506 953257
rect 674038 952021 674090 952073
rect 675478 952021 675530 952073
rect 42646 944621 42698 944673
rect 59542 944621 59594 944673
rect 42646 944251 42698 944303
rect 48886 944251 48938 944303
rect 42646 942697 42698 942749
rect 47542 942697 47594 942749
rect 39958 942179 40010 942231
rect 42646 942179 42698 942231
rect 44566 942179 44618 942231
rect 658102 939515 658154 939567
rect 674422 939515 674474 939567
rect 655318 939367 655370 939419
rect 674614 939367 674666 939419
rect 655222 939219 655274 939271
rect 676822 939219 676874 939271
rect 655126 939071 655178 939123
rect 676918 939071 676970 939123
rect 660886 937961 660938 938013
rect 674422 937961 674474 938013
rect 658006 936111 658058 936163
rect 676822 936111 676874 936163
rect 39958 933077 40010 933129
rect 40150 933077 40202 933129
rect 42646 932115 42698 932167
rect 53206 932115 53258 932167
rect 48886 930487 48938 930539
rect 59542 930487 59594 930539
rect 654454 927453 654506 927505
rect 666742 927453 666794 927505
rect 649654 927379 649706 927431
rect 677014 927379 677066 927431
rect 47446 915835 47498 915887
rect 59542 915835 59594 915887
rect 653974 915835 654026 915887
rect 660982 915835 661034 915887
rect 39862 907177 39914 907229
rect 40246 907177 40298 907229
rect 654454 904365 654506 904417
rect 663958 904365 664010 904417
rect 53302 901479 53354 901531
rect 59542 901479 59594 901531
rect 40246 892821 40298 892873
rect 40054 892747 40106 892799
rect 50518 887123 50570 887175
rect 59542 887123 59594 887175
rect 40054 886975 40106 887027
rect 40150 886975 40202 887027
rect 653974 881277 654026 881329
rect 660886 881277 660938 881329
rect 40150 872693 40202 872745
rect 41686 872619 41738 872671
rect 59542 872619 59594 872671
rect 40150 872471 40202 872523
rect 674614 872101 674666 872153
rect 675478 872101 675530 872153
rect 675094 871435 675146 871487
rect 675382 871435 675434 871487
rect 654454 869807 654506 869859
rect 663766 869807 663818 869859
rect 674422 868993 674474 869045
rect 675190 868993 675242 869045
rect 673366 866921 673418 866973
rect 675190 866921 675242 866973
rect 674518 866477 674570 866529
rect 675382 866477 675434 866529
rect 674326 864997 674378 865049
rect 675094 864997 675146 865049
rect 666646 864035 666698 864087
rect 675190 864035 675242 864087
rect 39862 863961 39914 864013
rect 40150 863961 40202 864013
rect 674422 862037 674474 862089
rect 674902 862037 674954 862089
rect 674998 861075 675050 861127
rect 675190 861075 675242 861127
rect 50326 858263 50378 858315
rect 58582 858263 58634 858315
rect 654166 858263 654218 858315
rect 661078 858263 661130 858315
rect 39862 843833 39914 843885
rect 40054 843833 40106 843885
rect 53398 843833 53450 843885
rect 59542 843833 59594 843885
rect 653974 835175 654026 835227
rect 666838 835175 666890 835227
rect 40054 832511 40106 832563
rect 40246 832215 40298 832267
rect 50614 829477 50666 829529
rect 59542 829477 59594 829529
rect 653974 823705 654026 823757
rect 669814 823705 669866 823757
rect 42646 819117 42698 819169
rect 50518 819117 50570 819169
rect 42646 818081 42698 818133
rect 53302 818081 53354 818133
rect 47542 815047 47594 815099
rect 59542 815047 59594 815099
rect 37366 814973 37418 815025
rect 40246 814973 40298 815025
rect 654454 812161 654506 812213
rect 664054 812161 664106 812213
rect 41974 802393 42026 802445
rect 42934 802393 42986 802445
rect 41782 802171 41834 802223
rect 41974 802171 42026 802223
rect 42742 800839 42794 800891
rect 43414 800839 43466 800891
rect 44662 800617 44714 800669
rect 59542 800617 59594 800669
rect 674998 800617 675050 800669
rect 675190 800617 675242 800669
rect 41878 800247 41930 800299
rect 42166 800247 42218 800299
rect 43510 800247 43562 800299
rect 41782 800173 41834 800225
rect 43318 800173 43370 800225
rect 41878 799951 41930 800003
rect 42166 798101 42218 798153
rect 42646 798101 42698 798153
rect 42550 797583 42602 797635
rect 43414 797583 43466 797635
rect 42070 797287 42122 797339
rect 45046 797287 45098 797339
rect 42166 796251 42218 796303
rect 43030 796251 43082 796303
rect 43030 796103 43082 796155
rect 43318 796103 43370 796155
rect 42166 794993 42218 795045
rect 42838 794993 42890 795045
rect 42070 794253 42122 794305
rect 42454 794253 42506 794305
rect 42166 793809 42218 793861
rect 43126 793809 43178 793861
rect 43126 793661 43178 793713
rect 43510 793661 43562 793713
rect 42166 793143 42218 793195
rect 42934 793143 42986 793195
rect 42550 792921 42602 792973
rect 43030 792921 43082 792973
rect 42166 790479 42218 790531
rect 42550 790479 42602 790531
rect 42166 789887 42218 789939
rect 43126 789887 43178 789939
rect 42166 789443 42218 789495
rect 42550 789443 42602 789495
rect 42166 788703 42218 788755
rect 42838 788703 42890 788755
rect 42166 787001 42218 787053
rect 43030 787001 43082 787053
rect 42166 786409 42218 786461
rect 42358 786409 42410 786461
rect 45046 786261 45098 786313
rect 59542 786261 59594 786313
rect 654070 786261 654122 786313
rect 669718 786261 669770 786313
rect 42070 785595 42122 785647
rect 42454 785595 42506 785647
rect 672502 783449 672554 783501
rect 675382 783449 675434 783501
rect 672982 783079 673034 783131
rect 675094 783079 675146 783131
rect 675478 783079 675530 783131
rect 673270 782931 673322 782983
rect 675382 782931 675434 782983
rect 674998 782487 675050 782539
rect 675478 782487 675530 782539
rect 663862 780489 663914 780541
rect 675094 780489 675146 780541
rect 673078 779749 673130 779801
rect 675382 779749 675434 779801
rect 672886 779305 672938 779357
rect 675478 779305 675530 779357
rect 673174 778565 673226 778617
rect 675382 778565 675434 778617
rect 672598 777603 672650 777655
rect 675478 777603 675530 777655
rect 675094 777011 675146 777063
rect 675382 777011 675434 777063
rect 42454 776049 42506 776101
rect 50614 776049 50666 776101
rect 674422 775457 674474 775509
rect 675382 775457 675434 775509
rect 42838 775309 42890 775361
rect 47542 775309 47594 775361
rect 42838 774791 42890 774843
rect 53398 774791 53450 774843
rect 654070 774717 654122 774769
rect 672406 774717 672458 774769
rect 674134 773607 674186 773659
rect 675478 773607 675530 773659
rect 53398 771831 53450 771883
rect 59542 771831 59594 771883
rect 653974 763247 654026 763299
rect 661174 763247 661226 763299
rect 660982 762877 661034 762929
rect 674326 762877 674378 762929
rect 666742 762285 666794 762337
rect 674326 762285 674378 762337
rect 663958 761989 664010 762041
rect 674614 761989 674666 762041
rect 672310 760435 672362 760487
rect 673846 760435 673898 760487
rect 42934 757549 42986 757601
rect 43606 757549 43658 757601
rect 44950 757475 45002 757527
rect 53590 757475 53642 757527
rect 59542 757475 59594 757527
rect 42934 757401 42986 757453
rect 41686 757253 41738 757305
rect 43510 757253 43562 757305
rect 41782 757031 41834 757083
rect 43318 757031 43370 757083
rect 42166 756735 42218 756787
rect 42358 756735 42410 756787
rect 42934 754219 42986 754271
rect 42166 754071 42218 754123
rect 42070 753035 42122 753087
rect 43126 753035 43178 753087
rect 42838 751629 42890 751681
rect 43510 751629 43562 751681
rect 42070 749779 42122 749831
rect 42838 749779 42890 749831
rect 649750 748817 649802 748869
rect 677014 748817 677066 748869
rect 42166 747263 42218 747315
rect 43126 747263 43178 747315
rect 42166 746893 42218 746945
rect 43606 746893 43658 746945
rect 42070 746227 42122 746279
rect 42742 746227 42794 746279
rect 672982 745931 673034 745983
rect 675094 745931 675146 745983
rect 42166 745487 42218 745539
rect 43030 745487 43082 745539
rect 674134 745413 674186 745465
rect 674518 745413 674570 745465
rect 42166 743785 42218 743837
rect 42838 743785 42890 743837
rect 42070 743193 42122 743245
rect 42742 743193 42794 743245
rect 53494 743045 53546 743097
rect 59542 743045 59594 743097
rect 42166 742379 42218 742431
rect 43126 742379 43178 742431
rect 653974 740159 654026 740211
rect 663958 740159 664010 740211
rect 672790 738087 672842 738139
rect 675094 738087 675146 738139
rect 675478 738087 675530 738139
rect 672694 737865 672746 737917
rect 675382 737865 675434 737917
rect 675190 737643 675242 737695
rect 675382 737643 675434 737695
rect 660982 737273 661034 737325
rect 675094 737273 675146 737325
rect 674230 735423 674282 735475
rect 675478 735423 675530 735475
rect 673366 734905 673418 734957
rect 675382 734905 675434 734957
rect 672982 733573 673034 733625
rect 675478 733573 675530 733625
rect 42742 732685 42794 732737
rect 53398 732685 53450 732737
rect 674902 732315 674954 732367
rect 675478 732315 675530 732367
rect 42742 732093 42794 732145
rect 53590 732093 53642 732145
rect 675094 732019 675146 732071
rect 675382 732019 675434 732071
rect 42358 731797 42410 731849
rect 45046 731797 45098 731849
rect 674614 730465 674666 730517
rect 675478 730465 675530 730517
rect 674230 728911 674282 728963
rect 674230 728689 674282 728741
rect 47542 728615 47594 728667
rect 59542 728615 59594 728667
rect 674326 728615 674378 728667
rect 675478 728615 675530 728667
rect 674998 725729 675050 725781
rect 675382 725729 675434 725781
rect 42742 720623 42794 720675
rect 42742 720401 42794 720453
rect 663766 717885 663818 717937
rect 674422 717885 674474 717937
rect 660886 717293 660938 717345
rect 674422 717293 674474 717345
rect 654262 717145 654314 717197
rect 666934 717145 666986 717197
rect 43126 717071 43178 717123
rect 44854 717071 44906 717123
rect 661078 716849 661130 716901
rect 674422 716849 674474 716901
rect 672310 716257 672362 716309
rect 674422 716257 674474 716309
rect 41680 714238 41732 714290
rect 44950 714259 45002 714311
rect 59542 714259 59594 714311
rect 43510 714037 43562 714089
rect 41782 713963 41834 714015
rect 43414 713963 43466 714015
rect 42070 713519 42122 713571
rect 42358 713519 42410 713571
rect 43414 711669 43466 711721
rect 43030 711521 43082 711573
rect 43030 711003 43082 711055
rect 43222 711003 43274 711055
rect 42166 710855 42218 710907
rect 43414 710855 43466 710907
rect 672502 709745 672554 709797
rect 674422 709745 674474 709797
rect 672598 709153 672650 709205
rect 674422 709153 674474 709205
rect 672886 708635 672938 708687
rect 674422 708635 674474 708687
rect 42070 708561 42122 708613
rect 43126 708561 43178 708613
rect 42166 708043 42218 708095
rect 42454 708043 42506 708095
rect 42166 706563 42218 706615
rect 43126 706563 43178 706615
rect 675190 705601 675242 705653
rect 675382 705601 675434 705653
rect 43030 704269 43082 704321
rect 42166 704047 42218 704099
rect 43030 704121 43082 704173
rect 43510 704121 43562 704173
rect 42070 703529 42122 703581
rect 42454 703529 42506 703581
rect 42166 702863 42218 702915
rect 43126 702863 43178 702915
rect 649846 702715 649898 702767
rect 677014 702715 677066 702767
rect 42166 702271 42218 702323
rect 43030 702271 43082 702323
rect 42166 700051 42218 700103
rect 42454 700051 42506 700103
rect 43126 699829 43178 699881
rect 59542 699829 59594 699881
rect 672790 699829 672842 699881
rect 673174 699829 673226 699881
rect 42166 699385 42218 699437
rect 42358 699385 42410 699437
rect 654454 694057 654506 694109
rect 672502 694057 672554 694109
rect 675094 693465 675146 693517
rect 675478 693465 675530 693517
rect 673174 692947 673226 692999
rect 675478 692947 675530 692999
rect 672790 692873 672842 692925
rect 675382 692873 675434 692925
rect 675190 692651 675242 692703
rect 675382 692651 675434 692703
rect 674998 690653 675050 690705
rect 675478 690653 675530 690705
rect 673270 689765 673322 689817
rect 675382 689765 675434 689817
rect 43222 689469 43274 689521
rect 44950 689469 45002 689521
rect 673078 688581 673130 688633
rect 675478 688581 675530 688633
rect 42838 688433 42890 688485
rect 47542 688433 47594 688485
rect 675094 687323 675146 687375
rect 675478 687323 675530 687375
rect 669622 686213 669674 686265
rect 675382 686213 675434 686265
rect 47542 685473 47594 685525
rect 59542 685473 59594 685525
rect 674326 685473 674378 685525
rect 675478 685473 675530 685525
rect 674902 684067 674954 684119
rect 674998 684067 675050 684119
rect 674998 683845 675050 683897
rect 674902 683771 674954 683823
rect 675094 683623 675146 683675
rect 675478 683623 675530 683675
rect 674998 680959 675050 681011
rect 675190 680959 675242 681011
rect 42166 674003 42218 674055
rect 43030 674003 43082 674055
rect 43414 673855 43466 673907
rect 44758 673855 44810 673907
rect 669814 672671 669866 672723
rect 674422 672671 674474 672723
rect 666838 672153 666890 672205
rect 674422 672153 674474 672205
rect 41878 672079 41930 672131
rect 42646 672079 42698 672131
rect 664054 671561 664106 671613
rect 674422 671561 674474 671613
rect 44854 671043 44906 671095
rect 59542 671043 59594 671095
rect 654454 671043 654506 671095
rect 661078 671043 661130 671095
rect 43222 670895 43274 670947
rect 43414 670821 43466 670873
rect 42646 670747 42698 670799
rect 42934 670747 42986 670799
rect 41974 670673 42026 670725
rect 43126 670673 43178 670725
rect 41782 670599 41834 670651
rect 42646 670599 42698 670651
rect 42166 670303 42218 670355
rect 42358 670303 42410 670355
rect 42166 668527 42218 668579
rect 42934 668527 42986 668579
rect 42934 668379 42986 668431
rect 43222 668379 43274 668431
rect 42166 667861 42218 667913
rect 43510 667861 43562 667913
rect 42166 666677 42218 666729
rect 42934 666677 42986 666729
rect 42934 665197 42986 665249
rect 43414 665197 43466 665249
rect 672694 665197 672746 665249
rect 673846 665197 673898 665249
rect 42070 664161 42122 664213
rect 42646 664161 42698 664213
rect 42166 663347 42218 663399
rect 43030 663347 43082 663399
rect 672982 662311 673034 662363
rect 673846 662311 673898 662363
rect 42070 661053 42122 661105
rect 43126 661053 43178 661105
rect 674422 660979 674474 661031
rect 675094 660979 675146 661031
rect 42070 660387 42122 660439
rect 42934 660387 42986 660439
rect 42166 659647 42218 659699
rect 42646 659647 42698 659699
rect 42646 659499 42698 659551
rect 43702 659499 43754 659551
rect 649942 659499 649994 659551
rect 674902 659499 674954 659551
rect 42070 659055 42122 659107
rect 42646 659055 42698 659107
rect 42070 657353 42122 657405
rect 42358 657353 42410 657405
rect 42934 656687 42986 656739
rect 59542 656687 59594 656739
rect 42166 656613 42218 656665
rect 43030 656613 43082 656665
rect 42166 656169 42218 656221
rect 43126 656169 43178 656221
rect 674614 655207 674666 655259
rect 675190 655207 675242 655259
rect 673174 653727 673226 653779
rect 675190 653727 675242 653779
rect 671734 648251 671786 648303
rect 675382 648251 675434 648303
rect 654262 648029 654314 648081
rect 664054 648029 664106 648081
rect 672310 648029 672362 648081
rect 675382 648029 675434 648081
rect 43222 647733 43274 647785
rect 44854 647733 44906 647785
rect 674518 647067 674570 647119
rect 675190 647067 675242 647119
rect 675382 647067 675434 647119
rect 674230 646401 674282 646453
rect 675094 646401 675146 646453
rect 675382 646401 675434 646453
rect 674614 645217 674666 645269
rect 674902 645217 674954 645269
rect 666742 645143 666794 645195
rect 675094 645143 675146 645195
rect 42358 645069 42410 645121
rect 59542 645069 59594 645121
rect 672214 644551 672266 644603
rect 675478 644551 675530 644603
rect 672598 644033 672650 644085
rect 675478 644033 675530 644085
rect 672886 643367 672938 643419
rect 675382 643367 675434 643419
rect 673366 642257 673418 642309
rect 675478 642257 675530 642309
rect 675094 641813 675146 641865
rect 675382 641813 675434 641865
rect 41782 631749 41834 631801
rect 42646 631749 42698 631801
rect 42646 628271 42698 628323
rect 42646 627975 42698 628027
rect 42454 627901 42506 627953
rect 47638 627901 47690 627953
rect 44758 627827 44810 627879
rect 59542 627827 59594 627879
rect 41014 627753 41066 627805
rect 43414 627753 43466 627805
rect 672406 627753 672458 627805
rect 673846 627753 673898 627805
rect 41590 627679 41642 627731
rect 43126 627679 43178 627731
rect 41878 627383 41930 627435
rect 669718 627309 669770 627361
rect 674614 627309 674666 627361
rect 41878 627161 41930 627213
rect 661174 626865 661226 626917
rect 674614 626865 674666 626917
rect 42166 625311 42218 625363
rect 42646 625311 42698 625363
rect 670966 625163 671018 625215
rect 674614 625163 674666 625215
rect 42166 624645 42218 624697
rect 42454 624645 42506 624697
rect 42166 623461 42218 623513
rect 43222 623461 43274 623513
rect 42166 622203 42218 622255
rect 42454 622203 42506 622255
rect 671926 622203 671978 622255
rect 677206 622203 677258 622255
rect 654070 622129 654122 622181
rect 672694 622129 672746 622181
rect 673750 622055 673802 622107
rect 676822 622055 676874 622107
rect 42166 621611 42218 621663
rect 42646 621611 42698 621663
rect 42070 620871 42122 620923
rect 43318 620871 43370 620923
rect 42166 620353 42218 620405
rect 43126 620353 43178 620405
rect 672790 619169 672842 619221
rect 673846 619169 673898 619221
rect 42070 617837 42122 617889
rect 42646 617837 42698 617889
rect 42166 617319 42218 617371
rect 42454 617319 42506 617371
rect 42166 616653 42218 616705
rect 42358 616653 42410 616705
rect 42166 615839 42218 615891
rect 43126 615839 43178 615891
rect 42166 614137 42218 614189
rect 43510 614137 43562 614189
rect 42166 613619 42218 613671
rect 42358 613619 42410 613671
rect 42358 613471 42410 613523
rect 59542 613471 59594 613523
rect 650038 613471 650090 613523
rect 677110 613471 677162 613523
rect 654358 613397 654410 613449
rect 669526 613397 669578 613449
rect 674230 613397 674282 613449
rect 675190 613397 675242 613449
rect 42070 612953 42122 613005
rect 42454 612953 42506 613005
rect 672118 604073 672170 604125
rect 675478 604073 675530 604125
rect 672022 603259 672074 603311
rect 675382 603259 675434 603311
rect 673270 602667 673322 602719
rect 675382 602667 675434 602719
rect 672406 602149 672458 602201
rect 675190 602149 675242 602201
rect 675382 602149 675434 602201
rect 673462 602075 673514 602127
rect 674518 602075 674570 602127
rect 675478 602075 675530 602127
rect 43222 601927 43274 601979
rect 46006 601927 46058 601979
rect 663766 601927 663818 601979
rect 675094 601927 675146 601979
rect 42454 601853 42506 601905
rect 59542 601853 59594 601905
rect 673174 601705 673226 601757
rect 673750 601705 673802 601757
rect 674614 600373 674666 600425
rect 675478 600373 675530 600425
rect 673078 599559 673130 599611
rect 675382 599559 675434 599611
rect 654454 599041 654506 599093
rect 669526 599041 669578 599093
rect 671830 599041 671882 599093
rect 675382 599041 675434 599093
rect 672982 598375 673034 598427
rect 675478 598375 675530 598427
rect 672790 597117 672842 597169
rect 675478 597117 675530 597169
rect 675094 596821 675146 596873
rect 675382 596821 675434 596873
rect 675094 590457 675146 590509
rect 675478 590457 675530 590509
rect 673174 590383 673226 590435
rect 673846 590383 673898 590435
rect 671926 588755 671978 588807
rect 676918 588755 676970 588807
rect 654454 587497 654506 587549
rect 666838 587497 666890 587549
rect 673846 587497 673898 587549
rect 676822 587497 676874 587549
rect 46006 584907 46058 584959
rect 58774 584907 58826 584959
rect 43126 584611 43178 584663
rect 43318 584611 43370 584663
rect 43414 584611 43466 584663
rect 43894 584611 43946 584663
rect 41590 584537 41642 584589
rect 43510 584537 43562 584589
rect 41686 584463 41738 584515
rect 43126 584463 43178 584515
rect 42934 584389 42986 584441
rect 43414 584389 43466 584441
rect 43030 584315 43082 584367
rect 43606 584315 43658 584367
rect 41782 584241 41834 584293
rect 42934 584241 42986 584293
rect 41878 584167 41930 584219
rect 42070 584167 42122 584219
rect 43030 584167 43082 584219
rect 42454 584093 42506 584145
rect 50422 584093 50474 584145
rect 41878 583945 41930 583997
rect 42166 582095 42218 582147
rect 43318 582095 43370 582147
rect 663958 582021 664010 582073
rect 674422 582021 674474 582073
rect 655222 581947 655274 581999
rect 674614 581947 674666 581999
rect 666934 581577 666986 581629
rect 674614 581577 674666 581629
rect 42070 581429 42122 581481
rect 42454 581429 42506 581481
rect 670966 580837 671018 580889
rect 674422 580837 674474 580889
rect 42070 580245 42122 580297
rect 43414 580245 43466 580297
rect 671926 580023 671978 580075
rect 674614 580023 674666 580075
rect 42070 578395 42122 578447
rect 43030 578395 43082 578447
rect 43030 578247 43082 578299
rect 43510 578247 43562 578299
rect 42166 577655 42218 577707
rect 43606 577655 43658 577707
rect 42070 577137 42122 577189
rect 42934 577137 42986 577189
rect 654454 576027 654506 576079
rect 669718 576027 669770 576079
rect 671734 574473 671786 574525
rect 674614 574473 674666 574525
rect 42166 573955 42218 574007
rect 43126 573955 43178 574007
rect 672598 573437 672650 573489
rect 674614 573437 674666 573489
rect 42070 573215 42122 573267
rect 42454 573215 42506 573267
rect 672214 573067 672266 573119
rect 673750 573067 673802 573119
rect 672310 572845 672362 572897
rect 674614 572845 674666 572897
rect 42166 572623 42218 572675
rect 43030 572623 43082 572675
rect 672886 571809 672938 571861
rect 674614 571809 674666 571861
rect 43510 571661 43562 571713
rect 43894 571661 43946 571713
rect 42166 570995 42218 571047
rect 42934 570995 42986 571047
rect 42166 570403 42218 570455
rect 42454 570403 42506 570455
rect 42934 570255 42986 570307
rect 59542 570255 59594 570307
rect 42070 569663 42122 569715
rect 43030 569663 43082 569715
rect 650134 567369 650186 567421
rect 677014 567369 677066 567421
rect 654454 567295 654506 567347
rect 666646 567295 666698 567347
rect 672406 564261 672458 564313
rect 675094 564261 675146 564313
rect 673462 563891 673514 563943
rect 675190 563891 675242 563943
rect 674614 559377 674666 559429
rect 675382 559377 675434 559429
rect 42454 559007 42506 559059
rect 50230 559007 50282 559059
rect 42550 558859 42602 558911
rect 59542 558859 59594 558911
rect 674902 558045 674954 558097
rect 675382 558045 675434 558097
rect 675190 557823 675242 557875
rect 675382 557823 675434 557875
rect 673462 557601 673514 557653
rect 675478 557601 675530 557653
rect 675094 557083 675146 557135
rect 675478 557083 675530 557135
rect 660886 555825 660938 555877
rect 675094 555825 675146 555877
rect 674422 555233 674474 555285
rect 675478 555233 675530 555285
rect 673174 553901 673226 553953
rect 675478 553901 675530 553953
rect 673366 553161 673418 553213
rect 675382 553161 675434 553213
rect 654454 552939 654506 552991
rect 666646 552939 666698 552991
rect 674326 551903 674378 551955
rect 675478 551903 675530 551955
rect 675094 551607 675146 551659
rect 675382 551607 675434 551659
rect 674902 550053 674954 550105
rect 675094 550053 675146 550105
rect 675478 550053 675530 550105
rect 41590 549831 41642 549883
rect 41782 549831 41834 549883
rect 674902 549831 674954 549883
rect 674518 548203 674570 548255
rect 675478 548203 675530 548255
rect 50230 544503 50282 544555
rect 59542 544503 59594 544555
rect 42166 542357 42218 542409
rect 43126 542357 43178 542409
rect 42934 541469 42986 541521
rect 53686 541469 53738 541521
rect 654454 541469 654506 541521
rect 672406 541469 672458 541521
rect 41590 541247 41642 541299
rect 43702 541247 43754 541299
rect 42838 541099 42890 541151
rect 43318 541099 43370 541151
rect 41974 540951 42026 541003
rect 42070 540951 42122 541003
rect 42838 540951 42890 541003
rect 42454 540359 42506 540411
rect 42070 538879 42122 538931
rect 42454 538879 42506 538931
rect 42454 538731 42506 538783
rect 43222 538731 43274 538783
rect 672502 538509 672554 538561
rect 673750 538509 673802 538561
rect 42166 538287 42218 538339
rect 42934 538287 42986 538339
rect 42934 538139 42986 538191
rect 43318 538139 43370 538191
rect 42070 537029 42122 537081
rect 42454 537029 42506 537081
rect 671926 536733 671978 536785
rect 673750 536733 673802 536785
rect 674614 536733 674666 536785
rect 674902 536733 674954 536785
rect 661078 536585 661130 536637
rect 674614 536585 674666 536637
rect 674518 536289 674570 536341
rect 675094 536289 675146 536341
rect 42070 535771 42122 535823
rect 43030 535771 43082 535823
rect 655126 535771 655178 535823
rect 676822 535771 676874 535823
rect 42166 535031 42218 535083
rect 43126 535031 43178 535083
rect 43126 534883 43178 534935
rect 43702 534883 43754 534935
rect 42166 534439 42218 534491
rect 42934 534439 42986 534491
rect 42070 533699 42122 533751
rect 43030 533699 43082 533751
rect 42166 531331 42218 531383
rect 42358 531331 42410 531383
rect 42166 530887 42218 530939
rect 42454 530887 42506 530939
rect 42454 530739 42506 530791
rect 42934 530739 42986 530791
rect 42070 530221 42122 530273
rect 42838 530221 42890 530273
rect 42838 529925 42890 529977
rect 59542 529925 59594 529977
rect 654070 529925 654122 529977
rect 672598 529925 672650 529977
rect 672118 529851 672170 529903
rect 673750 529851 673802 529903
rect 674902 529851 674954 529903
rect 675190 529851 675242 529903
rect 672790 529555 672842 529607
rect 673750 529555 673802 529607
rect 672022 529481 672074 529533
rect 674902 529481 674954 529533
rect 42166 529407 42218 529459
rect 43126 529407 43178 529459
rect 671830 528593 671882 528645
rect 673750 528593 673802 528645
rect 42166 527779 42218 527831
rect 42454 527779 42506 527831
rect 42070 527187 42122 527239
rect 42358 527187 42410 527239
rect 42166 526447 42218 526499
rect 42934 526447 42986 526499
rect 650230 524301 650282 524353
rect 677110 524301 677162 524353
rect 42358 524153 42410 524205
rect 42838 524153 42890 524205
rect 654454 519269 654506 519321
rect 663862 519269 663914 519321
rect 50518 515495 50570 515547
rect 59542 515495 59594 515547
rect 674902 514089 674954 514141
rect 675094 514089 675146 514141
rect 654454 506911 654506 506963
rect 663862 506911 663914 506963
rect 53878 501139 53930 501191
rect 59542 501139 59594 501191
rect 674614 499659 674666 499711
rect 674998 499659 675050 499711
rect 675094 495959 675146 496011
rect 675382 495959 675434 496011
rect 654358 495367 654410 495419
rect 661174 495367 661226 495419
rect 664054 492925 664106 492977
rect 674326 492925 674378 492977
rect 655318 492481 655370 492533
rect 674614 492481 674666 492533
rect 672694 492407 672746 492459
rect 673846 492407 673898 492459
rect 50422 486709 50474 486761
rect 58582 486709 58634 486761
rect 654262 483823 654314 483875
rect 666934 483823 666986 483875
rect 650326 479457 650378 479509
rect 677014 479457 677066 479509
rect 44950 472353 45002 472405
rect 59542 472353 59594 472405
rect 654454 472205 654506 472257
rect 660982 472205 661034 472257
rect 47830 457923 47882 457975
rect 59542 457923 59594 457975
rect 654454 457923 654506 457975
rect 660982 457923 661034 457975
rect 654358 446379 654410 446431
rect 672502 446379 672554 446431
rect 53686 443567 53738 443619
rect 59542 443567 59594 443619
rect 654454 434909 654506 434961
rect 663958 434909 664010 434961
rect 42838 432245 42890 432297
rect 50518 432245 50570 432297
rect 42838 431727 42890 431779
rect 53878 431727 53930 431779
rect 42838 429581 42890 429633
rect 43606 429581 43658 429633
rect 47638 429137 47690 429189
rect 59542 429137 59594 429189
rect 654454 426177 654506 426229
rect 669622 426177 669674 426229
rect 42358 417593 42410 417645
rect 56182 417593 56234 417645
rect 40246 416261 40298 416313
rect 42742 416261 42794 416313
rect 40054 415669 40106 415721
rect 43126 415669 43178 415721
rect 40150 415373 40202 415425
rect 43030 415373 43082 415425
rect 39958 414707 40010 414759
rect 43414 414707 43466 414759
rect 50518 414707 50570 414759
rect 58390 414707 58442 414759
rect 41878 413375 41930 413427
rect 41878 413153 41930 413205
rect 653878 411821 653930 411873
rect 669622 411821 669674 411873
rect 42166 411303 42218 411355
rect 42838 411303 42890 411355
rect 42070 410489 42122 410541
rect 47446 410489 47498 410541
rect 42166 409453 42218 409505
rect 42742 409453 42794 409505
rect 43030 409231 43082 409283
rect 42838 409157 42890 409209
rect 42934 409083 42986 409135
rect 43126 409083 43178 409135
rect 43126 408935 43178 408987
rect 43414 408935 43466 408987
rect 42166 408195 42218 408247
rect 42742 408195 42794 408247
rect 42070 407455 42122 407507
rect 43126 407455 43178 407507
rect 42166 407011 42218 407063
rect 42838 407011 42890 407063
rect 666838 405457 666890 405509
rect 674710 405457 674762 405509
rect 669526 404717 669578 404769
rect 674422 404717 674474 404769
rect 669718 404421 669770 404473
rect 674710 404421 674762 404473
rect 42166 403681 42218 403733
rect 42742 403681 42794 403733
rect 673462 400499 673514 400551
rect 677302 400499 677354 400551
rect 673366 400425 673418 400477
rect 677110 400425 677162 400477
rect 45046 400351 45098 400403
rect 58390 400351 58442 400403
rect 654454 400351 654506 400403
rect 666838 400351 666890 400403
rect 673654 400351 673706 400403
rect 673846 400351 673898 400403
rect 650422 391767 650474 391819
rect 677110 391767 677162 391819
rect 42358 389325 42410 389377
rect 44950 389325 45002 389377
rect 654454 388807 654506 388859
rect 669526 388807 669578 388859
rect 42358 388733 42410 388785
rect 47830 388733 47882 388785
rect 42742 387993 42794 388045
rect 50422 387993 50474 388045
rect 674998 386143 675050 386195
rect 675382 386143 675434 386195
rect 47734 385921 47786 385973
rect 59254 385921 59306 385973
rect 675190 385477 675242 385529
rect 675478 385403 675530 385455
rect 674710 385181 674762 385233
rect 674998 385181 675050 385233
rect 674902 384811 674954 384863
rect 675382 384811 675434 384863
rect 674518 383109 674570 383161
rect 675382 383109 675434 383161
rect 674422 382295 674474 382347
rect 675478 382295 675530 382347
rect 654454 380075 654506 380127
rect 666742 380075 666794 380127
rect 674806 378151 674858 378203
rect 675382 378151 675434 378203
rect 674614 377559 674666 377611
rect 675382 377559 675434 377611
rect 674230 376819 674282 376871
rect 675478 376819 675530 376871
rect 42646 376523 42698 376575
rect 44950 376523 45002 376575
rect 673942 375709 673994 375761
rect 675478 375709 675530 375761
rect 40246 373341 40298 373393
rect 43414 373341 43466 373393
rect 39958 372379 40010 372431
rect 43030 372379 43082 372431
rect 39862 371565 39914 371617
rect 43318 371565 43370 371617
rect 50422 371565 50474 371617
rect 59542 371565 59594 371617
rect 42166 370159 42218 370211
rect 42166 369937 42218 369989
rect 42358 369937 42410 369989
rect 42550 368827 42602 368879
rect 42070 368087 42122 368139
rect 42550 368087 42602 368139
rect 42934 367569 42986 367621
rect 43318 367569 43370 367621
rect 42070 367347 42122 367399
rect 50326 367347 50378 367399
rect 42070 366163 42122 366215
rect 43030 366163 43082 366215
rect 654454 365793 654506 365845
rect 661078 365793 661130 365845
rect 42166 364979 42218 365031
rect 43126 364979 43178 365031
rect 42070 364387 42122 364439
rect 42646 364387 42698 364439
rect 42166 363795 42218 363847
rect 43414 363795 43466 363847
rect 42166 360613 42218 360665
rect 42934 360613 42986 360665
rect 672406 360021 672458 360073
rect 674422 360021 674474 360073
rect 666646 359725 666698 359777
rect 674710 359725 674762 359777
rect 672598 358985 672650 359037
rect 674422 358985 674474 359037
rect 47446 357135 47498 357187
rect 59542 357135 59594 357187
rect 42454 346109 42506 346161
rect 47638 346109 47690 346161
rect 650518 345591 650570 345643
rect 677110 345591 677162 345643
rect 42454 345517 42506 345569
rect 50518 345517 50570 345569
rect 42934 344777 42986 344829
rect 53686 344777 53738 344829
rect 53878 342779 53930 342831
rect 58390 342779 58442 342831
rect 654454 342705 654506 342757
rect 666646 342705 666698 342757
rect 674806 341595 674858 341647
rect 675190 341595 675242 341647
rect 674902 341299 674954 341351
rect 675094 341299 675146 341351
rect 674614 339745 674666 339797
rect 675094 339745 675146 339797
rect 674422 339523 674474 339575
rect 675382 339523 675434 339575
rect 674518 337229 674570 337281
rect 675094 337229 675146 337281
rect 673942 333529 673994 333581
rect 675382 333529 675434 333581
rect 42838 333307 42890 333359
rect 47638 333307 47690 333359
rect 674230 332937 674282 332989
rect 675382 332937 675434 332989
rect 654454 332271 654506 332323
rect 663766 332271 663818 332323
rect 674326 332197 674378 332249
rect 675478 332197 675530 332249
rect 674038 331531 674090 331583
rect 675382 331531 675434 331583
rect 39862 329755 39914 329807
rect 43126 329755 43178 329807
rect 40054 329459 40106 329511
rect 42838 329459 42890 329511
rect 39958 329311 40010 329363
rect 42454 329311 42506 329363
rect 40246 329163 40298 329215
rect 42358 329163 42410 329215
rect 50326 328349 50378 328401
rect 57814 328349 57866 328401
rect 41878 327017 41930 327069
rect 41878 326721 41930 326773
rect 42454 325611 42506 325663
rect 42742 325315 42794 325367
rect 42070 324871 42122 324923
rect 42934 324871 42986 324923
rect 42166 324131 42218 324183
rect 44662 324131 44714 324183
rect 42166 323095 42218 323147
rect 42742 323095 42794 323147
rect 42838 322947 42890 322999
rect 42454 322725 42506 322777
rect 42070 321763 42122 321815
rect 43030 321763 43082 321815
rect 42166 321023 42218 321075
rect 42454 321023 42506 321075
rect 42166 320579 42218 320631
rect 43126 320579 43178 320631
rect 42166 317471 42218 317523
rect 42454 317471 42506 317523
rect 661174 315029 661226 315081
rect 674422 315029 674474 315081
rect 663862 314733 663914 314785
rect 674710 314733 674762 314785
rect 666934 313993 666986 314045
rect 674422 313993 674474 314045
rect 44662 313919 44714 313971
rect 58006 313919 58058 313971
rect 42550 302893 42602 302945
rect 47734 302893 47786 302945
rect 650614 302597 650666 302649
rect 674422 302597 674474 302649
rect 42550 302301 42602 302353
rect 50422 302301 50474 302353
rect 42550 301857 42602 301909
rect 45046 301857 45098 301909
rect 674518 300525 674570 300577
rect 674710 300525 674762 300577
rect 45142 299563 45194 299615
rect 59446 299563 59498 299615
rect 674518 295937 674570 295989
rect 675382 295937 675434 295989
rect 674902 295345 674954 295397
rect 675478 295345 675530 295397
rect 673942 294531 673994 294583
rect 675382 294531 675434 294583
rect 654550 293791 654602 293843
rect 663766 293791 663818 293843
rect 674326 292903 674378 292955
rect 675382 292903 675434 292955
rect 674806 291719 674858 291771
rect 675094 291719 675146 291771
rect 674614 291053 674666 291105
rect 675094 291053 675146 291105
rect 42550 289795 42602 289847
rect 47734 289795 47786 289847
rect 674998 288537 675050 288589
rect 675478 288537 675530 288589
rect 674422 287723 674474 287775
rect 675382 287723 675434 287775
rect 674038 287205 674090 287257
rect 675478 287205 675530 287257
rect 674230 286761 674282 286813
rect 675382 286761 675434 286813
rect 39862 285429 39914 285481
rect 43126 285429 43178 285481
rect 40054 285281 40106 285333
rect 43126 285281 43178 285333
rect 40150 285133 40202 285185
rect 43030 285133 43082 285185
rect 45046 285133 45098 285185
rect 58102 285133 58154 285185
rect 654070 284763 654122 284815
rect 660886 284763 660938 284815
rect 41206 284097 41258 284149
rect 41974 283801 42026 283853
rect 42454 283579 42506 283631
rect 41974 283505 42026 283557
rect 42166 281729 42218 281781
rect 42454 281729 42506 281781
rect 42166 281063 42218 281115
rect 53494 281063 53546 281115
rect 42166 279879 42218 279931
rect 43030 279879 43082 279931
rect 43126 279879 43178 279931
rect 43126 279657 43178 279709
rect 318166 278621 318218 278673
rect 42166 278547 42218 278599
rect 42934 278547 42986 278599
rect 64726 278547 64778 278599
rect 66646 278547 66698 278599
rect 295798 278547 295850 278599
rect 309046 278547 309098 278599
rect 370486 278547 370538 278599
rect 370966 278547 371018 278599
rect 379030 278547 379082 278599
rect 379126 278547 379178 278599
rect 379702 278547 379754 278599
rect 396214 278547 396266 278599
rect 403318 278547 403370 278599
rect 266038 278473 266090 278525
rect 334390 278473 334442 278525
rect 338326 278473 338378 278525
rect 358582 278473 358634 278525
rect 373174 278473 373226 278525
rect 387766 278473 387818 278525
rect 388342 278473 388394 278525
rect 490198 278473 490250 278525
rect 223126 278399 223178 278451
rect 329110 278399 329162 278451
rect 350326 278399 350378 278451
rect 393814 278399 393866 278451
rect 293782 278325 293834 278377
rect 389014 278325 389066 278377
rect 292054 278251 292106 278303
rect 374806 278251 374858 278303
rect 375478 278251 375530 278303
rect 385078 278251 385130 278303
rect 301846 278177 301898 278229
rect 453238 278177 453290 278229
rect 198166 278103 198218 278155
rect 325270 278103 325322 278155
rect 326614 278103 326666 278155
rect 635254 278103 635306 278155
rect 297526 278029 297578 278081
rect 417622 278029 417674 278081
rect 290806 277955 290858 278007
rect 309430 277955 309482 278007
rect 311830 277955 311882 278007
rect 328150 277955 328202 278007
rect 353494 277955 353546 278007
rect 64822 277881 64874 277933
rect 182230 277881 182282 277933
rect 301558 277881 301610 277933
rect 311926 277881 311978 277933
rect 312406 277881 312458 277933
rect 339958 277881 340010 277933
rect 355510 277881 355562 277933
rect 357430 277955 357482 278007
rect 415318 277955 415370 278007
rect 287254 277807 287306 277859
rect 335542 277807 335594 277859
rect 356854 277807 356906 277859
rect 422326 277881 422378 277933
rect 289942 277733 289994 277785
rect 357046 277733 357098 277785
rect 436630 277807 436682 277859
rect 450838 277733 450890 277785
rect 291478 277659 291530 277711
rect 356950 277659 357002 277711
rect 358870 277659 358922 277711
rect 465526 277659 465578 277711
rect 296470 277585 296522 277637
rect 410806 277585 410858 277637
rect 293206 277511 293258 277563
rect 382294 277511 382346 277563
rect 307990 277437 308042 277489
rect 318070 277437 318122 277489
rect 318358 277437 318410 277489
rect 331318 277437 331370 277489
rect 352918 277437 352970 277489
rect 357430 277437 357482 277489
rect 361558 277437 361610 277489
rect 486838 277437 486890 277489
rect 247894 277363 247946 277415
rect 292246 277363 292298 277415
rect 298198 277363 298250 277415
rect 425014 277363 425066 277415
rect 318454 277289 318506 277341
rect 327382 277289 327434 277341
rect 327670 277289 327722 277341
rect 460726 277289 460778 277341
rect 42070 277215 42122 277267
rect 43126 277215 43178 277267
rect 240694 277215 240746 277267
rect 290806 277215 290858 277267
rect 299062 277215 299114 277267
rect 432214 277215 432266 277267
rect 300214 277141 300266 277193
rect 439318 277141 439370 277193
rect 233494 277067 233546 277119
rect 330166 277067 330218 277119
rect 349078 277067 349130 277119
rect 386998 277067 387050 277119
rect 388438 277067 388490 277119
rect 402454 277067 402506 277119
rect 225238 276993 225290 277045
rect 273622 276993 273674 277045
rect 290806 276993 290858 277045
rect 364438 276993 364490 277045
rect 364822 276993 364874 277045
rect 300790 276919 300842 276971
rect 376630 276919 376682 276971
rect 289270 276845 289322 276897
rect 350038 276845 350090 276897
rect 365302 276845 365354 276897
rect 370966 276845 371018 276897
rect 377014 276993 377066 277045
rect 378550 276993 378602 277045
rect 378646 276993 378698 277045
rect 504694 276993 504746 277045
rect 376918 276919 376970 276971
rect 446518 276919 446570 276971
rect 515446 276845 515498 276897
rect 254902 276771 254954 276823
rect 332758 276771 332810 276823
rect 348886 276771 348938 276823
rect 383350 276771 383402 276823
rect 383734 276771 383786 276823
rect 523798 276771 523850 276823
rect 639382 276771 639434 276823
rect 649558 276771 649610 276823
rect 215734 276697 215786 276749
rect 311830 276697 311882 276749
rect 311926 276697 311978 276749
rect 338710 276697 338762 276749
rect 370966 276697 371018 276749
rect 518998 276697 519050 276749
rect 208534 276623 208586 276675
rect 309622 276623 309674 276675
rect 318166 276623 318218 276675
rect 338326 276623 338378 276675
rect 363766 276623 363818 276675
rect 368566 276623 368618 276675
rect 368758 276623 368810 276675
rect 378646 276623 378698 276675
rect 378742 276623 378794 276675
rect 611830 276623 611882 276675
rect 292246 276549 292298 276601
rect 307990 276549 308042 276601
rect 318070 276549 318122 276601
rect 332182 276549 332234 276601
rect 358582 276549 358634 276601
rect 379126 276549 379178 276601
rect 379798 276549 379850 276601
rect 636694 276549 636746 276601
rect 288406 276475 288458 276527
rect 342934 276475 342986 276527
rect 351094 276475 351146 276527
rect 401206 276475 401258 276527
rect 243766 276401 243818 276453
rect 434518 276401 434570 276453
rect 231958 276327 232010 276379
rect 338230 276327 338282 276379
rect 346774 276327 346826 276379
rect 365590 276327 365642 276379
rect 370966 276327 371018 276379
rect 375478 276327 375530 276379
rect 375574 276327 375626 276379
rect 380470 276327 380522 276379
rect 380566 276327 380618 276379
rect 232342 276253 232394 276305
rect 341782 276253 341834 276305
rect 348406 276253 348458 276305
rect 379510 276253 379562 276305
rect 379990 276253 380042 276305
rect 384886 276253 384938 276305
rect 385078 276327 385130 276379
rect 565462 276327 565514 276379
rect 572470 276253 572522 276305
rect 244726 276179 244778 276231
rect 441718 276179 441770 276231
rect 245398 276105 245450 276157
rect 448822 276105 448874 276157
rect 246358 276031 246410 276083
rect 455926 276031 455978 276083
rect 233494 275957 233546 276009
rect 348982 275957 349034 276009
rect 370390 275957 370442 276009
rect 384790 275957 384842 276009
rect 384886 275957 384938 276009
rect 579670 275957 579722 276009
rect 247414 275883 247466 275935
rect 463126 275883 463178 275935
rect 227446 275809 227498 275861
rect 298966 275809 299018 275861
rect 311542 275809 311594 275861
rect 532150 275809 532202 275861
rect 248086 275735 248138 275787
rect 470230 275735 470282 275787
rect 234070 275661 234122 275713
rect 356086 275661 356138 275713
rect 364246 275661 364298 275713
rect 380278 275661 380330 275713
rect 380470 275661 380522 275713
rect 601078 275661 601130 275713
rect 249142 275587 249194 275639
rect 477430 275587 477482 275639
rect 249814 275513 249866 275565
rect 484438 275513 484490 275565
rect 200182 275439 200234 275491
rect 270742 275439 270794 275491
rect 323254 275439 323306 275491
rect 564214 275439 564266 275491
rect 235030 275365 235082 275417
rect 363190 275365 363242 275417
rect 371830 275365 371882 275417
rect 235990 275291 236042 275343
rect 370294 275291 370346 275343
rect 372886 275291 372938 275343
rect 377590 275291 377642 275343
rect 377878 275365 377930 275417
rect 622486 275365 622538 275417
rect 379414 275291 379466 275343
rect 379510 275291 379562 275343
rect 633142 275291 633194 275343
rect 196726 275217 196778 275269
rect 270550 275217 270602 275269
rect 284950 275217 285002 275269
rect 314422 275217 314474 275269
rect 316054 275217 316106 275269
rect 571318 275217 571370 275269
rect 228022 275143 228074 275195
rect 306070 275143 306122 275195
rect 317302 275143 317354 275195
rect 578518 275143 578570 275195
rect 236758 275069 236810 275121
rect 377494 275069 377546 275121
rect 377590 275069 377642 275121
rect 379990 275069 380042 275121
rect 380086 275069 380138 275121
rect 380566 275069 380618 275121
rect 381430 275069 381482 275121
rect 647542 275069 647594 275121
rect 229078 274995 229130 275047
rect 313270 274995 313322 275047
rect 318070 274995 318122 275047
rect 585622 274995 585674 275047
rect 258550 274921 258602 274973
rect 333142 274921 333194 274973
rect 368086 274921 368138 274973
rect 378646 274921 378698 274973
rect 378742 274921 378794 274973
rect 384694 274921 384746 274973
rect 384790 274921 384842 274973
rect 558262 274921 558314 274973
rect 242998 274847 243050 274899
rect 427414 274847 427466 274899
rect 223030 274773 223082 274825
rect 263350 274773 263402 274825
rect 269206 274773 269258 274825
rect 334486 274773 334538 274825
rect 372310 274773 372362 274825
rect 384598 274773 384650 274825
rect 384694 274773 384746 274825
rect 551062 274773 551114 274825
rect 242230 274699 242282 274751
rect 420214 274699 420266 274751
rect 226294 274625 226346 274677
rect 291862 274625 291914 274677
rect 297814 274625 297866 274677
rect 337942 274625 337994 274677
rect 369526 274625 369578 274677
rect 378550 274625 378602 274677
rect 378646 274625 378698 274677
rect 540406 274625 540458 274677
rect 240502 274551 240554 274603
rect 406006 274551 406058 274603
rect 239350 274477 239402 274529
rect 398902 274477 398954 274529
rect 238486 274403 238538 274455
rect 391702 274403 391754 274455
rect 237814 274329 237866 274381
rect 372310 274329 372362 274381
rect 42166 274255 42218 274307
rect 43030 274255 43082 274307
rect 207382 274255 207434 274307
rect 271318 274255 271370 274307
rect 271414 274255 271466 274307
rect 214582 274181 214634 274233
rect 272470 274181 272522 274233
rect 276406 274255 276458 274307
rect 335638 274255 335690 274307
rect 358774 274255 358826 274307
rect 378742 274329 378794 274381
rect 378838 274329 378890 274381
rect 385558 274329 385610 274381
rect 385846 274329 385898 274381
rect 395350 274329 395402 274381
rect 225430 274107 225482 274159
rect 284662 274107 284714 274159
rect 225238 274033 225290 274085
rect 281110 274033 281162 274085
rect 239446 273959 239498 274011
rect 275254 273959 275306 274011
rect 287062 274181 287114 274233
rect 337558 274181 337610 274233
rect 352246 274181 352298 274233
rect 372406 274181 372458 274233
rect 286774 274107 286826 274159
rect 328726 274107 328778 274159
rect 364342 274107 364394 274159
rect 511894 274255 511946 274307
rect 374134 274181 374186 274233
rect 378454 274181 378506 274233
rect 378550 274181 378602 274233
rect 380182 274181 380234 274233
rect 380278 274181 380330 274233
rect 508342 274181 508394 274233
rect 374326 274107 374378 274159
rect 296662 274033 296714 274085
rect 297142 274033 297194 274085
rect 304918 274033 304970 274085
rect 338902 274033 338954 274085
rect 360502 274033 360554 274085
rect 378646 274033 378698 274085
rect 378838 274107 378890 274159
rect 479734 274107 479786 274159
rect 385750 274033 385802 274085
rect 388918 274033 388970 274085
rect 476182 274033 476234 274085
rect 378550 273959 378602 274011
rect 232438 273885 232490 273937
rect 274678 273885 274730 273937
rect 308854 273885 308906 273937
rect 230614 273811 230666 273863
rect 319702 273811 319754 273863
rect 229750 273737 229802 273789
rect 320086 273737 320138 273789
rect 322774 273885 322826 273937
rect 341302 273885 341354 273937
rect 360022 273885 360074 273937
rect 383062 273959 383114 274011
rect 378742 273885 378794 273937
rect 461974 273885 462026 273937
rect 325270 273811 325322 273863
rect 325942 273811 325994 273863
rect 356182 273811 356234 273863
rect 444118 273811 444170 273863
rect 377494 273737 377546 273789
rect 377590 273737 377642 273789
rect 392950 273737 393002 273789
rect 231766 273663 231818 273715
rect 325462 273663 325514 273715
rect 325654 273663 325706 273715
rect 327670 273663 327722 273715
rect 354454 273663 354506 273715
rect 429814 273663 429866 273715
rect 66646 273589 66698 273641
rect 236278 273589 236330 273641
rect 245494 273589 245546 273641
rect 262678 273589 262730 273641
rect 79222 273515 79274 273567
rect 106294 273515 106346 273567
rect 198742 273515 198794 273567
rect 91990 273441 92042 273493
rect 190582 273441 190634 273493
rect 190678 273441 190730 273493
rect 212374 273515 212426 273567
rect 227542 273515 227594 273567
rect 247606 273515 247658 273567
rect 262390 273515 262442 273567
rect 270358 273515 270410 273567
rect 270454 273515 270506 273567
rect 271414 273515 271466 273567
rect 271606 273515 271658 273567
rect 279478 273515 279530 273567
rect 284470 273515 284522 273567
rect 224086 273441 224138 273493
rect 274006 273441 274058 273493
rect 275158 273441 275210 273493
rect 279670 273441 279722 273493
rect 281206 273441 281258 273493
rect 285814 273441 285866 273493
rect 290902 273515 290954 273567
rect 293014 273515 293066 273567
rect 294742 273515 294794 273567
rect 309046 273515 309098 273567
rect 319798 273515 319850 273567
rect 321526 273515 321578 273567
rect 325462 273515 325514 273567
rect 334582 273515 334634 273567
rect 340630 273515 340682 273567
rect 343510 273515 343562 273567
rect 344662 273515 344714 273567
rect 347734 273515 347786 273567
rect 356950 273515 357002 273567
rect 367894 273515 367946 273567
rect 372406 273589 372458 273641
rect 411958 273589 412010 273641
rect 630742 273589 630794 273641
rect 639382 273589 639434 273641
rect 380278 273515 380330 273567
rect 380374 273515 380426 273567
rect 396214 273515 396266 273567
rect 396310 273515 396362 273567
rect 612982 273515 613034 273567
rect 642262 273515 642314 273567
rect 649462 273589 649514 273641
rect 310870 273441 310922 273493
rect 319702 273441 319754 273493
rect 327478 273441 327530 273493
rect 327574 273441 327626 273493
rect 557014 273441 557066 273493
rect 153814 273367 153866 273419
rect 160918 273367 160970 273419
rect 161014 273367 161066 273419
rect 404950 273367 405002 273419
rect 157462 273293 157514 273345
rect 404086 273293 404138 273345
rect 161302 273219 161354 273271
rect 147958 273145 148010 273197
rect 149686 273145 149738 273197
rect 151414 273145 151466 273197
rect 152566 273145 152618 273197
rect 152662 273145 152714 273197
rect 155350 273145 155402 273197
rect 156214 273145 156266 273197
rect 158326 273145 158378 273197
rect 162166 273145 162218 273197
rect 164086 273145 164138 273197
rect 164278 273219 164330 273271
rect 371542 273219 371594 273271
rect 374326 273219 374378 273271
rect 401302 273219 401354 273271
rect 403222 273145 403274 273197
rect 139606 273071 139658 273123
rect 142006 272997 142058 273049
rect 143926 272997 143978 273049
rect 146710 273071 146762 273123
rect 373846 273071 373898 273123
rect 374614 273071 374666 273123
rect 400630 273071 400682 273123
rect 399670 272997 399722 273049
rect 143158 272923 143210 272975
rect 374422 272923 374474 272975
rect 65878 272849 65930 272901
rect 190678 272849 190730 272901
rect 190774 272849 190826 272901
rect 192886 272849 192938 272901
rect 197110 272849 197162 272901
rect 213238 272849 213290 272901
rect 213334 272849 213386 272901
rect 216694 272849 216746 272901
rect 217558 272849 217610 272901
rect 220438 272849 220490 272901
rect 221014 272849 221066 272901
rect 249046 272849 249098 272901
rect 258358 272849 258410 272901
rect 374326 272849 374378 272901
rect 135958 272775 136010 272827
rect 396982 272923 397034 272975
rect 374614 272849 374666 272901
rect 378454 272849 378506 272901
rect 374806 272775 374858 272827
rect 376246 272775 376298 272827
rect 376342 272775 376394 272827
rect 377398 272775 377450 272827
rect 377494 272775 377546 272827
rect 378166 272775 378218 272827
rect 125302 272701 125354 272753
rect 128950 272627 129002 272679
rect 132502 272701 132554 272753
rect 146902 272701 146954 272753
rect 166966 272701 167018 272753
rect 227542 272701 227594 272753
rect 247606 272701 247658 272753
rect 378454 272701 378506 272753
rect 380374 272849 380426 272901
rect 380566 272849 380618 272901
rect 643894 272849 643946 272901
rect 127702 272553 127754 272605
rect 129526 272553 129578 272605
rect 322582 272553 322634 272605
rect 322966 272553 323018 272605
rect 397078 272775 397130 272827
rect 378838 272701 378890 272753
rect 398326 272701 398378 272753
rect 378742 272627 378794 272679
rect 392470 272627 392522 272679
rect 392566 272627 392618 272679
rect 407254 272627 407306 272679
rect 121750 272479 121802 272531
rect 378742 272479 378794 272531
rect 391702 272553 391754 272605
rect 379222 272479 379274 272531
rect 396790 272553 396842 272605
rect 397366 272553 397418 272605
rect 595126 272553 595178 272605
rect 394582 272479 394634 272531
rect 408118 272479 408170 272531
rect 64918 272405 64970 272457
rect 71926 272405 71978 272457
rect 84886 272405 84938 272457
rect 86326 272405 86378 272457
rect 105046 272405 105098 272457
rect 106486 272405 106538 272457
rect 118102 272405 118154 272457
rect 322582 272405 322634 272457
rect 322774 272405 322826 272457
rect 378454 272405 378506 272457
rect 378838 272405 378890 272457
rect 379126 272405 379178 272457
rect 394198 272405 394250 272457
rect 394486 272405 394538 272457
rect 591574 272405 591626 272457
rect 111094 272331 111146 272383
rect 378070 272331 378122 272383
rect 378934 272331 378986 272383
rect 389494 272331 389546 272383
rect 389590 272331 389642 272383
rect 408214 272331 408266 272383
rect 408310 272331 408362 272383
rect 587926 272331 587978 272383
rect 67030 272257 67082 272309
rect 197110 272257 197162 272309
rect 209782 272257 209834 272309
rect 216118 272257 216170 272309
rect 218230 272257 218282 272309
rect 223990 272257 224042 272309
rect 224566 272257 224618 272309
rect 277558 272257 277610 272309
rect 278806 272257 278858 272309
rect 280054 272257 280106 272309
rect 280726 272257 280778 272309
rect 282358 272257 282410 272309
rect 285526 272257 285578 272309
rect 319798 272257 319850 272309
rect 320374 272257 320426 272309
rect 607030 272257 607082 272309
rect 103894 272183 103946 272235
rect 107446 272109 107498 272161
rect 378358 272109 378410 272161
rect 379030 272183 379082 272235
rect 385270 272183 385322 272235
rect 385558 272183 385610 272235
rect 386806 272183 386858 272235
rect 383062 272109 383114 272161
rect 383254 272109 383306 272161
rect 396406 272109 396458 272161
rect 150262 272035 150314 272087
rect 164278 272035 164330 272087
rect 164566 272035 164618 272087
rect 382966 272035 383018 272087
rect 383350 272035 383402 272087
rect 392566 272035 392618 272087
rect 99190 271961 99242 272013
rect 197206 271961 197258 272013
rect 197302 271961 197354 272013
rect 207862 271961 207914 272013
rect 223702 271961 223754 272013
rect 262390 271961 262442 272013
rect 268054 271961 268106 272013
rect 278998 271961 279050 272013
rect 283798 271961 283850 272013
rect 307318 271961 307370 272013
rect 308470 271961 308522 272013
rect 331414 271961 331466 272013
rect 336982 271961 337034 272013
rect 343030 271961 343082 272013
rect 347926 271961 347978 272013
rect 374518 271961 374570 272013
rect 374710 271961 374762 272013
rect 378550 271961 378602 272013
rect 378646 271961 378698 272013
rect 389590 271961 389642 272013
rect 391606 271961 391658 272013
rect 566518 272183 566570 272235
rect 165814 271887 165866 271939
rect 166966 271887 167018 271939
rect 170518 271887 170570 271939
rect 172726 271887 172778 271939
rect 177622 271887 177674 271939
rect 178390 271887 178442 271939
rect 180022 271887 180074 271939
rect 181366 271887 181418 271939
rect 187030 271887 187082 271939
rect 207286 271887 207338 271939
rect 207382 271887 207434 271939
rect 296854 271887 296906 271939
rect 296950 271887 297002 271939
rect 322582 271887 322634 271939
rect 323062 271887 323114 271939
rect 383254 271887 383306 271939
rect 383446 271887 383498 271939
rect 95638 271813 95690 271865
rect 195862 271813 195914 271865
rect 208054 271813 208106 271865
rect 210262 271813 210314 271865
rect 210358 271813 210410 271865
rect 215446 271813 215498 271865
rect 220822 271813 220874 271865
rect 236182 271813 236234 271865
rect 250198 271813 250250 271865
rect 276790 271813 276842 271865
rect 283414 271813 283466 271865
rect 303670 271813 303722 271865
rect 313654 271813 313706 271865
rect 383350 271813 383402 271865
rect 385270 271887 385322 271939
rect 387478 271887 387530 271939
rect 394390 271887 394442 271939
rect 573718 272109 573770 272161
rect 396790 271961 396842 272013
rect 618838 271961 618890 272013
rect 396694 271887 396746 271939
rect 405718 271887 405770 271939
rect 549910 271813 549962 271865
rect 101494 271739 101546 271791
rect 103606 271739 103658 271791
rect 146902 271739 146954 271791
rect 166774 271739 166826 271791
rect 176470 271739 176522 271791
rect 178486 271739 178538 271791
rect 75382 271665 75434 271717
rect 77686 271665 77738 271717
rect 120982 271665 121034 271717
rect 141046 271665 141098 271717
rect 141334 271665 141386 271717
rect 161110 271665 161162 271717
rect 166582 271665 166634 271717
rect 166870 271665 166922 271717
rect 171670 271665 171722 271717
rect 186838 271739 186890 271791
rect 187030 271739 187082 271791
rect 259318 271739 259370 271791
rect 273526 271739 273578 271791
rect 296662 271739 296714 271791
rect 316726 271739 316778 271791
rect 334102 271739 334154 271791
rect 357046 271739 357098 271791
rect 377494 271739 377546 271791
rect 377782 271739 377834 271791
rect 378742 271739 378794 271791
rect 379030 271739 379082 271791
rect 383734 271739 383786 271791
rect 394102 271739 394154 271791
rect 406582 271739 406634 271791
rect 178870 271665 178922 271717
rect 382966 271665 383018 271717
rect 383254 271665 383306 271717
rect 409270 271665 409322 271717
rect 89590 271591 89642 271643
rect 92086 271591 92138 271643
rect 100822 271591 100874 271643
rect 120790 271591 120842 271643
rect 182422 271591 182474 271643
rect 296854 271591 296906 271643
rect 297046 271591 297098 271643
rect 383062 271591 383114 271643
rect 392758 271591 392810 271643
rect 409942 271591 409994 271643
rect 141142 271517 141194 271569
rect 141622 271517 141674 271569
rect 185974 271517 186026 271569
rect 156886 271443 156938 271495
rect 168118 271443 168170 271495
rect 175318 271443 175370 271495
rect 186838 271443 186890 271495
rect 410998 271517 411050 271569
rect 102646 271369 102698 271421
rect 197302 271443 197354 271495
rect 205846 271443 205898 271495
rect 411958 271443 412010 271495
rect 421846 271443 421898 271495
rect 431926 271443 431978 271495
rect 113494 271295 113546 271347
rect 211894 271369 211946 271421
rect 220342 271369 220394 271421
rect 241846 271369 241898 271421
rect 246646 271369 246698 271421
rect 257686 271369 257738 271421
rect 195958 271295 196010 271347
rect 206614 271295 206666 271347
rect 219766 271295 219818 271347
rect 238294 271295 238346 271347
rect 241558 271295 241610 271347
rect 242038 271295 242090 271347
rect 253750 271295 253802 271347
rect 277270 271369 277322 271421
rect 314326 271369 314378 271421
rect 327574 271369 327626 271421
rect 333430 271369 333482 271421
rect 342646 271369 342698 271421
rect 347446 271369 347498 271421
rect 372694 271369 372746 271421
rect 264502 271295 264554 271347
rect 278518 271295 278570 271347
rect 282934 271295 282986 271347
rect 300118 271295 300170 271347
rect 315382 271295 315434 271347
rect 322678 271295 322730 271347
rect 322774 271295 322826 271347
rect 325654 271295 325706 271347
rect 116950 271221 117002 271273
rect 156886 271221 156938 271273
rect 168118 271221 168170 271273
rect 211798 271221 211850 271273
rect 262198 271221 262250 271273
rect 282166 271221 282218 271273
rect 306262 271221 306314 271273
rect 315190 271221 315242 271273
rect 315670 271221 315722 271273
rect 322006 271221 322058 271273
rect 322102 271221 322154 271273
rect 327478 271295 327530 271347
rect 329974 271295 330026 271347
rect 341974 271295 342026 271347
rect 357334 271295 357386 271347
rect 326326 271221 326378 271273
rect 341494 271221 341546 271273
rect 345718 271221 345770 271273
rect 358102 271221 358154 271273
rect 120502 271147 120554 271199
rect 197110 271147 197162 271199
rect 202582 271147 202634 271199
rect 109846 271073 109898 271125
rect 184726 270999 184778 271051
rect 187030 270999 187082 271051
rect 188374 271073 188426 271125
rect 190006 271073 190058 271125
rect 190582 271073 190634 271125
rect 204502 271073 204554 271125
rect 219286 271147 219338 271199
rect 234646 271147 234698 271199
rect 269398 271147 269450 271199
rect 270454 271147 270506 271199
rect 282742 271147 282794 271199
rect 210358 271073 210410 271125
rect 210454 271073 210506 271125
rect 215542 271073 215594 271125
rect 218902 271073 218954 271125
rect 231190 271073 231242 271125
rect 260950 271073 261002 271125
rect 278134 271073 278186 271125
rect 282166 271073 282218 271125
rect 290902 271073 290954 271125
rect 195862 270999 195914 271051
rect 196246 270999 196298 271051
rect 269878 270999 269930 271051
rect 281686 270999 281738 271051
rect 289462 270999 289514 271051
rect 292534 271147 292586 271199
rect 315286 271147 315338 271199
rect 315478 271147 315530 271199
rect 327094 271147 327146 271199
rect 297142 271073 297194 271125
rect 302806 271073 302858 271125
rect 294262 270999 294314 271051
rect 319030 270999 319082 271051
rect 319318 271073 319370 271125
rect 322294 270999 322346 271051
rect 322774 271073 322826 271125
rect 327958 271147 328010 271199
rect 346390 271147 346442 271199
rect 362038 271147 362090 271199
rect 366454 271295 366506 271347
rect 380182 271369 380234 271421
rect 380374 271369 380426 271421
rect 367126 271221 367178 271273
rect 383158 271295 383210 271347
rect 383446 271369 383498 271421
rect 384118 271369 384170 271421
rect 384214 271369 384266 271421
rect 593974 271369 594026 271421
rect 590326 271295 590378 271347
rect 372982 271221 373034 271273
rect 421846 271221 421898 271273
rect 431926 271221 431978 271273
rect 480982 271221 481034 271273
rect 501046 271221 501098 271273
rect 543958 271221 544010 271273
rect 377110 271147 377162 271199
rect 377206 271147 377258 271199
rect 431638 271147 431690 271199
rect 431830 271147 431882 271199
rect 545206 271147 545258 271199
rect 340918 271073 340970 271125
rect 345238 271073 345290 271125
rect 354838 271073 354890 271125
rect 357718 271073 357770 271125
rect 371446 271073 371498 271125
rect 371542 271073 371594 271125
rect 327478 270999 327530 271051
rect 377014 270999 377066 271051
rect 377110 270999 377162 271051
rect 378646 270999 378698 271051
rect 378742 270999 378794 271051
rect 384214 270999 384266 271051
rect 385654 270999 385706 271051
rect 398806 270999 398858 271051
rect 398998 271073 399050 271125
rect 449302 271073 449354 271125
rect 449590 271073 449642 271125
rect 481078 271073 481130 271125
rect 481174 271073 481226 271125
rect 534454 271073 534506 271125
rect 402358 270999 402410 271051
rect 175606 270851 175658 270903
rect 130102 270777 130154 270829
rect 132406 270777 132458 270829
rect 144406 270777 144458 270829
rect 146806 270777 146858 270829
rect 168406 270777 168458 270829
rect 175510 270777 175562 270829
rect 189526 270851 189578 270903
rect 241846 270925 241898 270977
rect 241942 270925 241994 270977
rect 193078 270777 193130 270829
rect 195862 270777 195914 270829
rect 218710 270851 218762 270903
rect 227638 270851 227690 270903
rect 257686 270925 257738 270977
rect 276214 270925 276266 270977
rect 315190 270851 315242 270903
rect 316918 270851 316970 270903
rect 394102 270925 394154 270977
rect 394294 270925 394346 270977
rect 402838 270925 402890 270977
rect 402934 270925 402986 270977
rect 428182 270999 428234 271051
rect 446326 270999 446378 271051
rect 452182 270999 452234 271051
rect 469462 270999 469514 271051
rect 489526 270999 489578 271051
rect 489622 270925 489674 270977
rect 518422 270999 518474 271051
rect 518518 270999 518570 271051
rect 548566 270999 548618 271051
rect 558646 270999 558698 271051
rect 564502 270999 564554 271051
rect 322006 270851 322058 270903
rect 340438 270851 340490 270903
rect 344758 270851 344810 270903
rect 351286 270851 351338 270903
rect 205846 270777 205898 270829
rect 68182 270703 68234 270755
rect 69046 270703 69098 270755
rect 98038 270703 98090 270755
rect 100726 270703 100778 270755
rect 115798 270703 115850 270755
rect 118006 270703 118058 270755
rect 119350 270703 119402 270755
rect 120886 270703 120938 270755
rect 122902 270703 122954 270755
rect 123766 270703 123818 270755
rect 124150 270703 124202 270755
rect 126550 270703 126602 270755
rect 131254 270703 131306 270755
rect 132310 270703 132362 270755
rect 133558 270703 133610 270755
rect 135286 270703 135338 270755
rect 137206 270703 137258 270755
rect 138166 270703 138218 270755
rect 138358 270703 138410 270755
rect 140950 270703 141002 270755
rect 145558 270703 145610 270755
rect 146710 270703 146762 270755
rect 191926 270703 191978 270755
rect 195478 270703 195530 270755
rect 206230 270703 206282 270755
rect 210454 270703 210506 270755
rect 210646 270777 210698 270829
rect 212182 270777 212234 270829
rect 257302 270777 257354 270829
rect 277462 270777 277514 270829
rect 314806 270777 314858 270829
rect 319702 270777 319754 270829
rect 322966 270777 323018 270829
rect 324886 270777 324938 270829
rect 324982 270777 325034 270829
rect 328246 270777 328298 270829
rect 328342 270777 328394 270829
rect 331222 270777 331274 270829
rect 339862 270777 339914 270829
rect 345334 270777 345386 270829
rect 347830 270777 347882 270829
rect 369142 270851 369194 270903
rect 369238 270851 369290 270903
rect 380278 270851 380330 270903
rect 380950 270851 381002 270903
rect 381430 270851 381482 270903
rect 383062 270851 383114 270903
rect 392758 270851 392810 270903
rect 392854 270851 392906 270903
rect 452182 270851 452234 270903
rect 452470 270851 452522 270903
rect 541558 270851 541610 270903
rect 548566 270851 548618 270903
rect 558646 270851 558698 270903
rect 362038 270777 362090 270829
rect 369430 270777 369482 270829
rect 369910 270777 369962 270829
rect 374422 270777 374474 270829
rect 374518 270777 374570 270829
rect 380374 270777 380426 270829
rect 383158 270777 383210 270829
rect 386326 270777 386378 270829
rect 387478 270777 387530 270829
rect 510646 270777 510698 270829
rect 214486 270703 214538 270755
rect 251254 270703 251306 270755
rect 252214 270703 252266 270755
rect 268726 270703 268778 270755
rect 316726 270703 316778 270755
rect 317110 270703 317162 270755
rect 392086 270703 392138 270755
rect 394486 270703 394538 270755
rect 452182 270703 452234 270755
rect 452662 270703 452714 270755
rect 570166 270703 570218 270755
rect 213814 270629 213866 270681
rect 243286 270629 243338 270681
rect 431062 270629 431114 270681
rect 672502 270629 672554 270681
rect 673846 270629 673898 270681
rect 231286 270555 231338 270607
rect 328438 270555 328490 270607
rect 368470 270555 368522 270607
rect 368758 270555 368810 270607
rect 372502 270555 372554 270607
rect 387286 270555 387338 270607
rect 387382 270555 387434 270607
rect 561814 270555 561866 270607
rect 221974 270481 222026 270533
rect 256150 270481 256202 270533
rect 292150 270481 292202 270533
rect 304918 270481 304970 270533
rect 316726 270481 316778 270533
rect 370006 270481 370058 270533
rect 371446 270481 371498 270533
rect 454774 270481 454826 270533
rect 548566 270481 548618 270533
rect 575830 270481 575882 270533
rect 203830 270407 203882 270459
rect 270934 270407 270986 270459
rect 307798 270407 307850 270459
rect 503542 270407 503594 270459
rect 245302 270333 245354 270385
rect 445270 270333 445322 270385
rect 232822 270259 232874 270311
rect 328342 270259 328394 270311
rect 328438 270259 328490 270311
rect 331126 270259 331178 270311
rect 331222 270259 331274 270311
rect 339862 270259 339914 270311
rect 357622 270259 357674 270311
rect 366742 270259 366794 270311
rect 367030 270259 367082 270311
rect 371638 270259 371690 270311
rect 373366 270259 373418 270311
rect 387190 270259 387242 270311
rect 387382 270259 387434 270311
rect 568918 270259 568970 270311
rect 233974 270185 234026 270237
rect 352438 270185 352490 270237
rect 358486 270185 358538 270237
rect 373462 270185 373514 270237
rect 373558 270185 373610 270237
rect 387094 270185 387146 270237
rect 387286 270185 387338 270237
rect 576118 270185 576170 270237
rect 245878 270111 245930 270163
rect 452374 270111 452426 270163
rect 234550 270037 234602 270089
rect 359638 270037 359690 270089
rect 363094 270037 363146 270089
rect 386998 270037 387050 270089
rect 387190 270037 387242 270089
rect 583222 270037 583274 270089
rect 158614 269963 158666 270015
rect 161206 269963 161258 270015
rect 194326 269963 194378 270015
rect 318454 269963 318506 270015
rect 318550 269963 318602 270015
rect 323350 269963 323402 270015
rect 323446 269963 323498 270015
rect 366646 269963 366698 270015
rect 366742 269963 366794 270015
rect 373750 269963 373802 270015
rect 374038 269963 374090 270015
rect 374518 269963 374570 270015
rect 374902 269963 374954 270015
rect 379126 269963 379178 270015
rect 379222 269963 379274 270015
rect 386902 269963 386954 270015
rect 387094 269963 387146 270015
rect 586774 269963 586826 270015
rect 247030 269889 247082 269941
rect 459574 269889 459626 269941
rect 172918 269815 172970 269867
rect 175606 269815 175658 269867
rect 226966 269815 227018 269867
rect 295414 269815 295466 269867
rect 310390 269815 310442 269867
rect 524950 269815 525002 269867
rect 247606 269741 247658 269793
rect 466582 269741 466634 269793
rect 660982 269741 661034 269793
rect 674710 269741 674762 269793
rect 235702 269667 235754 269719
rect 357622 269667 357674 269719
rect 358582 269667 358634 269719
rect 375670 269667 375722 269719
rect 375766 269667 375818 269719
rect 379030 269667 379082 269719
rect 379126 269667 379178 269719
rect 597526 269667 597578 269719
rect 174070 269593 174122 269645
rect 175510 269593 175562 269645
rect 248566 269593 248618 269645
rect 473782 269593 473834 269645
rect 236278 269519 236330 269571
rect 358486 269519 358538 269571
rect 368470 269519 368522 269571
rect 372982 269519 373034 269571
rect 374422 269519 374474 269571
rect 378934 269519 378986 269571
rect 379030 269519 379082 269571
rect 604630 269519 604682 269571
rect 227542 269445 227594 269497
rect 302518 269445 302570 269497
rect 312598 269445 312650 269497
rect 542806 269445 542858 269497
rect 249622 269371 249674 269423
rect 481366 269371 481418 269423
rect 228502 269297 228554 269349
rect 309718 269297 309770 269349
rect 313846 269297 313898 269349
rect 553462 269297 553514 269349
rect 221494 269223 221546 269275
rect 251254 269223 251306 269275
rect 251350 269223 251402 269275
rect 495190 269223 495242 269275
rect 242614 269149 242666 269201
rect 423862 269149 423914 269201
rect 241558 269075 241610 269127
rect 416662 269075 416714 269127
rect 240886 269001 240938 269053
rect 409558 269001 409610 269053
rect 416278 269001 416330 269053
rect 486646 269149 486698 269201
rect 663958 269149 664010 269201
rect 674710 269149 674762 269201
rect 486646 269001 486698 269053
rect 230230 268927 230282 268979
rect 229558 268853 229610 268905
rect 316342 268853 316394 268905
rect 317974 268927 318026 268979
rect 337270 268927 337322 268979
rect 349078 268927 349130 268979
rect 369814 268927 369866 268979
rect 371350 268927 371402 268979
rect 378454 268927 378506 268979
rect 318262 268853 318314 268905
rect 318358 268853 318410 268905
rect 337846 268853 337898 268905
rect 351766 268853 351818 268905
rect 385558 268927 385610 268979
rect 386998 268927 387050 268979
rect 388534 268927 388586 268979
rect 388726 268927 388778 268979
rect 388822 268927 388874 268979
rect 489622 268927 489674 268979
rect 489718 268927 489770 268979
rect 518326 269001 518378 269053
rect 518422 268927 518474 268979
rect 536854 269001 536906 269053
rect 378646 268853 378698 268905
rect 529750 268853 529802 268905
rect 240022 268779 240074 268831
rect 378550 268779 378602 268831
rect 225814 268705 225866 268757
rect 288214 268705 288266 268757
rect 290614 268705 290666 268757
rect 317974 268705 318026 268757
rect 318262 268705 318314 268757
rect 334966 268705 335018 268757
rect 335062 268705 335114 268757
rect 348022 268705 348074 268757
rect 367510 268705 367562 268757
rect 416278 268779 416330 268831
rect 378742 268705 378794 268757
rect 526102 268705 526154 268757
rect 238870 268631 238922 268683
rect 378358 268631 378410 268683
rect 238294 268557 238346 268609
rect 366742 268557 366794 268609
rect 370774 268557 370826 268609
rect 376822 268557 376874 268609
rect 377014 268557 377066 268609
rect 378550 268557 378602 268609
rect 388438 268557 388490 268609
rect 237142 268483 237194 268535
rect 358582 268483 358634 268535
rect 366550 268483 366602 268535
rect 378646 268483 378698 268535
rect 378838 268483 378890 268535
rect 387286 268483 387338 268535
rect 388534 268483 388586 268535
rect 389206 268631 389258 268683
rect 415126 268631 415178 268683
rect 388918 268557 388970 268609
rect 389398 268557 389450 268609
rect 389494 268557 389546 268609
rect 395350 268557 395402 268609
rect 395446 268557 395498 268609
rect 399574 268557 399626 268609
rect 210934 268409 210986 268461
rect 271990 268409 272042 268461
rect 272758 268409 272810 268461
rect 228790 268335 228842 268387
rect 274198 268335 274250 268387
rect 287062 268335 287114 268387
rect 316918 268409 316970 268461
rect 336502 268409 336554 268461
rect 336598 268409 336650 268461
rect 337366 268409 337418 268461
rect 337750 268409 337802 268461
rect 366454 268409 366506 268461
rect 366646 268409 366698 268461
rect 377878 268409 377930 268461
rect 378934 268409 378986 268461
rect 388438 268409 388490 268461
rect 399286 268483 399338 268535
rect 403702 268483 403754 268535
rect 406102 268483 406154 268535
rect 501142 268409 501194 268461
rect 222550 268261 222602 268313
rect 259702 268261 259754 268313
rect 260086 268261 260138 268313
rect 292150 268261 292202 268313
rect 296662 268261 296714 268313
rect 312694 268261 312746 268313
rect 218038 268187 218090 268239
rect 272662 268187 272714 268239
rect 277654 268187 277706 268239
rect 282262 268187 282314 268239
rect 283510 268187 283562 268239
rect 316534 268187 316586 268239
rect 318262 268335 318314 268387
rect 318550 268335 318602 268387
rect 322966 268335 323018 268387
rect 323062 268335 323114 268387
rect 338326 268335 338378 268387
rect 360982 268335 361034 268387
rect 483286 268335 483338 268387
rect 317110 268261 317162 268313
rect 326710 268261 326762 268313
rect 326806 268261 326858 268313
rect 332278 268261 332330 268313
rect 332566 268261 332618 268313
rect 337462 268261 337514 268313
rect 348502 268261 348554 268313
rect 374326 268261 374378 268313
rect 374422 268261 374474 268313
rect 376342 268261 376394 268313
rect 376822 268261 376874 268313
rect 388726 268261 388778 268313
rect 388822 268261 388874 268313
rect 554710 268261 554762 268313
rect 322582 268187 322634 268239
rect 322870 268187 322922 268239
rect 323926 268187 323978 268239
rect 324022 268187 324074 268239
rect 324502 268187 324554 268239
rect 324598 268187 324650 268239
rect 347542 268187 347594 268239
rect 359446 268187 359498 268239
rect 468982 268187 469034 268239
rect 223222 268113 223274 268165
rect 266806 268113 266858 268165
rect 267382 268113 267434 268165
rect 268054 268113 268106 268165
rect 294550 268113 294602 268165
rect 318358 268113 318410 268165
rect 318454 268113 318506 268165
rect 325654 268113 325706 268165
rect 328438 268113 328490 268165
rect 336982 268113 337034 268165
rect 355702 268113 355754 268165
rect 440470 268113 440522 268165
rect 235894 268039 235946 268091
rect 274870 268039 274922 268091
rect 286006 268039 286058 268091
rect 316246 268039 316298 268091
rect 317110 268039 317162 268091
rect 326998 268039 327050 268091
rect 327766 268039 327818 268091
rect 336406 268039 336458 268091
rect 337366 268039 337418 268091
rect 348598 268039 348650 268091
rect 353974 268039 354026 268091
rect 426262 268039 426314 268091
rect 262006 267965 262058 268017
rect 324022 267965 324074 268017
rect 324118 267965 324170 268017
rect 326614 267965 326666 268017
rect 326710 267965 326762 268017
rect 328246 267965 328298 268017
rect 328342 267965 328394 268017
rect 438070 267965 438122 268017
rect 439126 267965 439178 268017
rect 449110 267965 449162 268017
rect 243094 267891 243146 267943
rect 275734 267891 275786 267943
rect 285046 267891 285098 267943
rect 316150 267891 316202 267943
rect 316246 267891 316298 267943
rect 212278 267817 212330 267869
rect 241078 267817 241130 267869
rect 258550 267817 258602 267869
rect 309622 267817 309674 267869
rect 318550 267891 318602 267943
rect 321334 267891 321386 267943
rect 336598 267891 336650 267943
rect 338326 267891 338378 267943
rect 377014 267891 377066 267943
rect 377878 267891 377930 267943
rect 378262 267891 378314 267943
rect 378550 267891 378602 267943
rect 385462 267891 385514 267943
rect 385558 267891 385610 267943
rect 317878 267817 317930 267869
rect 332566 267817 332618 267869
rect 334102 267817 334154 267869
rect 335062 267817 335114 267869
rect 337462 267817 337514 267869
rect 349078 267817 349130 267869
rect 366358 267817 366410 267869
rect 377974 267817 378026 267869
rect 378358 267817 378410 267869
rect 397270 267817 397322 267869
rect 397558 267891 397610 267943
rect 408790 267891 408842 267943
rect 408406 267817 408458 267869
rect 204982 267743 205034 267795
rect 221782 267743 221834 267795
rect 251926 267743 251978 267795
rect 258646 267743 258698 267795
rect 267478 267743 267530 267795
rect 269302 267743 269354 267795
rect 312022 267743 312074 267795
rect 312118 267743 312170 267795
rect 327766 267743 327818 267795
rect 327862 267743 327914 267795
rect 337750 267743 337802 267795
rect 338038 267743 338090 267795
rect 621238 267743 621290 267795
rect 219574 267669 219626 267721
rect 221782 267595 221834 267647
rect 197206 267521 197258 267573
rect 211510 267521 211562 267573
rect 251926 267595 251978 267647
rect 261814 267595 261866 267647
rect 241846 267521 241898 267573
rect 318262 267669 318314 267721
rect 267478 267595 267530 267647
rect 267766 267595 267818 267647
rect 287734 267595 287786 267647
rect 318454 267595 318506 267647
rect 279958 267521 280010 267573
rect 317110 267521 317162 267573
rect 317206 267521 317258 267573
rect 326902 267669 326954 267721
rect 326998 267669 327050 267721
rect 336118 267669 336170 267721
rect 336214 267669 336266 267721
rect 357334 267669 357386 267721
rect 357430 267669 357482 267721
rect 367798 267669 367850 267721
rect 368566 267669 368618 267721
rect 319222 267595 319274 267647
rect 326806 267595 326858 267647
rect 327094 267595 327146 267647
rect 344854 267595 344906 267647
rect 351286 267595 351338 267647
rect 322486 267521 322538 267573
rect 338038 267521 338090 267573
rect 353302 267521 353354 267573
rect 374998 267521 375050 267573
rect 256150 267447 256202 267499
rect 269014 267447 269066 267499
rect 241846 267373 241898 267425
rect 261814 267373 261866 267425
rect 269302 267373 269354 267425
rect 290326 267373 290378 267425
rect 338326 267447 338378 267499
rect 355030 267447 355082 267499
rect 297142 267373 297194 267425
rect 346582 267373 346634 267425
rect 347254 267373 347306 267425
rect 365206 267373 365258 267425
rect 367798 267447 367850 267499
rect 368758 267447 368810 267499
rect 369142 267447 369194 267499
rect 374806 267447 374858 267499
rect 375190 267595 375242 267647
rect 376822 267595 376874 267647
rect 376918 267595 376970 267647
rect 378358 267595 378410 267647
rect 378838 267669 378890 267721
rect 400054 267669 400106 267721
rect 401686 267669 401738 267721
rect 412822 267669 412874 267721
rect 397462 267595 397514 267647
rect 397558 267595 397610 267647
rect 404662 267595 404714 267647
rect 375382 267521 375434 267573
rect 419062 267521 419114 267573
rect 397558 267447 397610 267499
rect 397654 267447 397706 267499
rect 398806 267447 398858 267499
rect 398902 267447 398954 267499
rect 414358 267447 414410 267499
rect 433366 267373 433418 267425
rect 291670 267299 291722 267351
rect 367030 267299 367082 267351
rect 367126 267299 367178 267351
rect 378358 267299 378410 267351
rect 378454 267299 378506 267351
rect 385846 267299 385898 267351
rect 387478 267299 387530 267351
rect 608182 267299 608234 267351
rect 289462 267225 289514 267277
rect 353686 267225 353738 267277
rect 356566 267225 356618 267277
rect 369046 267225 369098 267277
rect 369334 267225 369386 267277
rect 447670 267225 447722 267277
rect 293590 267151 293642 267203
rect 367126 267151 367178 267203
rect 262102 267077 262154 267129
rect 309430 267077 309482 267129
rect 309622 267077 309674 267129
rect 317878 267077 317930 267129
rect 318262 267077 318314 267129
rect 328534 267077 328586 267129
rect 328630 267077 328682 267129
rect 348502 267077 348554 267129
rect 348598 267077 348650 267129
rect 377014 267151 377066 267203
rect 377206 267151 377258 267203
rect 387478 267151 387530 267203
rect 387574 267151 387626 267203
rect 398518 267151 398570 267203
rect 398806 267151 398858 267203
rect 421462 267151 421514 267203
rect 367318 267077 367370 267129
rect 375190 267077 375242 267129
rect 375958 267077 376010 267129
rect 458326 267077 458378 267129
rect 295318 267003 295370 267055
rect 378838 267003 378890 267055
rect 378934 267003 378986 267055
rect 398230 267003 398282 267055
rect 295990 266929 296042 266981
rect 397174 266929 397226 266981
rect 397270 266929 397322 266981
rect 398518 266929 398570 266981
rect 399190 266929 399242 266981
rect 413686 266929 413738 266981
rect 251638 266855 251690 266907
rect 332374 266855 332426 266907
rect 349558 266855 349610 266907
rect 357430 266855 357482 266907
rect 359830 266855 359882 266907
rect 472630 266855 472682 266907
rect 296854 266781 296906 266833
rect 398902 266781 398954 266833
rect 399094 266781 399146 266833
rect 407158 266781 407210 266833
rect 288790 266707 288842 266759
rect 297142 266707 297194 266759
rect 298006 266707 298058 266759
rect 398806 266707 398858 266759
rect 399286 266707 399338 266759
rect 408790 266707 408842 266759
rect 298582 266633 298634 266685
rect 428662 266633 428714 266685
rect 199126 266559 199178 266611
rect 214966 266559 215018 266611
rect 244246 266559 244298 266611
rect 331702 266559 331754 266611
rect 338326 266559 338378 266611
rect 360790 266559 360842 266611
rect 362230 266559 362282 266611
rect 494038 266559 494090 266611
rect 237430 266485 237482 266537
rect 330646 266485 330698 266537
rect 331414 266485 331466 266537
rect 339382 266485 339434 266537
rect 362710 266485 362762 266537
rect 497590 266485 497642 266537
rect 244150 266411 244202 266463
rect 261910 266411 261962 266463
rect 299734 266411 299786 266463
rect 435670 266411 435722 266463
rect 300310 266337 300362 266389
rect 442870 266337 442922 266389
rect 301270 266263 301322 266315
rect 449974 266263 450026 266315
rect 230038 266189 230090 266241
rect 329974 266189 330026 266241
rect 347254 266189 347306 266241
rect 347830 266189 347882 266241
rect 357814 266189 357866 266241
rect 375958 266189 376010 266241
rect 376918 266189 376970 266241
rect 522550 266189 522602 266241
rect 302326 266115 302378 266167
rect 457174 266115 457226 266167
rect 255094 266041 255146 266093
rect 258646 266041 258698 266093
rect 302998 266041 303050 266093
rect 464278 266041 464330 266093
rect 304054 265967 304106 266019
rect 471382 265967 471434 266019
rect 226390 265893 226442 265945
rect 318358 265893 318410 265945
rect 318454 265893 318506 265945
rect 339094 265893 339146 265945
rect 367030 265893 367082 265945
rect 378358 265893 378410 265945
rect 378454 265893 378506 265945
rect 397846 265893 397898 265945
rect 398230 265893 398282 265945
rect 533206 265893 533258 265945
rect 304726 265819 304778 265871
rect 478582 265819 478634 265871
rect 212470 265745 212522 265797
rect 318838 265745 318890 265797
rect 318934 265745 318986 265797
rect 327862 265745 327914 265797
rect 327958 265745 328010 265797
rect 348502 265745 348554 265797
rect 350710 265745 350762 265797
rect 368566 265745 368618 265797
rect 368758 265745 368810 265797
rect 378742 265745 378794 265797
rect 378838 265745 378890 265797
rect 399094 265745 399146 265797
rect 399190 265745 399242 265797
rect 547606 265745 547658 265797
rect 305590 265671 305642 265723
rect 485686 265671 485738 265723
rect 306742 265597 306794 265649
rect 318742 265597 318794 265649
rect 319030 265597 319082 265649
rect 492886 265597 492938 265649
rect 307318 265523 307370 265575
rect 499894 265523 499946 265575
rect 269014 265449 269066 265501
rect 288502 265449 288554 265501
rect 309334 265449 309386 265501
rect 309910 265375 309962 265427
rect 318550 265375 318602 265427
rect 319222 265375 319274 265427
rect 319702 265375 319754 265427
rect 321046 265375 321098 265427
rect 311638 265301 311690 265353
rect 318934 265301 318986 265353
rect 221686 265227 221738 265279
rect 273142 265227 273194 265279
rect 313270 265227 313322 265279
rect 318838 265227 318890 265279
rect 326470 265301 326522 265353
rect 326614 265301 326666 265353
rect 201430 265153 201482 265205
rect 79222 265005 79274 265057
rect 262102 265153 262154 265205
rect 282262 265153 282314 265205
rect 255670 265079 255722 265131
rect 267574 265079 267626 265131
rect 262102 265005 262154 265057
rect 282262 265005 282314 265057
rect 86422 264931 86474 264983
rect 211222 264931 211274 264983
rect 212278 264931 212330 264983
rect 256630 264931 256682 264983
rect 268246 264931 268298 264983
rect 287542 264931 287594 264983
rect 312022 265153 312074 265205
rect 316630 265153 316682 265205
rect 316534 265079 316586 265131
rect 317686 265153 317738 265205
rect 318742 265153 318794 265205
rect 319702 265227 319754 265279
rect 319318 265153 319370 265205
rect 329302 265153 329354 265205
rect 332278 265153 332330 265205
rect 367318 265153 367370 265205
rect 318550 265079 318602 265131
rect 318934 265079 318986 265131
rect 319222 265079 319274 265131
rect 326614 265079 326666 265131
rect 337078 265079 337130 265131
rect 337558 265079 337610 265131
rect 344854 265079 344906 265131
rect 374230 265079 374282 265131
rect 374806 265375 374858 265427
rect 376438 265375 376490 265427
rect 377206 265375 377258 265427
rect 378934 265375 378986 265427
rect 379126 265449 379178 265501
rect 387190 265449 387242 265501
rect 514294 265449 514346 265501
rect 399862 265375 399914 265427
rect 521398 265375 521450 265427
rect 378742 265301 378794 265353
rect 390550 265301 390602 265353
rect 392854 265301 392906 265353
rect 393622 265301 393674 265353
rect 398710 265301 398762 265353
rect 535606 265301 535658 265353
rect 398518 265153 398570 265205
rect 398998 265227 399050 265279
rect 546358 265227 546410 265279
rect 399862 265153 399914 265205
rect 406486 265153 406538 265205
rect 408118 265153 408170 265205
rect 411766 265153 411818 265205
rect 412054 265153 412106 265205
rect 309430 265005 309482 265057
rect 333622 265005 333674 265057
rect 365974 265005 366026 265057
rect 376726 265005 376778 265057
rect 377206 265005 377258 265057
rect 393334 265079 393386 265131
rect 615382 265079 615434 265131
rect 210646 264857 210698 264909
rect 212470 264857 212522 264909
rect 318742 264931 318794 264983
rect 318934 264931 318986 264983
rect 321046 264931 321098 264983
rect 348598 264931 348650 264983
rect 365206 264931 365258 264983
rect 385654 264931 385706 264983
rect 348502 264857 348554 264909
rect 382390 264857 382442 264909
rect 383446 264857 383498 264909
rect 392854 264931 392906 264983
rect 398998 265005 399050 265057
rect 399094 265005 399146 265057
rect 629686 265005 629738 265057
rect 393334 264931 393386 264983
rect 396982 264931 397034 264983
rect 398614 264931 398666 264983
rect 399574 264931 399626 264983
rect 412630 264931 412682 264983
rect 388983 264857 389035 264909
rect 412726 264857 412778 264909
rect 449398 264709 449450 264761
rect 469366 264709 469418 264761
rect 475798 264709 475850 264761
rect 489526 264709 489578 264761
rect 159862 263451 159914 263503
rect 161110 263451 161162 263503
rect 182230 262119 182282 262171
rect 192982 262045 193034 262097
rect 72022 260639 72074 260691
rect 84694 260639 84746 260691
rect 42454 259677 42506 259729
rect 53878 259677 53930 259729
rect 86422 259233 86474 259285
rect 632470 259233 632522 259285
rect 642166 259233 642218 259285
rect 92278 259159 92330 259211
rect 42838 258937 42890 258989
rect 50326 258937 50378 258989
rect 42454 258641 42506 258693
rect 47446 258641 47498 258693
rect 42454 257827 42506 257879
rect 43222 257827 43274 257879
rect 616342 257753 616394 257805
rect 630742 257753 630794 257805
rect 197110 257605 197162 257657
rect 212086 257605 212138 257657
rect 674614 256421 674666 256473
rect 674902 256421 674954 256473
rect 639286 256347 639338 256399
rect 677110 256347 677162 256399
rect 92278 254867 92330 254919
rect 104374 254867 104426 254919
rect 84694 253461 84746 253513
rect 92182 253387 92234 253439
rect 192982 253387 193034 253439
rect 198742 253387 198794 253439
rect 674614 253387 674666 253439
rect 675286 253387 675338 253439
rect 674518 252721 674570 252773
rect 675094 252721 675146 252773
rect 92182 250501 92234 250553
rect 97174 250501 97226 250553
rect 607702 250501 607754 250553
rect 616342 250575 616394 250627
rect 104374 250057 104426 250109
rect 106582 250057 106634 250109
rect 56182 249243 56234 249295
rect 205654 249243 205706 249295
rect 53782 249169 53834 249221
rect 210742 249169 210794 249221
rect 47638 249095 47690 249147
rect 206902 249095 206954 249147
rect 627862 248059 627914 248111
rect 632470 248059 632522 248111
rect 674422 247911 674474 247963
rect 675478 247911 675530 247963
rect 198742 247689 198794 247741
rect 211030 247689 211082 247741
rect 211318 247689 211370 247741
rect 209398 247615 209450 247667
rect 126550 247319 126602 247371
rect 129526 247245 129578 247297
rect 135190 247171 135242 247223
rect 132310 247097 132362 247149
rect 140950 247023 141002 247075
rect 65206 246727 65258 246779
rect 81142 246949 81194 247001
rect 143926 246949 143978 247001
rect 146710 246875 146762 246927
rect 181462 246801 181514 246853
rect 197590 246801 197642 246853
rect 211798 246801 211850 246853
rect 81142 246727 81194 246779
rect 205078 246727 205130 246779
rect 212278 246727 212330 246779
rect 227062 246727 227114 246779
rect 65014 246653 65066 246705
rect 80662 246653 80714 246705
rect 80950 246653 81002 246705
rect 210934 246653 210986 246705
rect 211894 246653 211946 246705
rect 385078 246727 385130 246779
rect 386998 246727 387050 246779
rect 388054 246727 388106 246779
rect 390262 246727 390314 246779
rect 237814 246653 237866 246705
rect 267478 246653 267530 246705
rect 267574 246653 267626 246705
rect 268630 246653 268682 246705
rect 56086 246579 56138 246631
rect 80758 246579 80810 246631
rect 81238 246579 81290 246631
rect 204886 246579 204938 246631
rect 276694 246653 276746 246705
rect 53206 246505 53258 246557
rect 204694 246505 204746 246557
rect 212182 246505 212234 246557
rect 269302 246579 269354 246631
rect 276886 246579 276938 246631
rect 232150 246505 232202 246557
rect 266614 246505 266666 246557
rect 266710 246505 266762 246557
rect 267574 246505 267626 246557
rect 267958 246505 268010 246557
rect 276598 246505 276650 246557
rect 276694 246505 276746 246557
rect 277366 246579 277418 246631
rect 278614 246579 278666 246631
rect 278806 246653 278858 246705
rect 288022 246653 288074 246705
rect 288886 246579 288938 246631
rect 297910 246579 297962 246631
rect 298006 246579 298058 246631
rect 302422 246579 302474 246631
rect 53398 246431 53450 246483
rect 204790 246431 204842 246483
rect 211702 246431 211754 246483
rect 226966 246431 227018 246483
rect 47734 246357 47786 246409
rect 210166 246357 210218 246409
rect 212086 246357 212138 246409
rect 221782 246357 221834 246409
rect 221878 246357 221930 246409
rect 276886 246431 276938 246483
rect 278710 246505 278762 246557
rect 308086 246579 308138 246631
rect 308470 246653 308522 246705
rect 350134 246653 350186 246705
rect 352342 246653 352394 246705
rect 362614 246653 362666 246705
rect 334870 246579 334922 246631
rect 334966 246579 335018 246631
rect 353206 246579 353258 246631
rect 353302 246579 353354 246631
rect 362806 246579 362858 246631
rect 368950 246579 369002 246631
rect 369142 246653 369194 246705
rect 389494 246653 389546 246705
rect 397654 246653 397706 246705
rect 402166 246727 402218 246779
rect 406102 246727 406154 246779
rect 406524 246778 406576 246830
rect 674326 247023 674378 247075
rect 675478 247023 675530 247075
rect 408982 246727 409034 246779
rect 409366 246727 409418 246779
rect 409462 246727 409514 246779
rect 412150 246727 412202 246779
rect 674710 246727 674762 246779
rect 675382 246727 675434 246779
rect 408790 246653 408842 246705
rect 402070 246579 402122 246631
rect 402166 246579 402218 246631
rect 406774 246579 406826 246631
rect 231862 246357 231914 246409
rect 304438 246431 304490 246483
rect 312406 246431 312458 246483
rect 44854 246283 44906 246335
rect 209686 246283 209738 246335
rect 209974 246283 210026 246335
rect 247222 246283 247274 246335
rect 267766 246283 267818 246335
rect 298006 246357 298058 246409
rect 298102 246357 298154 246409
rect 299254 246357 299306 246409
rect 302422 246357 302474 246409
rect 334966 246431 335018 246483
rect 335350 246505 335402 246557
rect 396790 246505 396842 246557
rect 397654 246505 397706 246557
rect 412054 246505 412106 246557
rect 322006 246357 322058 246409
rect 44950 246209 45002 246261
rect 80758 246209 80810 246261
rect 80950 246209 81002 246261
rect 209590 246209 209642 246261
rect 209878 246209 209930 246261
rect 237814 246209 237866 246261
rect 240502 246209 240554 246261
rect 277366 246209 277418 246261
rect 307990 246283 308042 246335
rect 308086 246283 308138 246335
rect 287638 246209 287690 246261
rect 118102 246135 118154 246187
rect 128086 246135 128138 246187
rect 46198 246061 46250 246113
rect 60502 246061 60554 246113
rect 66262 246061 66314 246113
rect 77782 246061 77834 246113
rect 97846 245987 97898 246039
rect 118102 245987 118154 246039
rect 128086 245987 128138 246039
rect 141142 245987 141194 246039
rect 151126 245987 151178 246039
rect 170902 246135 170954 246187
rect 211990 246135 212042 246187
rect 267766 246135 267818 246187
rect 267862 246135 267914 246187
rect 269302 246135 269354 246187
rect 272854 246135 272906 246187
rect 278038 246135 278090 246187
rect 278134 246135 278186 246187
rect 292246 246209 292298 246261
rect 292342 246209 292394 246261
rect 294166 246209 294218 246261
rect 294550 246209 294602 246261
rect 301270 246209 301322 246261
rect 301366 246209 301418 246261
rect 329686 246283 329738 246335
rect 288118 246135 288170 246187
rect 308470 246135 308522 246187
rect 308566 246135 308618 246187
rect 322006 246135 322058 246187
rect 334774 246209 334826 246261
rect 335158 246283 335210 246335
rect 352342 246283 352394 246335
rect 353206 246357 353258 246409
rect 378646 246357 378698 246409
rect 388534 246357 388586 246409
rect 389782 246357 389834 246409
rect 397366 246431 397418 246483
rect 407254 246431 407306 246483
rect 408598 246357 408650 246409
rect 387286 246283 387338 246335
rect 388918 246283 388970 246335
rect 407638 246283 407690 246335
rect 329686 246135 329738 246187
rect 330742 246135 330794 246187
rect 358006 246135 358058 246187
rect 181558 246061 181610 246113
rect 205846 246061 205898 246113
rect 170902 245987 170954 246039
rect 181462 245987 181514 246039
rect 205846 245913 205898 245965
rect 216022 246061 216074 246113
rect 237718 246061 237770 246113
rect 242518 246061 242570 246113
rect 227062 245987 227114 246039
rect 231862 245987 231914 246039
rect 240022 245987 240074 246039
rect 241750 245987 241802 246039
rect 236086 245913 236138 245965
rect 266518 246061 266570 246113
rect 266614 246061 266666 246113
rect 278614 246061 278666 246113
rect 278710 246061 278762 246113
rect 285910 246061 285962 246113
rect 286102 246061 286154 246113
rect 292630 246061 292682 246113
rect 292726 246061 292778 246113
rect 304438 246061 304490 246113
rect 304534 246061 304586 246113
rect 308950 246061 309002 246113
rect 312406 246061 312458 246113
rect 342742 246061 342794 246113
rect 350134 246061 350186 246113
rect 353302 246061 353354 246113
rect 378646 246209 378698 246261
rect 412246 246209 412298 246261
rect 389302 246135 389354 246187
rect 396790 246135 396842 246187
rect 406198 246135 406250 246187
rect 387382 246061 387434 246113
rect 388918 246061 388970 246113
rect 247222 245987 247274 246039
rect 252502 245987 252554 246039
rect 262582 245987 262634 246039
rect 277750 245987 277802 246039
rect 263830 245913 263882 245965
rect 367510 245987 367562 246039
rect 367702 245987 367754 246039
rect 505366 246061 505418 246113
rect 674806 246061 674858 246113
rect 675382 246061 675434 246113
rect 389302 245987 389354 246039
rect 409846 245987 409898 246039
rect 278038 245913 278090 245965
rect 368086 245913 368138 245965
rect 385078 245913 385130 245965
rect 409174 245913 409226 245965
rect 77782 245839 77834 245891
rect 97846 245839 97898 245891
rect 141142 245839 141194 245891
rect 151126 245839 151178 245891
rect 237046 245839 237098 245891
rect 252694 245839 252746 245891
rect 255094 245839 255146 245891
rect 338134 245839 338186 245891
rect 338230 245839 338282 245891
rect 357430 245839 357482 245891
rect 387286 245839 387338 245891
rect 409462 245839 409514 245891
rect 210838 245765 210890 245817
rect 227350 245765 227402 245817
rect 251350 245765 251402 245817
rect 356278 245765 356330 245817
rect 388054 245765 388106 245817
rect 397366 245765 397418 245817
rect 226966 245691 227018 245743
rect 232150 245691 232202 245743
rect 254134 245691 254186 245743
rect 330742 245691 330794 245743
rect 330838 245691 330890 245743
rect 357142 245691 357194 245743
rect 386998 245691 387050 245743
rect 390262 245691 390314 245743
rect 402070 245691 402122 245743
rect 407062 245691 407114 245743
rect 216022 245617 216074 245669
rect 236086 245617 236138 245669
rect 263062 245617 263114 245669
rect 210550 245543 210602 245595
rect 277750 245543 277802 245595
rect 277942 245617 277994 245669
rect 370966 245617 371018 245669
rect 369238 245543 369290 245595
rect 250294 245469 250346 245521
rect 338518 245469 338570 245521
rect 253366 245395 253418 245447
rect 338230 245395 338282 245447
rect 249622 245321 249674 245373
rect 355798 245395 355850 245447
rect 338422 245321 338474 245373
rect 358102 245321 358154 245373
rect 252406 245247 252458 245299
rect 330838 245247 330890 245299
rect 330934 245247 330986 245299
rect 358582 245395 358634 245447
rect 405910 245395 405962 245447
rect 412438 245395 412490 245447
rect 358486 245321 358538 245373
rect 362902 245321 362954 245373
rect 210166 245173 210218 245225
rect 214006 245173 214058 245225
rect 216598 245173 216650 245225
rect 358582 245173 358634 245225
rect 209590 245099 209642 245151
rect 213526 245099 213578 245151
rect 226390 245099 226442 245151
rect 251926 245099 251978 245151
rect 261814 245099 261866 245151
rect 372022 245173 372074 245225
rect 411478 245173 411530 245225
rect 405718 245099 405770 245151
rect 42454 245025 42506 245077
rect 214294 245025 214346 245077
rect 260854 245025 260906 245077
rect 374038 245025 374090 245077
rect 210070 244951 210122 245003
rect 252118 244951 252170 245003
rect 260758 244951 260810 245003
rect 374614 244951 374666 245003
rect 209686 244877 209738 244929
rect 213142 244877 213194 244929
rect 216502 244877 216554 244929
rect 106582 244803 106634 244855
rect 210070 244803 210122 244855
rect 149590 244729 149642 244781
rect 97174 244655 97226 244707
rect 142486 244655 142538 244707
rect 251926 244803 251978 244855
rect 319798 244803 319850 244855
rect 319990 244803 320042 244855
rect 330934 244803 330986 244855
rect 338518 244877 338570 244929
rect 355894 244877 355946 244929
rect 353590 244803 353642 244855
rect 252118 244729 252170 244781
rect 285718 244729 285770 244781
rect 285910 244729 285962 244781
rect 292726 244729 292778 244781
rect 292822 244729 292874 244781
rect 389302 244877 389354 244929
rect 268246 244655 268298 244707
rect 138166 244581 138218 244633
rect 206806 244581 206858 244633
rect 266518 244581 266570 244633
rect 277942 244655 277994 244707
rect 278038 244655 278090 244707
rect 277750 244581 277802 244633
rect 135286 244507 135338 244559
rect 204982 244507 205034 244559
rect 277366 244507 277418 244559
rect 282262 244507 282314 244559
rect 282454 244581 282506 244633
rect 288022 244581 288074 244633
rect 288214 244655 288266 244707
rect 408118 244803 408170 244855
rect 603094 244729 603146 244781
rect 607702 244803 607754 244855
rect 306646 244581 306698 244633
rect 306742 244581 306794 244633
rect 319702 244581 319754 244633
rect 342742 244581 342794 244633
rect 367702 244581 367754 244633
rect 291862 244507 291914 244559
rect 291958 244507 292010 244559
rect 301366 244507 301418 244559
rect 302326 244507 302378 244559
rect 304534 244507 304586 244559
rect 132406 244433 132458 244485
rect 205558 244433 205610 244485
rect 263446 244433 263498 244485
rect 272854 244433 272906 244485
rect 310774 244507 310826 244559
rect 312022 244507 312074 244559
rect 367606 244507 367658 244559
rect 126646 244359 126698 244411
rect 205366 244359 205418 244411
rect 264790 244359 264842 244411
rect 307894 244433 307946 244485
rect 308278 244433 308330 244485
rect 312214 244433 312266 244485
rect 319798 244433 319850 244485
rect 319894 244433 319946 244485
rect 321334 244433 321386 244485
rect 277846 244359 277898 244411
rect 310486 244359 310538 244411
rect 339862 244359 339914 244411
rect 368758 244433 368810 244485
rect 123766 244285 123818 244337
rect 205174 244285 205226 244337
rect 256534 244285 256586 244337
rect 276310 244285 276362 244337
rect 277942 244285 277994 244337
rect 306742 244285 306794 244337
rect 312406 244285 312458 244337
rect 339766 244285 339818 244337
rect 120886 244211 120938 244263
rect 205654 244211 205706 244263
rect 235126 244211 235178 244263
rect 267190 244211 267242 244263
rect 275926 244211 275978 244263
rect 276406 244211 276458 244263
rect 276598 244211 276650 244263
rect 318262 244211 318314 244263
rect 118006 244137 118058 244189
rect 204502 244137 204554 244189
rect 260086 244137 260138 244189
rect 318070 244137 318122 244189
rect 112246 244063 112298 244115
rect 206326 244063 206378 244115
rect 256342 244063 256394 244115
rect 335350 244063 335402 244115
rect 109366 243989 109418 244041
rect 206518 243989 206570 244041
rect 258358 243989 258410 244041
rect 336310 243989 336362 244041
rect 106486 243915 106538 243967
rect 205750 243915 205802 243967
rect 261142 243915 261194 243967
rect 318166 243915 318218 243967
rect 103606 243841 103658 243893
rect 206134 243841 206186 243893
rect 207190 243841 207242 243893
rect 268150 243841 268202 243893
rect 268246 243841 268298 243893
rect 287926 243841 287978 243893
rect 288022 243841 288074 243893
rect 292150 243841 292202 243893
rect 292246 243841 292298 243893
rect 307318 243841 307370 243893
rect 313366 243841 313418 243893
rect 370294 243841 370346 243893
rect 100726 243767 100778 243819
rect 206230 243767 206282 243819
rect 245398 243767 245450 243819
rect 353686 243767 353738 243819
rect 94966 243693 95018 243745
rect 205942 243693 205994 243745
rect 239350 243693 239402 243745
rect 350806 243693 350858 243745
rect 92086 243619 92138 243671
rect 206422 243619 206474 243671
rect 231766 243619 231818 243671
rect 347350 243619 347402 243671
rect 86326 243545 86378 243597
rect 206710 243545 206762 243597
rect 236278 243545 236330 243597
rect 349270 243545 349322 243597
rect 80566 243471 80618 243523
rect 206998 243471 207050 243523
rect 221206 243471 221258 243523
rect 227446 243471 227498 243523
rect 229750 243471 229802 243523
rect 346390 243471 346442 243523
rect 77686 243397 77738 243449
rect 204598 243397 204650 243449
rect 226774 243397 226826 243449
rect 345142 243397 345194 243449
rect 69046 243323 69098 243375
rect 206038 243323 206090 243375
rect 228502 243323 228554 243375
rect 345622 243323 345674 243375
rect 265942 243249 265994 243301
rect 277846 243249 277898 243301
rect 283702 243249 283754 243301
rect 298102 243249 298154 243301
rect 298294 243249 298346 243301
rect 299638 243249 299690 243301
rect 302422 243249 302474 243301
rect 312214 243249 312266 243301
rect 318262 243249 318314 243301
rect 340726 243249 340778 243301
rect 226006 243175 226058 243227
rect 236182 243175 236234 243227
rect 253366 243175 253418 243227
rect 256246 243175 256298 243227
rect 267382 243175 267434 243227
rect 262870 243101 262922 243153
rect 277942 243101 277994 243153
rect 284950 243101 285002 243153
rect 298006 243101 298058 243153
rect 318166 243175 318218 243227
rect 337558 243175 337610 243227
rect 305110 243101 305162 243153
rect 310486 243101 310538 243153
rect 339862 243101 339914 243153
rect 236182 243027 236234 243079
rect 253366 243027 253418 243079
rect 270838 243027 270890 243079
rect 291574 243027 291626 243079
rect 291766 243027 291818 243079
rect 294742 243027 294794 243079
rect 295318 243027 295370 243079
rect 303382 243027 303434 243079
rect 303478 243027 303530 243079
rect 320374 243027 320426 243079
rect 266038 242953 266090 243005
rect 277750 242953 277802 243005
rect 277846 242953 277898 243005
rect 279382 242953 279434 243005
rect 283222 242953 283274 243005
rect 302422 242953 302474 243005
rect 306454 242953 306506 243005
rect 316726 242953 316778 243005
rect 318070 242953 318122 243005
rect 337078 242953 337130 243005
rect 674998 242953 675050 243005
rect 675382 242953 675434 243005
rect 268150 242879 268202 242931
rect 287542 242879 287594 242931
rect 291382 242879 291434 242931
rect 292822 242879 292874 242931
rect 292918 242879 292970 242931
rect 302326 242879 302378 242931
rect 303094 242879 303146 242931
rect 312598 242879 312650 242931
rect 316534 242879 316586 242931
rect 266614 242805 266666 242857
rect 278038 242805 278090 242857
rect 285910 242805 285962 242857
rect 43414 242731 43466 242783
rect 46198 242731 46250 242783
rect 269206 242731 269258 242783
rect 294550 242731 294602 242783
rect 269686 242657 269738 242709
rect 285526 242657 285578 242709
rect 285718 242657 285770 242709
rect 291382 242657 291434 242709
rect 291574 242657 291626 242709
rect 293398 242657 293450 242709
rect 293494 242657 293546 242709
rect 294646 242657 294698 242709
rect 295126 242805 295178 242857
rect 297622 242805 297674 242857
rect 298006 242805 298058 242857
rect 317110 242805 317162 242857
rect 325078 242879 325130 242931
rect 339574 242879 339626 242931
rect 331126 242805 331178 242857
rect 295030 242731 295082 242783
rect 297814 242731 297866 242783
rect 298102 242731 298154 242783
rect 320086 242731 320138 242783
rect 314902 242657 314954 242709
rect 314998 242657 315050 242709
rect 316726 242657 316778 242709
rect 319702 242657 319754 242709
rect 338518 242657 338570 242709
rect 463702 242657 463754 242709
rect 483766 242657 483818 242709
rect 265270 242583 265322 242635
rect 277366 242583 277418 242635
rect 269878 242509 269930 242561
rect 277558 242509 277610 242561
rect 247510 242435 247562 242487
rect 221974 242361 222026 242413
rect 247606 242361 247658 242413
rect 267862 242435 267914 242487
rect 295318 242583 295370 242635
rect 299638 242583 299690 242635
rect 322582 242583 322634 242635
rect 277846 242509 277898 242561
rect 291766 242509 291818 242561
rect 285526 242435 285578 242487
rect 286294 242435 286346 242487
rect 286486 242435 286538 242487
rect 314326 242509 314378 242561
rect 317494 242509 317546 242561
rect 317974 242509 318026 242561
rect 328150 242509 328202 242561
rect 328534 242509 328586 242561
rect 443638 242509 443690 242561
rect 453622 242509 453674 242561
rect 292150 242435 292202 242487
rect 292918 242435 292970 242487
rect 293590 242435 293642 242487
rect 323446 242435 323498 242487
rect 273526 242361 273578 242413
rect 287734 242287 287786 242339
rect 287926 242361 287978 242413
rect 303478 242361 303530 242413
rect 308950 242361 309002 242413
rect 339766 242361 339818 242413
rect 430486 242361 430538 242413
rect 443446 242361 443498 242413
rect 504022 242361 504074 242413
rect 511126 242361 511178 242413
rect 355222 242287 355274 242339
rect 39958 242213 40010 242265
rect 42550 242213 42602 242265
rect 227350 242213 227402 242265
rect 227734 242213 227786 242265
rect 244150 242213 244202 242265
rect 353014 242213 353066 242265
rect 238294 242139 238346 242191
rect 350038 242139 350090 242191
rect 39862 242065 39914 242117
rect 42358 242065 42410 242117
rect 40054 241991 40106 242043
rect 42550 241991 42602 242043
rect 348694 242065 348746 242117
rect 40246 241917 40298 241969
rect 43126 241917 43178 241969
rect 50326 241917 50378 241969
rect 205846 241917 205898 241969
rect 218710 241843 218762 241895
rect 234358 241843 234410 241895
rect 234550 241843 234602 241895
rect 241462 241991 241514 242043
rect 351766 241991 351818 242043
rect 238966 241917 239018 241969
rect 347830 241917 347882 241969
rect 248566 241843 248618 241895
rect 273526 241843 273578 241895
rect 274006 241843 274058 241895
rect 281974 241843 282026 241895
rect 286870 241843 286922 241895
rect 297718 241843 297770 241895
rect 297814 241843 297866 241895
rect 305014 241843 305066 241895
rect 317878 241843 317930 241895
rect 327862 241843 327914 241895
rect 328054 241843 328106 241895
rect 375094 241843 375146 241895
rect 378166 241843 378218 241895
rect 215446 241769 215498 241821
rect 221398 241769 221450 241821
rect 233494 241769 233546 241821
rect 238966 241769 239018 241821
rect 239062 241769 239114 241821
rect 260662 241769 260714 241821
rect 327958 241769 328010 241821
rect 328726 241769 328778 241821
rect 333910 241769 333962 241821
rect 334486 241769 334538 241821
rect 365878 241769 365930 241821
rect 377206 241769 377258 241821
rect 395926 241769 395978 241821
rect 407542 241769 407594 241821
rect 219286 241695 219338 241747
rect 233782 241695 233834 241747
rect 262006 241695 262058 241747
rect 264310 241695 264362 241747
rect 271990 241695 272042 241747
rect 278134 241695 278186 241747
rect 221494 241621 221546 241673
rect 232918 241621 232970 241673
rect 236470 241621 236522 241673
rect 264406 241621 264458 241673
rect 213910 241547 213962 241599
rect 229174 241547 229226 241599
rect 252790 241547 252842 241599
rect 325174 241621 325226 241673
rect 325270 241621 325322 241673
rect 327862 241621 327914 241673
rect 329974 241695 330026 241747
rect 331030 241695 331082 241747
rect 358294 241695 358346 241747
rect 361558 241695 361610 241747
rect 396406 241695 396458 241747
rect 330070 241621 330122 241673
rect 348406 241621 348458 241673
rect 363190 241621 363242 241673
rect 400150 241621 400202 241673
rect 269302 241547 269354 241599
rect 317974 241547 318026 241599
rect 320470 241547 320522 241599
rect 336118 241547 336170 241599
rect 348502 241547 348554 241599
rect 356566 241547 356618 241599
rect 360982 241547 361034 241599
rect 395830 241547 395882 241599
rect 395926 241547 395978 241599
rect 405526 241547 405578 241599
rect 674038 241547 674090 241599
rect 675478 241547 675530 241599
rect 223222 241473 223274 241525
rect 232150 241473 232202 241525
rect 239158 241473 239210 241525
rect 258550 241473 258602 241525
rect 278230 241473 278282 241525
rect 318166 241473 318218 241525
rect 319510 241473 319562 241525
rect 329590 241473 329642 241525
rect 331510 241473 331562 241525
rect 359350 241473 359402 241525
rect 361942 241473 361994 241525
rect 397462 241473 397514 241525
rect 255958 241399 256010 241451
rect 318070 241399 318122 241451
rect 327382 241399 327434 241451
rect 332950 241399 333002 241451
rect 364534 241399 364586 241451
rect 402742 241399 402794 241451
rect 247414 241325 247466 241377
rect 250390 241325 250442 241377
rect 254998 241325 255050 241377
rect 318358 241325 318410 241377
rect 326710 241325 326762 241377
rect 328918 241325 328970 241377
rect 329014 241325 329066 241377
rect 347926 241325 347978 241377
rect 362326 241325 362378 241377
rect 398422 241325 398474 241377
rect 226294 241251 226346 241303
rect 230710 241251 230762 241303
rect 254230 241251 254282 241303
rect 337846 241251 337898 241303
rect 363766 241251 363818 241303
rect 400726 241251 400778 241303
rect 225430 241177 225482 241229
rect 230902 241177 230954 241229
rect 253750 241177 253802 241229
rect 339382 241177 339434 241229
rect 339478 241177 339530 241229
rect 360502 241177 360554 241229
rect 364150 241177 364202 241229
rect 401878 241177 401930 241229
rect 244726 241103 244778 241155
rect 326902 241103 326954 241155
rect 326998 241103 327050 241155
rect 330166 241103 330218 241155
rect 332278 241103 332330 241155
rect 361078 241103 361130 241155
rect 362422 241103 362474 241155
rect 398998 241103 399050 241155
rect 225238 241029 225290 241081
rect 231190 241029 231242 241081
rect 237526 241029 237578 241081
rect 254614 241029 254666 241081
rect 273142 241029 273194 241081
rect 280438 241029 280490 241081
rect 280534 241029 280586 241081
rect 290614 241029 290666 241081
rect 291958 241029 292010 241081
rect 376150 241029 376202 241081
rect 379606 241029 379658 241081
rect 409942 241029 409994 241081
rect 220438 240955 220490 241007
rect 233398 240955 233450 241007
rect 237622 240955 237674 241007
rect 252886 240955 252938 241007
rect 255094 240955 255146 241007
rect 317878 240955 317930 241007
rect 318166 240955 318218 241007
rect 331702 240955 331754 241007
rect 333718 240955 333770 241007
rect 364342 240955 364394 241007
rect 367222 240955 367274 241007
rect 408886 240955 408938 241007
rect 216694 240881 216746 240933
rect 236182 240881 236234 240933
rect 237430 240881 237482 240933
rect 248086 240881 248138 240933
rect 252310 240881 252362 240933
rect 342646 240881 342698 240933
rect 365398 240881 365450 240933
rect 405142 240881 405194 240933
rect 219286 240807 219338 240859
rect 250678 240807 250730 240859
rect 251542 240807 251594 240859
rect 344182 240807 344234 240859
rect 365974 240807 366026 240859
rect 406102 240807 406154 240859
rect 232342 240733 232394 240785
rect 238678 240733 238730 240785
rect 251830 240733 251882 240785
rect 274390 240733 274442 240785
rect 274486 240733 274538 240785
rect 281878 240733 281930 240785
rect 282262 240733 282314 240785
rect 375766 240733 375818 240785
rect 379222 240733 379274 240785
rect 409270 240733 409322 240785
rect 218806 240659 218858 240711
rect 252022 240659 252074 240711
rect 41878 240585 41930 240637
rect 212758 240585 212810 240637
rect 233302 240585 233354 240637
rect 250582 240585 250634 240637
rect 345718 240659 345770 240711
rect 366742 240659 366794 240711
rect 407734 240659 407786 240711
rect 257878 240585 257930 240637
rect 348022 240585 348074 240637
rect 365014 240585 365066 240637
rect 404470 240585 404522 240637
rect 221782 240511 221834 240563
rect 237526 240511 237578 240563
rect 250198 240511 250250 240563
rect 346294 240511 346346 240563
rect 364630 240511 364682 240563
rect 403414 240511 403466 240563
rect 674134 240511 674186 240563
rect 675478 240511 675530 240563
rect 220246 240437 220298 240489
rect 248662 240437 248714 240489
rect 249718 240437 249770 240489
rect 257686 240437 257738 240489
rect 257878 240437 257930 240489
rect 350230 240437 350282 240489
rect 366358 240437 366410 240489
rect 407158 240437 407210 240489
rect 607606 240437 607658 240489
rect 627862 240437 627914 240489
rect 41878 240363 41930 240415
rect 219670 240363 219722 240415
rect 249814 240363 249866 240415
rect 274678 240363 274730 240415
rect 283894 240363 283946 240415
rect 284086 240363 284138 240415
rect 297334 240363 297386 240415
rect 297718 240363 297770 240415
rect 313174 240363 313226 240415
rect 315190 240363 315242 240415
rect 374422 240363 374474 240415
rect 377014 240363 377066 240415
rect 404950 240363 405002 240415
rect 218422 240289 218474 240341
rect 237622 240289 237674 240341
rect 240886 240289 240938 240341
rect 255094 240289 255146 240341
rect 262102 240289 262154 240341
rect 278134 240289 278186 240341
rect 278326 240289 278378 240341
rect 283990 240289 284042 240341
rect 287254 240289 287306 240341
rect 303094 240289 303146 240341
rect 306550 240289 306602 240341
rect 308950 240289 309002 240341
rect 313654 240289 313706 240341
rect 371830 240289 371882 240341
rect 378262 240289 378314 240341
rect 408310 240289 408362 240341
rect 237910 240215 237962 240267
rect 261622 240215 261674 240267
rect 217558 240141 217610 240193
rect 234742 240141 234794 240193
rect 236950 240141 237002 240193
rect 263350 240141 263402 240193
rect 42358 240067 42410 240119
rect 43318 240067 43370 240119
rect 222550 240067 222602 240119
rect 232534 240067 232586 240119
rect 237334 240067 237386 240119
rect 262198 240067 262250 240119
rect 220630 239993 220682 240045
rect 237430 239993 237482 240045
rect 236566 239919 236618 239971
rect 263926 239993 263978 240045
rect 256438 239845 256490 239897
rect 269302 240215 269354 240267
rect 277462 240215 277514 240267
rect 295606 240215 295658 240267
rect 275734 240141 275786 240193
rect 281686 240141 281738 240193
rect 281878 240141 281930 240193
rect 289462 240141 289514 240193
rect 291094 240141 291146 240193
rect 293302 240141 293354 240193
rect 293782 240141 293834 240193
rect 312118 240215 312170 240267
rect 314614 240215 314666 240267
rect 373558 240215 373610 240267
rect 376438 240215 376490 240267
rect 404086 240215 404138 240267
rect 297142 240141 297194 240193
rect 304438 240141 304490 240193
rect 313750 240141 313802 240193
rect 371350 240141 371402 240193
rect 381814 240141 381866 240193
rect 389878 240141 389930 240193
rect 272470 240067 272522 240119
rect 285526 240067 285578 240119
rect 289558 240067 289610 240119
rect 275446 239993 275498 240045
rect 287446 239993 287498 240045
rect 288694 239993 288746 240045
rect 291862 239993 291914 240045
rect 279478 239919 279530 239971
rect 282166 239919 282218 239971
rect 284854 239919 284906 239971
rect 287830 239919 287882 239971
rect 290422 239919 290474 239971
rect 295222 239919 295274 239971
rect 314230 240067 314282 240119
rect 372406 240067 372458 240119
rect 376054 240067 376106 240119
rect 403222 240067 403274 240119
rect 296278 239993 296330 240045
rect 329110 239993 329162 240045
rect 329686 239993 329738 240045
rect 355702 239993 355754 240045
rect 360214 239993 360266 240045
rect 314806 239919 314858 239971
rect 317878 239919 317930 239971
rect 326998 239919 327050 239971
rect 328246 239919 328298 239971
rect 352438 239919 352490 239971
rect 268726 239845 268778 239897
rect 280150 239845 280202 239897
rect 280438 239845 280490 239897
rect 283030 239845 283082 239897
rect 283990 239845 284042 239897
rect 291670 239845 291722 239897
rect 149590 239771 149642 239823
rect 157750 239771 157802 239823
rect 248374 239771 248426 239823
rect 257878 239771 257930 239823
rect 274198 239771 274250 239823
rect 281494 239771 281546 239823
rect 214486 239697 214538 239749
rect 225142 239697 225194 239749
rect 228022 239697 228074 239749
rect 229942 239697 229994 239749
rect 268246 239697 268298 239749
rect 270934 239697 270986 239749
rect 275830 239697 275882 239749
rect 280534 239697 280586 239749
rect 215926 239623 215978 239675
rect 218902 239623 218954 239675
rect 229078 239623 229130 239675
rect 230230 239623 230282 239675
rect 257206 239623 257258 239675
rect 269302 239623 269354 239675
rect 270262 239623 270314 239675
rect 272278 239623 272330 239675
rect 273526 239623 273578 239675
rect 278326 239623 278378 239675
rect 278902 239623 278954 239675
rect 279670 239623 279722 239675
rect 279766 239623 279818 239675
rect 284086 239771 284138 239823
rect 289462 239771 289514 239823
rect 313846 239845 313898 239897
rect 324406 239845 324458 239897
rect 291862 239771 291914 239823
rect 293782 239771 293834 239823
rect 294262 239771 294314 239823
rect 303574 239771 303626 239823
rect 315574 239771 315626 239823
rect 325270 239771 325322 239823
rect 326230 239771 326282 239823
rect 329014 239771 329066 239823
rect 329302 239845 329354 239897
rect 354550 239845 354602 239897
rect 343702 239771 343754 239823
rect 282166 239697 282218 239749
rect 296566 239697 296618 239749
rect 297622 239697 297674 239749
rect 301078 239697 301130 239749
rect 301846 239697 301898 239749
rect 306646 239697 306698 239749
rect 281686 239623 281738 239675
rect 227254 239549 227306 239601
rect 230326 239549 230378 239601
rect 269398 239549 269450 239601
rect 276310 239549 276362 239601
rect 277654 239549 277706 239601
rect 282934 239549 282986 239601
rect 283030 239549 283082 239601
rect 292150 239549 292202 239601
rect 293206 239623 293258 239675
rect 302806 239623 302858 239675
rect 302998 239623 303050 239675
rect 307606 239623 307658 239675
rect 307894 239623 307946 239675
rect 312790 239697 312842 239749
rect 322678 239697 322730 239749
rect 309526 239623 309578 239675
rect 310294 239623 310346 239675
rect 320854 239623 320906 239675
rect 324694 239623 324746 239675
rect 326998 239697 327050 239749
rect 349558 239697 349610 239749
rect 340918 239623 340970 239675
rect 294742 239549 294794 239601
rect 295990 239549 296042 239601
rect 304150 239549 304202 239601
rect 308854 239549 308906 239601
rect 310198 239549 310250 239601
rect 323062 239549 323114 239601
rect 341302 239549 341354 239601
rect 277078 239475 277130 239527
rect 283798 239475 283850 239527
rect 283894 239475 283946 239527
rect 294358 239475 294410 239527
rect 322198 239475 322250 239527
rect 338902 239475 338954 239527
rect 271030 239401 271082 239453
rect 277942 239401 277994 239453
rect 278038 239401 278090 239453
rect 281782 239401 281834 239453
rect 281974 239401 282026 239453
rect 290806 239401 290858 239453
rect 290998 239401 291050 239453
rect 307894 239401 307946 239453
rect 323446 239401 323498 239453
rect 341974 239401 342026 239453
rect 240310 239327 240362 239379
rect 244150 239327 244202 239379
rect 276694 239327 276746 239379
rect 284470 239327 284522 239379
rect 285046 239327 285098 239379
rect 298870 239327 298922 239379
rect 307798 239327 307850 239379
rect 309814 239327 309866 239379
rect 321238 239327 321290 239379
rect 337174 239327 337226 239379
rect 377782 239993 377834 240045
rect 406678 239993 406730 240045
rect 375670 239919 375722 239971
rect 378646 239845 378698 239897
rect 383830 239845 383882 239897
rect 384022 239919 384074 239971
rect 398614 239919 398666 239971
rect 402358 239845 402410 239897
rect 380566 239771 380618 239823
rect 384886 239771 384938 239823
rect 383254 239697 383306 239749
rect 384406 239697 384458 239749
rect 387286 239697 387338 239749
rect 400630 239697 400682 239749
rect 374806 239623 374858 239675
rect 382678 239623 382730 239675
rect 383638 239623 383690 239675
rect 385558 239623 385610 239675
rect 380086 239549 380138 239601
rect 383734 239549 383786 239601
rect 380854 239475 380906 239527
rect 388150 239475 388202 239527
rect 375190 239401 375242 239453
rect 387286 239401 387338 239453
rect 392086 239327 392138 239379
rect 224086 239253 224138 239305
rect 231574 239253 231626 239305
rect 276214 239253 276266 239305
rect 286006 239253 286058 239305
rect 235510 239179 235562 239231
rect 238966 239179 239018 239231
rect 271798 239179 271850 239231
rect 290422 239253 290474 239305
rect 290518 239253 290570 239305
rect 316054 239253 316106 239305
rect 317974 239253 318026 239305
rect 332758 239253 332810 239305
rect 360598 239253 360650 239305
rect 394102 239253 394154 239305
rect 287350 239179 287402 239231
rect 237142 239105 237194 239157
rect 241654 239105 241706 239157
rect 244630 239105 244682 239157
rect 246262 239105 246314 239157
rect 272662 239105 272714 239157
rect 291094 239105 291146 239157
rect 291478 239179 291530 239231
rect 301846 239179 301898 239231
rect 302518 239179 302570 239231
rect 307222 239179 307274 239231
rect 326614 239179 326666 239231
rect 348598 239179 348650 239231
rect 380086 239179 380138 239231
rect 386614 239179 386666 239231
rect 596182 239179 596234 239231
rect 603094 239179 603146 239231
rect 300022 239105 300074 239157
rect 318070 239105 318122 239157
rect 334582 239105 334634 239157
rect 373366 239105 373418 239157
rect 396886 239105 396938 239157
rect 146614 239031 146666 239083
rect 174166 239031 174218 239083
rect 236182 239031 236234 239083
rect 238198 239031 238250 239083
rect 238486 239031 238538 239083
rect 241846 239031 241898 239083
rect 228502 238957 228554 239009
rect 230806 238957 230858 239009
rect 240502 238957 240554 239009
rect 255670 238957 255722 239009
rect 260374 238957 260426 239009
rect 228118 238883 228170 238935
rect 231958 238883 232010 238935
rect 239542 238883 239594 238935
rect 257398 238883 257450 238935
rect 259990 238883 260042 238935
rect 277846 238883 277898 238935
rect 278518 238883 278570 238935
rect 280726 238883 280778 238935
rect 283414 239031 283466 239083
rect 298390 239031 298442 239083
rect 318358 239031 318410 239083
rect 336502 239031 336554 239083
rect 373846 239031 373898 239083
rect 384022 239031 384074 239083
rect 280918 238957 280970 239009
rect 293974 238957 294026 239009
rect 294070 238957 294122 239009
rect 303190 238957 303242 239009
rect 304726 238957 304778 239009
rect 308182 238957 308234 239009
rect 311638 238957 311690 239009
rect 323638 238957 323690 239009
rect 323734 238957 323786 239009
rect 376630 238957 376682 239009
rect 380470 238957 380522 239009
rect 387574 238957 387626 239009
rect 282262 238883 282314 238935
rect 284374 238883 284426 238935
rect 288310 238883 288362 238935
rect 288406 238883 288458 238935
rect 300598 238883 300650 238935
rect 300790 238883 300842 238935
rect 306262 238883 306314 238935
rect 316438 238883 316490 238935
rect 377302 238883 377354 238935
rect 381430 238883 381482 238935
rect 389206 238883 389258 238935
rect 240118 238809 240170 238861
rect 256822 238809 256874 238861
rect 257110 238809 257162 238861
rect 318358 238809 318410 238861
rect 318646 238809 318698 238861
rect 332182 238809 332234 238861
rect 332470 238809 332522 238861
rect 347446 238809 347498 238861
rect 351382 238809 351434 238861
rect 358870 238809 358922 238861
rect 368182 238809 368234 238861
rect 384598 238809 384650 238861
rect 227254 238735 227306 238787
rect 234070 238735 234122 238787
rect 257782 238735 257834 238787
rect 318166 238735 318218 238787
rect 226294 238661 226346 238713
rect 235606 238661 235658 238713
rect 256246 238661 256298 238713
rect 318262 238661 318314 238713
rect 248950 238587 249002 238639
rect 315958 238587 316010 238639
rect 316054 238587 316106 238639
rect 323734 238735 323786 238787
rect 331222 238735 331274 238787
rect 358774 238735 358826 238787
rect 368662 238735 368714 238787
rect 381046 238735 381098 238787
rect 319030 238661 319082 238713
rect 332374 238661 332426 238713
rect 334102 238661 334154 238713
rect 365302 238661 365354 238713
rect 319606 238587 319658 238639
rect 333430 238587 333482 238639
rect 333622 238587 333674 238639
rect 363286 238587 363338 238639
rect 42166 238513 42218 238565
rect 43030 238513 43082 238565
rect 227734 238513 227786 238565
rect 232822 238513 232874 238565
rect 255574 238513 255626 238565
rect 318070 238513 318122 238565
rect 318358 238513 318410 238565
rect 324118 238513 324170 238565
rect 329782 238513 329834 238565
rect 332470 238513 332522 238565
rect 334870 238513 334922 238565
rect 367030 238513 367082 238565
rect 254614 238439 254666 238491
rect 42454 238365 42506 238417
rect 43030 238365 43082 238417
rect 221110 238365 221162 238417
rect 246550 238365 246602 238417
rect 254134 238365 254186 238417
rect 332854 238439 332906 238491
rect 362230 238439 362282 238491
rect 366838 238439 366890 238491
rect 383350 238661 383402 238713
rect 370486 238587 370538 238639
rect 382294 238587 382346 238639
rect 370006 238513 370058 238565
rect 380950 238513 381002 238565
rect 381046 238513 381098 238565
rect 385942 238513 385994 238565
rect 369430 238439 369482 238491
rect 388822 238439 388874 238491
rect 218038 238291 218090 238343
rect 253462 238291 253514 238343
rect 258550 238291 258602 238343
rect 280918 238291 280970 238343
rect 283318 238291 283370 238343
rect 284854 238291 284906 238343
rect 285814 238291 285866 238343
rect 298966 238291 299018 238343
rect 299062 238291 299114 238343
rect 305782 238291 305834 238343
rect 305878 238291 305930 238343
rect 332470 238291 332522 238343
rect 221878 238217 221930 238269
rect 244822 238217 244874 238269
rect 252406 238217 252458 238269
rect 336982 238365 337034 238417
rect 369814 238365 369866 238417
rect 389686 238365 389738 238417
rect 332758 238291 332810 238343
rect 385270 238291 385322 238343
rect 222838 238143 222890 238195
rect 243766 238143 243818 238195
rect 253366 238143 253418 238195
rect 332086 238143 332138 238195
rect 223222 238069 223274 238121
rect 242614 238069 242666 238121
rect 251158 238069 251210 238121
rect 338710 238217 338762 238269
rect 370390 238217 370442 238269
rect 390358 238217 390410 238269
rect 332566 238143 332618 238195
rect 340438 238143 340490 238195
rect 372022 238143 372074 238195
rect 394198 238143 394250 238195
rect 251926 237995 251978 238047
rect 341494 238069 341546 238121
rect 371638 238069 371690 238121
rect 393622 238069 393674 238121
rect 42934 237921 42986 237973
rect 43318 237921 43370 237973
rect 181462 237921 181514 237973
rect 201526 237921 201578 237973
rect 223318 237921 223370 237973
rect 242134 237921 242186 237973
rect 249814 237921 249866 237973
rect 329782 237921 329834 237973
rect 332278 237921 332330 237973
rect 332662 237995 332714 238047
rect 343510 237995 343562 238047
rect 371254 237995 371306 238047
rect 392470 237995 392522 238047
rect 345238 237921 345290 237973
rect 371158 237921 371210 237973
rect 391894 237921 391946 237973
rect 42166 237847 42218 237899
rect 47542 237847 47594 237899
rect 224086 237847 224138 237899
rect 240598 237847 240650 237899
rect 249334 237847 249386 237899
rect 349174 237847 349226 237899
rect 362806 237847 362858 237899
rect 370486 237847 370538 237899
rect 370582 237847 370634 237899
rect 379030 237847 379082 237899
rect 384406 237847 384458 237899
rect 410422 237847 410474 237899
rect 43318 237773 43370 237825
rect 43510 237773 43562 237825
rect 171286 237773 171338 237825
rect 181462 237773 181514 237825
rect 201526 237773 201578 237825
rect 207094 237773 207146 237825
rect 221974 237773 222026 237825
rect 225046 237773 225098 237825
rect 238870 237773 238922 237825
rect 247126 237773 247178 237825
rect 353974 237773 354026 237825
rect 375574 237773 375626 237825
rect 401206 237773 401258 237825
rect 221014 237699 221066 237751
rect 246934 237699 246986 237751
rect 247606 237699 247658 237751
rect 351958 237699 352010 237751
rect 359830 237699 359882 237751
rect 370006 237699 370058 237751
rect 370774 237699 370826 237751
rect 381142 237699 381194 237751
rect 384502 237699 384554 237751
rect 410998 237699 411050 237751
rect 549238 237699 549290 237751
rect 649366 237699 649418 237751
rect 245782 237625 245834 237677
rect 356182 237625 356234 237677
rect 373462 237625 373514 237677
rect 397942 237625 397994 237677
rect 497494 237625 497546 237677
rect 596182 237625 596234 237677
rect 148342 237551 148394 237603
rect 161302 237551 161354 237603
rect 246166 237551 246218 237603
rect 355030 237551 355082 237603
rect 355126 237551 355178 237603
rect 370582 237551 370634 237603
rect 374230 237551 374282 237603
rect 399670 237551 399722 237603
rect 420598 237551 420650 237603
rect 607606 237551 607658 237603
rect 275350 237477 275402 237529
rect 281110 237477 281162 237529
rect 288118 237477 288170 237529
rect 292342 237477 292394 237529
rect 293782 237477 293834 237529
rect 305878 237477 305930 237529
rect 305974 237477 306026 237529
rect 317590 237477 317642 237529
rect 317686 237477 317738 237529
rect 318454 237477 318506 237529
rect 318550 237477 318602 237529
rect 319702 237477 319754 237529
rect 161302 237403 161354 237455
rect 171286 237403 171338 237455
rect 227350 237403 227402 237455
rect 233590 237403 233642 237455
rect 238774 237403 238826 237455
rect 259414 237403 259466 237455
rect 275830 237403 275882 237455
rect 286582 237403 286634 237455
rect 288022 237403 288074 237455
rect 291958 237403 292010 237455
rect 294166 237403 294218 237455
rect 302230 237403 302282 237455
rect 316822 237403 316874 237455
rect 329782 237477 329834 237529
rect 331798 237477 331850 237529
rect 337942 237477 337994 237529
rect 372598 237477 372650 237529
rect 395350 237477 395402 237529
rect 319990 237403 320042 237455
rect 331318 237403 331370 237455
rect 339766 237403 339818 237455
rect 348406 237403 348458 237455
rect 348502 237403 348554 237455
rect 221494 237329 221546 237381
rect 245878 237329 245930 237381
rect 277846 237329 277898 237381
rect 287926 237329 287978 237381
rect 289366 237329 289418 237381
rect 300982 237329 301034 237381
rect 317398 237329 317450 237381
rect 338134 237329 338186 237381
rect 217078 237255 217130 237307
rect 255190 237255 255242 237307
rect 273238 237255 273290 237307
rect 287830 237255 287882 237307
rect 290134 237255 290186 237307
rect 301462 237255 301514 237307
rect 317782 237255 317834 237307
rect 319510 237255 319562 237307
rect 319894 237255 319946 237307
rect 321814 237255 321866 237307
rect 331798 237255 331850 237307
rect 331894 237255 331946 237307
rect 339478 237255 339530 237307
rect 353590 237329 353642 237381
rect 358774 237329 358826 237381
rect 355126 237255 355178 237307
rect 372982 237403 373034 237455
rect 396214 237403 396266 237455
rect 369046 237329 369098 237381
rect 387670 237329 387722 237381
rect 378358 237255 378410 237307
rect 379990 237255 380042 237307
rect 385366 237255 385418 237307
rect 274006 237181 274058 237233
rect 290230 237181 290282 237233
rect 291670 237181 291722 237233
rect 317686 237181 317738 237233
rect 318166 237181 318218 237233
rect 330550 237181 330602 237233
rect 330646 237181 330698 237233
rect 357238 237181 357290 237233
rect 288310 237107 288362 237159
rect 290422 237107 290474 237159
rect 290614 237107 290666 237159
rect 225910 237033 225962 237085
rect 236758 237033 236810 237085
rect 278806 237033 278858 237085
rect 295030 237033 295082 237085
rect 318262 237107 318314 237159
rect 328726 237107 328778 237159
rect 328822 237107 328874 237159
rect 353494 237107 353546 237159
rect 296950 237033 297002 237085
rect 315958 237033 316010 237085
rect 325846 237033 325898 237085
rect 327478 237033 327530 237085
rect 350710 237033 350762 237085
rect 224566 236959 224618 237011
rect 239638 236959 239690 237011
rect 276790 236959 276842 237011
rect 295126 236959 295178 237011
rect 295222 236959 295274 237011
rect 303670 236959 303722 237011
rect 327094 236959 327146 237011
rect 349750 236959 349802 237011
rect 223702 236885 223754 236937
rect 241558 236885 241610 236937
rect 286390 236885 286442 236937
rect 299638 236885 299690 236937
rect 327862 236885 327914 236937
rect 351478 236885 351530 236937
rect 277270 236811 277322 236863
rect 279766 236811 279818 236863
rect 288214 236811 288266 236863
rect 289942 236811 289994 236863
rect 291766 236811 291818 236863
rect 42166 236663 42218 236715
rect 43126 236663 43178 236715
rect 226870 236663 226922 236715
rect 235030 236663 235082 236715
rect 274102 236663 274154 236715
rect 288214 236663 288266 236715
rect 258166 236589 258218 236641
rect 262102 236589 262154 236641
rect 271894 236589 271946 236641
rect 291286 236737 291338 236789
rect 305974 236737 306026 236789
rect 324022 236811 324074 236863
rect 343030 236811 343082 236863
rect 319318 236737 319370 236789
rect 324790 236737 324842 236789
rect 344758 236737 344810 236789
rect 368950 236737 369002 236789
rect 387094 236737 387146 236789
rect 290422 236663 290474 236715
rect 298774 236663 298826 236715
rect 304054 236663 304106 236715
rect 307990 236663 308042 236715
rect 325654 236663 325706 236715
rect 346966 236663 347018 236715
rect 400342 236663 400394 236715
rect 420406 236663 420458 236715
rect 440662 236663 440714 236715
rect 460726 236663 460778 236715
rect 278422 236515 278474 236567
rect 281206 236515 281258 236567
rect 287350 236515 287402 236567
rect 291862 236515 291914 236567
rect 292054 236589 292106 236641
rect 311446 236589 311498 236641
rect 313654 236589 313706 236641
rect 313846 236589 313898 236641
rect 325270 236589 325322 236641
rect 345910 236589 345962 236641
rect 294454 236515 294506 236567
rect 300214 236515 300266 236567
rect 305878 236515 305930 236567
rect 322486 236515 322538 236567
rect 339958 236515 340010 236567
rect 638038 236515 638090 236567
rect 650518 236515 650570 236567
rect 275926 236441 275978 236493
rect 294838 236441 294890 236493
rect 295030 236441 295082 236493
rect 296182 236441 296234 236493
rect 320374 236441 320426 236493
rect 335254 236441 335306 236493
rect 637366 236441 637418 236493
rect 650230 236441 650282 236493
rect 225526 236367 225578 236419
rect 237238 236367 237290 236419
rect 273430 236367 273482 236419
rect 281590 236367 281642 236419
rect 268342 236293 268394 236345
rect 288118 236367 288170 236419
rect 289942 236367 289994 236419
rect 282742 236293 282794 236345
rect 297814 236293 297866 236345
rect 144118 236219 144170 236271
rect 168406 236219 168458 236271
rect 271414 236219 271466 236271
rect 288982 236219 289034 236271
rect 289078 236219 289130 236271
rect 290710 236219 290762 236271
rect 290806 236219 290858 236271
rect 293974 236219 294026 236271
rect 294070 236219 294122 236271
rect 296470 236219 296522 236271
rect 319990 236367 320042 236419
rect 334390 236367 334442 236419
rect 637942 236367 637994 236419
rect 650326 236367 650378 236419
rect 318070 236293 318122 236345
rect 335638 236293 335690 236345
rect 639190 236293 639242 236345
rect 649846 236293 649898 236345
rect 315382 236219 315434 236271
rect 315958 236219 316010 236271
rect 328438 236219 328490 236271
rect 638806 236219 638858 236271
rect 649654 236219 649706 236271
rect 144022 236145 144074 236197
rect 171286 236145 171338 236197
rect 210358 236145 210410 236197
rect 210742 236145 210794 236197
rect 213046 236145 213098 236197
rect 217462 236145 217514 236197
rect 221782 236145 221834 236197
rect 281686 236145 281738 236197
rect 297430 236145 297482 236197
rect 547126 236145 547178 236197
rect 549238 236145 549290 236197
rect 639766 236145 639818 236197
rect 650038 236145 650090 236197
rect 265654 236071 265706 236123
rect 308278 236071 308330 236123
rect 264886 235997 264938 236049
rect 309910 235997 309962 236049
rect 312982 235997 313034 236049
rect 369622 235997 369674 236049
rect 265078 235923 265130 235975
rect 339382 235923 339434 235975
rect 381910 235923 381962 235975
rect 390934 235923 390986 235975
rect 235702 235849 235754 235901
rect 266134 235849 266186 235901
rect 267094 235849 267146 235901
rect 340342 235849 340394 235901
rect 263734 235775 263786 235827
rect 338902 235775 338954 235827
rect 258934 235701 258986 235753
rect 336694 235701 336746 235753
rect 480982 235701 481034 235753
rect 497494 235701 497546 235753
rect 261910 235627 261962 235679
rect 338134 235627 338186 235679
rect 257302 235553 257354 235605
rect 335926 235553 335978 235605
rect 260566 235479 260618 235531
rect 337174 235479 337226 235531
rect 42166 235405 42218 235457
rect 43030 235405 43082 235457
rect 236086 235405 236138 235457
rect 265462 235405 265514 235457
rect 274390 235405 274442 235457
rect 356662 235405 356714 235457
rect 246262 235331 246314 235383
rect 353590 235331 353642 235383
rect 250390 235257 250442 235309
rect 354838 235257 354890 235309
rect 241654 235183 241706 235235
rect 349942 235183 349994 235235
rect 242038 235109 242090 235161
rect 352150 235109 352202 235161
rect 241846 235035 241898 235087
rect 350422 235035 350474 235087
rect 246454 234961 246506 235013
rect 354358 234961 354410 235013
rect 243286 234887 243338 234939
rect 352630 234887 352682 234939
rect 42166 234813 42218 234865
rect 42454 234813 42506 234865
rect 244150 234813 244202 234865
rect 351382 234813 351434 234865
rect 230614 234739 230666 234791
rect 346966 234739 347018 234791
rect 227830 234665 227882 234717
rect 345526 234665 345578 234717
rect 282454 234591 282506 234643
rect 322774 234591 322826 234643
rect 266998 234517 267050 234569
rect 305686 234517 305738 234569
rect 282838 234443 282890 234495
rect 321910 234443 321962 234495
rect 267478 234369 267530 234421
rect 304246 234369 304298 234421
rect 271606 234295 271658 234347
rect 309430 234295 309482 234347
rect 284662 234221 284714 234273
rect 317494 234221 317546 234273
rect 284278 234147 284330 234199
rect 319126 234147 319178 234199
rect 268822 234073 268874 234125
rect 301942 234073 301994 234125
rect 269590 233999 269642 234051
rect 300310 233999 300362 234051
rect 285142 233925 285194 233977
rect 316150 233925 316202 233977
rect 274870 233851 274922 233903
rect 288598 233851 288650 233903
rect 292534 233851 292586 233903
rect 320566 233851 320618 233903
rect 293110 233777 293162 233829
rect 321430 233777 321482 233829
rect 209782 233703 209834 233755
rect 212182 233703 212234 233755
rect 238054 233703 238106 233755
rect 239062 233703 239114 233755
rect 270070 233703 270122 233755
rect 298582 233703 298634 233755
rect 305590 233703 305642 233755
rect 308710 233703 308762 233755
rect 208150 233629 208202 233681
rect 213526 233629 213578 233681
rect 270646 233629 270698 233681
rect 298486 233629 298538 233681
rect 209974 233555 210026 233607
rect 213142 233555 213194 233607
rect 269110 233555 269162 233607
rect 297046 233555 297098 233607
rect 298198 233555 298250 233607
rect 210262 233481 210314 233533
rect 210934 233481 210986 233533
rect 211307 233474 211359 233526
rect 213910 233481 213962 233533
rect 316918 233629 316970 233681
rect 144022 233259 144074 233311
rect 165526 233259 165578 233311
rect 206518 233185 206570 233237
rect 206614 233185 206666 233237
rect 645718 233185 645770 233237
rect 649750 233185 649802 233237
rect 645814 233111 645866 233163
rect 649942 233111 649994 233163
rect 645142 233037 645194 233089
rect 650422 233037 650474 233089
rect 645334 232963 645386 233015
rect 650134 232963 650186 233015
rect 645238 232889 645290 232941
rect 650614 232889 650666 232941
rect 205078 232593 205130 232645
rect 205078 232445 205130 232497
rect 42070 231039 42122 231091
rect 42934 231039 42986 231091
rect 206902 230669 206954 230721
rect 207094 230669 207146 230721
rect 144022 230521 144074 230573
rect 151126 230521 151178 230573
rect 206326 230521 206378 230573
rect 206902 230521 206954 230573
rect 144118 230447 144170 230499
rect 202966 230447 203018 230499
rect 144022 227709 144074 227761
rect 188566 227709 188618 227761
rect 144118 227635 144170 227687
rect 194326 227635 194378 227687
rect 144214 227561 144266 227613
rect 197206 227561 197258 227613
rect 204886 227117 204938 227169
rect 205654 227117 205706 227169
rect 146806 225637 146858 225689
rect 156886 225637 156938 225689
rect 666838 225045 666890 225097
rect 674710 225045 674762 225097
rect 146806 224675 146858 224727
rect 200086 224675 200138 224727
rect 141046 224601 141098 224653
rect 199702 224601 199754 224653
rect 146422 224527 146474 224579
rect 201718 224527 201770 224579
rect 149686 224453 149738 224505
rect 201622 224453 201674 224505
rect 152566 224379 152618 224431
rect 201814 224379 201866 224431
rect 669622 224305 669674 224357
rect 674422 224305 674474 224357
rect 669526 224009 669578 224061
rect 674710 224009 674762 224061
rect 205750 223121 205802 223173
rect 206134 223121 206186 223173
rect 146710 221937 146762 221989
rect 177046 221937 177098 221989
rect 146806 221863 146858 221915
rect 179926 221863 179978 221915
rect 144406 221789 144458 221841
rect 182806 221789 182858 221841
rect 155446 221715 155498 221767
rect 198838 221715 198890 221767
rect 161206 221641 161258 221693
rect 210166 221641 210218 221693
rect 164086 221567 164138 221619
rect 201718 221567 201770 221619
rect 166966 221493 167018 221545
rect 201622 221493 201674 221545
rect 169846 221419 169898 221471
rect 196054 221419 196106 221471
rect 144406 218903 144458 218955
rect 174262 218903 174314 218955
rect 175606 218829 175658 218881
rect 200662 218829 200714 218881
rect 178486 218755 178538 218807
rect 201718 218755 201770 218807
rect 181366 218681 181418 218733
rect 210166 218681 210218 218733
rect 184246 218607 184298 218659
rect 201622 218607 201674 218659
rect 42454 216461 42506 216513
rect 45142 216461 45194 216513
rect 146806 216313 146858 216365
rect 154006 216313 154058 216365
rect 645430 216017 645482 216069
rect 645814 216017 645866 216069
rect 187126 215943 187178 215995
rect 210166 215943 210218 215995
rect 674134 215943 674186 215995
rect 674518 215943 674570 215995
rect 192886 215869 192938 215921
rect 201718 215869 201770 215921
rect 42838 215721 42890 215773
rect 45046 215721 45098 215773
rect 42838 215203 42890 215255
rect 44662 215203 44714 215255
rect 206038 213501 206090 213553
rect 206326 213501 206378 213553
rect 146806 213205 146858 213257
rect 168502 213205 168554 213257
rect 144214 213131 144266 213183
rect 171382 213131 171434 213183
rect 146806 210245 146858 210297
rect 148246 210245 148298 210297
rect 647926 210245 647978 210297
rect 677014 210245 677066 210297
rect 146710 207433 146762 207485
rect 165622 207433 165674 207485
rect 146806 207359 146858 207411
rect 203062 207359 203114 207411
rect 645430 207285 645482 207337
rect 645814 207285 645866 207337
rect 42454 204399 42506 204451
rect 50326 204399 50378 204451
rect 674998 204399 675050 204451
rect 675382 204399 675434 204451
rect 146806 201661 146858 201713
rect 159766 201661 159818 201713
rect 144982 201587 145034 201639
rect 162646 201587 162698 201639
rect 674134 201291 674186 201343
rect 675382 201291 675434 201343
rect 40054 200107 40106 200159
rect 43126 200107 43178 200159
rect 40150 198997 40202 199049
rect 42358 198997 42410 199049
rect 39958 198775 40010 198827
rect 43318 198775 43370 198827
rect 40246 198701 40298 198753
rect 41014 198701 41066 198753
rect 146806 198701 146858 198753
rect 191446 198701 191498 198753
rect 674710 197591 674762 197643
rect 675382 197591 675434 197643
rect 42070 197369 42122 197421
rect 42070 197147 42122 197199
rect 674518 196999 674570 197051
rect 675478 196999 675530 197051
rect 42358 196851 42410 196903
rect 43222 196851 43274 196903
rect 674614 196555 674666 196607
rect 675382 196555 675434 196607
rect 146806 195815 146858 195867
rect 185686 195815 185738 195867
rect 42454 195593 42506 195645
rect 42166 195297 42218 195349
rect 42934 194779 42986 194831
rect 43222 194779 43274 194831
rect 42838 194705 42890 194757
rect 43318 194705 43370 194757
rect 42070 194483 42122 194535
rect 44758 194483 44810 194535
rect 42070 193447 42122 193499
rect 43126 193447 43178 193499
rect 206902 192929 206954 192981
rect 206998 192929 207050 192981
rect 42166 192189 42218 192241
rect 43030 192189 43082 192241
rect 42070 191449 42122 191501
rect 42934 191449 42986 191501
rect 146710 190191 146762 190243
rect 151222 190191 151274 190243
rect 146806 190117 146858 190169
rect 148438 190117 148490 190169
rect 42166 187675 42218 187727
rect 42838 187675 42890 187727
rect 146806 187231 146858 187283
rect 197302 187231 197354 187283
rect 146806 184345 146858 184397
rect 194422 184345 194474 184397
rect 144502 181533 144554 181585
rect 148534 181533 148586 181585
rect 144022 181459 144074 181511
rect 188662 181459 188714 181511
rect 661078 179313 661130 179365
rect 674422 179313 674474 179365
rect 666646 178795 666698 178847
rect 674422 178795 674474 178847
rect 145270 178647 145322 178699
rect 148630 178647 148682 178699
rect 655222 178647 655274 178699
rect 674614 178647 674666 178699
rect 146806 178573 146858 178625
rect 191542 178573 191594 178625
rect 146806 175835 146858 175887
rect 148726 175835 148778 175887
rect 144118 175687 144170 175739
rect 185782 175687 185834 175739
rect 144790 172801 144842 172853
rect 162742 172801 162794 172853
rect 146806 169915 146858 169967
rect 159862 169915 159914 169967
rect 206710 169841 206762 169893
rect 206998 169841 207050 169893
rect 646870 167399 646922 167451
rect 674710 167399 674762 167451
rect 646294 167177 646346 167229
rect 674710 167177 674762 167229
rect 146806 167103 146858 167155
rect 156982 167103 157034 167155
rect 647926 167103 647978 167155
rect 674614 167103 674666 167155
rect 144790 167029 144842 167081
rect 148822 167029 148874 167081
rect 144790 164143 144842 164195
rect 148918 164143 148970 164195
rect 144982 162737 145034 162789
rect 146710 162737 146762 162789
rect 144886 161257 144938 161309
rect 149014 161257 149066 161309
rect 675478 160961 675530 161013
rect 675478 160739 675530 160791
rect 675094 159555 675146 159607
rect 675286 159555 675338 159607
rect 144886 158445 144938 158497
rect 149110 158445 149162 158497
rect 144886 155559 144938 155611
rect 200182 155559 200234 155611
rect 674038 153339 674090 153391
rect 675478 153339 675530 153391
rect 144886 152747 144938 152799
rect 180022 152747 180074 152799
rect 674230 152747 674282 152799
rect 675382 152747 675434 152799
rect 144790 152673 144842 152725
rect 182902 152673 182954 152725
rect 673942 152007 673994 152059
rect 675478 152007 675530 152059
rect 674134 151489 674186 151541
rect 675382 151489 675434 151541
rect 144886 149787 144938 149839
rect 177142 149787 177194 149839
rect 144886 146901 144938 146953
rect 174358 146901 174410 146953
rect 144502 146087 144554 146139
rect 144886 146087 144938 146139
rect 146134 144607 146186 144659
rect 146326 144607 146378 144659
rect 144310 144459 144362 144511
rect 146134 144459 146186 144511
rect 144502 144311 144554 144363
rect 154102 144311 154154 144363
rect 144310 144015 144362 144067
rect 208726 144015 208778 144067
rect 144310 141647 144362 141699
rect 171574 141647 171626 141699
rect 144310 141203 144362 141255
rect 149206 141203 149258 141255
rect 645430 141203 645482 141255
rect 645814 141203 645866 141255
rect 144502 141129 144554 141181
rect 208822 141129 208874 141181
rect 645142 141055 645194 141107
rect 645238 141055 645290 141107
rect 645430 141055 645482 141107
rect 645814 141055 645866 141107
rect 144502 140907 144554 140959
rect 146326 140907 146378 140959
rect 645238 140759 645290 140811
rect 645142 140537 645194 140589
rect 144310 138243 144362 138295
rect 168598 138243 168650 138295
rect 144886 137059 144938 137111
rect 144694 136911 144746 136963
rect 144886 136911 144938 136963
rect 144790 136689 144842 136741
rect 146902 135949 146954 136001
rect 149302 135949 149354 136001
rect 144310 135431 144362 135483
rect 208918 135357 208970 135409
rect 144502 134987 144554 135039
rect 146902 134987 146954 135039
rect 663766 133581 663818 133633
rect 674422 133581 674474 133633
rect 144310 132915 144362 132967
rect 165718 132915 165770 132967
rect 655318 132767 655370 132819
rect 676918 132767 676970 132819
rect 655126 132619 655178 132671
rect 676822 132619 676874 132671
rect 144310 132545 144362 132597
rect 209014 132545 209066 132597
rect 144502 132471 144554 132523
rect 209110 132471 209162 132523
rect 647638 132471 647690 132523
rect 674422 132471 674474 132523
rect 144502 129659 144554 129711
rect 151414 129659 151466 129711
rect 144310 129585 144362 129637
rect 208630 129585 208682 129637
rect 144502 129511 144554 129563
rect 144886 129511 144938 129563
rect 144886 129363 144938 129415
rect 146134 129363 146186 129415
rect 146134 128475 146186 128527
rect 146518 128475 146570 128527
rect 144022 126995 144074 127047
rect 144118 126995 144170 127047
rect 144214 126995 144266 127047
rect 144310 126921 144362 126973
rect 144022 126773 144074 126825
rect 144118 126773 144170 126825
rect 144214 126773 144266 126825
rect 146326 126773 146378 126825
rect 146998 126847 147050 126899
rect 149398 126847 149450 126899
rect 203158 126773 203210 126825
rect 143926 126699 143978 126751
rect 146518 126699 146570 126751
rect 208534 126699 208586 126751
rect 145078 126625 145130 126677
rect 146326 126625 146378 126677
rect 645526 126625 645578 126677
rect 645814 126625 645866 126677
rect 143926 126477 143978 126529
rect 145078 126477 145130 126529
rect 144598 125367 144650 125419
rect 146518 125367 146570 125419
rect 39862 125293 39914 125345
rect 42934 125293 42986 125345
rect 144406 125219 144458 125271
rect 144598 125219 144650 125271
rect 146326 124997 146378 125049
rect 146134 124849 146186 124901
rect 146326 124849 146378 124901
rect 146134 124701 146186 124753
rect 144310 123961 144362 124013
rect 197398 123961 197450 124013
rect 144406 123887 144458 123939
rect 200278 123887 200330 123939
rect 645814 121223 645866 121275
rect 676822 121223 676874 121275
rect 645910 121149 645962 121201
rect 674710 121149 674762 121201
rect 144406 121075 144458 121127
rect 149494 121075 149546 121127
rect 646006 121075 646058 121127
rect 676918 121075 676970 121127
rect 144310 121001 144362 121053
rect 149590 121001 149642 121053
rect 144406 120927 144458 120979
rect 144598 120927 144650 120979
rect 207094 120927 207146 120979
rect 207190 120927 207242 120979
rect 144310 118411 144362 118463
rect 144406 118263 144458 118315
rect 171478 118263 171530 118315
rect 144310 118189 144362 118241
rect 188758 118189 188810 118241
rect 144598 118115 144650 118167
rect 194518 118115 194570 118167
rect 144598 117967 144650 118019
rect 144310 116191 144362 116243
rect 149686 116191 149738 116243
rect 144310 115525 144362 115577
rect 148150 115525 148202 115577
rect 144310 115377 144362 115429
rect 146134 115377 146186 115429
rect 146134 115007 146186 115059
rect 146902 115007 146954 115059
rect 674518 114119 674570 114171
rect 675382 114119 675434 114171
rect 674326 113601 674378 113653
rect 675094 113601 675146 113653
rect 144310 112639 144362 112691
rect 147958 112639 148010 112691
rect 144310 112417 144362 112469
rect 148054 112417 148106 112469
rect 144406 112343 144458 112395
rect 191638 112343 191690 112395
rect 674230 111825 674282 111877
rect 675094 111825 675146 111877
rect 674710 111307 674762 111359
rect 675382 111307 675434 111359
rect 674806 111233 674858 111285
rect 675094 111233 675146 111285
rect 144406 109531 144458 109583
rect 147862 109531 147914 109583
rect 144310 109457 144362 109509
rect 185878 109457 185930 109509
rect 144406 109383 144458 109435
rect 144598 109383 144650 109435
rect 674902 107533 674954 107585
rect 675382 107533 675434 107585
rect 143830 106941 143882 106993
rect 144406 106941 144458 106993
rect 144310 106867 144362 106919
rect 162838 106867 162890 106919
rect 673942 106867 673994 106919
rect 675478 106867 675530 106919
rect 143926 106793 143978 106845
rect 146518 106793 146570 106845
rect 144310 106719 144362 106771
rect 145078 106719 145130 106771
rect 144598 106571 144650 106623
rect 147766 106571 147818 106623
rect 645526 106497 645578 106549
rect 645910 106497 645962 106549
rect 668182 106497 668234 106549
rect 675094 106497 675146 106549
rect 143926 106423 143978 106475
rect 144598 106423 144650 106475
rect 146518 106423 146570 106475
rect 159958 106423 160010 106475
rect 674422 106349 674474 106401
rect 675382 106349 675434 106401
rect 146326 104795 146378 104847
rect 146902 104795 146954 104847
rect 645430 104499 645482 104551
rect 665206 104499 665258 104551
rect 659542 104425 659594 104477
rect 665302 104425 665354 104477
rect 146518 104351 146570 104403
rect 160054 104351 160106 104403
rect 146326 103685 146378 103737
rect 208438 103685 208490 103737
rect 146134 103611 146186 103663
rect 204598 103611 204650 103663
rect 145078 103537 145130 103589
rect 204694 103537 204746 103589
rect 146902 103463 146954 103515
rect 204502 103463 204554 103515
rect 143830 103389 143882 103441
rect 145078 103389 145130 103441
rect 146518 101539 146570 101591
rect 157078 101539 157130 101591
rect 146326 100799 146378 100851
rect 151318 100799 151370 100851
rect 145078 100725 145130 100777
rect 194710 100725 194762 100777
rect 144406 100651 144458 100703
rect 201718 100651 201770 100703
rect 144598 100577 144650 100629
rect 204598 100577 204650 100629
rect 151126 100503 151178 100555
rect 198358 100503 198410 100555
rect 159766 100429 159818 100481
rect 210166 100429 210218 100481
rect 146518 98061 146570 98113
rect 180118 98061 180170 98113
rect 146326 97987 146378 98039
rect 182998 97987 183050 98039
rect 146134 97913 146186 97965
rect 208342 97913 208394 97965
rect 154006 97839 154058 97891
rect 200758 97839 200810 97891
rect 156886 97765 156938 97817
rect 200566 97765 200618 97817
rect 171382 97691 171434 97743
rect 201718 97691 201770 97743
rect 174262 97617 174314 97669
rect 210166 97617 210218 97669
rect 182806 97543 182858 97595
rect 201046 97543 201098 97595
rect 146518 95101 146570 95153
rect 174454 95101 174506 95153
rect 146326 95027 146378 95079
rect 177238 95027 177290 95079
rect 144214 94879 144266 94931
rect 201622 94879 201674 94931
rect 151222 94805 151274 94857
rect 195478 94805 195530 94857
rect 165622 94731 165674 94783
rect 201718 94731 201770 94783
rect 168502 94657 168554 94709
rect 210166 94657 210218 94709
rect 144022 94583 144074 94635
rect 194806 94583 194858 94635
rect 651286 93695 651338 93747
rect 659542 93695 659594 93747
rect 646390 92659 646442 92711
rect 659830 92659 659882 92711
rect 647446 92585 647498 92637
rect 661750 92585 661802 92637
rect 646198 92511 646250 92563
rect 660694 92511 660746 92563
rect 647830 92363 647882 92415
rect 663094 92363 663146 92415
rect 647254 92289 647306 92341
rect 661174 92289 661226 92341
rect 146326 92215 146378 92267
rect 154006 92215 154058 92267
rect 647734 92215 647786 92267
rect 662518 92215 662570 92267
rect 146518 92141 146570 92193
rect 171382 92141 171434 92193
rect 646678 92141 646730 92193
rect 658870 92141 658922 92193
rect 144118 92067 144170 92119
rect 210166 92067 210218 92119
rect 188662 91771 188714 91823
rect 201718 91771 201770 91823
rect 146134 89403 146186 89455
rect 151126 89403 151178 89455
rect 146518 89329 146570 89381
rect 165622 89329 165674 89381
rect 146326 89255 146378 89307
rect 168502 89255 168554 89307
rect 156982 89181 157034 89233
rect 197878 89181 197930 89233
rect 159862 89107 159914 89159
rect 201814 89107 201866 89159
rect 162742 89033 162794 89085
rect 201622 89033 201674 89085
rect 185782 88959 185834 89011
rect 201334 88959 201386 89011
rect 191542 88885 191594 88937
rect 201718 88885 201770 88937
rect 650614 87331 650666 87383
rect 659350 87331 659402 87383
rect 658006 87257 658058 87309
rect 657046 87109 657098 87161
rect 645430 87035 645482 87087
rect 663286 87035 663338 87087
rect 645814 86961 645866 87013
rect 650998 86961 651050 87013
rect 645430 86887 645482 86939
rect 645910 86887 645962 86939
rect 645814 86443 645866 86495
rect 651094 86443 651146 86495
rect 154102 86369 154154 86421
rect 196054 86369 196106 86421
rect 645430 86369 645482 86421
rect 646102 86369 646154 86421
rect 174358 86295 174410 86347
rect 201814 86295 201866 86347
rect 177142 86221 177194 86273
rect 198742 86221 198794 86273
rect 180022 86147 180074 86199
rect 201718 86147 201770 86199
rect 182902 86073 182954 86125
rect 201622 86073 201674 86125
rect 645430 85185 645482 85237
rect 650902 85185 650954 85237
rect 146518 84963 146570 85015
rect 197782 84963 197834 85015
rect 151414 83483 151466 83535
rect 201526 83483 201578 83535
rect 165718 83409 165770 83461
rect 201814 83409 201866 83461
rect 645430 83409 645482 83461
rect 657046 83409 657098 83461
rect 168598 83335 168650 83387
rect 201622 83335 201674 83387
rect 171574 83261 171626 83313
rect 201718 83261 201770 83313
rect 146518 82077 146570 82129
rect 201718 82077 201770 82129
rect 645430 81855 645482 81907
rect 663286 81855 663338 81907
rect 645814 81781 645866 81833
rect 663382 81781 663434 81833
rect 647542 81633 647594 81685
rect 661078 81633 661130 81685
rect 645430 81263 645482 81315
rect 657526 81263 657578 81315
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 188758 80301 188810 80353
rect 210166 80301 210218 80353
rect 645430 80153 645482 80205
rect 656950 80153 657002 80205
rect 645910 79043 645962 79095
rect 651190 79043 651242 79095
rect 645430 78895 645482 78947
rect 658870 78895 658922 78947
rect 645814 78377 645866 78429
rect 662518 78377 662570 78429
rect 646006 78007 646058 78059
rect 660694 78007 660746 78059
rect 146326 77859 146378 77911
rect 190006 77859 190058 77911
rect 146518 77785 146570 77837
rect 208246 77785 208298 77837
rect 157078 77711 157130 77763
rect 196918 77711 196970 77763
rect 647638 77711 647690 77763
rect 659446 77711 659498 77763
rect 160054 77637 160106 77689
rect 201622 77637 201674 77689
rect 645430 77637 645482 77689
rect 650998 77637 651050 77689
rect 162838 77563 162890 77615
rect 200278 77563 200330 77615
rect 185878 77489 185930 77541
rect 210166 77489 210218 77541
rect 191638 77415 191690 77467
rect 201718 77415 201770 77467
rect 645430 77267 645482 77319
rect 662902 77267 662954 77319
rect 190006 77193 190058 77245
rect 201718 77193 201770 77245
rect 645910 76971 645962 77023
rect 661750 76971 661802 77023
rect 645430 76897 645482 76949
rect 658294 76897 658346 76949
rect 645814 76675 645866 76727
rect 650902 76675 650954 76727
rect 640726 76231 640778 76283
rect 651286 76231 651338 76283
rect 645430 75491 645482 75543
rect 656854 75491 656906 75543
rect 146326 75269 146378 75321
rect 146134 75195 146186 75247
rect 146518 75195 146570 75247
rect 144022 75121 144074 75173
rect 144214 75047 144266 75099
rect 146134 75047 146186 75099
rect 144118 74973 144170 75025
rect 146326 74973 146378 75025
rect 160054 75047 160106 75099
rect 156406 74973 156458 75025
rect 144406 74899 144458 74951
rect 161494 74899 161546 74951
rect 154006 74825 154058 74877
rect 201526 74825 201578 74877
rect 174454 74751 174506 74803
rect 201814 74751 201866 74803
rect 177238 74677 177290 74729
rect 210166 74677 210218 74729
rect 180118 74603 180170 74655
rect 201622 74603 201674 74655
rect 182998 74529 183050 74581
rect 201718 74529 201770 74581
rect 144406 74455 144458 74507
rect 148342 74455 148394 74507
rect 144214 74011 144266 74063
rect 146710 74011 146762 74063
rect 645430 72975 645482 73027
rect 663382 72975 663434 73027
rect 645814 72309 645866 72361
rect 660118 72309 660170 72361
rect 645430 72087 645482 72139
rect 663190 72087 663242 72139
rect 146710 72013 146762 72065
rect 153910 72013 153962 72065
rect 151126 71939 151178 71991
rect 200374 71939 200426 71991
rect 209782 71939 209834 71991
rect 210166 71939 210218 71991
rect 161494 71865 161546 71917
rect 201814 71865 201866 71917
rect 165622 71791 165674 71843
rect 201622 71791 201674 71843
rect 209782 71791 209834 71843
rect 209974 71791 210026 71843
rect 168502 71717 168554 71769
rect 201718 71717 201770 71769
rect 171382 71643 171434 71695
rect 209974 71643 210026 71695
rect 146710 70903 146762 70955
rect 149782 70903 149834 70955
rect 144118 69497 144170 69549
rect 145654 69497 145706 69549
rect 145462 69349 145514 69401
rect 145654 69349 145706 69401
rect 145462 69201 145514 69253
rect 145846 69201 145898 69253
rect 144022 69127 144074 69179
rect 201814 69053 201866 69105
rect 149782 68979 149834 69031
rect 201622 68979 201674 69031
rect 153910 68905 153962 68957
rect 201718 68905 201770 68957
rect 156406 68831 156458 68883
rect 196246 68831 196298 68883
rect 160054 68757 160106 68809
rect 195478 68757 195530 68809
rect 146710 67351 146762 67403
rect 152662 67351 152714 67403
rect 145846 66389 145898 66441
rect 158326 66389 158378 66441
rect 146806 66241 146858 66293
rect 645526 66241 645578 66293
rect 646102 66241 646154 66293
rect 201718 66167 201770 66219
rect 152662 66093 152714 66145
rect 198550 66093 198602 66145
rect 158326 66019 158378 66071
rect 193654 66019 193706 66071
rect 145654 64835 145706 64887
rect 146710 64835 146762 64887
rect 201718 64835 201770 64887
rect 144502 64613 144554 64665
rect 144694 64613 144746 64665
rect 144790 64613 144842 64665
rect 145558 64613 145610 64665
rect 144694 64465 144746 64517
rect 146806 64761 146858 64813
rect 201814 64761 201866 64813
rect 144214 64391 144266 64443
rect 145942 64391 145994 64443
rect 146902 63355 146954 63407
rect 195478 63355 195530 63407
rect 209398 62763 209450 62815
rect 210262 62763 210314 62815
rect 209494 62615 209546 62667
rect 210262 62615 210314 62667
rect 146806 62467 146858 62519
rect 149782 62467 149834 62519
rect 160534 60765 160586 60817
rect 201718 60765 201770 60817
rect 156310 60691 156362 60743
rect 201622 60691 201674 60743
rect 152662 60617 152714 60669
rect 195478 60617 195530 60669
rect 151126 60543 151178 60595
rect 201526 60543 201578 60595
rect 148342 60469 148394 60521
rect 201814 60469 201866 60521
rect 146902 60395 146954 60447
rect 209974 60395 210026 60447
rect 149782 60321 149834 60373
rect 198358 60321 198410 60373
rect 146806 59581 146858 59633
rect 160534 59581 160586 59633
rect 146806 58989 146858 59041
rect 201718 58989 201770 59041
rect 146806 57065 146858 57117
rect 156310 57065 156362 57117
rect 144118 56917 144170 56969
rect 146806 56917 146858 56969
rect 144022 56473 144074 56525
rect 152662 56473 152714 56525
rect 144790 54623 144842 54675
rect 151126 54623 151178 54675
rect 144214 54327 144266 54379
rect 144598 54327 144650 54379
rect 210262 54327 210314 54379
rect 209302 54253 209354 54305
rect 217462 54253 217514 54305
rect 219382 54253 219434 54305
rect 209782 54179 209834 54231
rect 219190 54179 219242 54231
rect 144502 54105 144554 54157
rect 148342 54105 148394 54157
rect 209686 54105 209738 54157
rect 213766 54105 213818 54157
rect 205654 53957 205706 54009
rect 218182 53957 218234 54009
rect 208342 53883 208394 53935
rect 214966 53883 215018 53935
rect 210358 53809 210410 53861
rect 221398 53809 221450 53861
rect 231766 53809 231818 53861
rect 261910 53883 261962 53935
rect 262006 53809 262058 53861
rect 209974 53735 210026 53787
rect 219190 53735 219242 53787
rect 282166 53883 282218 53935
rect 210166 53661 210218 53713
rect 207958 53587 208010 53639
rect 231766 53587 231818 53639
rect 209398 53513 209450 53565
rect 215254 53513 215306 53565
rect 216358 53513 216410 53565
rect 209494 53439 209546 53491
rect 218902 53439 218954 53491
rect 210646 53365 210698 53417
rect 351286 53513 351338 53565
rect 219190 53439 219242 53491
rect 384406 53439 384458 53491
rect 219382 53365 219434 53417
rect 467446 53365 467498 53417
rect 469366 53365 469418 53417
rect 501046 53365 501098 53417
rect 210262 53291 210314 53343
rect 219670 53291 219722 53343
rect 221398 53291 221450 53343
rect 501142 53291 501194 53343
rect 204886 53217 204938 53269
rect 215638 53217 215690 53269
rect 210454 53143 210506 53195
rect 213430 53143 213482 53195
rect 251926 53143 251978 53195
rect 208054 53069 208106 53121
rect 220342 53069 220394 53121
rect 315670 53217 315722 53269
rect 368566 53217 368618 53269
rect 388822 53217 388874 53269
rect 408982 53217 409034 53269
rect 368662 53143 368714 53195
rect 388726 53143 388778 53195
rect 216982 52995 217034 53047
rect 315670 52995 315722 53047
rect 409078 52995 409130 53047
rect 469366 53143 469418 53195
rect 501046 53143 501098 53195
rect 509686 53143 509738 53195
rect 251926 52921 251978 52973
rect 159958 52847 160010 52899
rect 217270 52847 217322 52899
rect 211606 52773 211658 52825
rect 219958 52773 220010 52825
rect 151318 52699 151370 52751
rect 216502 52699 216554 52751
rect 212278 52477 212330 52529
rect 213430 52477 213482 52529
rect 211222 52403 211274 52455
rect 213814 52403 213866 52455
rect 203062 52329 203114 52381
rect 226582 52329 226634 52381
rect 146518 52255 146570 52307
rect 225718 52255 225770 52307
rect 171478 52181 171530 52233
rect 219862 52181 219914 52233
rect 146326 52107 146378 52159
rect 226966 52107 227018 52159
rect 144214 52033 144266 52085
rect 220918 52033 220970 52085
rect 145078 51959 145130 52011
rect 203062 51959 203114 52011
rect 146134 51885 146186 51937
rect 227542 51885 227594 51937
rect 213430 51811 213482 51863
rect 213814 51737 213866 51789
rect 219958 51811 220010 51863
rect 645526 51811 645578 51863
rect 209878 51663 209930 51715
rect 214102 51663 214154 51715
rect 645718 51737 645770 51789
rect 639670 51663 639722 51715
rect 209590 51589 209642 51641
rect 214486 51589 214538 51641
rect 144982 51441 145034 51493
rect 233590 51441 233642 51493
rect 145174 51367 145226 51419
rect 234550 51367 234602 51419
rect 145366 51293 145418 51345
rect 235798 51293 235850 51345
rect 145654 51219 145706 51271
rect 235318 51219 235370 51271
rect 146038 51145 146090 51197
rect 232342 51145 232394 51197
rect 146230 51071 146282 51123
rect 231382 51071 231434 51123
rect 146422 50997 146474 51049
rect 231958 50997 232010 51049
rect 146614 50923 146666 50975
rect 230902 50923 230954 50975
rect 144886 50849 144938 50901
rect 230134 50849 230186 50901
rect 145270 50775 145322 50827
rect 228790 50775 228842 50827
rect 146710 50701 146762 50753
rect 228694 50701 228746 50753
rect 145942 50627 145994 50679
rect 229174 50627 229226 50679
rect 144406 50553 144458 50605
rect 208054 50553 208106 50605
rect 208246 50553 208298 50605
rect 216118 50553 216170 50605
rect 144694 50479 144746 50531
rect 208342 50479 208394 50531
rect 208438 50479 208490 50531
rect 216886 50479 216938 50531
rect 145558 50405 145610 50457
rect 211510 50405 211562 50457
rect 144310 50331 144362 50383
rect 209110 50331 209162 50383
rect 209398 50331 209450 50383
rect 221494 50331 221546 50383
rect 144790 50257 144842 50309
rect 235414 50257 235466 50309
rect 145750 50183 145802 50235
rect 234934 50183 234986 50235
rect 145846 50109 145898 50161
rect 232726 50109 232778 50161
rect 209110 50035 209162 50087
rect 223894 50035 223946 50087
rect 208054 49961 208106 50013
rect 225334 49961 225386 50013
rect 146806 49887 146858 49939
rect 241174 49887 241226 49939
rect 145366 49813 145418 49865
rect 244150 49813 244202 49865
rect 208342 49739 208394 49791
rect 226102 49739 226154 49791
rect 145462 49665 145514 49717
rect 237142 49665 237194 49717
rect 211510 49591 211562 49643
rect 226486 49591 226538 49643
rect 208918 48925 208970 48977
rect 220246 48999 220298 49051
rect 509686 48999 509738 49051
rect 525910 48999 525962 49051
rect 218614 48925 218666 48977
rect 645622 48925 645674 48977
rect 210070 48851 210122 48903
rect 220726 48851 220778 48903
rect 501142 48851 501194 48903
rect 507094 48851 507146 48903
rect 208150 48777 208202 48829
rect 220054 48777 220106 48829
rect 220246 48777 220298 48829
rect 223510 48777 223562 48829
rect 208534 48703 208586 48755
rect 221686 48703 221738 48755
rect 222262 48703 222314 48755
rect 645238 48703 645290 48755
rect 209014 48629 209066 48681
rect 222454 48629 222506 48681
rect 222934 48629 222986 48681
rect 645142 48629 645194 48681
rect 188566 48555 188618 48607
rect 239350 48555 239402 48607
rect 185686 48481 185738 48533
rect 240214 48481 240266 48533
rect 194326 48407 194378 48459
rect 239734 48407 239786 48459
rect 197206 48333 197258 48385
rect 239830 48333 239882 48385
rect 162646 48259 162698 48311
rect 241558 48259 241610 48311
rect 149302 48185 149354 48237
rect 209206 48185 209258 48237
rect 209302 48185 209354 48237
rect 222742 48185 222794 48237
rect 224086 48185 224138 48237
rect 645334 48185 645386 48237
rect 149206 48111 149258 48163
rect 208534 48111 208586 48163
rect 208630 48111 208682 48163
rect 222070 48111 222122 48163
rect 148150 48037 148202 48089
rect 219094 48037 219146 48089
rect 149398 47963 149450 48015
rect 221302 47963 221354 48015
rect 149494 47889 149546 47941
rect 220534 47889 220586 47941
rect 149686 47815 149738 47867
rect 219478 47815 219530 47867
rect 149590 47741 149642 47793
rect 220150 47741 220202 47793
rect 147862 47667 147914 47719
rect 218038 47667 218090 47719
rect 147766 47593 147818 47645
rect 217654 47593 217706 47645
rect 148054 47519 148106 47571
rect 218326 47519 218378 47571
rect 623446 47519 623498 47571
rect 640726 47519 640778 47571
rect 147958 47445 148010 47497
rect 218710 47445 218762 47497
rect 177046 47371 177098 47423
rect 238006 47371 238058 47423
rect 179926 47297 179978 47349
rect 238582 47297 238634 47349
rect 200086 47223 200138 47275
rect 238966 47223 239018 47275
rect 148534 47149 148586 47201
rect 230998 47149 231050 47201
rect 148246 47075 148298 47127
rect 236374 47075 236426 47127
rect 149110 47001 149162 47053
rect 233302 47001 233354 47053
rect 149014 46927 149066 46979
rect 234166 46927 234218 46979
rect 148726 46853 148778 46905
rect 229750 46853 229802 46905
rect 148630 46779 148682 46831
rect 230518 46779 230570 46831
rect 148822 46705 148874 46757
rect 228310 46705 228362 46757
rect 209206 46631 209258 46683
rect 223126 46631 223178 46683
rect 148918 46557 148970 46609
rect 227926 46557 227978 46609
rect 148438 46483 148490 46535
rect 233110 46483 233162 46535
rect 208822 46409 208874 46461
rect 224662 46409 224714 46461
rect 208726 46335 208778 46387
rect 224950 46335 225002 46387
rect 208534 46261 208586 46313
rect 224278 46261 224330 46313
rect 191446 46187 191498 46239
rect 240790 46187 240842 46239
rect 206998 46039 207050 46091
rect 465814 46039 465866 46091
rect 384406 45373 384458 45425
rect 388822 45373 388874 45425
rect 212086 45003 212138 45055
rect 297238 45003 297290 45055
rect 211414 44929 211466 44981
rect 361750 44929 361802 44981
rect 213910 44855 213962 44907
rect 455734 44855 455786 44907
rect 211702 44781 211754 44833
rect 362806 44781 362858 44833
rect 212470 44633 212522 44685
rect 310102 44633 310154 44685
rect 507094 43301 507146 43353
rect 215062 43227 215114 43279
rect 518710 43227 518762 43279
rect 520342 43153 520394 43205
rect 206902 42265 206954 42317
rect 405526 42265 405578 42317
rect 213622 42191 213674 42243
rect 460054 42191 460106 42243
rect 214294 42117 214346 42169
rect 514870 42117 514922 42169
rect 404374 41525 404426 41577
rect 334102 40859 334154 40911
rect 344182 40859 344234 40911
rect 388822 40267 388874 40319
rect 394582 40267 394634 40319
rect 394582 37381 394634 37433
rect 404374 37381 404426 37433
<< metal2 >>
rect 92276 1016714 92332 1016723
rect 92276 1016649 92332 1016658
rect 81044 995846 81100 995855
rect 80784 995804 81044 995832
rect 82032 995813 82334 995832
rect 91248 995813 91550 995832
rect 92290 995813 92318 1016649
rect 148532 1015974 148588 1015983
rect 148532 1015909 148588 1015918
rect 353396 1015974 353452 1015983
rect 353396 1015909 353452 1015918
rect 148546 1007991 148574 1015909
rect 145364 1007982 145420 1007991
rect 145364 1007917 145420 1007926
rect 148532 1007982 148588 1007991
rect 148532 1007917 148588 1007926
rect 143734 1002393 143786 1002399
rect 143650 1002341 143734 1002344
rect 143650 1002335 143786 1002341
rect 143650 1002316 143774 1002335
rect 143926 1002319 143978 1002325
rect 92566 999507 92618 999513
rect 92566 999449 92618 999455
rect 92374 999433 92426 999439
rect 92374 999375 92426 999381
rect 82032 995807 82346 995813
rect 82032 995804 82294 995807
rect 81044 995781 81100 995790
rect 91248 995807 91562 995813
rect 91248 995804 91510 995807
rect 82294 995749 82346 995755
rect 91510 995749 91562 995755
rect 92278 995807 92330 995813
rect 92278 995749 92330 995755
rect 92386 995739 92414 999375
rect 89782 995733 89834 995739
rect 85940 995698 85996 995707
rect 85728 995656 85940 995684
rect 89424 995681 89782 995684
rect 89424 995675 89834 995681
rect 92374 995733 92426 995739
rect 92374 995675 92426 995681
rect 89424 995656 89822 995675
rect 85940 995633 85996 995642
rect 77088 995508 77342 995536
rect 66838 995141 66890 995147
rect 66838 995083 66890 995089
rect 61846 993587 61898 993593
rect 61846 993529 61898 993535
rect 50422 988333 50474 988339
rect 50422 988275 50474 988281
rect 47638 988259 47690 988265
rect 47638 988201 47690 988207
rect 44758 988185 44810 988191
rect 44758 988127 44810 988133
rect 43126 987889 43178 987895
rect 43126 987831 43178 987837
rect 42082 968771 42110 969252
rect 42068 968762 42124 968771
rect 42068 968697 42124 968706
rect 41794 967143 41822 967402
rect 43138 967323 43166 987831
rect 44566 986557 44618 986563
rect 44566 986499 44618 986505
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 43126 967317 43178 967323
rect 43126 967259 43178 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 42082 965071 42110 965552
rect 42068 965062 42124 965071
rect 42068 964997 42124 965006
rect 41794 964035 41822 964368
rect 41780 964026 41836 964035
rect 41780 963961 41836 963970
rect 41794 963295 41822 963702
rect 41780 963286 41836 963295
rect 41780 963221 41836 963230
rect 42836 963286 42892 963295
rect 42836 963221 42892 963230
rect 41794 962703 41822 963081
rect 41780 962694 41836 962703
rect 41780 962629 41836 962638
rect 41890 962111 41918 962518
rect 41876 962102 41932 962111
rect 41876 962037 41932 962046
rect 42178 960959 42206 961260
rect 42850 960959 42878 963221
rect 42166 960953 42218 960959
rect 42166 960895 42218 960901
rect 42838 960953 42890 960959
rect 42838 960895 42890 960901
rect 42178 960483 42206 960594
rect 42164 960474 42220 960483
rect 42164 960409 42220 960418
rect 41794 959743 41822 960045
rect 41780 959734 41836 959743
rect 41780 959669 41836 959678
rect 41794 959151 41822 959410
rect 41780 959142 41836 959151
rect 41780 959077 41836 959086
rect 42742 959103 42794 959109
rect 42742 959045 42794 959051
rect 41794 958559 41822 958744
rect 41780 958550 41836 958559
rect 41780 958485 41836 958494
rect 41890 957819 41918 958226
rect 41876 957810 41932 957819
rect 41876 957745 41932 957754
rect 42178 955895 42206 956376
rect 42164 955886 42220 955895
rect 42164 955821 42220 955830
rect 42192 955696 42494 955724
rect 42192 955063 42398 955091
rect 42166 953257 42218 953263
rect 42166 953199 42218 953205
rect 40340 943010 40396 943019
rect 40340 942945 40396 942954
rect 39958 942231 40010 942237
rect 39958 942173 40010 942179
rect 39970 933135 39998 942173
rect 39958 933129 40010 933135
rect 39958 933071 40010 933077
rect 40150 933129 40202 933135
rect 40150 933071 40202 933077
rect 35156 932650 35212 932659
rect 35156 932585 35212 932594
rect 35170 932215 35198 932585
rect 35156 932206 35212 932215
rect 35156 932141 35212 932150
rect 40162 927331 40190 933071
rect 40148 927322 40204 927331
rect 40148 927257 40204 927266
rect 39860 927174 39916 927183
rect 39860 927109 39916 927118
rect 39874 907235 39902 927109
rect 39862 907229 39914 907235
rect 39862 907171 39914 907177
rect 40246 907229 40298 907235
rect 40246 907171 40298 907177
rect 40258 892879 40286 907171
rect 40246 892873 40298 892879
rect 40246 892815 40298 892821
rect 40054 892799 40106 892805
rect 40054 892741 40106 892747
rect 40066 887033 40094 892741
rect 40054 887027 40106 887033
rect 40054 886969 40106 886975
rect 40150 887027 40202 887033
rect 40150 886969 40202 886975
rect 40162 872751 40190 886969
rect 40150 872745 40202 872751
rect 40150 872687 40202 872693
rect 40150 872523 40202 872529
rect 40150 872465 40202 872471
rect 40162 864019 40190 872465
rect 39862 864013 39914 864019
rect 39862 863955 39914 863961
rect 40150 864013 40202 864019
rect 40150 863955 40202 863961
rect 39874 843891 39902 863955
rect 39862 843885 39914 843891
rect 39862 843827 39914 843833
rect 40054 843885 40106 843891
rect 40054 843827 40106 843833
rect 40066 832569 40094 843827
rect 40054 832563 40106 832569
rect 40054 832505 40106 832511
rect 40246 832267 40298 832273
rect 40246 832209 40298 832215
rect 40258 816775 40286 832209
rect 40354 817219 40382 942945
rect 42178 938135 42206 953199
rect 42370 940355 42398 955063
rect 42466 953263 42494 955696
rect 42454 953257 42506 953263
rect 42454 953199 42506 953205
rect 42434 950148 42494 950157
rect 42434 950079 42494 950088
rect 42450 950040 42494 950079
rect 42356 940346 42412 940355
rect 42356 940281 42412 940290
rect 42164 938126 42220 938135
rect 42164 938061 42220 938070
rect 41686 872671 41738 872677
rect 41686 872613 41738 872619
rect 41698 818847 41726 872613
rect 41684 818838 41740 818847
rect 41684 818773 41740 818782
rect 40340 817210 40396 817219
rect 40340 817145 40396 817154
rect 40244 816766 40300 816775
rect 40244 816701 40300 816710
rect 40258 815031 40286 816701
rect 37366 815025 37418 815031
rect 37366 814967 37418 814973
rect 40246 815025 40298 815031
rect 40246 814967 40298 814973
rect 41780 814990 41836 814999
rect 35156 806850 35212 806859
rect 35156 806785 35212 806794
rect 35170 806415 35198 806785
rect 35156 806406 35212 806415
rect 35156 806341 35212 806350
rect 37378 802123 37406 814967
rect 41780 814925 41836 814934
rect 41684 813362 41740 813371
rect 41684 813297 41740 813306
rect 37364 802114 37420 802123
rect 41698 802100 41726 813297
rect 41794 802229 41822 814925
rect 41972 812770 42028 812779
rect 41972 812705 42028 812714
rect 41876 812326 41932 812335
rect 41876 812261 41932 812270
rect 41782 802223 41834 802229
rect 41782 802165 41834 802171
rect 41698 802072 41822 802100
rect 37364 802049 37420 802058
rect 41794 800231 41822 802072
rect 41890 800305 41918 812261
rect 41986 802451 42014 812705
rect 42068 811142 42124 811151
rect 42068 811077 42124 811086
rect 41974 802445 42026 802451
rect 41974 802387 42026 802393
rect 41974 802223 42026 802229
rect 41974 802165 42026 802171
rect 41986 800347 42014 802165
rect 42082 800495 42110 811077
rect 42164 810550 42220 810559
rect 42164 810485 42220 810494
rect 42068 800486 42124 800495
rect 42068 800421 42124 800430
rect 41972 800338 42028 800347
rect 41878 800299 41930 800305
rect 42178 800305 42206 810485
rect 42356 809514 42412 809523
rect 42356 809449 42412 809458
rect 41972 800273 42028 800282
rect 42166 800299 42218 800305
rect 41878 800241 41930 800247
rect 42166 800241 42218 800247
rect 41782 800225 41834 800231
rect 41782 800167 41834 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 42370 799755 42398 809449
rect 42356 799746 42412 799755
rect 42356 799681 42412 799690
rect 42166 798153 42218 798159
rect 42166 798095 42218 798101
rect 42178 797605 42206 798095
rect 42466 797683 42494 950040
rect 42644 944934 42700 944943
rect 42644 944869 42700 944878
rect 42658 944679 42686 944869
rect 42646 944673 42698 944679
rect 42646 944615 42698 944621
rect 42644 944342 42700 944351
rect 42644 944277 42646 944286
rect 42698 944277 42700 944286
rect 42646 944245 42698 944251
rect 42754 943833 42782 959045
rect 42850 950159 42878 960895
rect 42834 950150 42894 950159
rect 42834 950081 42894 950090
rect 42740 943824 42796 943833
rect 42740 943759 42796 943768
rect 42646 942749 42698 942755
rect 42644 942714 42646 942723
rect 42698 942714 42700 942723
rect 42644 942649 42700 942658
rect 44578 942237 44606 986499
rect 42646 942231 42698 942237
rect 42644 942196 42646 942205
rect 44566 942231 44618 942237
rect 42698 942196 42700 942205
rect 44566 942173 44618 942179
rect 42644 942131 42700 942140
rect 42644 932206 42700 932215
rect 42644 932141 42646 932150
rect 42698 932141 42700 932150
rect 42646 932109 42698 932115
rect 42646 819169 42698 819175
rect 42644 819134 42646 819143
rect 42698 819134 42700 819143
rect 42644 819069 42700 819078
rect 42646 818133 42698 818139
rect 42644 818098 42646 818107
rect 42698 818098 42700 818107
rect 42644 818033 42700 818042
rect 43220 817506 43276 817515
rect 43220 817441 43276 817450
rect 42644 814398 42700 814407
rect 42644 814333 42700 814342
rect 42658 798159 42686 814333
rect 43028 810402 43084 810411
rect 43028 810337 43084 810346
rect 42740 809292 42796 809301
rect 42740 809227 42796 809236
rect 42754 800897 42782 809227
rect 42836 808182 42892 808191
rect 42836 808117 42892 808126
rect 42742 800891 42794 800897
rect 42742 800833 42794 800839
rect 42646 798153 42698 798159
rect 42646 798095 42698 798101
rect 42452 797674 42508 797683
rect 42452 797609 42508 797618
rect 42550 797635 42602 797641
rect 42550 797577 42602 797583
rect 42452 797526 42508 797535
rect 42562 797512 42590 797577
rect 42562 797484 42686 797512
rect 42452 797461 42508 797470
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 42466 794311 42494 797461
rect 42548 797082 42604 797091
rect 42548 797017 42604 797026
rect 42070 794305 42122 794311
rect 42070 794247 42122 794253
rect 42454 794305 42506 794311
rect 42454 794247 42506 794253
rect 42082 793946 42110 794247
rect 42166 793861 42218 793867
rect 42166 793803 42218 793809
rect 42178 793280 42206 793803
rect 42166 793195 42218 793201
rect 42166 793137 42218 793143
rect 42178 792729 42206 793137
rect 42562 792979 42590 797017
rect 42550 792973 42602 792979
rect 42550 792915 42602 792921
rect 42658 792776 42686 797484
rect 42850 795051 42878 808117
rect 42934 802445 42986 802451
rect 42934 802387 42986 802393
rect 42838 795045 42890 795051
rect 42838 794987 42890 794993
rect 42946 793201 42974 802387
rect 43042 796309 43070 810337
rect 43124 808774 43180 808783
rect 43124 808709 43180 808718
rect 43030 796303 43082 796309
rect 43030 796245 43082 796251
rect 43030 796155 43082 796161
rect 43030 796097 43082 796103
rect 42934 793195 42986 793201
rect 42934 793137 42986 793143
rect 43042 793072 43070 796097
rect 43138 793867 43166 808709
rect 43126 793861 43178 793867
rect 43126 793803 43178 793809
rect 43126 793713 43178 793719
rect 43126 793655 43178 793661
rect 42946 793044 43070 793072
rect 42946 792924 42974 793044
rect 42466 792748 42686 792776
rect 42850 792896 42974 792924
rect 43030 792973 43082 792979
rect 43030 792915 43082 792921
rect 42466 792480 42494 792748
rect 42548 792642 42604 792651
rect 42604 792600 42686 792628
rect 42548 792577 42604 792586
rect 42466 792452 42590 792480
rect 42356 791902 42412 791911
rect 42356 791837 42412 791846
rect 42082 791319 42110 791430
rect 42068 791310 42124 791319
rect 42068 791245 42124 791254
rect 42164 791162 42220 791171
rect 42164 791097 42220 791106
rect 42178 790797 42206 791097
rect 42166 790531 42218 790537
rect 42166 790473 42218 790479
rect 42178 790246 42206 790473
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42166 788755 42218 788761
rect 42166 788697 42218 788703
rect 42178 788396 42206 788697
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42370 786467 42398 791837
rect 42452 791754 42508 791763
rect 42452 791689 42508 791698
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42358 786461 42410 786467
rect 42358 786403 42410 786409
rect 42178 785921 42206 786403
rect 42466 785653 42494 791689
rect 42562 790537 42590 792452
rect 42550 790531 42602 790537
rect 42550 790473 42602 790479
rect 42658 789520 42686 792600
rect 42562 789501 42686 789520
rect 42550 789495 42686 789501
rect 42602 789492 42686 789495
rect 42550 789437 42602 789443
rect 42850 788761 42878 792896
rect 42838 788755 42890 788761
rect 42838 788697 42890 788703
rect 43042 787059 43070 792915
rect 43138 789945 43166 793655
rect 43126 789939 43178 789945
rect 43126 789881 43178 789887
rect 43030 787053 43082 787059
rect 43030 786995 43082 787001
rect 42070 785647 42122 785653
rect 42070 785589 42122 785595
rect 42454 785647 42506 785653
rect 42454 785589 42506 785595
rect 42082 785288 42110 785589
rect 42454 776101 42506 776107
rect 42452 776066 42454 776075
rect 42506 776066 42508 776075
rect 42452 776001 42508 776010
rect 42838 775361 42890 775367
rect 42836 775326 42838 775335
rect 42890 775326 42892 775335
rect 42836 775261 42892 775270
rect 42838 774843 42890 774849
rect 42836 774808 42838 774817
rect 42890 774808 42892 774817
rect 42836 774743 42892 774752
rect 43234 773707 43262 817441
rect 44564 806554 44620 806563
rect 44564 806489 44620 806498
rect 43414 800891 43466 800897
rect 43414 800833 43466 800839
rect 43318 800225 43370 800231
rect 43318 800167 43370 800173
rect 43330 796161 43358 800167
rect 43426 797641 43454 800833
rect 43510 800299 43562 800305
rect 43510 800241 43562 800247
rect 43414 797635 43466 797641
rect 43414 797577 43466 797583
rect 43318 796155 43370 796161
rect 43318 796097 43370 796103
rect 43522 793719 43550 800241
rect 43510 793713 43562 793719
rect 43510 793655 43562 793661
rect 43412 774290 43468 774299
rect 43412 774225 43468 774234
rect 43220 773698 43276 773707
rect 43220 773633 43276 773642
rect 43028 772070 43084 772079
rect 43028 772005 43084 772014
rect 42068 771182 42124 771191
rect 42068 771117 42124 771126
rect 40244 770738 40300 770747
rect 40244 770673 40300 770682
rect 35156 763634 35212 763643
rect 35156 763569 35212 763578
rect 35170 763199 35198 763569
rect 35156 763190 35212 763199
rect 35156 763125 35212 763134
rect 40258 760239 40286 770673
rect 41684 769554 41740 769563
rect 41684 769489 41740 769498
rect 41588 764818 41644 764827
rect 41588 764753 41644 764762
rect 40244 760230 40300 760239
rect 40244 760165 40300 760174
rect 41602 757427 41630 764753
rect 41588 757418 41644 757427
rect 41588 757353 41644 757362
rect 41698 757311 41726 769489
rect 41876 766298 41932 766307
rect 41876 766233 41932 766242
rect 41780 765854 41836 765863
rect 41780 765789 41836 765798
rect 41686 757305 41738 757311
rect 41686 757247 41738 757253
rect 41794 757089 41822 765789
rect 41890 757131 41918 766233
rect 42082 760239 42110 771117
rect 42836 770442 42892 770451
rect 42836 770377 42892 770386
rect 42356 769110 42412 769119
rect 42356 769045 42412 769054
rect 42164 767926 42220 767935
rect 42164 767861 42220 767870
rect 42068 760230 42124 760239
rect 42068 760165 42124 760174
rect 42178 757131 42206 767861
rect 41876 757122 41932 757131
rect 41782 757083 41834 757089
rect 41876 757057 41932 757066
rect 42164 757122 42220 757131
rect 42164 757057 42220 757066
rect 41782 757025 41834 757031
rect 42370 756793 42398 769045
rect 42850 759203 42878 770377
rect 42932 767778 42988 767787
rect 42932 767713 42988 767722
rect 42836 759194 42892 759203
rect 42836 759129 42892 759138
rect 42946 757607 42974 767713
rect 42934 757601 42986 757607
rect 42934 757543 42986 757549
rect 42934 757453 42986 757459
rect 42934 757395 42986 757401
rect 42166 756787 42218 756793
rect 42166 756729 42218 756735
rect 42358 756787 42410 756793
rect 42358 756729 42410 756735
rect 42178 756245 42206 756729
rect 42068 754902 42124 754911
rect 42068 754837 42124 754846
rect 42082 754430 42110 754837
rect 42946 754277 42974 757395
rect 42934 754271 42986 754277
rect 42934 754213 42986 754219
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42082 752580 42110 753029
rect 43042 751951 43070 772005
rect 43124 767186 43180 767195
rect 43124 767121 43180 767130
rect 43138 753093 43166 767121
rect 43318 757083 43370 757089
rect 43318 757025 43370 757031
rect 43126 753087 43178 753093
rect 43126 753029 43178 753035
rect 43330 752964 43358 757025
rect 43138 752936 43358 752964
rect 43028 751942 43084 751951
rect 43028 751877 43084 751886
rect 42068 751794 42124 751803
rect 42068 751729 42124 751738
rect 42082 751396 42110 751729
rect 42838 751681 42890 751687
rect 42740 751646 42796 751655
rect 42838 751623 42890 751629
rect 42740 751581 42796 751590
rect 41876 751054 41932 751063
rect 41876 750989 41932 750998
rect 41890 750730 41918 750989
rect 42164 750610 42220 750619
rect 42164 750545 42220 750554
rect 42178 750064 42206 750545
rect 42070 749831 42122 749837
rect 42070 749773 42122 749779
rect 42082 749546 42110 749773
rect 41972 748686 42028 748695
rect 41972 748621 42028 748630
rect 41986 748214 42014 748621
rect 41794 747215 41822 747622
rect 42166 747315 42218 747321
rect 42166 747257 42218 747263
rect 41780 747206 41836 747215
rect 41780 747141 41836 747150
rect 42178 747030 42206 747257
rect 42166 746945 42218 746951
rect 42166 746887 42218 746893
rect 42178 746401 42206 746887
rect 42754 746285 42782 751581
rect 42850 749837 42878 751623
rect 43028 750314 43084 750323
rect 43028 750249 43084 750258
rect 42838 749831 42890 749837
rect 42838 749773 42890 749779
rect 42836 749722 42892 749731
rect 42836 749657 42892 749666
rect 42070 746279 42122 746285
rect 42070 746221 42122 746227
rect 42742 746279 42794 746285
rect 42742 746221 42794 746227
rect 42082 745772 42110 746221
rect 42740 746170 42796 746179
rect 42740 746105 42796 746114
rect 42166 745539 42218 745545
rect 42166 745481 42218 745487
rect 42178 745180 42206 745481
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42178 743365 42206 743779
rect 42754 743251 42782 746105
rect 42850 743843 42878 749657
rect 43042 745545 43070 750249
rect 43138 747321 43166 752936
rect 43126 747315 43178 747321
rect 43126 747257 43178 747263
rect 43124 746910 43180 746919
rect 43124 746845 43180 746854
rect 43030 745539 43082 745545
rect 43030 745481 43082 745487
rect 42838 743837 42890 743843
rect 42838 743779 42890 743785
rect 42070 743245 42122 743251
rect 42070 743187 42122 743193
rect 42742 743245 42794 743251
rect 42742 743187 42794 743193
rect 42082 742738 42110 743187
rect 43138 742437 43166 746845
rect 42166 742431 42218 742437
rect 42166 742373 42218 742379
rect 43126 742431 43178 742437
rect 43126 742373 43178 742379
rect 42178 742072 42206 742373
rect 42742 732737 42794 732743
rect 42740 732702 42742 732711
rect 42794 732702 42796 732711
rect 42740 732637 42796 732646
rect 42742 732145 42794 732151
rect 42740 732110 42742 732119
rect 42794 732110 42796 732119
rect 42740 732045 42796 732054
rect 42358 731849 42410 731855
rect 42356 731814 42358 731823
rect 42410 731814 42412 731823
rect 42356 731749 42412 731758
rect 43426 730491 43454 774225
rect 43606 757601 43658 757607
rect 43606 757543 43658 757549
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43522 751687 43550 757247
rect 43510 751681 43562 751687
rect 43510 751623 43562 751629
rect 43618 746951 43646 757543
rect 43606 746945 43658 746951
rect 43606 746887 43658 746893
rect 43700 731074 43756 731083
rect 43700 731009 43756 731018
rect 43412 730482 43468 730491
rect 43412 730417 43468 730426
rect 41588 728706 41644 728715
rect 41588 728641 41644 728650
rect 40724 724266 40780 724275
rect 40724 724201 40780 724210
rect 35156 720418 35212 720427
rect 35156 720353 35212 720362
rect 35170 719983 35198 720353
rect 35156 719974 35212 719983
rect 35156 719909 35212 719918
rect 40738 714211 40766 724201
rect 41492 723082 41548 723091
rect 41492 723017 41548 723026
rect 41506 714211 41534 723017
rect 41602 714359 41630 728641
rect 41876 727966 41932 727975
rect 41876 727901 41932 727910
rect 41684 726930 41740 726939
rect 41684 726865 41740 726874
rect 41588 714350 41644 714359
rect 41588 714285 41644 714294
rect 41698 714290 41726 726865
rect 41780 726338 41836 726347
rect 41780 726273 41836 726282
rect 41674 714238 41680 714290
rect 41732 714238 41738 714290
rect 40724 714202 40780 714211
rect 40724 714137 40780 714146
rect 41492 714202 41548 714211
rect 41492 714137 41548 714146
rect 41794 714021 41822 726273
rect 41782 714015 41834 714021
rect 41782 713957 41834 713963
rect 41890 713915 41918 727901
rect 42356 725894 42412 725903
rect 42356 725829 42412 725838
rect 42164 723674 42220 723683
rect 42164 723609 42220 723618
rect 42178 713915 42206 723609
rect 41876 713906 41932 713915
rect 41876 713841 41932 713850
rect 42164 713906 42220 713915
rect 42164 713841 42220 713850
rect 42370 713577 42398 725829
rect 43028 722934 43084 722943
rect 43028 722869 43084 722878
rect 42740 721824 42796 721833
rect 42740 721759 42796 721768
rect 42754 720681 42782 721759
rect 42742 720675 42794 720681
rect 42742 720617 42794 720623
rect 42742 720453 42794 720459
rect 42742 720395 42794 720401
rect 42070 713571 42122 713577
rect 42070 713513 42122 713519
rect 42358 713571 42410 713577
rect 42358 713513 42410 713519
rect 42082 713064 42110 713513
rect 42068 711686 42124 711695
rect 42068 711621 42124 711630
rect 42082 711214 42110 711621
rect 42754 711547 42782 720395
rect 43042 711695 43070 722869
rect 43126 717123 43178 717129
rect 43126 717065 43178 717071
rect 43028 711686 43084 711695
rect 43028 711621 43084 711630
rect 43030 711573 43082 711579
rect 42740 711538 42796 711547
rect 43030 711515 43082 711521
rect 43138 711524 43166 717065
rect 43510 714089 43562 714095
rect 43510 714031 43562 714037
rect 43414 714015 43466 714021
rect 43414 713957 43466 713963
rect 43426 711727 43454 713957
rect 43414 711721 43466 711727
rect 43414 711663 43466 711669
rect 42740 711473 42796 711482
rect 42452 711242 42508 711251
rect 42452 711177 42508 711186
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42164 709910 42220 709919
rect 42164 709845 42220 709854
rect 42178 709364 42206 709845
rect 42070 708613 42122 708619
rect 42070 708555 42122 708561
rect 42082 708180 42110 708555
rect 42466 708101 42494 711177
rect 43042 711061 43070 711515
rect 43138 711496 43454 711524
rect 43220 711390 43276 711399
rect 43220 711325 43276 711334
rect 43234 711228 43262 711325
rect 43138 711200 43262 711228
rect 43030 711055 43082 711061
rect 43030 710997 43082 711003
rect 43028 710946 43084 710955
rect 43028 710881 43084 710890
rect 42166 708095 42218 708101
rect 42166 708037 42218 708043
rect 42454 708095 42506 708101
rect 42454 708037 42506 708043
rect 42178 707514 42206 708037
rect 41780 707394 41836 707403
rect 41780 707329 41836 707338
rect 41794 706881 41822 707329
rect 42452 707246 42508 707255
rect 42452 707181 42508 707190
rect 42166 706615 42218 706621
rect 42166 706557 42218 706563
rect 42178 706330 42206 706557
rect 42356 705174 42412 705183
rect 42356 705109 42412 705118
rect 42178 704591 42206 705041
rect 42164 704582 42220 704591
rect 42164 704517 42220 704526
rect 41794 704147 41822 704406
rect 41780 704138 41836 704147
rect 41780 704073 41836 704082
rect 42166 704099 42218 704105
rect 42166 704041 42218 704047
rect 42178 703845 42206 704041
rect 42070 703581 42122 703587
rect 42070 703523 42122 703529
rect 42082 703222 42110 703523
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42178 702556 42206 702857
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42068 700586 42124 700595
rect 42068 700521 42124 700530
rect 42082 700188 42110 700521
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42178 699522 42206 700045
rect 42370 699443 42398 705109
rect 42466 703587 42494 707181
rect 43042 704327 43070 710881
rect 43138 708619 43166 711200
rect 43222 711055 43274 711061
rect 43222 710997 43274 711003
rect 43126 708613 43178 708619
rect 43126 708555 43178 708561
rect 43234 708416 43262 710997
rect 43426 710913 43454 711496
rect 43414 710907 43466 710913
rect 43414 710849 43466 710855
rect 43138 708388 43262 708416
rect 43138 706621 43166 708388
rect 43126 706615 43178 706621
rect 43126 706557 43178 706563
rect 43124 706506 43180 706515
rect 43124 706441 43180 706450
rect 43030 704321 43082 704327
rect 43030 704263 43082 704269
rect 43030 704173 43082 704179
rect 43030 704115 43082 704121
rect 42454 703581 42506 703587
rect 42454 703523 42506 703529
rect 42452 703398 42508 703407
rect 42452 703333 42508 703342
rect 42466 700109 42494 703333
rect 43042 702329 43070 704115
rect 43138 702921 43166 706441
rect 43522 704179 43550 714031
rect 43510 704173 43562 704179
rect 43510 704115 43562 704121
rect 43126 702915 43178 702921
rect 43126 702857 43178 702863
rect 43030 702323 43082 702329
rect 43030 702265 43082 702271
rect 43714 701312 43742 731009
rect 43522 701284 43742 701312
rect 42454 700103 42506 700109
rect 42454 700045 42506 700051
rect 43126 699881 43178 699887
rect 43126 699823 43178 699829
rect 42166 699437 42218 699443
rect 42166 699379 42218 699385
rect 42358 699437 42410 699443
rect 42358 699379 42410 699385
rect 42178 698856 42206 699379
rect 43138 689051 43166 699823
rect 43222 689521 43274 689527
rect 43220 689486 43222 689495
rect 43274 689486 43276 689495
rect 43220 689421 43276 689430
rect 43124 689042 43180 689051
rect 43124 688977 43180 688986
rect 42838 688485 42890 688491
rect 42836 688450 42838 688459
rect 42890 688450 42892 688459
rect 42836 688385 42892 688394
rect 43412 687858 43468 687867
rect 43412 687793 43468 687802
rect 42068 685490 42124 685499
rect 42068 685425 42124 685434
rect 41876 684898 41932 684907
rect 41876 684833 41932 684842
rect 41012 681494 41068 681503
rect 41012 681429 41068 681438
rect 35156 677202 35212 677211
rect 35156 677137 35212 677146
rect 35170 676767 35198 677137
rect 35156 676758 35212 676767
rect 35156 676693 35212 676702
rect 41026 670995 41054 681429
rect 41780 678830 41836 678839
rect 41780 678765 41836 678774
rect 41684 675574 41740 675583
rect 41684 675509 41740 675518
rect 41698 670995 41726 675509
rect 41012 670986 41068 670995
rect 41012 670921 41068 670930
rect 41684 670986 41740 670995
rect 41684 670921 41740 670930
rect 41794 670657 41822 678765
rect 41890 672137 41918 684833
rect 41972 679866 42028 679875
rect 41972 679801 42028 679810
rect 41878 672131 41930 672137
rect 41878 672073 41930 672079
rect 41986 670731 42014 679801
rect 41974 670725 42026 670731
rect 42082 670699 42110 685425
rect 42356 682678 42412 682687
rect 42356 682613 42412 682622
rect 42164 680458 42220 680467
rect 42164 680393 42220 680402
rect 42178 674061 42206 680393
rect 42166 674055 42218 674061
rect 42166 673997 42218 674003
rect 41974 670667 42026 670673
rect 42068 670690 42124 670699
rect 41782 670651 41834 670657
rect 42068 670625 42124 670634
rect 41782 670593 41834 670599
rect 42370 670361 42398 682613
rect 43220 681346 43276 681355
rect 43220 681281 43276 681290
rect 43124 679866 43180 679875
rect 43124 679801 43180 679810
rect 43138 675708 43166 679801
rect 42946 675680 43166 675708
rect 42646 672131 42698 672137
rect 42646 672073 42698 672079
rect 42658 670805 42686 672073
rect 42946 670995 42974 675680
rect 43030 674055 43082 674061
rect 43030 673997 43082 674003
rect 42932 670986 42988 670995
rect 42932 670921 42988 670930
rect 43042 670824 43070 673997
rect 43234 670953 43262 681281
rect 43426 679408 43454 687793
rect 43522 687719 43550 701284
rect 43508 687710 43564 687719
rect 43508 687645 43564 687654
rect 43700 683714 43756 683723
rect 43700 683649 43756 683658
rect 43330 679380 43454 679408
rect 43222 670947 43274 670953
rect 43222 670889 43274 670895
rect 42646 670799 42698 670805
rect 42646 670741 42698 670747
rect 42934 670799 42986 670805
rect 43042 670796 43262 670824
rect 42934 670741 42986 670747
rect 42646 670651 42698 670657
rect 42646 670593 42698 670599
rect 42166 670355 42218 670361
rect 42166 670297 42218 670303
rect 42358 670355 42410 670361
rect 42358 670297 42410 670303
rect 42178 669848 42206 670297
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42164 665362 42220 665371
rect 42164 665297 42220 665306
rect 42178 664964 42206 665297
rect 42164 664770 42220 664779
rect 42164 664705 42220 664714
rect 42178 664298 42206 664705
rect 42658 664219 42686 670593
rect 42946 668585 42974 670741
rect 43126 670725 43178 670731
rect 43028 670690 43084 670699
rect 43126 670667 43178 670673
rect 43028 670625 43084 670634
rect 42934 668579 42986 668585
rect 42934 668521 42986 668527
rect 42934 668431 42986 668437
rect 42934 668373 42986 668379
rect 42946 666735 42974 668373
rect 42934 666729 42986 666735
rect 42934 666671 42986 666677
rect 42934 665249 42986 665255
rect 42934 665191 42986 665197
rect 42070 664213 42122 664219
rect 42070 664155 42122 664161
rect 42646 664213 42698 664219
rect 42646 664155 42698 664161
rect 42082 663706 42110 664155
rect 42644 664030 42700 664039
rect 42644 663965 42700 663974
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42178 663114 42206 663341
rect 42356 662846 42412 662855
rect 42356 662781 42412 662790
rect 42068 662254 42124 662263
rect 42068 662189 42124 662198
rect 42082 661856 42110 662189
rect 41890 661079 41918 661190
rect 42070 661105 42122 661111
rect 41876 661070 41932 661079
rect 42070 661047 42122 661053
rect 41876 661005 41932 661014
rect 42082 660672 42110 661047
rect 42070 660439 42122 660445
rect 42070 660381 42122 660387
rect 42082 660006 42110 660381
rect 42166 659699 42218 659705
rect 42166 659641 42218 659647
rect 42178 659340 42206 659641
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42082 658822 42110 659049
rect 42370 657411 42398 662781
rect 42658 659705 42686 663965
rect 42946 660445 42974 665191
rect 43042 663405 43070 670625
rect 43030 663399 43082 663405
rect 43030 663341 43082 663347
rect 43028 662402 43084 662411
rect 43028 662337 43084 662346
rect 42934 660439 42986 660445
rect 42934 660381 42986 660387
rect 42646 659699 42698 659705
rect 42646 659641 42698 659647
rect 42658 659557 42782 659576
rect 42646 659551 42782 659557
rect 42698 659548 42782 659551
rect 42646 659493 42698 659499
rect 42754 659132 42782 659548
rect 42658 659113 42782 659132
rect 42646 659107 42782 659113
rect 42698 659104 42782 659107
rect 42646 659049 42698 659055
rect 42070 657405 42122 657411
rect 42070 657347 42122 657353
rect 42358 657405 42410 657411
rect 42358 657347 42410 657353
rect 42082 656972 42110 657347
rect 42934 656739 42986 656745
rect 42934 656681 42986 656687
rect 42166 656665 42218 656671
rect 42166 656607 42218 656613
rect 42178 656306 42206 656607
rect 42166 656221 42218 656227
rect 42166 656163 42218 656169
rect 42178 655677 42206 656163
rect 42946 646279 42974 656681
rect 43042 656671 43070 662337
rect 43138 661111 43166 670667
rect 43234 668437 43262 670796
rect 43222 668431 43274 668437
rect 43222 668373 43274 668379
rect 43126 661105 43178 661111
rect 43126 661047 43178 661053
rect 43124 660922 43180 660931
rect 43124 660857 43180 660866
rect 43030 656665 43082 656671
rect 43030 656607 43082 656613
rect 43138 656227 43166 660857
rect 43126 656221 43178 656227
rect 43126 656163 43178 656169
rect 43222 647785 43274 647791
rect 43222 647727 43274 647733
rect 42932 646270 42988 646279
rect 42932 646205 42988 646214
rect 42356 645530 42412 645539
rect 42356 645465 42412 645474
rect 42370 645127 42398 645465
rect 43234 645243 43262 647727
rect 43220 645234 43276 645243
rect 43220 645169 43276 645178
rect 42358 645121 42410 645127
rect 42358 645063 42410 645069
rect 43330 644503 43358 679380
rect 43414 673907 43466 673913
rect 43414 673849 43466 673855
rect 43426 670972 43454 673849
rect 43426 670944 43550 670972
rect 43414 670873 43466 670879
rect 43414 670815 43466 670821
rect 43426 665255 43454 670815
rect 43522 667919 43550 670944
rect 43510 667913 43562 667919
rect 43510 667855 43562 667861
rect 43414 665249 43466 665255
rect 43414 665191 43466 665197
rect 43714 659557 43742 683649
rect 43702 659551 43754 659557
rect 43702 659493 43754 659499
rect 43796 647158 43852 647167
rect 43796 647093 43852 647102
rect 43604 647010 43660 647019
rect 43604 646945 43660 646954
rect 43316 644494 43372 644503
rect 43316 644429 43372 644438
rect 43618 643023 43646 646945
rect 43810 643615 43838 647093
rect 43988 644642 44044 644651
rect 43988 644577 44044 644586
rect 43796 643606 43852 643615
rect 43796 643541 43852 643550
rect 43604 643014 43660 643023
rect 43604 642949 43660 642958
rect 43508 642126 43564 642135
rect 43508 642061 43564 642070
rect 41780 641682 41836 641691
rect 41780 641617 41836 641626
rect 41012 640498 41068 640507
rect 41012 640433 41068 640442
rect 35156 633986 35212 633995
rect 35156 633921 35212 633930
rect 35170 633551 35198 633921
rect 35156 633542 35212 633551
rect 35156 633477 35212 633486
rect 41026 627811 41054 640433
rect 41588 640054 41644 640063
rect 41588 639989 41644 639998
rect 41492 638426 41548 638435
rect 41492 638361 41548 638370
rect 41014 627805 41066 627811
rect 41506 627779 41534 638361
rect 41014 627747 41066 627753
rect 41492 627770 41548 627779
rect 41602 627737 41630 639989
rect 41794 631807 41822 641617
rect 41876 639462 41932 639471
rect 41876 639397 41932 639406
rect 41782 631801 41834 631807
rect 41782 631743 41834 631749
rect 41492 627705 41548 627714
rect 41590 627731 41642 627737
rect 41590 627673 41642 627679
rect 41890 627441 41918 639397
rect 41972 637834 42028 637843
rect 41972 637769 42028 637778
rect 41986 627483 42014 637769
rect 43220 637242 43276 637251
rect 43220 637177 43276 637186
rect 42164 636798 42220 636807
rect 42164 636733 42220 636742
rect 42068 636206 42124 636215
rect 42068 636141 42124 636150
rect 42082 627631 42110 636141
rect 42178 628223 42206 636733
rect 42356 635170 42412 635179
rect 42356 635105 42412 635114
rect 42164 628214 42220 628223
rect 42164 628149 42220 628158
rect 42068 627622 42124 627631
rect 42068 627557 42124 627566
rect 41972 627474 42028 627483
rect 41878 627435 41930 627441
rect 41972 627409 42028 627418
rect 41878 627377 41930 627383
rect 41878 627213 41930 627219
rect 41878 627155 41930 627161
rect 41890 626632 41918 627155
rect 42370 627039 42398 635105
rect 42646 631801 42698 631807
rect 42646 631743 42698 631749
rect 42658 628329 42686 631743
rect 42646 628323 42698 628329
rect 42646 628265 42698 628271
rect 42644 628214 42700 628223
rect 42700 628172 42782 628200
rect 42644 628149 42700 628158
rect 42646 628027 42698 628033
rect 42646 627969 42698 627975
rect 42454 627953 42506 627959
rect 42454 627895 42506 627901
rect 42356 627030 42412 627039
rect 42356 626965 42412 626974
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42178 624782 42206 625305
rect 42466 624703 42494 627895
rect 42658 625369 42686 627969
rect 42646 625363 42698 625369
rect 42646 625305 42698 625311
rect 42754 625240 42782 628172
rect 43126 627731 43178 627737
rect 43126 627673 43178 627679
rect 42658 625212 42782 625240
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42454 624697 42506 624703
rect 42454 624639 42506 624645
rect 42178 624161 42206 624639
rect 42452 624514 42508 624523
rect 42452 624449 42508 624458
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42466 622261 42494 624449
rect 42166 622255 42218 622261
rect 42166 622197 42218 622203
rect 42454 622255 42506 622261
rect 42454 622197 42506 622203
rect 42178 621748 42206 622197
rect 42452 622146 42508 622155
rect 42452 622081 42508 622090
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42070 620923 42122 620929
rect 42070 620865 42122 620871
rect 42082 620490 42110 620865
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 42178 619929 42206 620347
rect 42356 619630 42412 619639
rect 42356 619565 42412 619574
rect 42178 618307 42206 618640
rect 42164 618298 42220 618307
rect 42164 618233 42220 618242
rect 41986 617715 42014 617974
rect 42070 617889 42122 617895
rect 42070 617831 42122 617837
rect 41972 617706 42028 617715
rect 41972 617641 42028 617650
rect 42082 617456 42110 617831
rect 42166 617371 42218 617377
rect 42166 617313 42218 617319
rect 42178 616790 42206 617313
rect 42370 616711 42398 619565
rect 42466 617377 42494 622081
rect 42658 621669 42686 625212
rect 42646 621663 42698 621669
rect 42646 621605 42698 621611
rect 42644 621554 42700 621563
rect 42644 621489 42700 621498
rect 42658 617895 42686 621489
rect 43138 620411 43166 627673
rect 43234 623519 43262 637177
rect 43316 635614 43372 635623
rect 43316 635549 43372 635558
rect 43222 623513 43274 623519
rect 43222 623455 43274 623461
rect 43330 620929 43358 635549
rect 43414 627805 43466 627811
rect 43414 627747 43466 627753
rect 43318 620923 43370 620929
rect 43318 620865 43370 620871
rect 43126 620405 43178 620411
rect 43126 620347 43178 620353
rect 43426 620208 43454 627747
rect 43138 620180 43454 620208
rect 42646 617889 42698 617895
rect 42646 617831 42698 617837
rect 42454 617371 42506 617377
rect 42454 617313 42506 617319
rect 42452 617262 42508 617271
rect 42452 617197 42508 617206
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42358 616705 42410 616711
rect 42358 616647 42410 616653
rect 42178 616157 42206 616647
rect 42356 616522 42412 616531
rect 42356 616457 42412 616466
rect 42166 615891 42218 615897
rect 42166 615833 42218 615839
rect 42178 615606 42206 615833
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 42178 613756 42206 614131
rect 42370 613677 42398 616457
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42358 613671 42410 613677
rect 42358 613613 42410 613619
rect 42178 613121 42206 613613
rect 42358 613523 42410 613529
rect 42358 613465 42410 613471
rect 42070 613005 42122 613011
rect 42070 612947 42122 612953
rect 42082 612498 42110 612947
rect 42370 602175 42398 613465
rect 42466 613011 42494 617197
rect 43138 615897 43166 620180
rect 43126 615891 43178 615897
rect 43126 615833 43178 615839
rect 43522 614195 43550 642061
rect 43510 614189 43562 614195
rect 43510 614131 43562 614137
rect 42454 613005 42506 613011
rect 42454 612947 42506 612953
rect 42452 602906 42508 602915
rect 42452 602841 42508 602850
rect 42356 602166 42412 602175
rect 42356 602101 42412 602110
rect 42466 601911 42494 602841
rect 43220 602462 43276 602471
rect 43220 602397 43276 602406
rect 43234 601985 43262 602397
rect 43222 601979 43274 601985
rect 43222 601921 43274 601927
rect 42454 601905 42506 601911
rect 42454 601847 42506 601853
rect 43220 601426 43276 601435
rect 43220 601361 43276 601370
rect 43124 598762 43180 598771
rect 43124 598697 43180 598706
rect 41588 597282 41644 597291
rect 41588 597217 41644 597226
rect 41602 584595 41630 597217
rect 41780 596838 41836 596847
rect 41780 596773 41836 596782
rect 41684 594618 41740 594627
rect 41684 594553 41740 594562
rect 41590 584589 41642 584595
rect 41590 584531 41642 584537
rect 41698 584521 41726 594553
rect 41686 584515 41738 584521
rect 41686 584457 41738 584463
rect 41794 584299 41822 596773
rect 41876 596246 41932 596255
rect 41876 596181 41932 596190
rect 41782 584293 41834 584299
rect 41782 584235 41834 584241
rect 41890 584225 41918 596181
rect 41972 595210 42028 595219
rect 41972 595145 42028 595154
rect 41986 584267 42014 595145
rect 42932 594396 42988 594405
rect 42932 594331 42988 594340
rect 42068 593582 42124 593591
rect 42068 593517 42124 593526
rect 41972 584258 42028 584267
rect 41878 584219 41930 584225
rect 42082 584225 42110 593517
rect 42946 584447 42974 594331
rect 43028 592768 43084 592777
rect 43028 592703 43084 592712
rect 42934 584441 42986 584447
rect 42934 584383 42986 584389
rect 43042 584373 43070 592703
rect 43138 584669 43166 598697
rect 43126 584663 43178 584669
rect 43126 584605 43178 584611
rect 43126 584515 43178 584521
rect 43126 584457 43178 584463
rect 43030 584367 43082 584373
rect 43030 584309 43082 584315
rect 42934 584293 42986 584299
rect 42934 584235 42986 584241
rect 41972 584193 42028 584202
rect 42070 584219 42122 584225
rect 41878 584161 41930 584167
rect 42070 584161 42122 584167
rect 42454 584145 42506 584151
rect 42454 584087 42506 584093
rect 41878 583997 41930 584003
rect 41878 583939 41930 583945
rect 41890 583445 41918 583939
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42178 581605 42206 582089
rect 42466 581487 42494 584087
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42454 581481 42506 581487
rect 42454 581423 42506 581429
rect 42082 580974 42110 581423
rect 42452 581298 42508 581307
rect 42452 581233 42508 581242
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42082 579790 42110 580239
rect 42164 578930 42220 578939
rect 42164 578865 42220 578874
rect 42178 578569 42206 578865
rect 42070 578447 42122 578453
rect 42070 578389 42122 578395
rect 42082 577940 42110 578389
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 42070 577189 42122 577195
rect 42070 577131 42122 577137
rect 42082 576756 42110 577131
rect 41972 575970 42028 575979
rect 41972 575905 42028 575914
rect 41986 575424 42014 575905
rect 41794 574499 41822 574797
rect 42068 574638 42124 574647
rect 42068 574573 42124 574582
rect 41780 574490 41836 574499
rect 41780 574425 41836 574434
rect 42082 574240 42110 574573
rect 42166 574007 42218 574013
rect 42166 573949 42218 573955
rect 42178 573574 42206 573949
rect 42466 573273 42494 581233
rect 42946 577195 42974 584235
rect 43030 584219 43082 584225
rect 43030 584161 43082 584167
rect 43042 578453 43070 584161
rect 43030 578447 43082 578453
rect 43030 578389 43082 578395
rect 43030 578299 43082 578305
rect 43030 578241 43082 578247
rect 42934 577189 42986 577195
rect 42934 577131 42986 577137
rect 42932 577006 42988 577015
rect 42932 576941 42988 576950
rect 42070 573267 42122 573273
rect 42070 573209 42122 573215
rect 42454 573267 42506 573273
rect 42454 573209 42506 573215
rect 42082 572982 42110 573209
rect 42452 573158 42508 573167
rect 42452 573093 42508 573102
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42178 572390 42206 572617
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 42178 570540 42206 570989
rect 42466 570461 42494 573093
rect 42946 571053 42974 576941
rect 43042 572681 43070 578241
rect 43138 574013 43166 584457
rect 43126 574007 43178 574013
rect 43126 573949 43178 573955
rect 43124 573898 43180 573907
rect 43124 573833 43180 573842
rect 43030 572675 43082 572681
rect 43030 572617 43082 572623
rect 43138 572552 43166 573833
rect 43042 572524 43166 572552
rect 42934 571047 42986 571053
rect 42934 570989 42986 570995
rect 42166 570455 42218 570461
rect 42166 570397 42218 570403
rect 42454 570455 42506 570461
rect 42454 570397 42506 570403
rect 42178 570332 42206 570397
rect 42082 570304 42206 570332
rect 42934 570307 42986 570313
rect 42082 569948 42110 570304
rect 42934 570249 42986 570255
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42082 569282 42110 569657
rect 42548 559542 42604 559551
rect 42548 559477 42604 559486
rect 42452 559098 42508 559107
rect 42452 559033 42454 559042
rect 42506 559033 42508 559042
rect 42454 559001 42506 559007
rect 42562 558917 42590 559477
rect 42550 558911 42602 558917
rect 42550 558853 42602 558859
rect 42946 558811 42974 570249
rect 43042 569721 43070 572524
rect 43030 569715 43082 569721
rect 43030 569657 43082 569663
rect 42932 558802 42988 558811
rect 42932 558737 42988 558746
rect 43234 558071 43262 601361
rect 43618 600103 43646 642949
rect 43810 600399 43838 643541
rect 44002 601287 44030 644577
rect 43988 601278 44044 601287
rect 43988 601213 44044 601222
rect 43796 600390 43852 600399
rect 43796 600325 43852 600334
rect 43412 600094 43468 600103
rect 43412 600029 43468 600038
rect 43604 600094 43660 600103
rect 43604 600029 43660 600038
rect 43426 584669 43454 600029
rect 43318 584663 43370 584669
rect 43318 584605 43370 584611
rect 43414 584663 43466 584669
rect 43414 584605 43466 584611
rect 43330 582153 43358 584605
rect 43510 584589 43562 584595
rect 43510 584531 43562 584537
rect 43414 584441 43466 584447
rect 43414 584383 43466 584389
rect 43318 582147 43370 582153
rect 43318 582089 43370 582095
rect 43426 580303 43454 584383
rect 43414 580297 43466 580303
rect 43414 580239 43466 580245
rect 43522 578305 43550 584531
rect 43606 584367 43658 584373
rect 43606 584309 43658 584315
rect 43510 578299 43562 578305
rect 43510 578241 43562 578247
rect 43618 577713 43646 584309
rect 43606 577707 43658 577713
rect 43606 577649 43658 577655
rect 43510 571713 43562 571719
rect 43510 571655 43562 571661
rect 43522 560587 43550 571655
rect 43810 570355 43838 600325
rect 43894 584663 43946 584669
rect 43894 584605 43946 584611
rect 43906 571719 43934 584605
rect 43894 571713 43946 571719
rect 43894 571655 43946 571661
rect 43796 570346 43852 570355
rect 43796 570281 43852 570290
rect 43796 570198 43852 570207
rect 43796 570133 43852 570142
rect 43508 560578 43564 560587
rect 43508 560513 43564 560522
rect 43412 558506 43468 558515
rect 43412 558441 43468 558450
rect 43220 558062 43276 558071
rect 43220 557997 43276 558006
rect 41684 555842 41740 555851
rect 41684 555777 41740 555786
rect 41590 549883 41642 549889
rect 41590 549825 41642 549831
rect 35156 547554 35212 547563
rect 35156 547489 35212 547498
rect 35170 547119 35198 547489
rect 35156 547110 35212 547119
rect 35156 547045 35212 547054
rect 41602 541305 41630 549825
rect 41698 541347 41726 555777
rect 41972 555250 42028 555259
rect 41972 555185 42028 555194
rect 41780 554066 41836 554075
rect 41780 554001 41836 554010
rect 41794 549889 41822 554001
rect 41876 551402 41932 551411
rect 41876 551337 41932 551346
rect 41782 549883 41834 549889
rect 41782 549825 41834 549831
rect 41780 549774 41836 549783
rect 41780 549709 41836 549718
rect 41684 541338 41740 541347
rect 41590 541299 41642 541305
rect 41684 541273 41740 541282
rect 41590 541241 41642 541247
rect 41794 541199 41822 549709
rect 41780 541190 41836 541199
rect 41780 541125 41836 541134
rect 41890 541051 41918 551337
rect 41876 541042 41932 541051
rect 41986 541009 42014 555185
rect 42932 553918 42988 553927
rect 42932 553853 42988 553862
rect 42452 553030 42508 553039
rect 42452 552965 42508 552974
rect 42068 551994 42124 552003
rect 42068 551929 42124 551938
rect 42082 541009 42110 551929
rect 42164 550366 42220 550375
rect 42164 550301 42220 550310
rect 42178 542415 42206 550301
rect 42166 542409 42218 542415
rect 42166 542351 42218 542357
rect 41876 540977 41932 540986
rect 41974 541003 42026 541009
rect 41974 540945 42026 540951
rect 42070 541003 42122 541009
rect 42070 540945 42122 540951
rect 42466 540755 42494 552965
rect 42836 549552 42892 549561
rect 42836 549487 42892 549496
rect 42850 541157 42878 549487
rect 42946 541643 42974 553853
rect 43028 551180 43084 551189
rect 43028 551115 43084 551124
rect 43042 549168 43070 551115
rect 43042 549140 43166 549168
rect 43028 549034 43084 549043
rect 43028 548969 43084 548978
rect 42932 541634 42988 541643
rect 42932 541569 42988 541578
rect 42934 541521 42986 541527
rect 42934 541463 42986 541469
rect 42838 541151 42890 541157
rect 42838 541093 42890 541099
rect 42838 541003 42890 541009
rect 42838 540945 42890 540951
rect 42164 540746 42220 540755
rect 42164 540681 42220 540690
rect 42452 540746 42508 540755
rect 42452 540681 42508 540690
rect 42178 540245 42206 540681
rect 42454 540411 42506 540417
rect 42454 540353 42506 540359
rect 42466 538937 42494 540353
rect 42070 538931 42122 538937
rect 42070 538873 42122 538879
rect 42454 538931 42506 538937
rect 42454 538873 42506 538879
rect 42082 538424 42110 538873
rect 42454 538783 42506 538789
rect 42454 538725 42506 538731
rect 42166 538339 42218 538345
rect 42166 538281 42218 538287
rect 42178 537758 42206 538281
rect 42466 537087 42494 538725
rect 42070 537081 42122 537087
rect 42070 537023 42122 537029
rect 42454 537081 42506 537087
rect 42454 537023 42506 537029
rect 42082 536574 42110 537023
rect 42452 536898 42508 536907
rect 42452 536833 42508 536842
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42082 535390 42110 535765
rect 42166 535083 42218 535089
rect 42166 535025 42218 535031
rect 42178 534724 42206 535025
rect 42166 534491 42218 534497
rect 42166 534433 42218 534439
rect 42178 534058 42206 534433
rect 42070 533751 42122 533757
rect 42070 533693 42122 533699
rect 42082 533540 42110 533693
rect 42356 533346 42412 533355
rect 42356 533281 42412 533290
rect 42164 532754 42220 532763
rect 42164 532689 42220 532698
rect 42178 531875 42206 532689
rect 42164 531866 42220 531875
rect 42164 531801 42220 531810
rect 41780 531718 41836 531727
rect 41780 531653 41836 531662
rect 41794 531616 41822 531653
rect 42370 531389 42398 533281
rect 42166 531383 42218 531389
rect 42166 531325 42218 531331
rect 42358 531383 42410 531389
rect 42358 531325 42410 531331
rect 42178 531024 42206 531325
rect 42356 531274 42412 531283
rect 42356 531209 42412 531218
rect 42166 530939 42218 530945
rect 42166 530881 42218 530887
rect 42178 530401 42206 530881
rect 42070 530273 42122 530279
rect 42070 530215 42122 530221
rect 42082 529766 42110 530215
rect 42166 529459 42218 529465
rect 42166 529401 42218 529407
rect 42178 529205 42206 529401
rect 42166 527831 42218 527837
rect 42166 527773 42218 527779
rect 42178 527365 42206 527773
rect 42370 527245 42398 531209
rect 42466 530945 42494 536833
rect 42454 530939 42506 530945
rect 42454 530881 42506 530887
rect 42454 530791 42506 530797
rect 42454 530733 42506 530739
rect 42466 527837 42494 530733
rect 42850 530279 42878 540945
rect 42946 538345 42974 541463
rect 42934 538339 42986 538345
rect 42934 538281 42986 538287
rect 42934 538191 42986 538197
rect 42934 538133 42986 538139
rect 42946 534497 42974 538133
rect 43042 535829 43070 548969
rect 43138 542508 43166 549140
rect 43138 542480 43262 542508
rect 43126 542409 43178 542415
rect 43126 542351 43178 542357
rect 43030 535823 43082 535829
rect 43030 535765 43082 535771
rect 43028 535714 43084 535723
rect 43028 535649 43084 535658
rect 42934 534491 42986 534497
rect 42934 534433 42986 534439
rect 42932 534382 42988 534391
rect 42932 534317 42988 534326
rect 42946 530797 42974 534317
rect 43042 533757 43070 535649
rect 43138 535089 43166 542351
rect 43234 538789 43262 542480
rect 43318 541151 43370 541157
rect 43318 541093 43370 541099
rect 43222 538783 43274 538789
rect 43222 538725 43274 538731
rect 43330 538197 43358 541093
rect 43318 538191 43370 538197
rect 43318 538133 43370 538139
rect 43126 535083 43178 535089
rect 43126 535025 43178 535031
rect 43126 534935 43178 534941
rect 43126 534877 43178 534883
rect 43030 533751 43082 533757
rect 43030 533693 43082 533699
rect 42934 530791 42986 530797
rect 42934 530733 42986 530739
rect 42932 530682 42988 530691
rect 42932 530617 42988 530626
rect 42838 530273 42890 530279
rect 42838 530215 42890 530221
rect 42838 529977 42890 529983
rect 42838 529919 42890 529925
rect 42454 527831 42506 527837
rect 42454 527773 42506 527779
rect 42070 527239 42122 527245
rect 42070 527181 42122 527187
rect 42358 527239 42410 527245
rect 42358 527181 42410 527187
rect 42082 526732 42110 527181
rect 42166 526499 42218 526505
rect 42166 526441 42218 526447
rect 42178 526066 42206 526441
rect 42850 524211 42878 529919
rect 42946 526505 42974 530617
rect 43138 529465 43166 534877
rect 43126 529459 43178 529465
rect 43126 529401 43178 529407
rect 42934 526499 42986 526505
rect 42934 526441 42986 526447
rect 42358 524205 42410 524211
rect 42358 524147 42410 524153
rect 42838 524205 42890 524211
rect 42838 524147 42890 524153
rect 42370 431383 42398 524147
rect 42838 432297 42890 432303
rect 42836 432262 42838 432271
rect 42890 432262 42892 432271
rect 42836 432197 42892 432206
rect 42838 431779 42890 431785
rect 42836 431744 42838 431753
rect 42890 431744 42892 431753
rect 42836 431679 42892 431688
rect 42356 431374 42412 431383
rect 42356 431309 42412 431318
rect 43220 430634 43276 430643
rect 43220 430569 43276 430578
rect 42838 429633 42890 429639
rect 42836 429598 42838 429607
rect 42890 429598 42892 429607
rect 42836 429533 42892 429542
rect 42836 427970 42892 427979
rect 42836 427905 42892 427914
rect 41876 425454 41932 425463
rect 41876 425389 41932 425398
rect 40244 423382 40300 423391
rect 40244 423317 40300 423326
rect 39956 422790 40012 422799
rect 39956 422725 40012 422734
rect 35156 419978 35212 419987
rect 35156 419913 35212 419922
rect 35170 419543 35198 419913
rect 35156 419534 35212 419543
rect 35156 419469 35212 419478
rect 39970 414765 39998 422725
rect 40052 422198 40108 422207
rect 40052 422133 40108 422142
rect 40066 415727 40094 422133
rect 40148 421606 40204 421615
rect 40148 421541 40204 421550
rect 40054 415721 40106 415727
rect 40054 415663 40106 415669
rect 40162 415431 40190 421541
rect 40258 416319 40286 423317
rect 40246 416313 40298 416319
rect 40246 416255 40298 416261
rect 40150 415425 40202 415431
rect 40150 415367 40202 415373
rect 39958 414759 40010 414765
rect 39958 414701 40010 414707
rect 41890 413433 41918 425389
rect 42356 420570 42412 420579
rect 42356 420505 42412 420514
rect 42370 419543 42398 420505
rect 42356 419534 42412 419543
rect 42356 419469 42412 419478
rect 42370 417651 42398 419469
rect 42358 417645 42410 417651
rect 42358 417587 42410 417593
rect 42742 416313 42794 416319
rect 42742 416255 42794 416261
rect 41878 413427 41930 413433
rect 41878 413369 41930 413375
rect 41878 413205 41930 413211
rect 41878 413147 41930 413153
rect 41890 412624 41918 413147
rect 42166 411355 42218 411361
rect 42166 411297 42218 411303
rect 42178 410805 42206 411297
rect 42070 410541 42122 410547
rect 42070 410483 42122 410489
rect 42082 410182 42110 410483
rect 42754 409511 42782 416255
rect 42850 411361 42878 427905
rect 42932 421458 42988 421467
rect 42932 421393 42988 421402
rect 42838 411355 42890 411361
rect 42838 411297 42890 411303
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42742 409505 42794 409511
rect 42742 409447 42794 409453
rect 42178 408965 42206 409447
rect 42946 409308 42974 421393
rect 43126 415721 43178 415727
rect 43126 415663 43178 415669
rect 43030 415425 43082 415431
rect 43030 415367 43082 415373
rect 42754 409280 42974 409308
rect 43042 409289 43070 415367
rect 43030 409283 43082 409289
rect 42754 408253 42782 409280
rect 43030 409225 43082 409231
rect 42838 409209 42890 409215
rect 42838 409151 42890 409157
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42742 408247 42794 408253
rect 42742 408189 42794 408195
rect 42178 407769 42206 408189
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42850 407069 42878 409151
rect 43138 409141 43166 415663
rect 42934 409135 42986 409141
rect 42934 409077 42986 409083
rect 43126 409135 43178 409141
rect 43126 409077 43178 409083
rect 42166 407063 42218 407069
rect 42166 407005 42218 407011
rect 42838 407063 42890 407069
rect 42838 407005 42890 407011
rect 42178 406482 42206 407005
rect 42946 406940 42974 409077
rect 43126 408987 43178 408993
rect 43126 408929 43178 408935
rect 43138 407513 43166 408929
rect 43126 407507 43178 407513
rect 43126 407449 43178 407455
rect 42754 406912 42974 406940
rect 41780 406066 41836 406075
rect 41780 406001 41836 406010
rect 41794 405929 41822 406001
rect 41876 405178 41932 405187
rect 41876 405113 41932 405122
rect 41890 404632 41918 405113
rect 41780 404438 41836 404447
rect 41780 404373 41836 404382
rect 41794 403997 41822 404373
rect 42754 403739 42782 406912
rect 42166 403733 42218 403739
rect 42166 403675 42218 403681
rect 42742 403733 42794 403739
rect 42742 403675 42794 403681
rect 42178 403448 42206 403675
rect 42164 403106 42220 403115
rect 42164 403041 42220 403050
rect 42178 402782 42206 403041
rect 42164 402662 42220 402671
rect 42164 402597 42220 402606
rect 42178 402157 42206 402597
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42358 389377 42410 389383
rect 42356 389342 42358 389351
rect 42410 389342 42412 389351
rect 42356 389277 42412 389286
rect 42358 388785 42410 388791
rect 42356 388750 42358 388759
rect 42410 388750 42412 388759
rect 42356 388685 42412 388694
rect 42742 388045 42794 388051
rect 42740 388010 42742 388019
rect 42794 388010 42796 388019
rect 42740 387945 42796 387954
rect 43234 387131 43262 430569
rect 43426 430199 43454 558441
rect 43412 430190 43468 430199
rect 43412 430125 43468 430134
rect 43522 429015 43550 560513
rect 43604 556878 43660 556887
rect 43810 556864 43838 570133
rect 43660 556836 43838 556864
rect 43604 556813 43660 556822
rect 43618 429639 43646 556813
rect 43702 541299 43754 541305
rect 43702 541241 43754 541247
rect 43714 534941 43742 541241
rect 43702 534935 43754 534941
rect 43702 534877 43754 534883
rect 43606 429633 43658 429639
rect 43606 429575 43658 429581
rect 43508 429006 43564 429015
rect 43508 428941 43564 428950
rect 43414 414759 43466 414765
rect 43414 414701 43466 414707
rect 43426 408993 43454 414701
rect 43414 408987 43466 408993
rect 43414 408929 43466 408935
rect 43316 387270 43372 387279
rect 43316 387205 43372 387214
rect 43220 387122 43276 387131
rect 43220 387057 43276 387066
rect 42164 384458 42220 384467
rect 42164 384393 42220 384402
rect 40052 381202 40108 381211
rect 40052 381137 40108 381146
rect 39956 380166 40012 380175
rect 39956 380101 40012 380110
rect 39860 378982 39916 378991
rect 39860 378917 39916 378926
rect 35156 376762 35212 376771
rect 35156 376697 35212 376706
rect 35170 376327 35198 376697
rect 35156 376318 35212 376327
rect 35156 376253 35212 376262
rect 39874 371623 39902 378917
rect 39970 372437 39998 380101
rect 40066 375143 40094 381137
rect 40148 380610 40204 380619
rect 40148 380545 40204 380554
rect 40052 375134 40108 375143
rect 40052 375069 40108 375078
rect 40162 372923 40190 380545
rect 40244 378390 40300 378399
rect 40244 378325 40300 378334
rect 40258 373399 40286 378325
rect 40246 373393 40298 373399
rect 40246 373335 40298 373341
rect 40148 372914 40204 372923
rect 40148 372849 40204 372858
rect 39958 372431 40010 372437
rect 39958 372373 40010 372379
rect 39862 371617 39914 371623
rect 39862 371559 39914 371565
rect 42178 370217 42206 384393
rect 42356 382238 42412 382247
rect 42356 382173 42412 382182
rect 42166 370211 42218 370217
rect 42166 370153 42218 370159
rect 42370 369995 42398 382173
rect 42548 379574 42604 379583
rect 42548 379509 42604 379518
rect 42562 372308 42590 379509
rect 43124 378242 43180 378251
rect 43124 378177 43180 378186
rect 42644 377650 42700 377659
rect 42644 377585 42700 377594
rect 42658 376623 42686 377585
rect 42644 376614 42700 376623
rect 42644 376549 42646 376558
rect 42698 376549 42700 376558
rect 42646 376517 42698 376523
rect 43030 372431 43082 372437
rect 43030 372373 43082 372379
rect 42562 372280 42686 372308
rect 42166 369989 42218 369995
rect 42166 369931 42218 369937
rect 42358 369989 42410 369995
rect 42358 369931 42410 369937
rect 42178 369445 42206 369931
rect 42550 368879 42602 368885
rect 42550 368821 42602 368827
rect 42562 368145 42590 368821
rect 42070 368139 42122 368145
rect 42070 368081 42122 368087
rect 42550 368139 42602 368145
rect 42550 368081 42602 368087
rect 42082 367632 42110 368081
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42070 366215 42122 366221
rect 42070 366157 42122 366163
rect 42082 365782 42110 366157
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42178 364569 42206 364973
rect 42658 364445 42686 372280
rect 42934 367621 42986 367627
rect 42934 367563 42986 367569
rect 42070 364439 42122 364445
rect 42070 364381 42122 364387
rect 42646 364439 42698 364445
rect 42646 364381 42698 364387
rect 42082 363932 42110 364381
rect 42166 363847 42218 363853
rect 42166 363789 42218 363795
rect 42178 363266 42206 363789
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 42082 360935 42110 361416
rect 42068 360926 42124 360935
rect 42068 360861 42124 360870
rect 41986 360639 42014 360824
rect 42946 360671 42974 367563
rect 43042 366221 43070 372373
rect 43030 366215 43082 366221
rect 43030 366157 43082 366163
rect 43138 365037 43166 378177
rect 43330 378080 43358 387205
rect 43234 378052 43358 378080
rect 43126 365031 43178 365037
rect 43126 364973 43178 364979
rect 42166 360665 42218 360671
rect 41972 360630 42028 360639
rect 42166 360607 42218 360613
rect 42934 360665 42986 360671
rect 42934 360607 42986 360613
rect 41972 360565 42028 360574
rect 42178 360232 42206 360607
rect 42164 359890 42220 359899
rect 42164 359825 42220 359834
rect 42178 359601 42206 359825
rect 42068 359446 42124 359455
rect 42068 359381 42124 359390
rect 42082 358974 42110 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41780 356930 41836 356939
rect 41780 356865 41836 356874
rect 41794 356565 41822 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42454 346161 42506 346167
rect 42452 346126 42454 346135
rect 42506 346126 42508 346135
rect 42452 346061 42508 346070
rect 42454 345569 42506 345575
rect 42452 345534 42454 345543
rect 42506 345534 42508 345543
rect 42452 345469 42508 345478
rect 42934 344829 42986 344835
rect 42932 344794 42934 344803
rect 42986 344794 42988 344803
rect 42932 344729 42988 344738
rect 43124 344054 43180 344063
rect 43124 343989 43180 343998
rect 43138 343596 43166 343989
rect 43234 343767 43262 378052
rect 43414 373393 43466 373399
rect 43414 373335 43466 373341
rect 43318 371617 43370 371623
rect 43318 371559 43370 371565
rect 43330 367627 43358 371559
rect 43318 367621 43370 367627
rect 43318 367563 43370 367569
rect 43426 363853 43454 373335
rect 43414 363847 43466 363853
rect 43414 363789 43466 363795
rect 43220 343758 43276 343767
rect 43220 343693 43276 343702
rect 43138 343568 43262 343596
rect 42932 341538 42988 341547
rect 42932 341473 42988 341482
rect 41876 339022 41932 339031
rect 41876 338957 41932 338966
rect 40148 337394 40204 337403
rect 40148 337329 40204 337338
rect 39956 336950 40012 336959
rect 39956 336885 40012 336894
rect 39860 335174 39916 335183
rect 39860 335109 39916 335118
rect 35156 333546 35212 333555
rect 35156 333481 35212 333490
rect 35170 333111 35198 333481
rect 35156 333102 35212 333111
rect 35156 333037 35212 333046
rect 39874 329813 39902 335109
rect 39862 329807 39914 329813
rect 39862 329749 39914 329755
rect 39970 329369 39998 336885
rect 40052 336358 40108 336367
rect 40052 336293 40108 336302
rect 40066 329517 40094 336293
rect 40162 329855 40190 337329
rect 40244 335766 40300 335775
rect 40244 335701 40300 335710
rect 40148 329846 40204 329855
rect 40148 329781 40204 329790
rect 40054 329511 40106 329517
rect 40054 329453 40106 329459
rect 39958 329363 40010 329369
rect 39958 329305 40010 329311
rect 40258 329221 40286 335701
rect 40246 329215 40298 329221
rect 40246 329157 40298 329163
rect 41890 327075 41918 338957
rect 42836 333398 42892 333407
rect 42836 333333 42838 333342
rect 42890 333333 42892 333342
rect 42838 333301 42890 333307
rect 42838 329511 42890 329517
rect 42838 329453 42890 329459
rect 42454 329363 42506 329369
rect 42454 329305 42506 329311
rect 42358 329215 42410 329221
rect 42358 329157 42410 329163
rect 41878 327069 41930 327075
rect 41878 327011 41930 327017
rect 41878 326773 41930 326779
rect 41878 326715 41930 326721
rect 41890 326266 41918 326715
rect 42370 326599 42398 329157
rect 42356 326590 42412 326599
rect 42356 326525 42412 326534
rect 42466 325669 42494 329305
rect 42454 325663 42506 325669
rect 42454 325605 42506 325611
rect 42742 325367 42794 325373
rect 42742 325309 42794 325315
rect 42070 324923 42122 324929
rect 42070 324865 42122 324871
rect 42082 324416 42110 324865
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42754 323153 42782 325309
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42742 323147 42794 323153
rect 42742 323089 42794 323095
rect 42178 322566 42206 323089
rect 42850 323005 42878 329453
rect 42946 324929 42974 341473
rect 43028 335026 43084 335035
rect 43028 334961 43084 334970
rect 42934 324923 42986 324929
rect 42934 324865 42986 324871
rect 42838 322999 42890 323005
rect 42838 322941 42890 322947
rect 42454 322777 42506 322783
rect 42454 322719 42506 322725
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42082 321382 42110 321757
rect 42466 321081 42494 322719
rect 43042 321821 43070 334961
rect 43126 329807 43178 329813
rect 43126 329749 43178 329755
rect 43030 321815 43082 321821
rect 43030 321757 43082 321763
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42454 321075 42506 321081
rect 42454 321017 42506 321023
rect 42178 320716 42206 321017
rect 42452 320966 42508 320975
rect 42452 320901 42508 320910
rect 42166 320631 42218 320637
rect 42166 320573 42218 320579
rect 42178 320081 42206 320573
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 41972 318746 42028 318755
rect 41972 318681 42028 318690
rect 41986 318241 42014 318681
rect 41972 317858 42028 317867
rect 41972 317793 42028 317802
rect 41986 317608 42014 317793
rect 42466 317529 42494 320901
rect 43138 320637 43166 329749
rect 43126 320631 43178 320637
rect 43126 320573 43178 320579
rect 42166 317523 42218 317529
rect 42166 317465 42218 317471
rect 42454 317523 42506 317529
rect 42454 317465 42506 317471
rect 42178 317045 42206 317465
rect 42068 316674 42124 316683
rect 42068 316609 42124 316618
rect 42082 316424 42110 316609
rect 42068 316082 42124 316091
rect 42068 316017 42124 316026
rect 42082 315758 42110 316017
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41876 313714 41932 313723
rect 41876 313649 41932 313658
rect 41890 313390 41918 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42550 302945 42602 302951
rect 42548 302910 42550 302919
rect 42602 302910 42604 302919
rect 42548 302845 42604 302854
rect 42550 302353 42602 302359
rect 42548 302318 42550 302327
rect 42602 302318 42604 302327
rect 42548 302253 42604 302262
rect 42550 301909 42602 301915
rect 42548 301874 42550 301883
rect 42602 301874 42604 301883
rect 42548 301809 42604 301818
rect 43234 300551 43262 343568
rect 43316 300986 43372 300995
rect 43316 300921 43372 300930
rect 43220 300542 43276 300551
rect 43220 300477 43276 300486
rect 41204 298026 41260 298035
rect 41204 297961 41260 297970
rect 40244 294178 40300 294187
rect 40244 294113 40300 294122
rect 40148 293734 40204 293743
rect 40148 293669 40204 293678
rect 39860 292550 39916 292559
rect 39860 292485 39916 292494
rect 35156 290478 35212 290487
rect 35156 290413 35212 290422
rect 35170 289895 35198 290413
rect 35156 289886 35212 289895
rect 35156 289821 35212 289830
rect 39874 285487 39902 292485
rect 40052 292106 40108 292115
rect 40052 292041 40108 292050
rect 39862 285481 39914 285487
rect 39862 285423 39914 285429
rect 40066 285339 40094 292041
rect 40054 285333 40106 285339
rect 40054 285275 40106 285281
rect 40162 285191 40190 293669
rect 40150 285185 40202 285191
rect 40258 285159 40286 294113
rect 40150 285127 40202 285133
rect 40244 285150 40300 285159
rect 40244 285085 40300 285094
rect 41218 284155 41246 297961
rect 41972 295806 42028 295815
rect 41972 295741 42028 295750
rect 41206 284149 41258 284155
rect 41206 284091 41258 284097
rect 41986 283859 42014 295741
rect 42932 291810 42988 291819
rect 42932 291745 42988 291754
rect 42548 289886 42604 289895
rect 42548 289821 42550 289830
rect 42602 289821 42604 289830
rect 42550 289789 42602 289795
rect 41974 283853 42026 283859
rect 41974 283795 42026 283801
rect 42454 283631 42506 283637
rect 42454 283573 42506 283579
rect 41974 283557 42026 283563
rect 41974 283499 42026 283505
rect 41986 283050 42014 283499
rect 42466 281787 42494 283573
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42454 281781 42506 281787
rect 42454 281723 42506 281729
rect 42178 281200 42206 281723
rect 42166 281115 42218 281121
rect 42166 281057 42218 281063
rect 42178 280534 42206 281057
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42946 278605 42974 291745
rect 43126 285481 43178 285487
rect 43178 285429 43262 285432
rect 43126 285423 43262 285429
rect 43138 285404 43262 285423
rect 43126 285333 43178 285339
rect 43126 285275 43178 285281
rect 43030 285185 43082 285191
rect 43030 285127 43082 285133
rect 43042 279937 43070 285127
rect 43138 279937 43166 285275
rect 43030 279931 43082 279937
rect 43030 279873 43082 279879
rect 43126 279931 43178 279937
rect 43126 279873 43178 279879
rect 43234 279808 43262 285404
rect 43042 279780 43262 279808
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42934 278599 42986 278605
rect 42934 278541 42986 278547
rect 42178 278166 42206 278541
rect 42164 278046 42220 278055
rect 42164 277981 42220 277990
rect 42178 277500 42206 277981
rect 42070 277267 42122 277273
rect 42070 277209 42122 277215
rect 42082 276908 42110 277209
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 41972 275530 42028 275539
rect 41972 275465 42028 275474
rect 41986 275058 42014 275465
rect 42164 274790 42220 274799
rect 42164 274725 42220 274734
rect 42178 274392 42206 274725
rect 43042 274313 43070 279780
rect 43126 279709 43178 279715
rect 43126 279651 43178 279657
rect 43138 277273 43166 279651
rect 43330 277884 43358 300921
rect 43234 277856 43358 277884
rect 43126 277267 43178 277273
rect 43126 277209 43178 277215
rect 43124 274790 43180 274799
rect 43124 274725 43180 274734
rect 42166 274307 42218 274313
rect 42166 274249 42218 274255
rect 43030 274307 43082 274313
rect 43030 274249 43082 274255
rect 42178 273845 42206 274249
rect 41780 273606 41836 273615
rect 41780 273541 41836 273550
rect 41794 273208 41822 273541
rect 42068 273014 42124 273023
rect 42068 272949 42124 272958
rect 42082 272542 42110 272949
rect 41780 272274 41836 272283
rect 41780 272209 41836 272218
rect 41794 272024 41822 272209
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 42454 259729 42506 259735
rect 42452 259694 42454 259703
rect 42506 259694 42508 259703
rect 42452 259629 42508 259638
rect 42838 258989 42890 258995
rect 42836 258954 42838 258963
rect 42890 258954 42892 258963
rect 42836 258889 42892 258898
rect 42454 258693 42506 258699
rect 42452 258658 42454 258667
rect 42506 258658 42508 258667
rect 42452 258593 42508 258602
rect 42454 257879 42506 257885
rect 42454 257821 42506 257827
rect 42466 257483 42494 257821
rect 42452 257474 42508 257483
rect 42452 257409 42508 257418
rect 42164 255994 42220 256003
rect 42164 255929 42220 255938
rect 41876 252590 41932 252599
rect 41876 252525 41932 252534
rect 40148 250962 40204 250971
rect 40148 250897 40204 250906
rect 39956 249926 40012 249935
rect 39956 249861 40012 249870
rect 39860 249334 39916 249343
rect 39860 249269 39916 249278
rect 35156 247262 35212 247271
rect 35156 247197 35212 247206
rect 35170 246827 35198 247197
rect 35156 246818 35212 246827
rect 35156 246753 35212 246762
rect 39874 242123 39902 249269
rect 39970 242271 39998 249861
rect 40052 248890 40108 248899
rect 40052 248825 40108 248834
rect 39958 242265 40010 242271
rect 39958 242207 40010 242213
rect 39862 242117 39914 242123
rect 39862 242059 39914 242065
rect 40066 242049 40094 248825
rect 40162 244903 40190 250897
rect 40244 250518 40300 250527
rect 40244 250453 40300 250462
rect 40148 244894 40204 244903
rect 40148 244829 40204 244838
rect 40054 242043 40106 242049
rect 40054 241985 40106 241991
rect 40258 241975 40286 250453
rect 40246 241969 40298 241975
rect 40246 241911 40298 241917
rect 41890 240643 41918 252525
rect 42068 248298 42124 248307
rect 42068 248233 42124 248242
rect 42082 242091 42110 248233
rect 42178 242535 42206 255929
rect 43028 255106 43084 255115
rect 43028 255041 43084 255050
rect 42452 246818 42508 246827
rect 42452 246753 42508 246762
rect 42466 245083 42494 246753
rect 42454 245077 42506 245083
rect 42454 245019 42506 245025
rect 42164 242526 42220 242535
rect 42164 242461 42220 242470
rect 42550 242265 42602 242271
rect 42602 242213 42686 242216
rect 42550 242207 42686 242213
rect 42562 242188 42686 242207
rect 42358 242117 42410 242123
rect 42068 242082 42124 242091
rect 42358 242059 42410 242065
rect 42452 242082 42508 242091
rect 42068 242017 42124 242026
rect 41878 240637 41930 240643
rect 41878 240579 41930 240585
rect 41878 240415 41930 240421
rect 41878 240357 41930 240363
rect 41890 239834 41918 240357
rect 42370 240125 42398 242059
rect 42452 242017 42508 242026
rect 42550 242043 42602 242049
rect 42358 240119 42410 240125
rect 42358 240061 42410 240067
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42178 237984 42206 238507
rect 42466 238423 42494 242017
rect 42550 241985 42602 241991
rect 42454 238417 42506 238423
rect 42562 238391 42590 241985
rect 42454 238359 42506 238365
rect 42548 238382 42604 238391
rect 42548 238317 42604 238326
rect 42658 238220 42686 242188
rect 43042 238571 43070 255041
rect 43138 243867 43166 274725
rect 43234 257885 43262 277856
rect 43222 257879 43274 257885
rect 43222 257821 43274 257827
rect 43220 257622 43276 257631
rect 43220 257557 43276 257566
rect 43124 243858 43180 243867
rect 43124 243793 43180 243802
rect 43126 241969 43178 241975
rect 43126 241911 43178 241917
rect 43030 238565 43082 238571
rect 43030 238507 43082 238513
rect 43030 238417 43082 238423
rect 43030 238359 43082 238365
rect 42466 238192 42686 238220
rect 42466 237961 42494 238192
rect 42934 237973 42986 237979
rect 42466 237933 42590 237961
rect 42166 237899 42218 237905
rect 42166 237841 42218 237847
rect 42178 237361 42206 237841
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42178 236165 42206 236657
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42454 234865 42506 234871
rect 42562 234853 42590 237933
rect 42934 237915 42986 237921
rect 42506 234825 42590 234853
rect 42454 234807 42506 234813
rect 42178 234325 42206 234807
rect 42068 234090 42124 234099
rect 42068 234025 42124 234034
rect 42082 233692 42110 234025
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41794 231731 41822 231842
rect 41780 231722 41836 231731
rect 41780 231657 41836 231666
rect 41986 231139 42014 231176
rect 41972 231130 42028 231139
rect 42946 231097 42974 237915
rect 43042 235463 43070 238359
rect 43138 236721 43166 241911
rect 43126 236715 43178 236721
rect 43126 236657 43178 236663
rect 43030 235457 43082 235463
rect 43030 235399 43082 235405
rect 41972 231065 42028 231074
rect 42070 231091 42122 231097
rect 42070 231033 42122 231039
rect 42934 231091 42986 231097
rect 42934 231033 42986 231039
rect 42082 230658 42110 231033
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227282 41836 227291
rect 41780 227217 41836 227226
rect 41794 226958 41822 227217
rect 41780 226690 41836 226699
rect 41780 226625 41836 226634
rect 41794 226321 41822 226625
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42454 216513 42506 216519
rect 42452 216478 42454 216487
rect 42506 216478 42508 216487
rect 42452 216413 42508 216422
rect 42838 215773 42890 215779
rect 42836 215738 42838 215747
rect 42890 215738 42892 215747
rect 42836 215673 42892 215682
rect 42838 215255 42890 215261
rect 42836 215220 42838 215229
rect 42890 215220 42892 215229
rect 42836 215155 42892 215164
rect 43234 214119 43262 257557
rect 44578 246235 44606 806489
rect 44662 800669 44714 800675
rect 44662 800611 44714 800617
rect 44674 324189 44702 800611
rect 44770 673913 44798 988127
rect 44854 988111 44906 988117
rect 44854 988053 44906 988059
rect 44866 717129 44894 988053
rect 44950 988037 45002 988043
rect 44950 987979 45002 987985
rect 44962 757533 44990 987979
rect 45046 987963 45098 987969
rect 45046 987905 45098 987911
rect 45058 797345 45086 987905
rect 47542 986705 47594 986711
rect 47542 986647 47594 986653
rect 47446 986631 47498 986637
rect 47446 986573 47498 986579
rect 47458 941687 47486 986573
rect 47554 942755 47582 986647
rect 47542 942749 47594 942755
rect 47542 942691 47594 942697
rect 47444 941678 47500 941687
rect 47444 941613 47500 941622
rect 47446 915887 47498 915893
rect 47446 915829 47498 915835
rect 45046 797339 45098 797345
rect 45046 797281 45098 797287
rect 45046 786313 45098 786319
rect 45046 786255 45098 786261
rect 44950 757527 45002 757533
rect 44950 757469 45002 757475
rect 45058 731855 45086 786255
rect 45046 731849 45098 731855
rect 45046 731791 45098 731797
rect 44854 717123 44906 717129
rect 44854 717065 44906 717071
rect 44950 714311 45002 714317
rect 44950 714253 45002 714259
rect 44962 689527 44990 714253
rect 44950 689521 45002 689527
rect 44950 689463 45002 689469
rect 44758 673907 44810 673913
rect 44758 673849 44810 673855
rect 44854 671095 44906 671101
rect 44854 671037 44906 671043
rect 44866 647791 44894 671037
rect 44854 647785 44906 647791
rect 44854 647727 44906 647733
rect 44758 627879 44810 627885
rect 44758 627821 44810 627827
rect 44662 324183 44714 324189
rect 44662 324125 44714 324131
rect 44662 313971 44714 313977
rect 44662 313913 44714 313919
rect 44564 246226 44620 246235
rect 44564 246161 44620 246170
rect 43414 242783 43466 242789
rect 43414 242725 43466 242731
rect 43318 240119 43370 240125
rect 43318 240061 43370 240067
rect 43330 237979 43358 240061
rect 43318 237973 43370 237979
rect 43318 237915 43370 237921
rect 43318 237825 43370 237831
rect 43318 237767 43370 237773
rect 43220 214110 43276 214119
rect 43220 214045 43276 214054
rect 43330 213083 43358 237767
rect 43426 213675 43454 242725
rect 43508 242526 43564 242535
rect 43508 242461 43564 242470
rect 43522 237831 43550 242461
rect 43510 237825 43562 237831
rect 43510 237767 43562 237773
rect 44674 215261 44702 313913
rect 44662 215255 44714 215261
rect 44662 215197 44714 215203
rect 43412 213666 43468 213675
rect 43412 213601 43468 213610
rect 43316 213074 43372 213083
rect 43316 213009 43372 213018
rect 42452 211742 42508 211751
rect 42508 211700 42590 211728
rect 42452 211677 42508 211686
rect 42068 209522 42124 209531
rect 42068 209457 42124 209466
rect 40052 207302 40108 207311
rect 40052 207237 40108 207246
rect 39956 206118 40012 206127
rect 39956 206053 40012 206062
rect 35156 204046 35212 204055
rect 35156 203981 35212 203990
rect 35170 203611 35198 203981
rect 35156 203602 35212 203611
rect 35156 203537 35212 203546
rect 39970 198833 39998 206053
rect 40066 200165 40094 207237
rect 40148 206710 40204 206719
rect 40148 206645 40204 206654
rect 40054 200159 40106 200165
rect 40054 200101 40106 200107
rect 40162 199055 40190 206645
rect 40244 205674 40300 205683
rect 40244 205609 40300 205618
rect 40150 199049 40202 199055
rect 40150 198991 40202 198997
rect 39958 198827 40010 198833
rect 39958 198769 40010 198775
rect 40258 198759 40286 205609
rect 40246 198753 40298 198759
rect 40246 198695 40298 198701
rect 41014 198753 41066 198759
rect 41014 198695 41066 198701
rect 41026 197811 41054 198695
rect 41112 197811 41121 197827
rect 41026 197783 41121 197811
rect 41112 197767 41121 197783
rect 41181 197767 41190 197827
rect 42082 197427 42110 209457
rect 42452 204490 42508 204499
rect 42452 204425 42454 204434
rect 42506 204425 42508 204434
rect 42454 204393 42506 204399
rect 42466 204055 42494 204393
rect 42452 204046 42508 204055
rect 42452 203981 42508 203990
rect 42358 199049 42410 199055
rect 42358 198991 42410 198997
rect 42070 197421 42122 197427
rect 42070 197363 42122 197369
rect 42070 197199 42122 197205
rect 42070 197141 42122 197147
rect 42082 196618 42110 197141
rect 42370 196909 42398 198991
rect 42358 196903 42410 196909
rect 42358 196845 42410 196851
rect 42562 195892 42590 211700
rect 43028 205378 43084 205387
rect 43028 205313 43084 205322
rect 42466 195864 42590 195892
rect 42466 195651 42494 195864
rect 42454 195645 42506 195651
rect 42454 195587 42506 195593
rect 42166 195349 42218 195355
rect 42166 195291 42218 195297
rect 42178 194805 42206 195291
rect 42934 194831 42986 194837
rect 42934 194773 42986 194779
rect 42838 194757 42890 194763
rect 42838 194699 42890 194705
rect 42070 194535 42122 194541
rect 42070 194477 42122 194483
rect 42082 194176 42110 194477
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42178 191769 42206 192183
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42082 191142 42110 191443
rect 42164 191022 42220 191031
rect 42164 190957 42220 190966
rect 42178 190476 42206 190957
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 41780 189098 41836 189107
rect 41780 189033 41836 189042
rect 41794 188626 41822 189033
rect 41972 188358 42028 188367
rect 41972 188293 42028 188302
rect 41986 187997 42014 188293
rect 42850 187733 42878 194699
rect 42946 191507 42974 194773
rect 43042 192247 43070 205313
rect 43126 200159 43178 200165
rect 43126 200101 43178 200107
rect 43138 193505 43166 200101
rect 43318 198827 43370 198833
rect 43318 198769 43370 198775
rect 43222 196903 43274 196909
rect 43222 196845 43274 196851
rect 43234 194837 43262 196845
rect 43222 194831 43274 194837
rect 43222 194773 43274 194779
rect 43330 194763 43358 198769
rect 43318 194757 43370 194763
rect 43318 194699 43370 194705
rect 44770 194541 44798 627821
rect 46006 601979 46058 601985
rect 46006 601921 46058 601927
rect 46018 584965 46046 601921
rect 46006 584959 46058 584965
rect 46006 584901 46058 584907
rect 44852 547406 44908 547415
rect 44852 547341 44908 547350
rect 44866 246341 44894 547341
rect 44950 472405 45002 472411
rect 44950 472347 45002 472353
rect 44962 389383 44990 472347
rect 47458 410547 47486 915829
rect 47542 815099 47594 815105
rect 47542 815041 47594 815047
rect 47554 775367 47582 815041
rect 47542 775361 47594 775367
rect 47542 775303 47594 775309
rect 47542 728667 47594 728673
rect 47542 728609 47594 728615
rect 47554 688491 47582 728609
rect 47542 688485 47594 688491
rect 47542 688427 47594 688433
rect 47542 685525 47594 685531
rect 47542 685467 47594 685473
rect 47446 410541 47498 410547
rect 47446 410483 47498 410489
rect 45046 400403 45098 400409
rect 45046 400345 45098 400351
rect 44950 389377 45002 389383
rect 44950 389319 45002 389325
rect 44950 376575 45002 376581
rect 44950 376517 45002 376523
rect 44854 246335 44906 246341
rect 44854 246277 44906 246283
rect 44962 246267 44990 376517
rect 45058 301915 45086 400345
rect 47446 357187 47498 357193
rect 47446 357129 47498 357135
rect 45046 301909 45098 301915
rect 45046 301851 45098 301857
rect 45142 299615 45194 299621
rect 45142 299557 45194 299563
rect 45046 285185 45098 285191
rect 45046 285127 45098 285133
rect 44950 246261 45002 246267
rect 44950 246203 45002 246209
rect 45058 215779 45086 285127
rect 45154 216519 45182 299557
rect 47458 258699 47486 357129
rect 47446 258693 47498 258699
rect 47446 258635 47498 258641
rect 46196 256734 46252 256743
rect 46196 256669 46252 256678
rect 46210 246119 46238 256669
rect 46198 246113 46250 246119
rect 46198 246055 46250 246061
rect 46210 242789 46238 246055
rect 46198 242783 46250 242789
rect 46198 242725 46250 242731
rect 47554 237905 47582 685467
rect 47650 627959 47678 988201
rect 48886 944303 48938 944309
rect 48886 944245 48938 944251
rect 48898 930545 48926 944245
rect 48886 930539 48938 930545
rect 48886 930481 48938 930487
rect 50326 858315 50378 858321
rect 50326 858257 50378 858263
rect 47638 627953 47690 627959
rect 47638 627895 47690 627901
rect 50230 559059 50282 559065
rect 50230 559001 50282 559007
rect 50242 544561 50270 559001
rect 50230 544555 50282 544561
rect 50230 544497 50282 544503
rect 47830 457975 47882 457981
rect 47830 457917 47882 457923
rect 47638 429189 47690 429195
rect 47638 429131 47690 429137
rect 47650 346167 47678 429131
rect 47842 388791 47870 457917
rect 47830 388785 47882 388791
rect 47830 388727 47882 388733
rect 47734 385973 47786 385979
rect 47734 385915 47786 385921
rect 47638 346161 47690 346167
rect 47638 346103 47690 346109
rect 47638 333359 47690 333365
rect 47638 333301 47690 333307
rect 47650 249153 47678 333301
rect 47746 302951 47774 385915
rect 50338 367405 50366 858257
rect 50434 584151 50462 988275
rect 59444 975422 59500 975431
rect 59444 975357 59500 975366
rect 59458 973539 59486 975357
rect 53686 973533 53738 973539
rect 53686 973475 53738 973481
rect 59446 973533 59498 973539
rect 59446 973475 59498 973481
rect 53206 932167 53258 932173
rect 53206 932109 53258 932115
rect 50518 887175 50570 887181
rect 50518 887117 50570 887123
rect 50530 819175 50558 887117
rect 50614 829529 50666 829535
rect 50614 829471 50666 829477
rect 50518 819169 50570 819175
rect 50518 819111 50570 819117
rect 50626 776107 50654 829471
rect 50614 776101 50666 776107
rect 50614 776043 50666 776049
rect 50422 584145 50474 584151
rect 50422 584087 50474 584093
rect 50518 515547 50570 515553
rect 50518 515489 50570 515495
rect 50422 486761 50474 486767
rect 50422 486703 50474 486709
rect 50434 388051 50462 486703
rect 50530 432303 50558 515489
rect 50518 432297 50570 432303
rect 50518 432239 50570 432245
rect 50518 414759 50570 414765
rect 50518 414701 50570 414707
rect 50422 388045 50474 388051
rect 50422 387987 50474 387993
rect 50422 371617 50474 371623
rect 50422 371559 50474 371565
rect 50326 367399 50378 367405
rect 50326 367341 50378 367347
rect 50326 328401 50378 328407
rect 50326 328343 50378 328349
rect 47734 302945 47786 302951
rect 47734 302887 47786 302893
rect 47734 289847 47786 289853
rect 47734 289789 47786 289795
rect 47638 249147 47690 249153
rect 47638 249089 47690 249095
rect 47746 246415 47774 289789
rect 50338 258995 50366 328343
rect 50434 302359 50462 371559
rect 50530 345575 50558 414701
rect 50518 345569 50570 345575
rect 50518 345511 50570 345517
rect 50422 302353 50474 302359
rect 50422 302295 50474 302301
rect 50326 258989 50378 258995
rect 50326 258931 50378 258937
rect 53218 246563 53246 932109
rect 53302 901531 53354 901537
rect 53302 901473 53354 901479
rect 53314 818139 53342 901473
rect 53398 843885 53450 843891
rect 53398 843827 53450 843833
rect 53302 818133 53354 818139
rect 53302 818075 53354 818081
rect 53410 774849 53438 843827
rect 53398 774843 53450 774849
rect 53398 774785 53450 774791
rect 53398 771883 53450 771889
rect 53398 771825 53450 771831
rect 53300 763338 53356 763347
rect 53300 763273 53356 763282
rect 53314 247715 53342 763273
rect 53410 732743 53438 771825
rect 53590 757527 53642 757533
rect 53590 757469 53642 757475
rect 53494 743097 53546 743103
rect 53494 743039 53546 743045
rect 53398 732737 53450 732743
rect 53398 732679 53450 732685
rect 53396 720122 53452 720131
rect 53396 720057 53452 720066
rect 53300 247706 53356 247715
rect 53300 247641 53356 247650
rect 53206 246557 53258 246563
rect 53206 246499 53258 246505
rect 53410 246489 53438 720057
rect 53506 281121 53534 743039
rect 53602 732151 53630 757469
rect 53590 732145 53642 732151
rect 53590 732087 53642 732093
rect 53588 676906 53644 676915
rect 53588 676841 53644 676850
rect 53494 281115 53546 281121
rect 53494 281057 53546 281063
rect 53602 246531 53630 676841
rect 53698 541527 53726 973475
rect 61858 961963 61886 993529
rect 62038 993513 62090 993519
rect 62038 993455 62090 993461
rect 62050 963295 62078 993455
rect 66850 988561 66878 995083
rect 77314 993667 77342 995508
rect 77698 993889 77726 995522
rect 77686 993883 77738 993889
rect 77686 993825 77738 993831
rect 78370 993741 78398 995522
rect 80194 993815 80222 995522
rect 81408 995517 81662 995536
rect 81408 995511 81674 995517
rect 81408 995508 81622 995511
rect 81622 995453 81674 995459
rect 80182 993809 80234 993815
rect 80182 993751 80234 993757
rect 78358 993735 78410 993741
rect 78358 993677 78410 993683
rect 77302 993661 77354 993667
rect 77302 993603 77354 993609
rect 82594 993593 82622 995522
rect 83232 995508 83486 995536
rect 82582 993587 82634 993593
rect 82582 993529 82634 993535
rect 83458 993519 83486 995508
rect 84514 993783 84542 995522
rect 85104 995508 85406 995536
rect 86352 995508 86462 995536
rect 87552 995508 87806 995536
rect 85378 995411 85406 995508
rect 85364 995402 85420 995411
rect 85364 995337 85420 995346
rect 86434 995263 86462 995508
rect 86420 995254 86476 995263
rect 86420 995189 86476 995198
rect 87778 995115 87806 995508
rect 87764 995106 87820 995115
rect 87764 995041 87820 995050
rect 88738 993931 88766 995522
rect 88724 993922 88780 993931
rect 88724 993857 88780 993866
rect 84500 993774 84556 993783
rect 84500 993709 84556 993718
rect 92578 993519 92606 999449
rect 106294 999433 106346 999439
rect 106292 999398 106294 999407
rect 126646 999433 126698 999439
rect 106346 999398 106348 999407
rect 126646 999375 126698 999381
rect 106292 999333 106348 999342
rect 107926 996177 107978 996183
rect 107926 996119 107978 996125
rect 107542 996103 107594 996109
rect 107542 996045 107594 996051
rect 99572 995994 99628 996003
rect 94966 995955 95018 995961
rect 99572 995929 99628 995938
rect 102932 995994 102988 996003
rect 102932 995929 102934 995938
rect 94966 995897 95018 995903
rect 94978 995855 95006 995897
rect 97846 995881 97898 995887
rect 94964 995846 95020 995855
rect 93526 995807 93578 995813
rect 97846 995823 97898 995829
rect 97940 995846 97996 995855
rect 94964 995781 95020 995790
rect 93526 995749 93578 995755
rect 83446 993513 83498 993519
rect 83446 993455 83498 993461
rect 92566 993513 92618 993519
rect 92566 993455 92618 993461
rect 73462 992181 73514 992187
rect 73462 992123 73514 992129
rect 64822 988555 64874 988561
rect 64822 988497 64874 988503
rect 66838 988555 66890 988561
rect 66838 988497 66890 988503
rect 64726 983597 64778 983603
rect 64726 983539 64778 983545
rect 62036 963286 62092 963295
rect 62036 963221 62092 963230
rect 61844 961954 61900 961963
rect 61844 961889 61900 961898
rect 59540 960918 59596 960927
rect 59540 960853 59596 960862
rect 59554 959109 59582 960853
rect 59542 959103 59594 959109
rect 59542 959045 59594 959051
rect 59540 946710 59596 946719
rect 59540 946645 59596 946654
rect 59554 944679 59582 946645
rect 59542 944673 59594 944679
rect 59542 944615 59594 944621
rect 59540 932206 59596 932215
rect 59540 932141 59596 932150
rect 59554 930545 59582 932141
rect 59542 930539 59594 930545
rect 59542 930481 59594 930487
rect 59540 917850 59596 917859
rect 59540 917785 59596 917794
rect 59554 915893 59582 917785
rect 59542 915887 59594 915893
rect 59542 915829 59594 915835
rect 59540 903494 59596 903503
rect 59540 903429 59596 903438
rect 59554 901537 59582 903429
rect 59542 901531 59594 901537
rect 59542 901473 59594 901479
rect 59540 889138 59596 889147
rect 59540 889073 59596 889082
rect 59554 887181 59582 889073
rect 59542 887175 59594 887181
rect 59542 887117 59594 887123
rect 59540 874782 59596 874791
rect 59540 874717 59596 874726
rect 59554 872677 59582 874717
rect 59542 872671 59594 872677
rect 59542 872613 59594 872619
rect 58580 860426 58636 860435
rect 58580 860361 58636 860370
rect 58594 858321 58622 860361
rect 58582 858315 58634 858321
rect 58582 858257 58634 858263
rect 59540 846070 59596 846079
rect 59540 846005 59596 846014
rect 59554 843891 59582 846005
rect 59542 843885 59594 843891
rect 59542 843827 59594 843833
rect 59540 831714 59596 831723
rect 59540 831649 59596 831658
rect 59554 829535 59582 831649
rect 59542 829529 59594 829535
rect 59542 829471 59594 829477
rect 59540 817358 59596 817367
rect 59540 817293 59596 817302
rect 59554 815105 59582 817293
rect 59542 815099 59594 815105
rect 59542 815041 59594 815047
rect 59540 802854 59596 802863
rect 59540 802789 59596 802798
rect 59554 800675 59582 802789
rect 59542 800669 59594 800675
rect 59542 800611 59594 800617
rect 59540 788646 59596 788655
rect 59540 788581 59596 788590
rect 59554 786319 59582 788581
rect 59542 786313 59594 786319
rect 59542 786255 59594 786261
rect 59540 774142 59596 774151
rect 59540 774077 59596 774086
rect 59554 771889 59582 774077
rect 59542 771883 59594 771889
rect 59542 771825 59594 771831
rect 59540 759786 59596 759795
rect 59540 759721 59596 759730
rect 59554 757533 59582 759721
rect 59542 757527 59594 757533
rect 59542 757469 59594 757475
rect 59540 745578 59596 745587
rect 59540 745513 59596 745522
rect 59554 743103 59582 745513
rect 59542 743097 59594 743103
rect 59542 743039 59594 743045
rect 59540 731074 59596 731083
rect 59540 731009 59596 731018
rect 59554 728673 59582 731009
rect 59542 728667 59594 728673
rect 59542 728609 59594 728615
rect 59540 716718 59596 716727
rect 59540 716653 59596 716662
rect 59554 714317 59582 716653
rect 59542 714311 59594 714317
rect 59542 714253 59594 714259
rect 59540 702362 59596 702371
rect 59540 702297 59596 702306
rect 59554 699887 59582 702297
rect 59542 699881 59594 699887
rect 59542 699823 59594 699829
rect 59540 688006 59596 688015
rect 59540 687941 59596 687950
rect 59554 685531 59582 687941
rect 59542 685525 59594 685531
rect 59542 685467 59594 685473
rect 59540 673650 59596 673659
rect 59540 673585 59596 673594
rect 59554 671101 59582 673585
rect 59542 671095 59594 671101
rect 59542 671037 59594 671043
rect 59540 659294 59596 659303
rect 59540 659229 59596 659238
rect 59554 656745 59582 659229
rect 59542 656739 59594 656745
rect 59542 656681 59594 656687
rect 59542 645121 59594 645127
rect 59542 645063 59594 645069
rect 59554 644947 59582 645063
rect 59540 644938 59596 644947
rect 59540 644873 59596 644882
rect 56084 633986 56140 633995
rect 56084 633921 56140 633930
rect 53780 590622 53836 590631
rect 53780 590557 53836 590566
rect 53686 541521 53738 541527
rect 53686 541463 53738 541469
rect 53686 443619 53738 443625
rect 53686 443561 53738 443567
rect 53698 344835 53726 443561
rect 53686 344829 53738 344835
rect 53686 344771 53738 344777
rect 53794 249227 53822 590557
rect 53878 501191 53930 501197
rect 53878 501133 53930 501139
rect 53890 431785 53918 501133
rect 53878 431779 53930 431785
rect 53878 431721 53930 431727
rect 53878 342831 53930 342837
rect 53878 342773 53930 342779
rect 53890 259735 53918 342773
rect 53878 259729 53930 259735
rect 53878 259671 53930 259677
rect 53782 249221 53834 249227
rect 53782 249163 53834 249169
rect 56098 246637 56126 633921
rect 59540 630582 59596 630591
rect 59540 630517 59596 630526
rect 59554 627885 59582 630517
rect 59542 627879 59594 627885
rect 59542 627821 59594 627827
rect 59540 616226 59596 616235
rect 59540 616161 59596 616170
rect 59554 613529 59582 616161
rect 59542 613523 59594 613529
rect 59542 613465 59594 613471
rect 59542 601905 59594 601911
rect 59540 601870 59542 601879
rect 59594 601870 59596 601879
rect 59540 601805 59596 601814
rect 58772 587514 58828 587523
rect 58772 587449 58828 587458
rect 58786 584965 58814 587449
rect 58774 584959 58826 584965
rect 58774 584901 58826 584907
rect 59540 573010 59596 573019
rect 59540 572945 59596 572954
rect 59554 570313 59582 572945
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 59540 558950 59596 558959
rect 59540 558885 59542 558894
rect 59594 558885 59596 558894
rect 59542 558853 59594 558859
rect 59542 544555 59594 544561
rect 59542 544497 59594 544503
rect 59554 544455 59582 544497
rect 59540 544446 59596 544455
rect 59540 544381 59596 544390
rect 59540 530090 59596 530099
rect 59540 530025 59596 530034
rect 59554 529983 59582 530025
rect 59542 529977 59594 529983
rect 59542 529919 59594 529925
rect 59540 515734 59596 515743
rect 59540 515669 59596 515678
rect 59554 515553 59582 515669
rect 59542 515547 59594 515553
rect 59542 515489 59594 515495
rect 59540 501230 59596 501239
rect 59540 501165 59542 501174
rect 59594 501165 59596 501174
rect 59542 501133 59594 501139
rect 58580 486874 58636 486883
rect 58580 486809 58636 486818
rect 58594 486767 58622 486809
rect 58582 486761 58634 486767
rect 58582 486703 58634 486709
rect 59540 472518 59596 472527
rect 59540 472453 59596 472462
rect 59554 472411 59582 472453
rect 59542 472405 59594 472411
rect 59542 472347 59594 472353
rect 59540 458162 59596 458171
rect 59540 458097 59596 458106
rect 59554 457981 59582 458097
rect 59542 457975 59594 457981
rect 59542 457917 59594 457923
rect 59540 443806 59596 443815
rect 59540 443741 59596 443750
rect 59554 443625 59582 443741
rect 59542 443619 59594 443625
rect 59542 443561 59594 443567
rect 59540 429450 59596 429459
rect 59540 429385 59596 429394
rect 59554 429195 59582 429385
rect 59542 429189 59594 429195
rect 59542 429131 59594 429137
rect 56182 417645 56234 417651
rect 56182 417587 56234 417593
rect 56194 249301 56222 417587
rect 58388 415094 58444 415103
rect 58388 415029 58444 415038
rect 58402 414765 58430 415029
rect 58390 414759 58442 414765
rect 58390 414701 58442 414707
rect 58388 400738 58444 400747
rect 58388 400673 58444 400682
rect 58402 400409 58430 400673
rect 58390 400403 58442 400409
rect 58390 400345 58442 400351
rect 59252 386382 59308 386391
rect 59252 386317 59308 386326
rect 59266 385979 59294 386317
rect 59254 385973 59306 385979
rect 59254 385915 59306 385921
rect 59540 371878 59596 371887
rect 59540 371813 59596 371822
rect 59554 371623 59582 371813
rect 59542 371617 59594 371623
rect 59542 371559 59594 371565
rect 59540 357670 59596 357679
rect 59540 357605 59596 357614
rect 59554 357193 59582 357605
rect 59542 357187 59594 357193
rect 59542 357129 59594 357135
rect 58388 343166 58444 343175
rect 58388 343101 58444 343110
rect 58402 342837 58430 343101
rect 58390 342831 58442 342837
rect 58390 342773 58442 342779
rect 57812 328810 57868 328819
rect 57812 328745 57868 328754
rect 57826 328407 57854 328745
rect 57814 328401 57866 328407
rect 57814 328343 57866 328349
rect 58004 314602 58060 314611
rect 58004 314537 58060 314546
rect 58018 313977 58046 314537
rect 58006 313971 58058 313977
rect 58006 313913 58058 313919
rect 59444 300098 59500 300107
rect 59444 300033 59500 300042
rect 59458 299621 59486 300033
rect 59446 299615 59498 299621
rect 59446 299557 59498 299563
rect 58100 285890 58156 285899
rect 58100 285825 58156 285834
rect 58114 285191 58142 285825
rect 58102 285185 58154 285191
rect 58102 285127 58154 285133
rect 64738 278605 64766 983539
rect 64726 278599 64778 278605
rect 64726 278541 64778 278547
rect 64834 277939 64862 988497
rect 65110 986779 65162 986785
rect 65110 986721 65162 986727
rect 65014 986409 65066 986415
rect 65014 986351 65066 986357
rect 64918 983523 64970 983529
rect 64918 983465 64970 983471
rect 64822 277933 64874 277939
rect 64822 277875 64874 277881
rect 64930 272463 64958 983465
rect 64918 272457 64970 272463
rect 64918 272399 64970 272405
rect 56182 249295 56234 249301
rect 56182 249237 56234 249243
rect 65026 246711 65054 986351
rect 65014 246705 65066 246711
rect 65014 246647 65066 246653
rect 56086 246631 56138 246637
rect 56086 246573 56138 246579
rect 53588 246522 53644 246531
rect 53398 246483 53450 246489
rect 53588 246457 53644 246466
rect 53398 246425 53450 246431
rect 47734 246409 47786 246415
rect 65122 246383 65150 986721
rect 65206 986483 65258 986489
rect 65206 986425 65258 986431
rect 65218 246785 65246 986425
rect 73474 983534 73502 992123
rect 89590 989295 89642 989301
rect 89590 989237 89642 989243
rect 89602 983534 89630 989237
rect 93538 986785 93566 995749
rect 93814 995659 93866 995665
rect 93814 995601 93866 995607
rect 93826 995411 93854 995601
rect 97858 995559 97886 995823
rect 97940 995781 97942 995790
rect 97994 995781 97996 995790
rect 97942 995749 97994 995755
rect 98996 995698 99052 995707
rect 98996 995633 98998 995642
rect 99050 995633 99052 995642
rect 98998 995601 99050 995607
rect 97844 995550 97900 995559
rect 97844 995485 97900 995494
rect 93812 995402 93868 995411
rect 93812 995337 93868 995346
rect 99586 995263 99614 995929
rect 102986 995929 102988 995938
rect 102934 995897 102986 995903
rect 102452 995846 102508 995855
rect 102452 995781 102508 995790
rect 104468 995846 104524 995855
rect 104468 995781 104524 995790
rect 102466 995517 102494 995781
rect 102454 995511 102506 995517
rect 102454 995453 102506 995459
rect 99572 995254 99628 995263
rect 99572 995189 99628 995198
rect 97844 994958 97900 994967
rect 97844 994893 97900 994902
rect 97858 993889 97886 994893
rect 97846 993883 97898 993889
rect 97846 993825 97898 993831
rect 104482 993783 104510 995781
rect 107554 995559 107582 996045
rect 107938 995855 107966 996119
rect 108982 996029 109034 996035
rect 108980 995994 108982 996003
rect 109034 995994 109036 996003
rect 108980 995929 109036 995938
rect 109556 995994 109612 996003
rect 109556 995929 109612 995938
rect 107924 995846 107980 995855
rect 107924 995781 107980 995790
rect 107540 995550 107596 995559
rect 107540 995485 107596 995494
rect 105908 995402 105964 995411
rect 105908 995337 105964 995346
rect 105332 995254 105388 995263
rect 105332 995189 105388 995198
rect 105346 993815 105374 995189
rect 105334 993809 105386 993815
rect 104468 993774 104524 993783
rect 105334 993751 105386 993757
rect 104468 993709 104524 993718
rect 105922 993667 105950 995337
rect 106964 995254 107020 995263
rect 106964 995189 107020 995198
rect 106978 993741 107006 995189
rect 106966 993735 107018 993741
rect 106966 993677 107018 993683
rect 105910 993661 105962 993667
rect 105910 993603 105962 993609
rect 105814 990479 105866 990485
rect 105814 990421 105866 990427
rect 93526 986779 93578 986785
rect 93526 986721 93578 986727
rect 105826 983534 105854 990421
rect 107554 986637 107582 995485
rect 107542 986631 107594 986637
rect 107542 986573 107594 986579
rect 107938 986563 107966 995781
rect 109172 995550 109228 995559
rect 109172 995485 109228 995494
rect 109186 986711 109214 995485
rect 109364 995106 109420 995115
rect 109364 995041 109420 995050
rect 109378 989301 109406 995041
rect 109570 990485 109598 995929
rect 126658 995855 126686 999375
rect 126644 995846 126700 995855
rect 126644 995781 126700 995790
rect 134324 995846 134380 995855
rect 136148 995846 136204 995855
rect 134380 995804 135134 995832
rect 135936 995804 136148 995832
rect 134324 995781 134380 995790
rect 110228 995254 110284 995263
rect 110228 995189 110284 995198
rect 110242 992187 110270 995189
rect 128482 993741 128510 995522
rect 129120 995508 129374 995536
rect 129346 993815 129374 995508
rect 129334 993809 129386 993815
rect 129334 993751 129386 993757
rect 128470 993735 128522 993741
rect 128470 993677 128522 993683
rect 129730 993667 129758 995522
rect 131616 995508 131870 995536
rect 131842 994227 131870 995508
rect 131828 994218 131884 994227
rect 131828 994153 131884 994162
rect 132130 993889 132158 995522
rect 132802 994375 132830 995522
rect 133440 995508 133694 995536
rect 133666 994523 133694 995508
rect 133954 995508 134016 995536
rect 133652 994514 133708 994523
rect 133652 994449 133708 994458
rect 132788 994366 132844 994375
rect 132788 994301 132844 994310
rect 132118 993883 132170 993889
rect 132118 993825 132170 993831
rect 129718 993661 129770 993667
rect 129718 993603 129770 993609
rect 133954 993593 133982 995508
rect 135106 994056 135134 995804
rect 137136 995813 137438 995832
rect 137760 995813 138014 995832
rect 143650 995813 143678 1002316
rect 143926 1002261 143978 1002267
rect 143830 1000839 143882 1000845
rect 143830 1000781 143882 1000787
rect 143734 999507 143786 999513
rect 143734 999449 143786 999455
rect 137136 995807 137450 995813
rect 137136 995804 137398 995807
rect 136148 995781 136204 995790
rect 137760 995807 138026 995813
rect 137760 995804 137974 995807
rect 137398 995749 137450 995755
rect 137974 995749 138026 995755
rect 143638 995807 143690 995813
rect 143638 995749 143690 995755
rect 136726 995733 136778 995739
rect 136464 995681 136726 995684
rect 136464 995675 136778 995681
rect 136464 995656 136766 995675
rect 142656 995665 143006 995684
rect 143746 995665 143774 999449
rect 142656 995659 143018 995665
rect 142656 995656 142966 995659
rect 142966 995601 143018 995607
rect 143734 995659 143786 995665
rect 143734 995601 143786 995607
rect 143842 995591 143870 1000781
rect 141046 995585 141098 995591
rect 139220 995550 139276 995559
rect 138960 995508 139220 995536
rect 140160 995508 140414 995536
rect 140784 995533 141046 995536
rect 140784 995527 141098 995533
rect 143830 995585 143882 995591
rect 143830 995527 143882 995533
rect 140784 995508 141086 995527
rect 139220 995485 139276 995494
rect 135188 994070 135244 994079
rect 135106 994028 135188 994056
rect 135188 994005 135244 994014
rect 140386 993783 140414 995508
rect 140372 993774 140428 993783
rect 140372 993709 140428 993718
rect 143938 993593 143966 1002261
rect 144022 999433 144074 999439
rect 144022 999375 144074 999381
rect 144034 995887 144062 999375
rect 144118 996547 144170 996553
rect 144118 996489 144170 996495
rect 144022 995881 144074 995887
rect 144130 995855 144158 996489
rect 144022 995823 144074 995829
rect 144116 995846 144172 995855
rect 144116 995781 144172 995790
rect 144692 995402 144748 995411
rect 144692 995337 144748 995346
rect 144706 994375 144734 995337
rect 144692 994366 144748 994375
rect 144692 994301 144748 994310
rect 133942 993587 133994 993593
rect 133942 993529 133994 993535
rect 143926 993587 143978 993593
rect 143926 993529 143978 993535
rect 110230 992181 110282 992187
rect 110230 992123 110282 992129
rect 109558 990479 109610 990485
rect 109558 990421 109610 990427
rect 109366 989295 109418 989301
rect 109366 989237 109418 989243
rect 138262 989295 138314 989301
rect 138262 989237 138314 989243
rect 122038 988333 122090 988339
rect 122038 988275 122090 988281
rect 109174 986705 109226 986711
rect 109174 986647 109226 986653
rect 107926 986557 107978 986563
rect 107926 986499 107978 986505
rect 122050 983534 122078 988275
rect 138274 983534 138302 989237
rect 145378 986489 145406 1007917
rect 349652 1007834 349708 1007843
rect 349652 1007769 349708 1007778
rect 353300 1007834 353356 1007843
rect 353410 1007820 353438 1015909
rect 434998 1008091 435050 1008097
rect 434998 1008033 435050 1008039
rect 470806 1008091 470858 1008097
rect 470806 1008033 470858 1008039
rect 353356 1007792 353438 1007820
rect 353300 1007769 353356 1007778
rect 299156 1005910 299212 1005919
rect 299156 1005845 299212 1005854
rect 302996 1005910 303052 1005919
rect 302996 1005845 303052 1005854
rect 164278 1005279 164330 1005285
rect 164278 1005221 164330 1005227
rect 172822 1005279 172874 1005285
rect 172822 1005221 172874 1005227
rect 160436 1003246 160492 1003255
rect 160436 1003181 160438 1003190
rect 160490 1003181 160492 1003190
rect 161492 1003209 161548 1003218
rect 164290 1003213 164318 1005221
rect 160438 1003149 160490 1003155
rect 161492 1003144 161548 1003153
rect 164278 1003207 164330 1003213
rect 164278 1003149 164330 1003155
rect 161506 1002843 161534 1003144
rect 161494 1002837 161546 1002843
rect 161494 1002779 161546 1002785
rect 169942 1002837 169994 1002843
rect 169942 1002779 169994 1002785
rect 151124 1002506 151180 1002515
rect 151124 1002441 151126 1002450
rect 151178 1002441 151180 1002450
rect 151126 1002409 151178 1002415
rect 146806 1002393 146858 1002399
rect 152758 1002393 152810 1002399
rect 146806 1002335 146858 1002341
rect 152756 1002358 152758 1002367
rect 152810 1002358 152812 1002367
rect 146818 999439 146846 1002335
rect 152756 1002293 152812 1002302
rect 157652 1000878 157708 1000887
rect 157652 1000813 157654 1000822
rect 157706 1000813 157708 1000822
rect 157654 1000781 157706 1000787
rect 155540 999546 155596 999555
rect 155540 999481 155542 999490
rect 155594 999481 155596 999490
rect 155542 999449 155594 999455
rect 146806 999433 146858 999439
rect 146806 999375 146858 999381
rect 156020 996586 156076 996595
rect 156020 996521 156022 996530
rect 156074 996521 156076 996530
rect 156022 996489 156074 996495
rect 159766 996177 159818 996183
rect 159188 996142 159244 996151
rect 159188 996077 159190 996086
rect 159242 996077 159244 996086
rect 159764 996142 159766 996151
rect 159818 996142 159820 996151
rect 159764 996077 159820 996086
rect 159190 996045 159242 996051
rect 160438 996029 160490 996035
rect 152084 995994 152140 996003
rect 146806 995955 146858 995961
rect 152084 995929 152086 995938
rect 146806 995897 146858 995903
rect 152138 995929 152140 995938
rect 160436 995994 160438 996003
rect 160490 995994 160492 996003
rect 160436 995929 160492 995938
rect 152086 995897 152138 995903
rect 146818 994523 146846 995897
rect 151700 995846 151756 995855
rect 149590 995807 149642 995813
rect 151700 995781 151756 995790
rect 154868 995846 154924 995855
rect 154868 995781 154870 995790
rect 149590 995749 149642 995755
rect 146804 994514 146860 994523
rect 146804 994449 146860 994458
rect 146900 994366 146956 994375
rect 146900 994301 146956 994310
rect 146914 994079 146942 994301
rect 146900 994070 146956 994079
rect 146900 994005 146956 994014
rect 149602 993815 149630 995749
rect 151714 995739 151742 995781
rect 154922 995781 154924 995790
rect 158228 995846 158284 995855
rect 158228 995781 158284 995790
rect 161492 995846 161548 995855
rect 161492 995781 161548 995790
rect 154870 995749 154922 995755
rect 151702 995733 151754 995739
rect 151702 995675 151754 995681
rect 154772 995402 154828 995411
rect 154772 995337 154828 995346
rect 149684 995254 149740 995263
rect 149684 995189 149740 995198
rect 149698 993889 149726 995189
rect 154786 994227 154814 995337
rect 157268 995254 157324 995263
rect 157268 995189 157324 995198
rect 154772 994218 154828 994227
rect 154772 994153 154828 994162
rect 149686 993883 149738 993889
rect 149686 993825 149738 993831
rect 149590 993809 149642 993815
rect 149590 993751 149642 993757
rect 157282 993741 157310 995189
rect 157270 993735 157322 993741
rect 157270 993677 157322 993683
rect 158242 993667 158270 995781
rect 158230 993661 158282 993667
rect 158230 993603 158282 993609
rect 154486 989369 154538 989375
rect 154486 989311 154538 989317
rect 145366 986483 145418 986489
rect 145366 986425 145418 986431
rect 154498 983534 154526 989311
rect 161506 989301 161534 995781
rect 161684 995254 161740 995263
rect 161684 995189 161740 995198
rect 161698 989375 161726 995189
rect 161686 989369 161738 989375
rect 161686 989311 161738 989317
rect 161494 989295 161546 989301
rect 161494 989237 161546 989243
rect 169954 983548 169982 1002779
rect 172834 995961 172862 1005221
rect 218806 1005205 218858 1005211
rect 213812 1005170 213868 1005179
rect 213812 1005105 213868 1005114
rect 218804 1005170 218806 1005179
rect 222742 1005205 222794 1005211
rect 218858 1005170 218860 1005179
rect 222742 1005147 222794 1005153
rect 218804 1005105 218860 1005114
rect 211796 1003246 211852 1003255
rect 213826 1003213 213854 1005105
rect 211796 1003181 211798 1003190
rect 211850 1003181 211852 1003190
rect 213814 1003207 213866 1003213
rect 211798 1003149 211850 1003155
rect 213814 1003149 213866 1003155
rect 175702 1002319 175754 1002325
rect 175702 1002261 175754 1002267
rect 172822 995955 172874 995961
rect 172822 995897 172874 995903
rect 175714 995739 175742 1002261
rect 209108 1000878 209164 1000887
rect 195190 1000839 195242 1000845
rect 209108 1000813 209110 1000822
rect 195190 1000781 195242 1000787
rect 209162 1000813 209164 1000822
rect 209110 1000781 209162 1000787
rect 195094 999433 195146 999439
rect 195094 999375 195146 999381
rect 178486 996177 178538 996183
rect 178486 996119 178538 996125
rect 178498 996035 178526 996119
rect 178486 996029 178538 996035
rect 178486 995971 178538 995977
rect 188756 995846 188812 995855
rect 183552 995813 183806 995832
rect 183552 995807 183818 995813
rect 183552 995804 183766 995807
rect 188544 995804 188756 995832
rect 189428 995846 189484 995855
rect 189168 995804 189428 995832
rect 188756 995781 188812 995790
rect 189428 995781 189484 995790
rect 183766 995749 183818 995755
rect 195106 995739 195134 999375
rect 175702 995733 175754 995739
rect 175702 995675 175754 995681
rect 185206 995733 185258 995739
rect 194422 995733 194474 995739
rect 185258 995681 185424 995684
rect 185206 995675 185424 995681
rect 185218 995670 185424 995675
rect 185218 995656 185438 995670
rect 192192 995665 192542 995684
rect 194064 995681 194422 995684
rect 194064 995675 194474 995681
rect 195094 995733 195146 995739
rect 195094 995675 195146 995681
rect 192192 995659 192554 995665
rect 192192 995656 192502 995659
rect 185110 995585 185162 995591
rect 179842 993741 179870 995522
rect 180514 993963 180542 995522
rect 181152 995508 181406 995536
rect 180502 993957 180554 993963
rect 180502 993899 180554 993905
rect 181378 993815 181406 995508
rect 183010 993889 183038 995522
rect 184066 995517 184176 995536
rect 184054 995511 184176 995517
rect 184106 995508 184176 995511
rect 184848 995533 185110 995536
rect 184848 995527 185162 995533
rect 184848 995508 185150 995527
rect 184054 995453 184106 995459
rect 182998 993883 183050 993889
rect 182998 993825 183050 993831
rect 181366 993809 181418 993815
rect 181366 993751 181418 993757
rect 179830 993735 179882 993741
rect 179830 993677 179882 993683
rect 185410 993667 185438 995656
rect 194064 995656 194462 995675
rect 195202 995665 195230 1000781
rect 206902 999433 206954 999439
rect 206900 999398 206902 999407
rect 206954 999398 206956 999407
rect 206900 999333 206956 999342
rect 205268 996586 205324 996595
rect 195766 996547 195818 996553
rect 205268 996521 205270 996530
rect 195766 996489 195818 996495
rect 205322 996521 205324 996530
rect 205270 996489 205322 996495
rect 195190 995659 195242 995665
rect 192502 995601 192554 995607
rect 195190 995601 195242 995607
rect 188084 995550 188140 995559
rect 185794 995508 186048 995536
rect 185794 994375 185822 995508
rect 187330 994375 187358 995522
rect 187872 995508 188084 995536
rect 190368 995508 190622 995536
rect 188084 995485 188140 995494
rect 190594 995411 190622 995508
rect 190580 995402 190636 995411
rect 190580 995337 190636 995346
rect 185780 994366 185836 994375
rect 185780 994301 185836 994310
rect 187316 994366 187372 994375
rect 187316 994301 187372 994310
rect 191554 994079 191582 995522
rect 195778 995517 195806 996489
rect 210166 996473 210218 996479
rect 210166 996415 210218 996421
rect 198646 996177 198698 996183
rect 204022 996177 204074 996183
rect 198646 996119 198698 996125
rect 204020 996142 204022 996151
rect 210178 996151 210206 996415
rect 204074 996142 204076 996151
rect 198658 996003 198686 996119
rect 204020 996077 204076 996086
rect 210164 996142 210220 996151
rect 210164 996077 210166 996086
rect 210218 996077 210220 996086
rect 210166 996045 210218 996051
rect 222754 996035 222782 1005147
rect 255478 1002393 255530 1002399
rect 253844 1002358 253900 1002367
rect 246646 1002319 246698 1002325
rect 253844 1002293 253846 1002302
rect 246646 1002261 246698 1002267
rect 253898 1002293 253900 1002302
rect 255476 1002358 255478 1002367
rect 255530 1002358 255532 1002367
rect 255476 1002293 255532 1002302
rect 253846 1002261 253898 1002267
rect 246550 1002245 246602 1002251
rect 246550 1002187 246602 1002193
rect 225430 996473 225482 996479
rect 225430 996415 225482 996421
rect 225442 996109 225470 996415
rect 225430 996103 225482 996109
rect 225430 996045 225482 996051
rect 210646 996029 210698 996035
rect 198644 995994 198700 996003
rect 198644 995929 198700 995938
rect 207380 995994 207436 996003
rect 207380 995929 207436 995938
rect 210644 995994 210646 996003
rect 222742 996029 222794 996035
rect 210698 995994 210700 996003
rect 210644 995929 210700 995938
rect 211796 995994 211852 996003
rect 211796 995929 211798 995938
rect 198646 995881 198698 995887
rect 198644 995846 198646 995855
rect 202486 995881 202538 995887
rect 198698 995846 198700 995855
rect 198644 995781 198700 995790
rect 202484 995846 202486 995855
rect 202538 995846 202540 995855
rect 202484 995781 202540 995790
rect 202964 995846 203020 995855
rect 202964 995781 203020 995790
rect 205652 995846 205708 995855
rect 205652 995781 205654 995790
rect 202978 995739 203006 995781
rect 205706 995781 205708 995790
rect 205654 995749 205706 995755
rect 198454 995733 198506 995739
rect 197204 995698 197260 995707
rect 198454 995675 198506 995681
rect 202966 995733 203018 995739
rect 202966 995675 203018 995681
rect 197204 995633 197260 995642
rect 195766 995511 195818 995517
rect 195766 995453 195818 995459
rect 191540 994070 191596 994079
rect 191540 994005 191596 994014
rect 185398 993661 185450 993667
rect 185398 993603 185450 993609
rect 186934 988259 186986 988265
rect 186934 988201 186986 988207
rect 169954 983520 170736 983548
rect 186946 983534 186974 988201
rect 197218 986415 197246 995633
rect 198466 995559 198494 995675
rect 198646 995585 198698 995591
rect 198452 995550 198508 995559
rect 198452 995485 198508 995494
rect 198644 995550 198646 995559
rect 198698 995550 198700 995559
rect 198644 995485 198700 995494
rect 198644 995254 198700 995263
rect 198644 995189 198700 995198
rect 198658 993963 198686 995189
rect 207394 994375 207422 995929
rect 211850 995929 211852 995938
rect 219092 995994 219148 996003
rect 222742 995971 222794 995977
rect 219092 995929 219148 995938
rect 211798 995897 211850 995903
rect 213332 995846 213388 995855
rect 213332 995781 213388 995790
rect 208148 995254 208204 995263
rect 208148 995189 208204 995198
rect 208724 995254 208780 995263
rect 208724 995189 208780 995198
rect 209780 995254 209836 995263
rect 209780 995189 209836 995198
rect 207380 994366 207436 994375
rect 207380 994301 207436 994310
rect 198646 993957 198698 993963
rect 198646 993899 198698 993905
rect 208162 993889 208190 995189
rect 208150 993883 208202 993889
rect 208150 993825 208202 993831
rect 208738 993741 208766 995189
rect 209794 993815 209822 995189
rect 209782 993809 209834 993815
rect 209782 993751 209834 993757
rect 208726 993735 208778 993741
rect 208726 993677 208778 993683
rect 213346 989375 213374 995781
rect 216020 995698 216076 995707
rect 216020 995633 216076 995642
rect 203158 989369 203210 989375
rect 203158 989311 203210 989317
rect 213334 989369 213386 989375
rect 213334 989311 213386 989317
rect 197206 986409 197258 986415
rect 197206 986351 197258 986357
rect 203170 983534 203198 989311
rect 216034 989301 216062 995633
rect 216022 989295 216074 989301
rect 216022 989237 216074 989243
rect 219106 983548 219134 995929
rect 243188 995846 243244 995855
rect 239280 995813 239582 995832
rect 240576 995813 240926 995832
rect 239280 995807 239594 995813
rect 239280 995804 239542 995807
rect 240576 995807 240938 995813
rect 240576 995804 240886 995807
rect 239542 995749 239594 995755
rect 242976 995804 243188 995832
rect 243956 995846 244012 995855
rect 243600 995804 243956 995832
rect 243188 995781 243244 995790
rect 243956 995781 244012 995790
rect 240886 995749 240938 995755
rect 246562 995739 246590 1002187
rect 246658 995813 246686 1002261
rect 258836 999694 258892 999703
rect 247030 999655 247082 999661
rect 258836 999629 258838 999638
rect 247030 999597 247082 999603
rect 258890 999629 258892 999638
rect 258838 999597 258890 999603
rect 246742 999581 246794 999587
rect 246742 999523 246794 999529
rect 246646 995807 246698 995813
rect 246646 995749 246698 995755
rect 240310 995733 240362 995739
rect 239952 995681 240310 995684
rect 246550 995733 246602 995739
rect 241844 995698 241900 995707
rect 239952 995675 240362 995681
rect 239952 995656 240350 995675
rect 241776 995656 241844 995684
rect 246550 995675 246602 995681
rect 241844 995633 241900 995642
rect 236468 995550 236524 995559
rect 231264 995508 231518 995536
rect 231936 995508 232190 995536
rect 231490 993815 231518 995508
rect 232162 993889 232190 995508
rect 232546 994375 232574 995522
rect 233302 995067 233354 995073
rect 233302 995009 233354 995015
rect 232532 994366 232588 994375
rect 232532 994301 232588 994310
rect 232150 993883 232202 993889
rect 232150 993825 232202 993831
rect 231478 993809 231530 993815
rect 231478 993751 231530 993757
rect 233314 988876 233342 995009
rect 234370 993741 234398 995522
rect 234946 993963 234974 995522
rect 235584 995508 235838 995536
rect 236256 995508 236468 995536
rect 235810 994037 235838 995508
rect 236468 995485 236524 995494
rect 235798 994031 235850 994037
rect 235798 993973 235850 993979
rect 234934 993957 234986 993963
rect 234934 993899 234986 993905
rect 234358 993735 234410 993741
rect 234358 993677 234410 993683
rect 236770 993667 236798 995522
rect 237456 995508 237566 995536
rect 238704 995508 239006 995536
rect 245424 995517 245726 995536
rect 246754 995517 246782 999523
rect 246838 999507 246890 999513
rect 246838 999449 246890 999455
rect 246850 995855 246878 999449
rect 246934 999433 246986 999439
rect 246934 999375 246986 999381
rect 246946 996003 246974 999375
rect 246932 995994 246988 996003
rect 246932 995929 246988 995938
rect 246836 995846 246892 995855
rect 246836 995781 246892 995790
rect 246934 995807 246986 995813
rect 246934 995749 246986 995755
rect 245424 995511 245738 995517
rect 245424 995508 245686 995511
rect 237538 994227 237566 995508
rect 238978 995411 239006 995508
rect 245686 995453 245738 995459
rect 246742 995511 246794 995517
rect 246742 995453 246794 995459
rect 238964 995402 239020 995411
rect 238964 995337 239020 995346
rect 237524 994218 237580 994227
rect 237524 994153 237580 994162
rect 246946 993889 246974 995749
rect 247042 995411 247070 999597
rect 258358 999581 258410 999587
rect 258356 999546 258358 999555
rect 298294 999581 298346 999587
rect 258410 999546 258412 999555
rect 258356 999481 258412 999490
rect 260468 999546 260524 999555
rect 298294 999523 298346 999529
rect 260468 999481 260470 999490
rect 260522 999481 260524 999490
rect 260470 999449 260522 999455
rect 279286 999433 279338 999439
rect 279286 999375 279338 999381
rect 298102 999433 298154 999439
rect 298102 999375 298154 999381
rect 259988 996586 260044 996595
rect 247126 996547 247178 996553
rect 259988 996521 259990 996530
rect 247126 996489 247178 996495
rect 260042 996521 260044 996530
rect 259990 996489 260042 996495
rect 247028 995402 247084 995411
rect 247028 995337 247084 995346
rect 246934 993883 246986 993889
rect 246934 993825 246986 993831
rect 247138 993815 247166 996489
rect 262100 996290 262156 996299
rect 262100 996225 262156 996234
rect 262114 996183 262142 996225
rect 262102 996177 262154 996183
rect 262004 996142 262060 996151
rect 263062 996177 263114 996183
rect 262102 996119 262154 996125
rect 263060 996142 263062 996151
rect 263114 996142 263116 996151
rect 262004 996077 262006 996086
rect 262058 996077 262060 996086
rect 263060 996077 263116 996086
rect 262006 996045 262058 996051
rect 263254 996029 263306 996035
rect 254516 995994 254572 996003
rect 254516 995929 254572 995938
rect 257684 995994 257740 996003
rect 257684 995929 257740 995938
rect 263252 995994 263254 996003
rect 263306 995994 263308 996003
rect 263252 995929 263308 995938
rect 254530 995887 254558 995929
rect 254518 995881 254570 995887
rect 254518 995823 254570 995829
rect 256148 995846 256204 995855
rect 257698 995813 257726 995929
rect 259412 995846 259468 995855
rect 256148 995781 256204 995790
rect 257686 995807 257738 995813
rect 256162 995739 256190 995781
rect 259412 995781 259468 995790
rect 270740 995846 270796 995855
rect 270740 995781 270796 995790
rect 257686 995749 257738 995755
rect 247606 995733 247658 995739
rect 247604 995698 247606 995707
rect 256150 995733 256202 995739
rect 247658 995698 247660 995707
rect 247604 995633 247660 995642
rect 247796 995698 247852 995707
rect 256150 995675 256202 995681
rect 247796 995633 247852 995642
rect 247604 995402 247660 995411
rect 247604 995337 247660 995346
rect 247618 994037 247646 995337
rect 247810 995073 247838 995633
rect 250484 995254 250540 995263
rect 250484 995189 250540 995198
rect 247798 995067 247850 995073
rect 247798 995009 247850 995015
rect 247606 994031 247658 994037
rect 247606 993973 247658 993979
rect 250498 993963 250526 995189
rect 250486 993957 250538 993963
rect 250486 993899 250538 993905
rect 247126 993809 247178 993815
rect 247126 993751 247178 993757
rect 259426 993741 259454 995781
rect 267956 995698 268012 995707
rect 267956 995633 268012 995642
rect 267860 995550 267916 995559
rect 267860 995485 267916 995494
rect 259414 993735 259466 993741
rect 259414 993677 259466 993683
rect 236758 993661 236810 993667
rect 236758 993603 236810 993609
rect 267874 989301 267902 995485
rect 235606 989295 235658 989301
rect 235606 989237 235658 989243
rect 267862 989295 267914 989301
rect 267862 989237 267914 989243
rect 233218 988848 233342 988876
rect 233218 985009 233246 988848
rect 225526 985003 225578 985009
rect 225526 984945 225578 984951
rect 233206 985003 233258 985009
rect 233206 984945 233258 984951
rect 225538 983603 225566 984945
rect 225526 983597 225578 983603
rect 219106 983520 219408 983548
rect 225526 983539 225578 983545
rect 235618 983534 235646 989237
rect 251830 988185 251882 988191
rect 251830 988127 251882 988133
rect 251842 983534 251870 988127
rect 267862 986409 267914 986415
rect 267862 986351 267914 986357
rect 267874 983529 267902 986351
rect 267970 983548 267998 995633
rect 270754 989375 270782 995781
rect 279298 995073 279326 999375
rect 298114 997578 298142 999375
rect 298114 997528 298236 997578
rect 298114 997468 298162 997528
rect 298222 997468 298236 997528
rect 298114 997402 298236 997468
rect 298114 997400 298142 997402
rect 280244 997178 280300 997187
rect 280244 997113 280300 997122
rect 298100 997178 298156 997187
rect 298100 997113 298102 997122
rect 280258 996257 280286 997113
rect 298154 997113 298156 997122
rect 298102 997081 298154 997087
rect 298120 996740 298240 996766
rect 298120 996680 298164 996740
rect 298224 996680 298240 996740
rect 298120 996664 298240 996680
rect 280246 996251 280298 996257
rect 280246 996193 280298 996199
rect 298166 995930 298194 996664
rect 298018 995902 298194 995930
rect 290516 995846 290572 995855
rect 283536 995813 283838 995832
rect 283536 995807 283850 995813
rect 283536 995804 283798 995807
rect 290352 995804 290516 995832
rect 290880 995813 291230 995832
rect 290516 995781 290572 995790
rect 290710 995807 290762 995813
rect 283798 995749 283850 995755
rect 290880 995807 291242 995813
rect 290880 995804 291190 995807
rect 290710 995749 290762 995755
rect 291190 995749 291242 995755
rect 288994 995656 289056 995684
rect 286774 995585 286826 995591
rect 279286 995067 279338 995073
rect 279286 995009 279338 995015
rect 282850 993741 282878 995522
rect 284160 995508 284414 995536
rect 286560 995533 286774 995536
rect 286560 995527 286826 995533
rect 282838 993735 282890 993741
rect 282838 993677 282890 993683
rect 284386 993667 284414 995508
rect 286018 994523 286046 995522
rect 286560 995508 286814 995527
rect 287184 995517 287486 995536
rect 287184 995511 287498 995517
rect 287184 995508 287446 995511
rect 287856 995508 287966 995536
rect 287446 995453 287498 995459
rect 287938 995443 287966 995508
rect 288130 995508 288384 995536
rect 287926 995437 287978 995443
rect 287926 995379 287978 995385
rect 288020 994662 288076 994671
rect 288020 994597 288076 994606
rect 286004 994514 286060 994523
rect 286004 994449 286060 994458
rect 288034 994227 288062 994597
rect 288020 994218 288076 994227
rect 288020 994153 288076 994162
rect 284374 993661 284426 993667
rect 284374 993603 284426 993609
rect 288130 993445 288158 995508
rect 288994 994671 289022 995656
rect 290722 995517 290750 995749
rect 291766 995733 291818 995739
rect 291504 995681 291766 995684
rect 292532 995698 292588 995707
rect 291504 995675 291818 995681
rect 291504 995656 291806 995675
rect 292176 995656 292532 995684
rect 297072 995665 297374 995684
rect 298018 995665 298046 995902
rect 297072 995659 297386 995665
rect 297072 995656 297334 995659
rect 292532 995633 292588 995642
rect 297334 995601 297386 995607
rect 298006 995659 298058 995665
rect 298006 995601 298058 995607
rect 298306 995591 298334 999523
rect 298390 999507 298442 999513
rect 298390 999449 298442 999455
rect 298402 995855 298430 999449
rect 298388 995846 298444 995855
rect 298388 995781 298444 995790
rect 295414 995585 295466 995591
rect 293588 995550 293644 995559
rect 290710 995511 290762 995517
rect 293376 995508 293588 995536
rect 295200 995533 295414 995536
rect 295200 995527 295466 995533
rect 298294 995585 298346 995591
rect 298294 995527 298346 995533
rect 293588 995485 293644 995494
rect 290710 995453 290762 995459
rect 288980 994662 289036 994671
rect 288980 994597 289036 994606
rect 290902 994327 290954 994333
rect 290902 994269 290954 994275
rect 288118 993439 288170 993445
rect 288118 993381 288170 993387
rect 270742 989369 270794 989375
rect 270742 989311 270794 989317
rect 284278 989369 284330 989375
rect 284278 989311 284330 989317
rect 267862 983523 267914 983529
rect 267970 983520 268080 983548
rect 284290 983534 284318 989311
rect 290914 986415 290942 994269
rect 294562 994227 294590 995522
rect 295200 995508 295454 995527
rect 299170 994333 299198 1005845
rect 299350 1002911 299402 1002917
rect 299350 1002853 299402 1002859
rect 299254 1002763 299306 1002769
rect 299254 1002705 299306 1002711
rect 299266 995887 299294 1002705
rect 299254 995881 299306 995887
rect 299254 995823 299306 995829
rect 299362 995517 299390 1002853
rect 299446 1002837 299498 1002843
rect 299446 1002779 299498 1002785
rect 299458 996035 299486 1002779
rect 303010 999291 303038 1005845
rect 316822 1005279 316874 1005285
rect 316822 1005221 316874 1005227
rect 331222 1005279 331274 1005285
rect 331222 1005221 331274 1005227
rect 316436 1003246 316492 1003255
rect 316834 1003232 316862 1005221
rect 316492 1003204 316862 1003232
rect 316436 1003181 316492 1003190
rect 308852 1002950 308908 1002959
rect 308852 1002885 308854 1002894
rect 308906 1002885 308908 1002894
rect 308854 1002853 308906 1002859
rect 309334 1002837 309386 1002843
rect 308276 1002802 308332 1002811
rect 308276 1002737 308278 1002746
rect 308330 1002737 308332 1002746
rect 309332 1002802 309334 1002811
rect 309386 1002802 309388 1002811
rect 309332 1002737 309388 1002746
rect 308278 1002705 308330 1002711
rect 312118 999581 312170 999587
rect 310484 999546 310540 999555
rect 310484 999481 310486 999490
rect 310538 999481 310540 999490
rect 312116 999546 312118 999555
rect 312170 999546 312172 999555
rect 312116 999481 312172 999490
rect 310486 999449 310538 999455
rect 309910 999433 309962 999439
rect 309908 999398 309910 999407
rect 309962 999398 309964 999407
rect 309908 999333 309964 999342
rect 313750 999359 313802 999365
rect 313750 999301 313802 999307
rect 331126 999359 331178 999365
rect 331126 999301 331178 999307
rect 302998 999285 303050 999291
rect 304342 999285 304394 999291
rect 302998 999227 303050 999233
rect 304340 999250 304342 999259
rect 304918 999285 304970 999291
rect 304394 999250 304396 999259
rect 304340 999185 304396 999194
rect 304916 999250 304918 999259
rect 304970 999250 304972 999259
rect 304916 999185 304972 999194
rect 313762 997187 313790 999301
rect 314804 997770 314860 997779
rect 314804 997705 314806 997714
rect 314858 997705 314860 997714
rect 314806 997673 314858 997679
rect 331138 997663 331166 999301
rect 331126 997657 331178 997663
rect 331126 997599 331178 997605
rect 313748 997178 313804 997187
rect 313748 997113 313750 997122
rect 313802 997113 313804 997122
rect 313750 997081 313802 997087
rect 313174 996473 313226 996479
rect 313174 996415 313226 996421
rect 313186 996151 313214 996415
rect 314806 996177 314858 996183
rect 313172 996142 313228 996151
rect 313172 996077 313174 996086
rect 313226 996077 313228 996086
rect 314804 996142 314806 996151
rect 314858 996142 314860 996151
rect 314804 996077 314860 996086
rect 313174 996045 313226 996051
rect 299446 996029 299498 996035
rect 299446 995971 299498 995977
rect 303956 995994 304012 996003
rect 304340 995994 304396 996003
rect 304012 995952 304340 995980
rect 303956 995929 304012 995938
rect 304340 995929 304396 995938
rect 311540 995994 311596 996003
rect 311540 995929 311596 995938
rect 319604 995994 319660 996003
rect 319604 995929 319660 995938
rect 306068 995846 306124 995855
rect 306068 995781 306070 995790
rect 306122 995781 306124 995790
rect 306548 995846 306604 995855
rect 306548 995781 306604 995790
rect 306070 995749 306122 995755
rect 306454 995733 306506 995739
rect 306452 995698 306454 995707
rect 306506 995698 306508 995707
rect 306452 995633 306508 995642
rect 299350 995511 299402 995517
rect 299350 995453 299402 995459
rect 306562 995443 306590 995781
rect 306550 995437 306602 995443
rect 306550 995379 306602 995385
rect 308084 994662 308140 994671
rect 308084 994597 308140 994606
rect 308098 994375 308126 994597
rect 308084 994366 308140 994375
rect 299158 994327 299210 994333
rect 308084 994301 308140 994310
rect 299158 994269 299210 994275
rect 294548 994218 294604 994227
rect 294548 994153 294604 994162
rect 311554 993741 311582 995929
rect 312788 995402 312844 995411
rect 312788 995337 312844 995346
rect 311542 993735 311594 993741
rect 311542 993677 311594 993683
rect 312802 993667 312830 995337
rect 312790 993661 312842 993667
rect 312790 993603 312842 993609
rect 319618 989375 319646 995929
rect 319700 995698 319756 995707
rect 319700 995633 319756 995642
rect 319606 989369 319658 989375
rect 319606 989311 319658 989317
rect 319714 989301 319742 995633
rect 328246 993587 328298 993593
rect 328246 993529 328298 993535
rect 328258 993464 328286 993529
rect 328258 993445 328478 993464
rect 328258 993439 328490 993445
rect 328258 993436 328438 993439
rect 328438 993381 328490 993387
rect 300502 989295 300554 989301
rect 300502 989237 300554 989243
rect 319702 989295 319754 989301
rect 319702 989237 319754 989243
rect 290902 986409 290954 986415
rect 290902 986351 290954 986357
rect 300514 983534 300542 989237
rect 331234 988339 331262 1005221
rect 349666 995147 349694 1007769
rect 434710 1005575 434762 1005581
rect 434710 1005517 434762 1005523
rect 367222 1005427 367274 1005433
rect 367222 1005369 367274 1005375
rect 383638 1005427 383690 1005433
rect 383638 1005369 383690 1005375
rect 359060 1003246 359116 1003255
rect 359060 1003181 359062 1003190
rect 359114 1003181 359116 1003190
rect 362516 1003246 362572 1003255
rect 367234 1003213 367262 1005369
rect 377686 1003281 377738 1003287
rect 377686 1003223 377738 1003229
rect 362516 1003181 362518 1003190
rect 359062 1003149 359114 1003155
rect 362570 1003181 362572 1003190
rect 367222 1003207 367274 1003213
rect 362518 1003149 362570 1003155
rect 367222 1003149 367274 1003155
rect 361268 1002654 361324 1002663
rect 361268 1002589 361270 1002598
rect 361322 1002589 361324 1002598
rect 368854 1002615 368906 1002621
rect 361270 1002557 361322 1002563
rect 368854 1002557 368906 1002563
rect 361846 1002541 361898 1002547
rect 361844 1002506 361846 1002515
rect 368662 1002541 368714 1002547
rect 361898 1002506 361900 1002515
rect 368662 1002483 368714 1002489
rect 361844 1002441 361900 1002450
rect 363478 1002393 363530 1002399
rect 362900 1002358 362956 1002367
rect 362900 1002293 362902 1002302
rect 362954 1002293 362956 1002302
rect 363476 1002358 363478 1002367
rect 363530 1002358 363532 1002367
rect 363476 1002293 363532 1002302
rect 362902 1002261 362954 1002267
rect 356374 1000913 356426 1000919
rect 356372 1000878 356374 1000887
rect 356426 1000878 356428 1000887
rect 356372 1000813 356428 1000822
rect 360212 1000878 360268 1000887
rect 360212 1000813 360214 1000822
rect 360266 1000813 360268 1000822
rect 360214 1000781 360266 1000787
rect 357142 999433 357194 999439
rect 357044 999398 357100 999407
rect 357100 999381 357142 999384
rect 357100 999375 357194 999381
rect 357100 999356 357182 999375
rect 357044 999333 357100 999342
rect 364532 999250 364588 999259
rect 364532 999185 364534 999194
rect 364586 999185 364588 999194
rect 364534 999153 364586 999159
rect 364546 997663 364574 999153
rect 365204 997770 365260 997779
rect 365204 997705 365206 997714
rect 365258 997705 365260 997714
rect 365206 997673 365258 997679
rect 364534 997657 364586 997663
rect 364534 997599 364586 997605
rect 368674 996553 368702 1002483
rect 368758 1002319 368810 1002325
rect 368758 1002261 368810 1002267
rect 368770 997145 368798 1002261
rect 368866 998699 368894 1002557
rect 377110 1002393 377162 1002399
rect 377110 1002335 377162 1002341
rect 377122 999439 377150 1002335
rect 377698 1002325 377726 1003223
rect 377686 1002319 377738 1002325
rect 377686 1002261 377738 1002267
rect 383446 1002319 383498 1002325
rect 383446 1002261 383498 1002267
rect 377206 1000913 377258 1000919
rect 377206 1000855 377258 1000861
rect 377110 999433 377162 999439
rect 377110 999375 377162 999381
rect 368854 998693 368906 998699
rect 368854 998635 368906 998641
rect 374518 998693 374570 998699
rect 374518 998635 374570 998641
rect 368758 997139 368810 997145
rect 368758 997081 368810 997087
rect 368662 996547 368714 996553
rect 368662 996489 368714 996495
rect 363958 996473 364010 996479
rect 363958 996415 364010 996421
rect 363970 996035 363998 996415
rect 368662 996177 368714 996183
rect 368662 996119 368714 996125
rect 363958 996029 364010 996035
rect 363956 995994 363958 996003
rect 364010 995994 364012 996003
rect 363956 995929 364012 995938
rect 358100 995846 358156 995855
rect 358100 995781 358156 995790
rect 366164 995846 366220 995855
rect 366164 995781 366220 995790
rect 366740 995846 366796 995855
rect 366740 995781 366742 995790
rect 349654 995141 349706 995147
rect 349654 995083 349706 995089
rect 358114 994523 358142 995781
rect 366178 995739 366206 995781
rect 366794 995781 366796 995790
rect 366742 995749 366794 995755
rect 366166 995733 366218 995739
rect 358196 995698 358252 995707
rect 358252 995656 358526 995684
rect 368674 995707 368702 996119
rect 371540 995846 371596 995855
rect 371540 995781 371596 995790
rect 371638 995807 371690 995813
rect 366166 995675 366218 995681
rect 368660 995698 368716 995707
rect 358196 995633 358252 995642
rect 358498 994819 358526 995656
rect 368660 995633 368716 995642
rect 365780 995550 365836 995559
rect 365780 995485 365836 995494
rect 358484 994810 358540 994819
rect 358484 994745 358540 994754
rect 358100 994514 358156 994523
rect 358100 994449 358156 994458
rect 365794 993667 365822 995485
rect 365782 993661 365834 993667
rect 365782 993603 365834 993609
rect 348406 993513 348458 993519
rect 348458 993461 348542 993464
rect 348406 993455 348542 993461
rect 348418 993445 348542 993455
rect 348418 993439 348554 993445
rect 348418 993436 348502 993439
rect 348502 993381 348554 993387
rect 362902 993365 362954 993371
rect 362900 993330 362902 993339
rect 362954 993330 362956 993339
rect 362900 993265 362956 993274
rect 371554 989375 371582 995781
rect 371638 995749 371690 995755
rect 371650 989449 371678 995749
rect 371734 995733 371786 995739
rect 371734 995675 371786 995681
rect 371638 989443 371690 989449
rect 371638 989385 371690 989391
rect 349174 989369 349226 989375
rect 349174 989311 349226 989317
rect 371542 989369 371594 989375
rect 371542 989311 371594 989317
rect 331222 988333 331274 988339
rect 331222 988275 331274 988281
rect 332566 988333 332618 988339
rect 332566 988275 332618 988281
rect 316726 988111 316778 988117
rect 316726 988053 316778 988059
rect 316738 983534 316766 988053
rect 332578 983548 332606 988275
rect 332578 983520 332976 983548
rect 349186 983534 349214 989311
rect 371746 989301 371774 995675
rect 374530 993741 374558 998635
rect 377218 997885 377246 1000855
rect 383158 999359 383210 999365
rect 383158 999301 383210 999307
rect 380182 999211 380234 999217
rect 380182 999153 380234 999159
rect 377206 997879 377258 997885
rect 377206 997821 377258 997827
rect 377110 997139 377162 997145
rect 377110 997081 377162 997087
rect 377122 995115 377150 997081
rect 377206 996547 377258 996553
rect 377206 996489 377258 996495
rect 377218 995707 377246 996489
rect 380194 996109 380222 999153
rect 383062 997879 383114 997885
rect 383062 997821 383114 997827
rect 380182 996103 380234 996109
rect 380182 996045 380234 996051
rect 383074 995855 383102 997821
rect 383060 995846 383116 995855
rect 383060 995781 383116 995790
rect 377204 995698 377260 995707
rect 377204 995633 377260 995642
rect 383170 995591 383198 999301
rect 383458 995887 383486 1002261
rect 383650 1001012 383678 1005369
rect 434614 1005279 434666 1005285
rect 434614 1005221 434666 1005227
rect 426068 1003246 426124 1003255
rect 426068 1003181 426070 1003190
rect 426122 1003181 426124 1003190
rect 429236 1003246 429292 1003255
rect 434626 1003213 434654 1005221
rect 429236 1003181 429238 1003190
rect 426070 1003149 426122 1003155
rect 429290 1003181 429292 1003190
rect 434614 1003207 434666 1003213
rect 429238 1003149 429290 1003155
rect 434614 1003149 434666 1003155
rect 425396 1003098 425452 1003107
rect 430292 1003098 430348 1003107
rect 425396 1003033 425398 1003042
rect 425450 1003033 425452 1003042
rect 430198 1003059 430250 1003065
rect 425398 1003001 425450 1003007
rect 430292 1003033 430294 1003042
rect 430198 1003001 430250 1003007
rect 430346 1003033 430348 1003042
rect 430294 1003001 430346 1003007
rect 424342 1002985 424394 1002991
rect 424340 1002950 424342 1002959
rect 424394 1002950 424396 1002959
rect 424340 1002885 424396 1002894
rect 428756 1002950 428812 1002959
rect 428756 1002885 428758 1002894
rect 428810 1002885 428812 1002894
rect 428758 1002853 428810 1002859
rect 428278 1002837 428330 1002843
rect 423764 1002802 423820 1002811
rect 423764 1002737 423766 1002746
rect 423818 1002737 423820 1002746
rect 428276 1002802 428278 1002811
rect 428330 1002802 428332 1002811
rect 428276 1002737 428332 1002746
rect 423766 1002705 423818 1002711
rect 424822 1002689 424874 1002695
rect 424820 1002654 424822 1002663
rect 424874 1002654 424876 1002663
rect 424820 1002589 424876 1002598
rect 427700 1002654 427756 1002663
rect 427700 1002589 427702 1002598
rect 427754 1002589 427756 1002598
rect 427702 1002557 427754 1002563
rect 426646 1002541 426698 1002547
rect 426644 1002506 426646 1002515
rect 426698 1002506 426700 1002515
rect 426644 1002441 426700 1002450
rect 427124 1002506 427180 1002515
rect 427124 1002441 427126 1002450
rect 427178 1002441 427180 1002450
rect 427126 1002409 427178 1002415
rect 430210 1002325 430238 1003001
rect 434722 1002917 434750 1005517
rect 434902 1005427 434954 1005433
rect 434902 1005369 434954 1005375
rect 434806 1005205 434858 1005211
rect 434806 1005147 434858 1005153
rect 434710 1002911 434762 1002917
rect 434710 1002853 434762 1002859
rect 434818 1002843 434846 1005147
rect 434914 1003065 434942 1005369
rect 434902 1003059 434954 1003065
rect 434902 1003001 434954 1003007
rect 434806 1002837 434858 1002843
rect 434806 1002779 434858 1002785
rect 435010 1002399 435038 1008033
rect 435188 1005910 435244 1005919
rect 435188 1005845 435244 1005854
rect 465716 1005910 465772 1005919
rect 465716 1005845 465772 1005854
rect 435092 1005170 435148 1005179
rect 435092 1005105 435148 1005114
rect 435106 1002547 435134 1005105
rect 435202 1002621 435230 1005845
rect 459286 1005427 459338 1005433
rect 459286 1005369 459338 1005375
rect 436918 1005353 436970 1005359
rect 436918 1005295 436970 1005301
rect 435190 1002615 435242 1002621
rect 435190 1002557 435242 1002563
rect 435094 1002541 435146 1002547
rect 435094 1002483 435146 1002489
rect 431926 1002393 431978 1002399
rect 431924 1002358 431926 1002367
rect 434998 1002393 435050 1002399
rect 431978 1002358 431980 1002367
rect 430198 1002319 430250 1002325
rect 434998 1002335 435050 1002341
rect 431924 1002293 431980 1002302
rect 430198 1002261 430250 1002267
rect 383650 1000984 383774 1001012
rect 383638 1000839 383690 1000845
rect 383638 1000781 383690 1000787
rect 383542 999433 383594 999439
rect 383542 999375 383594 999381
rect 383446 995881 383498 995887
rect 383446 995823 383498 995829
rect 383554 995739 383582 999375
rect 383650 995813 383678 1000781
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 383542 995733 383594 995739
rect 383542 995675 383594 995681
rect 383746 995665 383774 1000984
rect 429910 1000913 429962 1000919
rect 429908 1000878 429910 1000887
rect 429962 1000878 429964 1000887
rect 429908 1000813 429964 1000822
rect 430964 1000878 431020 1000887
rect 430964 1000813 430966 1000822
rect 431018 1000813 431020 1000822
rect 430966 1000781 431018 1000787
rect 432596 996290 432652 996299
rect 432596 996225 432598 996234
rect 432650 996225 432652 996234
rect 432598 996193 432650 996199
rect 432502 996177 432554 996183
rect 432500 996142 432502 996151
rect 432554 996142 432556 996151
rect 435010 996109 435038 1002335
rect 432500 996077 432556 996086
rect 434998 996103 435050 996109
rect 434998 996045 435050 996051
rect 436930 996035 436958 1005295
rect 443734 1005205 443786 1005211
rect 443540 1005170 443596 1005179
rect 443734 1005147 443786 1005153
rect 443540 1005105 443596 1005114
rect 443554 1003731 443582 1005105
rect 443542 1003725 443594 1003731
rect 443542 1003667 443594 1003673
rect 439222 1003207 439274 1003213
rect 439222 1003149 439274 1003155
rect 439126 1003059 439178 1003065
rect 439126 1003001 439178 1003007
rect 439138 1002769 439166 1003001
rect 439126 1002763 439178 1002769
rect 439126 1002705 439178 1002711
rect 439234 1002695 439262 1003149
rect 439222 1002689 439274 1002695
rect 439222 1002631 439274 1002637
rect 443638 1002467 443690 1002473
rect 443638 1002409 443690 1002415
rect 443650 1000993 443678 1002409
rect 443638 1000987 443690 1000993
rect 443638 1000929 443690 1000935
rect 430966 996029 431018 996035
rect 430964 995994 430966 996003
rect 436918 996029 436970 996035
rect 431018 995994 431020 996003
rect 436918 995971 436970 995977
rect 437876 995994 437932 996003
rect 430964 995929 431020 995938
rect 437876 995929 437932 995938
rect 393716 995846 393772 995855
rect 384994 995813 385296 995832
rect 388834 995813 388992 995832
rect 384982 995807 385296 995813
rect 385034 995804 385296 995807
rect 388822 995807 388992 995813
rect 384982 995749 385034 995755
rect 388874 995804 388992 995807
rect 422132 995846 422188 995855
rect 393772 995804 393984 995832
rect 393716 995781 393772 995790
rect 422132 995781 422188 995790
rect 388822 995749 388874 995755
rect 386038 995733 386090 995739
rect 384418 995665 384672 995684
rect 383734 995659 383786 995665
rect 383734 995601 383786 995607
rect 384406 995659 384672 995665
rect 384458 995656 384672 995659
rect 385968 995681 386038 995684
rect 385968 995675 386090 995681
rect 387476 995698 387532 995707
rect 385968 995656 386078 995675
rect 387532 995656 387792 995684
rect 390192 995656 390494 995684
rect 387476 995633 387532 995642
rect 384406 995601 384458 995607
rect 383158 995585 383210 995591
rect 383158 995527 383210 995533
rect 383158 995437 383210 995443
rect 383158 995379 383210 995385
rect 377108 995106 377164 995115
rect 377108 995041 377164 995050
rect 374518 993735 374570 993741
rect 374518 993677 374570 993683
rect 382966 993365 383018 993371
rect 382964 993330 382966 993339
rect 383018 993330 383020 993339
rect 383170 993316 383198 995379
rect 388354 994967 388382 995522
rect 389410 995508 389664 995536
rect 388340 994958 388396 994967
rect 388340 994893 388396 994902
rect 389410 994819 389438 995508
rect 390466 995443 390494 995656
rect 392374 995585 392426 995591
rect 390864 995522 391166 995536
rect 392426 995533 392688 995536
rect 392374 995527 392688 995533
rect 390850 995508 391166 995522
rect 390454 995437 390506 995443
rect 390454 995379 390506 995385
rect 389396 994810 389452 994819
rect 389396 994745 389452 994754
rect 390850 994375 390878 995508
rect 391138 995411 391166 995508
rect 391124 995402 391180 995411
rect 391124 995337 391180 995346
rect 390836 994366 390892 994375
rect 390836 994301 390892 994310
rect 392098 993741 392126 995522
rect 392386 995508 392688 995527
rect 393058 995508 393312 995536
rect 393058 994523 393086 995508
rect 395170 994671 395198 995522
rect 395156 994662 395212 994671
rect 395156 994597 395212 994606
rect 393044 994514 393100 994523
rect 393044 994449 393100 994458
rect 396322 994375 396350 995522
rect 396994 995115 397022 995522
rect 396980 995106 397036 995115
rect 396980 995041 397036 995050
rect 396308 994366 396364 994375
rect 396308 994301 396364 994310
rect 392086 993735 392138 993741
rect 392086 993677 392138 993683
rect 398818 993667 398846 995522
rect 403126 995437 403178 995443
rect 403126 995379 403178 995385
rect 398806 993661 398858 993667
rect 398806 993603 398858 993609
rect 403138 993445 403166 995379
rect 408982 993513 409034 993519
rect 408898 993461 408982 993464
rect 408898 993455 409034 993461
rect 408898 993445 409022 993455
rect 403126 993439 403178 993445
rect 403126 993381 403178 993387
rect 408886 993439 409022 993445
rect 408938 993436 409022 993439
rect 408886 993381 408938 993387
rect 383074 993297 383198 993316
rect 382964 993265 383020 993274
rect 383062 993291 383198 993297
rect 383114 993288 383198 993291
rect 383062 993233 383114 993239
rect 422146 992779 422174 995781
rect 437780 995698 437836 995707
rect 437780 995633 437836 995642
rect 423380 993626 423436 993635
rect 423380 993561 423382 993570
rect 423434 993561 423436 993570
rect 423382 993529 423434 993535
rect 422134 992773 422186 992779
rect 422134 992715 422186 992721
rect 426262 992773 426314 992779
rect 426262 992715 426314 992721
rect 397846 989443 397898 989449
rect 397846 989385 397898 989391
rect 365398 989295 365450 989301
rect 365398 989237 365450 989243
rect 371734 989295 371786 989301
rect 371734 989237 371786 989243
rect 365410 983534 365438 989237
rect 381622 988037 381674 988043
rect 381622 987979 381674 987985
rect 381634 983534 381662 987979
rect 397858 983534 397886 989385
rect 414070 989369 414122 989375
rect 414070 989311 414122 989317
rect 414082 983534 414110 989311
rect 426274 983529 426302 992715
rect 437794 989449 437822 995633
rect 437782 989443 437834 989449
rect 437782 989385 437834 989391
rect 437890 989375 437918 995929
rect 437972 995550 438028 995559
rect 437972 995485 438028 995494
rect 437878 989369 437930 989375
rect 437878 989311 437930 989317
rect 437986 989301 438014 995485
rect 443746 993667 443774 1005147
rect 449206 1003133 449258 1003139
rect 449206 1003075 449258 1003081
rect 449218 1002325 449246 1003075
rect 449206 1002319 449258 1002325
rect 449206 1002261 449258 1002267
rect 459298 999439 459326 1005369
rect 463798 1003725 463850 1003731
rect 463798 1003667 463850 1003673
rect 463510 1003059 463562 1003065
rect 463510 1003001 463562 1003007
rect 459286 999433 459338 999439
rect 459286 999375 459338 999381
rect 463522 997219 463550 1003001
rect 463606 1002985 463658 1002991
rect 463606 1002927 463658 1002933
rect 463510 997213 463562 997219
rect 463510 997155 463562 997161
rect 463618 996572 463646 1002927
rect 463618 996544 463742 996572
rect 463714 996151 463742 996544
rect 463700 996142 463756 996151
rect 463700 996077 463756 996086
rect 463810 995707 463838 1003667
rect 465730 1001067 465758 1005845
rect 467062 1003281 467114 1003287
rect 467062 1003223 467114 1003229
rect 466582 1003207 466634 1003213
rect 466582 1003149 466634 1003155
rect 465718 1001061 465770 1001067
rect 465718 1001003 465770 1001009
rect 464758 999359 464810 999365
rect 464758 999301 464810 999307
rect 463796 995698 463852 995707
rect 463796 995633 463852 995642
rect 464770 994819 464798 999301
rect 465334 997213 465386 997219
rect 465334 997155 465386 997161
rect 465346 995559 465374 997155
rect 466594 995591 466622 1003149
rect 466582 995585 466634 995591
rect 465332 995550 465388 995559
rect 466582 995527 466634 995533
rect 465332 995485 465388 995494
rect 467074 994967 467102 1003223
rect 467830 1003133 467882 1003139
rect 467830 1003075 467882 1003081
rect 467842 996003 467870 1003075
rect 470818 996109 470846 1008033
rect 472150 1005575 472202 1005581
rect 472150 1005517 472202 1005523
rect 471382 1005353 471434 1005359
rect 471382 1005295 471434 1005301
rect 470806 996103 470858 996109
rect 470806 996045 470858 996051
rect 467828 995994 467884 996003
rect 471394 995961 471422 1005295
rect 467828 995929 467884 995938
rect 471382 995955 471434 995961
rect 471382 995897 471434 995903
rect 472162 995115 472190 1005517
rect 472246 1005279 472298 1005285
rect 472246 1005221 472298 1005227
rect 472258 995855 472286 1005221
rect 518614 1003281 518666 1003287
rect 518614 1003223 518666 1003229
rect 502390 1003133 502442 1003139
rect 501332 1003098 501388 1003107
rect 501332 1003033 501334 1003042
rect 501386 1003033 501388 1003042
rect 502388 1003098 502390 1003107
rect 502966 1003133 503018 1003139
rect 502442 1003098 502444 1003107
rect 502388 1003033 502444 1003042
rect 502964 1003098 502966 1003107
rect 503018 1003098 503020 1003107
rect 502964 1003033 503020 1003042
rect 504020 1003098 504076 1003107
rect 504020 1003033 504022 1003042
rect 501334 1003001 501386 1003007
rect 504074 1003033 504076 1003042
rect 518422 1003059 518474 1003065
rect 504022 1003001 504074 1003007
rect 518422 1003001 518474 1003007
rect 503446 1002393 503498 1002399
rect 503444 1002358 503446 1002367
rect 514006 1002393 514058 1002399
rect 503498 1002358 503500 1002367
rect 489526 1002319 489578 1002325
rect 514006 1002335 514058 1002341
rect 503444 1002293 503500 1002302
rect 489526 1002261 489578 1002267
rect 472630 1001061 472682 1001067
rect 472682 1001009 472766 1001012
rect 472630 1001003 472766 1001009
rect 472438 1000987 472490 1000993
rect 472642 1000984 472766 1001003
rect 472438 1000929 472490 1000935
rect 472450 995887 472478 1000929
rect 472630 1000913 472682 1000919
rect 472630 1000855 472682 1000861
rect 472534 1000839 472586 1000845
rect 472534 1000781 472586 1000787
rect 472438 995881 472490 995887
rect 472244 995846 472300 995855
rect 472438 995823 472490 995829
rect 472244 995781 472300 995790
rect 472546 995739 472574 1000781
rect 472642 995813 472670 1000855
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 472738 995665 472766 1000984
rect 476468 995846 476524 995855
rect 473314 995813 473664 995832
rect 473302 995807 473664 995813
rect 473354 995804 473664 995807
rect 481460 995846 481516 995855
rect 476524 995804 476784 995832
rect 476962 995813 477360 995832
rect 476950 995807 477360 995813
rect 476468 995781 476524 995790
rect 473302 995749 473354 995755
rect 477002 995804 477360 995807
rect 482036 995846 482092 995855
rect 481516 995804 481680 995832
rect 481460 995781 481516 995790
rect 482092 995804 482352 995832
rect 482036 995781 482092 995790
rect 476950 995749 477002 995755
rect 474646 995733 474698 995739
rect 474082 995665 474336 995684
rect 477716 995698 477772 995707
rect 474698 995681 474960 995684
rect 474646 995675 474960 995681
rect 472726 995659 472778 995665
rect 472726 995601 472778 995607
rect 474070 995659 474336 995665
rect 474122 995656 474336 995659
rect 474658 995656 474960 995675
rect 482708 995698 482764 995707
rect 477772 995656 477984 995684
rect 478402 995665 478656 995684
rect 478390 995659 478656 995665
rect 477716 995633 477772 995642
rect 474070 995601 474122 995607
rect 478442 995656 478656 995659
rect 482764 995656 482976 995684
rect 482708 995633 482764 995642
rect 478390 995601 478442 995607
rect 478100 995254 478156 995263
rect 478100 995189 478156 995198
rect 472148 995106 472204 995115
rect 472148 995041 472204 995050
rect 467060 994958 467116 994967
rect 467060 994893 467116 994902
rect 464756 994810 464812 994819
rect 464756 994745 464812 994754
rect 478114 994671 478142 995189
rect 478100 994662 478156 994671
rect 478100 994597 478156 994606
rect 479170 994185 479198 995522
rect 479842 994671 479870 995522
rect 481090 995115 481118 995522
rect 481076 995106 481132 995115
rect 481076 995041 481132 995050
rect 484162 994967 484190 995522
rect 485376 995508 485630 995536
rect 484148 994958 484204 994967
rect 484148 994893 484204 994902
rect 479828 994662 479884 994671
rect 479828 994597 479884 994606
rect 485602 994523 485630 995508
rect 485986 994819 486014 995522
rect 485972 994810 486028 994819
rect 485972 994745 486028 994754
rect 485588 994514 485644 994523
rect 485588 994449 485644 994458
rect 463702 994179 463754 994185
rect 463702 994121 463754 994127
rect 479158 994179 479210 994185
rect 479158 994121 479210 994127
rect 443734 993661 443786 993667
rect 443444 993626 443500 993635
rect 443734 993603 443786 993609
rect 443444 993561 443500 993570
rect 443458 993519 443486 993561
rect 443446 993513 443498 993519
rect 443446 993455 443498 993461
rect 449206 993513 449258 993519
rect 449258 993461 449438 993464
rect 449206 993455 449438 993461
rect 449218 993445 449438 993455
rect 463714 993445 463742 994121
rect 479170 993445 479198 994121
rect 487810 993667 487838 995522
rect 487798 993661 487850 993667
rect 487798 993603 487850 993609
rect 489538 993445 489566 1002261
rect 506230 1001505 506282 1001511
rect 506228 1001470 506230 1001479
rect 506282 1001470 506284 1001479
rect 506228 1001405 506284 1001414
rect 507860 1001026 507916 1001035
rect 507860 1000961 507862 1000970
rect 507914 1000961 507916 1000970
rect 512660 1001026 512716 1001035
rect 512660 1000961 512662 1000970
rect 507862 1000929 507914 1000935
rect 512714 1000961 512716 1000970
rect 512662 1000929 512714 1000935
rect 514018 1000887 514046 1002335
rect 500756 1000878 500812 1000887
rect 500756 1000813 500758 1000822
rect 500810 1000813 500812 1000822
rect 514004 1000878 514060 1000887
rect 514004 1000813 514060 1000822
rect 500758 1000781 500810 1000787
rect 506900 1000730 506956 1000739
rect 506900 1000665 506902 1000674
rect 506954 1000665 506956 1000674
rect 512084 1000730 512140 1000739
rect 512084 1000665 512086 1000674
rect 506902 1000633 506954 1000639
rect 512138 1000665 512140 1000674
rect 512086 1000633 512138 1000639
rect 518434 999851 518462 1003001
rect 518518 1001505 518570 1001511
rect 518518 1001447 518570 1001453
rect 518420 999842 518476 999851
rect 518420 999777 518476 999786
rect 502006 999729 502058 999735
rect 502004 999694 502006 999703
rect 512086 999729 512138 999735
rect 502058 999694 502060 999703
rect 502004 999629 502060 999638
rect 512084 999694 512086 999703
rect 512138 999694 512140 999703
rect 512084 999629 512140 999638
rect 504694 999581 504746 999587
rect 504692 999546 504694 999555
rect 512086 999581 512138 999587
rect 504746 999546 504748 999555
rect 504692 999481 504748 999490
rect 512084 999546 512086 999555
rect 512138 999546 512140 999555
rect 512084 999481 512140 999490
rect 500182 999433 500234 999439
rect 500180 999398 500182 999407
rect 515830 999433 515882 999439
rect 500234 999398 500236 999407
rect 518530 999407 518558 1001447
rect 515830 999375 515882 999381
rect 518516 999398 518572 999407
rect 500180 999333 500236 999342
rect 507286 996621 507338 996627
rect 505652 996586 505708 996595
rect 505652 996521 505654 996530
rect 505706 996521 505708 996530
rect 507284 996586 507286 996595
rect 507338 996586 507340 996595
rect 507284 996521 507340 996530
rect 505654 996489 505706 996495
rect 508340 996290 508396 996299
rect 508340 996225 508342 996234
rect 508394 996225 508396 996234
rect 508342 996193 508394 996199
rect 508354 995961 508382 996193
rect 509590 996177 509642 996183
rect 508532 996142 508588 996151
rect 508532 996077 508534 996086
rect 508586 996077 508588 996086
rect 509588 996142 509590 996151
rect 509642 996142 509644 996151
rect 509588 996077 509644 996086
rect 508534 996045 508586 996051
rect 510548 995994 510604 996003
rect 508342 995955 508394 995961
rect 510548 995929 510550 995938
rect 508342 995897 508394 995903
rect 510602 995929 510604 995938
rect 515540 995994 515596 996003
rect 515540 995929 515596 995938
rect 515734 995955 515786 995961
rect 510550 995897 510602 995903
rect 511124 995846 511180 995855
rect 511124 995781 511126 995790
rect 511178 995781 511180 995790
rect 511126 995749 511178 995755
rect 449218 993439 449450 993445
rect 449218 993436 449398 993439
rect 449398 993381 449450 993387
rect 463702 993439 463754 993445
rect 463702 993381 463754 993387
rect 479158 993439 479210 993445
rect 479158 993381 479210 993387
rect 489526 993439 489578 993445
rect 489526 993381 489578 993387
rect 462742 989443 462794 989449
rect 462742 989385 462794 989391
rect 430294 989295 430346 989301
rect 430294 989237 430346 989243
rect 437974 989295 438026 989301
rect 437974 989237 438026 989243
rect 430306 983534 430334 989237
rect 446518 987963 446570 987969
rect 446518 987905 446570 987911
rect 446530 983534 446558 987905
rect 462754 983534 462782 989385
rect 515554 989375 515582 995929
rect 515734 995897 515786 995903
rect 515638 995807 515690 995813
rect 515638 995749 515690 995755
rect 515650 989449 515678 995749
rect 515638 989443 515690 989449
rect 515638 989385 515690 989391
rect 478966 989369 479018 989375
rect 478966 989311 479018 989317
rect 515542 989369 515594 989375
rect 515542 989311 515594 989317
rect 478978 983534 479006 989311
rect 515746 989301 515774 995897
rect 495190 989295 495242 989301
rect 495190 989237 495242 989243
rect 515734 989295 515786 989301
rect 515734 989237 515786 989243
rect 495202 983534 495230 989237
rect 511414 987889 511466 987895
rect 511414 987831 511466 987837
rect 511426 983534 511454 987831
rect 515842 983603 515870 999375
rect 518516 999333 518572 999342
rect 518422 996177 518474 996183
rect 518422 996119 518474 996125
rect 518434 995707 518462 996119
rect 518420 995698 518476 995707
rect 518420 995633 518476 995642
rect 518626 995443 518654 1003223
rect 518806 1003207 518858 1003213
rect 518806 1003149 518858 1003155
rect 518710 1003133 518762 1003139
rect 518710 1003075 518762 1003081
rect 518614 995437 518666 995443
rect 518614 995379 518666 995385
rect 518722 995369 518750 1003075
rect 518818 995517 518846 1003149
rect 554902 1002985 554954 1002991
rect 554900 1002950 554902 1002959
rect 573046 1002985 573098 1002991
rect 554954 1002950 554956 1002959
rect 573046 1002927 573098 1002933
rect 554900 1002885 554956 1002894
rect 554326 1002837 554378 1002843
rect 554324 1002802 554326 1002811
rect 572854 1002837 572906 1002843
rect 554378 1002802 554380 1002811
rect 572854 1002779 572906 1002785
rect 554324 1002737 554380 1002746
rect 553748 1002654 553804 1002663
rect 553748 1002589 553750 1002598
rect 553802 1002589 553804 1002598
rect 553750 1002557 553802 1002563
rect 553270 1002393 553322 1002399
rect 553268 1002358 553270 1002367
rect 567478 1002393 567530 1002399
rect 553322 1002358 553324 1002367
rect 519862 1002319 519914 1002325
rect 553268 1002293 553324 1002302
rect 555380 1002358 555436 1002367
rect 567478 1002335 567530 1002341
rect 555380 1002293 555382 1002302
rect 519862 1002261 519914 1002267
rect 555434 1002293 555436 1002302
rect 567382 1002319 567434 1002325
rect 555382 1002261 555434 1002267
rect 567382 1002261 567434 1002267
rect 518806 995511 518858 995517
rect 518806 995453 518858 995459
rect 518710 995363 518762 995369
rect 518710 995305 518762 995311
rect 519874 995147 519902 1002261
rect 557782 1001357 557834 1001363
rect 557780 1001322 557782 1001331
rect 557834 1001322 557836 1001331
rect 557780 1001257 557836 1001266
rect 523796 1001026 523852 1001035
rect 523796 1000961 523852 1000970
rect 523508 1000878 523564 1000887
rect 523318 1000839 523370 1000845
rect 523508 1000813 523564 1000822
rect 523318 1000781 523370 1000787
rect 521206 996547 521258 996553
rect 521206 996489 521258 996495
rect 521218 995855 521246 996489
rect 521204 995846 521260 995855
rect 521204 995781 521260 995790
rect 521300 995550 521356 995559
rect 521300 995485 521356 995494
rect 519862 995141 519914 995147
rect 519862 995083 519914 995089
rect 521314 993815 521342 995485
rect 523330 995221 523358 1000781
rect 523414 996621 523466 996627
rect 523414 996563 523466 996569
rect 523426 995295 523454 996563
rect 523522 995707 523550 1000813
rect 523700 999694 523756 999703
rect 523700 999629 523756 999638
rect 523604 999398 523660 999407
rect 523604 999333 523660 999342
rect 523508 995698 523564 995707
rect 523508 995633 523564 995642
rect 523618 995591 523646 999333
rect 523714 995961 523742 999629
rect 523702 995955 523754 995961
rect 523702 995897 523754 995903
rect 523810 995665 523838 1000961
rect 552310 1000913 552362 1000919
rect 552308 1000878 552310 1000887
rect 552362 1000878 552364 1000887
rect 552308 1000813 552364 1000822
rect 552884 1000878 552940 1000887
rect 552940 1000845 553022 1000864
rect 552940 1000839 553034 1000845
rect 552940 1000836 552982 1000839
rect 552884 1000813 552940 1000822
rect 552982 1000781 553034 1000787
rect 523988 1000730 524044 1000739
rect 523988 1000665 524044 1000674
rect 523892 999842 523948 999851
rect 523892 999777 523948 999786
rect 523906 995887 523934 999777
rect 523894 995881 523946 995887
rect 523894 995823 523946 995829
rect 524002 995739 524030 1000665
rect 524084 999546 524140 999555
rect 524084 999481 524140 999490
rect 524098 995832 524126 999481
rect 557206 999137 557258 999143
rect 557204 999102 557206 999111
rect 557258 999102 557260 999111
rect 557204 999037 557260 999046
rect 558838 998989 558890 998995
rect 558836 998954 558838 998963
rect 558890 998954 558892 998963
rect 558836 998889 558892 998898
rect 555956 997770 556012 997779
rect 555956 997705 555958 997714
rect 556010 997705 556012 997714
rect 555958 997673 556010 997679
rect 567394 997589 567422 1002261
rect 567490 997663 567518 1002335
rect 571030 1001357 571082 1001363
rect 571030 1001299 571082 1001305
rect 567478 997657 567530 997663
rect 567478 997599 567530 997605
rect 567382 997583 567434 997589
rect 567382 997525 567434 997531
rect 571042 997515 571070 1001299
rect 571030 997509 571082 997515
rect 558164 997474 558220 997483
rect 571030 997451 571082 997457
rect 558164 997409 558166 997418
rect 558218 997409 558220 997418
rect 558166 997377 558218 997383
rect 559414 997361 559466 997367
rect 559412 997326 559414 997335
rect 559466 997326 559468 997335
rect 559412 997261 559468 997270
rect 561046 996177 561098 996183
rect 561044 996142 561046 996151
rect 561098 996142 561100 996151
rect 559798 996103 559850 996109
rect 561044 996077 561100 996086
rect 559798 996045 559850 996051
rect 559810 995855 559838 996045
rect 560182 996029 560234 996035
rect 560182 995971 560234 995977
rect 561908 995994 561964 996003
rect 532244 995846 532300 995855
rect 524098 995813 524222 995832
rect 525346 995813 525744 995832
rect 528418 995813 528768 995832
rect 529858 995813 530064 995832
rect 524098 995807 524234 995813
rect 524098 995804 524182 995807
rect 524182 995749 524234 995755
rect 525334 995807 525744 995813
rect 525386 995804 525744 995807
rect 528406 995807 528768 995813
rect 525334 995749 525386 995755
rect 528458 995804 528768 995807
rect 529846 995807 530064 995813
rect 528406 995749 528458 995755
rect 529898 995804 530064 995807
rect 530592 995804 530750 995832
rect 529846 995749 529898 995755
rect 523990 995733 524042 995739
rect 523990 995675 524042 995681
rect 524758 995733 524810 995739
rect 529076 995698 529132 995707
rect 524810 995681 525072 995684
rect 524758 995675 525072 995681
rect 523798 995659 523850 995665
rect 524770 995656 525072 995675
rect 526114 995665 526368 995684
rect 526102 995659 526368 995665
rect 523798 995601 523850 995607
rect 526154 995656 526368 995659
rect 529132 995656 529392 995684
rect 529076 995633 529132 995642
rect 526102 995601 526154 995607
rect 523606 995585 523658 995591
rect 523606 995527 523658 995533
rect 527830 995585 527882 995591
rect 527882 995533 528192 995536
rect 527830 995527 528192 995533
rect 527842 995508 528192 995527
rect 523414 995289 523466 995295
rect 523414 995231 523466 995237
rect 523318 995215 523370 995221
rect 523318 995157 523370 995163
rect 530722 995147 530750 995804
rect 550484 995846 550540 995855
rect 532300 995804 532512 995832
rect 532244 995781 532300 995790
rect 550484 995781 550540 995790
rect 559796 995846 559852 995855
rect 559796 995781 559798 995790
rect 550498 995559 550526 995781
rect 559850 995781 559852 995790
rect 559798 995749 559850 995755
rect 560194 995707 560222 995971
rect 561908 995929 561910 995938
rect 561962 995929 561964 995938
rect 569782 995955 569834 995961
rect 561910 995897 561962 995903
rect 569782 995897 569834 995903
rect 564598 995807 564650 995813
rect 564598 995749 564650 995755
rect 555380 995698 555436 995707
rect 555380 995633 555436 995642
rect 560180 995698 560236 995707
rect 560180 995633 560182 995642
rect 550484 995550 550540 995559
rect 530710 995141 530762 995147
rect 530710 995083 530762 995089
rect 531202 994703 531230 995522
rect 532834 995517 533088 995536
rect 532822 995511 533088 995517
rect 532874 995508 533088 995511
rect 533410 995508 533712 995536
rect 532822 995453 532874 995459
rect 533410 995443 533438 995508
rect 533398 995437 533450 995443
rect 533398 995379 533450 995385
rect 534370 995221 534398 995522
rect 535570 995369 535598 995522
rect 535558 995363 535610 995369
rect 535558 995305 535610 995311
rect 534358 995215 534410 995221
rect 534358 995157 534410 995163
rect 532726 995141 532778 995147
rect 532726 995083 532778 995089
rect 524086 994697 524138 994703
rect 524084 994662 524086 994671
rect 531190 994697 531242 994703
rect 524138 994662 524140 994671
rect 531190 994639 531242 994645
rect 524084 994597 524140 994606
rect 521302 993809 521354 993815
rect 521302 993751 521354 993757
rect 531202 993667 531230 994639
rect 532738 993741 532766 995083
rect 536770 994671 536798 995522
rect 537394 995295 537422 995522
rect 538978 995508 539232 995536
rect 537382 995289 537434 995295
rect 537382 995231 537434 995237
rect 536756 994662 536812 994671
rect 536756 994597 536812 994606
rect 538978 993815 539006 995508
rect 550484 995485 550540 995494
rect 555394 995147 555422 995633
rect 560234 995633 560236 995642
rect 564502 995659 564554 995665
rect 560182 995601 560234 995607
rect 564502 995601 564554 995607
rect 561620 995402 561676 995411
rect 561620 995337 561676 995346
rect 555382 995141 555434 995147
rect 555382 995083 555434 995089
rect 561634 993889 561662 995337
rect 561622 993883 561674 993889
rect 561622 993825 561674 993831
rect 538966 993809 539018 993815
rect 538966 993751 539018 993757
rect 532726 993735 532778 993741
rect 532726 993677 532778 993683
rect 531190 993661 531242 993667
rect 531190 993603 531242 993609
rect 527638 989443 527690 989449
rect 527638 989385 527690 989391
rect 515830 983597 515882 983603
rect 515830 983539 515882 983545
rect 527650 983534 527678 989385
rect 543766 989369 543818 989375
rect 543766 989311 543818 989317
rect 543778 983534 543806 989311
rect 560086 989295 560138 989301
rect 560086 989237 560138 989243
rect 560098 983534 560126 989237
rect 564514 986563 564542 995601
rect 564502 986557 564554 986563
rect 564502 986499 564554 986505
rect 564610 986415 564638 995749
rect 569684 995698 569740 995707
rect 569684 995633 569740 995642
rect 565844 995550 565900 995559
rect 565844 995485 565900 995494
rect 565858 986489 565886 995485
rect 569698 989449 569726 995633
rect 569686 989443 569738 989449
rect 569686 989385 569738 989391
rect 569794 989301 569822 995897
rect 569876 995846 569932 995855
rect 569876 995781 569932 995790
rect 569890 989375 569918 995781
rect 572866 994819 572894 1002779
rect 572950 1002615 573002 1002621
rect 572950 1002557 573002 1002563
rect 572962 994967 572990 1002557
rect 573058 995559 573086 1002927
rect 573238 1000913 573290 1000919
rect 573238 1000855 573290 1000861
rect 573044 995550 573100 995559
rect 573044 995485 573100 995494
rect 573250 995263 573278 1000855
rect 575158 1000839 575210 1000845
rect 575158 1000781 575210 1000787
rect 573814 999137 573866 999143
rect 573814 999079 573866 999085
rect 573526 998989 573578 998995
rect 573526 998931 573578 998937
rect 573236 995254 573292 995263
rect 573236 995189 573292 995198
rect 573538 995115 573566 998931
rect 573826 995707 573854 999079
rect 573812 995698 573868 995707
rect 573812 995633 573868 995642
rect 575170 995411 575198 1000781
rect 610678 999803 610730 999809
rect 610678 999745 610730 999751
rect 625846 999803 625898 999809
rect 625846 999745 625898 999751
rect 609046 999729 609098 999735
rect 609046 999671 609098 999677
rect 596278 999581 596330 999587
rect 596278 999523 596330 999529
rect 593302 999507 593354 999513
rect 593302 999449 593354 999455
rect 593314 997737 593342 999449
rect 596182 999433 596234 999439
rect 596182 999375 596234 999381
rect 593302 997731 593354 997737
rect 593302 997673 593354 997679
rect 596194 997663 596222 999375
rect 596182 997657 596234 997663
rect 596182 997599 596234 997605
rect 596290 997589 596318 999523
rect 596278 997583 596330 997589
rect 596278 997525 596330 997531
rect 609058 997441 609086 999671
rect 610582 999655 610634 999661
rect 610582 999597 610634 999603
rect 610594 997515 610622 999597
rect 610582 997509 610634 997515
rect 610582 997451 610634 997457
rect 609046 997435 609098 997441
rect 609046 997377 609098 997383
rect 610690 997367 610718 999745
rect 625750 999729 625802 999735
rect 625750 999671 625802 999677
rect 625858 999680 625886 999745
rect 625654 999655 625706 999661
rect 625654 999597 625706 999603
rect 625558 999581 625610 999587
rect 625558 999523 625610 999529
rect 625462 999433 625514 999439
rect 625462 999375 625514 999381
rect 610678 997361 610730 997367
rect 610678 997303 610730 997309
rect 625474 995961 625502 999375
rect 625462 995955 625514 995961
rect 625462 995897 625514 995903
rect 625570 995665 625598 999523
rect 625666 995887 625694 999597
rect 625654 995881 625706 995887
rect 625654 995823 625706 995829
rect 625762 995739 625790 999671
rect 625858 999652 625982 999680
rect 625846 999507 625898 999513
rect 625846 999449 625898 999455
rect 625858 995813 625886 999449
rect 625846 995807 625898 995813
rect 625846 995749 625898 995755
rect 625750 995733 625802 995739
rect 625750 995675 625802 995681
rect 625558 995659 625610 995665
rect 625558 995601 625610 995607
rect 625954 995591 625982 999652
rect 627106 995813 627504 995832
rect 629602 995813 630000 995832
rect 631522 995813 631824 995832
rect 627094 995807 627504 995813
rect 627146 995804 627504 995807
rect 629590 995807 630000 995813
rect 627094 995749 627146 995755
rect 629642 995804 630000 995807
rect 631510 995807 631824 995813
rect 629590 995749 629642 995755
rect 631562 995804 631824 995807
rect 631510 995749 631562 995755
rect 626518 995733 626570 995739
rect 634004 995698 634060 995707
rect 626570 995681 626880 995684
rect 626518 995675 626880 995681
rect 626530 995656 626880 995675
rect 630178 995665 630576 995684
rect 630166 995659 630576 995665
rect 630218 995656 630576 995659
rect 634060 995656 634320 995684
rect 634004 995633 634060 995642
rect 630166 995601 630218 995607
rect 625942 995585 625994 995591
rect 625942 995527 625994 995533
rect 627862 995585 627914 995591
rect 630932 995550 630988 995559
rect 627914 995533 628176 995536
rect 627862 995527 628176 995533
rect 627874 995508 628176 995527
rect 630988 995508 631200 995536
rect 630932 995485 630988 995494
rect 575156 995402 575212 995411
rect 575156 995337 575212 995346
rect 573524 995106 573580 995115
rect 573524 995041 573580 995050
rect 609046 995067 609098 995073
rect 609046 995009 609098 995015
rect 572948 994958 573004 994967
rect 572948 994893 573004 994902
rect 572852 994810 572908 994819
rect 572852 994745 572908 994754
rect 604628 994366 604684 994375
rect 604628 994301 604684 994310
rect 576308 993922 576364 993931
rect 576308 993857 576364 993866
rect 569878 989369 569930 989375
rect 569878 989311 569930 989317
rect 569782 989295 569834 989301
rect 569782 989237 569834 989243
rect 565846 986483 565898 986489
rect 565846 986425 565898 986431
rect 564598 986409 564650 986415
rect 564598 986351 564650 986357
rect 576322 983534 576350 993857
rect 604642 991873 604670 994301
rect 604726 991959 604778 991965
rect 604726 991901 604778 991907
rect 605782 991959 605834 991965
rect 605782 991901 605834 991907
rect 604738 991873 604766 991901
rect 604642 991845 604766 991873
rect 605794 991669 605822 991901
rect 605782 991663 605834 991669
rect 605782 991605 605834 991611
rect 592438 989443 592490 989449
rect 592438 989385 592490 989391
rect 592450 983534 592478 989385
rect 608758 989369 608810 989375
rect 608758 989311 608810 989317
rect 608770 983534 608798 989311
rect 609058 986637 609086 995009
rect 632386 993741 632414 995522
rect 633024 995508 633086 995536
rect 632374 993735 632426 993741
rect 632374 993677 632426 993683
rect 619798 991663 619850 991669
rect 619798 991605 619850 991611
rect 619810 986711 619838 991605
rect 624982 989295 625034 989301
rect 624982 989237 625034 989243
rect 619798 986705 619850 986711
rect 619798 986647 619850 986653
rect 609046 986631 609098 986637
rect 609046 986573 609098 986579
rect 624994 983534 625022 989237
rect 632386 983751 632414 993677
rect 633058 993667 633086 995508
rect 634594 995508 634896 995536
rect 635266 995508 635520 995536
rect 634594 995411 634622 995508
rect 634580 995402 634636 995411
rect 634580 995337 634636 995346
rect 635266 994967 635294 995508
rect 636130 995263 636158 995522
rect 636116 995254 636172 995263
rect 636116 995189 636172 995198
rect 635252 994958 635308 994967
rect 635252 994893 635308 994902
rect 637378 994819 637406 995522
rect 637364 994810 637420 994819
rect 637364 994745 637420 994754
rect 634292 994662 634348 994671
rect 634292 994597 634348 994606
rect 633046 993661 633098 993667
rect 633046 993603 633098 993609
rect 632374 983745 632426 983751
rect 632374 983687 632426 983693
rect 633058 983677 633086 993603
rect 634306 989301 634334 994597
rect 638530 993931 638558 995522
rect 639202 995115 639230 995522
rect 639188 995106 639244 995115
rect 639188 995041 639244 995050
rect 638516 993922 638572 993931
rect 641026 993889 641054 995522
rect 649366 995141 649418 995147
rect 649366 995083 649418 995089
rect 642260 993922 642316 993931
rect 638516 993857 638572 993866
rect 641014 993883 641066 993889
rect 642260 993857 642316 993866
rect 641014 993825 641066 993831
rect 641108 993774 641164 993783
rect 641108 993709 641164 993718
rect 634294 989295 634346 989301
rect 634294 989237 634346 989243
rect 633046 983671 633098 983677
rect 633046 983613 633098 983619
rect 641122 983534 641150 993709
rect 642274 993519 642302 993857
rect 642262 993513 642314 993519
rect 642262 993455 642314 993461
rect 426262 983523 426314 983529
rect 267862 983465 267914 983471
rect 426262 983465 426314 983471
rect 318166 278673 318218 278679
rect 318166 278615 318218 278621
rect 373172 278638 373228 278647
rect 66646 278599 66698 278605
rect 66646 278541 66698 278547
rect 295798 278599 295850 278605
rect 295798 278541 295850 278547
rect 309046 278599 309098 278605
rect 309046 278541 309098 278547
rect 65890 272907 65918 277870
rect 66658 273647 66686 278541
rect 266038 278525 266090 278531
rect 204500 278490 204556 278499
rect 263732 278490 263788 278499
rect 222864 278457 223166 278476
rect 222864 278451 223178 278457
rect 222864 278448 223126 278451
rect 204500 278425 204556 278434
rect 197904 278161 198206 278180
rect 197904 278155 198218 278161
rect 197904 278152 198166 278155
rect 198166 278097 198218 278103
rect 166594 278004 166896 278032
rect 66646 273641 66698 273647
rect 66646 273583 66698 273589
rect 65878 272901 65930 272907
rect 65878 272843 65930 272849
rect 67042 272315 67070 277870
rect 67030 272309 67082 272315
rect 67030 272251 67082 272257
rect 68194 270761 68222 277870
rect 69442 272431 69470 277870
rect 70594 272727 70622 277870
rect 70580 272718 70636 272727
rect 70580 272653 70636 272662
rect 69428 272422 69484 272431
rect 69428 272357 69484 272366
rect 71746 272135 71774 277870
rect 71926 272457 71978 272463
rect 71926 272399 71978 272405
rect 71732 272126 71788 272135
rect 71732 272061 71788 272070
rect 68182 270755 68234 270761
rect 68182 270697 68234 270703
rect 69046 270755 69098 270761
rect 69046 270697 69098 270703
rect 65206 246779 65258 246785
rect 65206 246721 65258 246727
rect 47734 246351 47786 246357
rect 65108 246374 65164 246383
rect 65108 246309 65164 246318
rect 60502 246113 60554 246119
rect 60500 246078 60502 246087
rect 66262 246113 66314 246119
rect 60554 246078 60556 246087
rect 60500 246013 60556 246022
rect 66260 246078 66262 246087
rect 66314 246078 66316 246087
rect 66260 246013 66316 246022
rect 69058 243381 69086 270697
rect 71938 270632 71966 272399
rect 72994 271395 73022 277870
rect 74146 272283 74174 277870
rect 74900 273162 74956 273171
rect 74900 273097 74956 273106
rect 74914 272431 74942 273097
rect 74900 272422 74956 272431
rect 74900 272357 74956 272366
rect 74132 272274 74188 272283
rect 74132 272209 74188 272218
rect 75394 271723 75422 277870
rect 76546 272727 76574 277870
rect 76340 272718 76396 272727
rect 76340 272653 76396 272662
rect 76532 272718 76588 272727
rect 76532 272653 76588 272662
rect 75382 271717 75434 271723
rect 76354 271691 76382 272653
rect 77686 271717 77738 271723
rect 75382 271659 75434 271665
rect 76340 271682 76396 271691
rect 77686 271659 77738 271665
rect 76340 271617 76396 271626
rect 72980 271386 73036 271395
rect 72980 271321 73036 271330
rect 71938 270604 72062 270632
rect 72034 260697 72062 270604
rect 72022 260691 72074 260697
rect 72022 260633 72074 260639
rect 77698 243455 77726 271659
rect 77794 270951 77822 277870
rect 78946 272875 78974 277870
rect 80208 277856 80606 277884
rect 79222 273567 79274 273573
rect 79222 273509 79274 273515
rect 78932 272866 78988 272875
rect 78932 272801 78988 272810
rect 77780 270942 77836 270951
rect 77780 270877 77836 270886
rect 79234 265063 79262 273509
rect 79222 265057 79274 265063
rect 79222 264999 79274 265005
rect 77782 246113 77834 246119
rect 77782 246055 77834 246061
rect 77794 245897 77822 246055
rect 77782 245891 77834 245897
rect 77782 245833 77834 245839
rect 80578 243529 80606 277856
rect 81346 273023 81374 277870
rect 81332 273014 81388 273023
rect 81332 272949 81388 272958
rect 82594 271247 82622 277870
rect 83650 273615 83678 277870
rect 83636 273606 83692 273615
rect 83636 273541 83692 273550
rect 84898 272463 84926 277870
rect 86050 273319 86078 277870
rect 86036 273310 86092 273319
rect 86036 273245 86092 273254
rect 84886 272457 84938 272463
rect 84886 272399 84938 272405
rect 86326 272457 86378 272463
rect 86326 272399 86378 272405
rect 82580 271238 82636 271247
rect 82580 271173 82636 271182
rect 84694 260691 84746 260697
rect 84694 260633 84746 260639
rect 84706 253519 84734 260633
rect 84694 253513 84746 253519
rect 84694 253455 84746 253461
rect 81142 247001 81194 247007
rect 80674 246924 80990 246952
rect 81142 246943 81194 246949
rect 80674 246711 80702 246924
rect 80962 246711 80990 246924
rect 81154 246785 81182 246943
rect 81142 246779 81194 246785
rect 81142 246721 81194 246727
rect 80662 246705 80714 246711
rect 80662 246647 80714 246653
rect 80950 246705 81002 246711
rect 80950 246647 81002 246653
rect 80758 246631 80810 246637
rect 80758 246573 80810 246579
rect 81238 246631 81290 246637
rect 81238 246573 81290 246579
rect 80770 246508 80798 246573
rect 80770 246480 80894 246508
rect 80866 246360 80894 246480
rect 80866 246332 81086 246360
rect 80758 246261 80810 246267
rect 80950 246261 81002 246267
rect 80810 246209 80950 246212
rect 80758 246203 81002 246209
rect 81058 246212 81086 246332
rect 81250 246212 81278 246573
rect 80770 246184 80990 246203
rect 81058 246184 81278 246212
rect 86338 243603 86366 272399
rect 87202 271099 87230 277870
rect 88450 273467 88478 277870
rect 88436 273458 88492 273467
rect 88436 273393 88492 273402
rect 89602 271649 89630 277870
rect 90850 271987 90878 277870
rect 92002 273499 92030 277870
rect 91990 273493 92042 273499
rect 91990 273435 92042 273441
rect 90836 271978 90892 271987
rect 90836 271913 90892 271922
rect 93250 271839 93278 277870
rect 94416 277856 95006 277884
rect 94868 273162 94924 273171
rect 94868 273097 94924 273106
rect 94772 272570 94828 272579
rect 94772 272505 94828 272514
rect 93236 271830 93292 271839
rect 93236 271765 93292 271774
rect 94786 271691 94814 272505
rect 94882 272431 94910 273097
rect 94868 272422 94924 272431
rect 94868 272357 94924 272366
rect 94772 271682 94828 271691
rect 89590 271643 89642 271649
rect 89590 271585 89642 271591
rect 92086 271643 92138 271649
rect 94772 271617 94828 271626
rect 92086 271585 92138 271591
rect 87188 271090 87244 271099
rect 87188 271025 87244 271034
rect 86422 264983 86474 264989
rect 86422 264925 86474 264931
rect 86434 259291 86462 264925
rect 86422 259285 86474 259291
rect 86422 259227 86474 259233
rect 92098 243677 92126 271585
rect 92278 259211 92330 259217
rect 92278 259153 92330 259159
rect 92290 254925 92318 259153
rect 92278 254919 92330 254925
rect 92278 254861 92330 254867
rect 92182 253439 92234 253445
rect 92182 253381 92234 253387
rect 92194 250559 92222 253381
rect 92182 250553 92234 250559
rect 92182 250495 92234 250501
rect 94978 243751 95006 277856
rect 95650 271871 95678 277870
rect 95638 271865 95690 271871
rect 95638 271807 95690 271813
rect 96802 271691 96830 277870
rect 96788 271682 96844 271691
rect 96788 271617 96844 271626
rect 98050 270761 98078 277870
rect 99202 272019 99230 277870
rect 100368 277856 100670 277884
rect 99190 272013 99242 272019
rect 99190 271955 99242 271961
rect 100642 271520 100670 277856
rect 101506 271797 101534 277870
rect 101494 271791 101546 271797
rect 101494 271733 101546 271739
rect 100820 271682 100876 271691
rect 100820 271617 100822 271626
rect 100874 271617 100876 271626
rect 100822 271585 100874 271591
rect 100724 271534 100780 271543
rect 100642 271492 100724 271520
rect 100724 271469 100780 271478
rect 102658 271427 102686 277870
rect 103906 272241 103934 277870
rect 105058 272463 105086 277870
rect 106306 273573 106334 277870
rect 106294 273567 106346 273573
rect 106294 273509 106346 273515
rect 105046 272457 105098 272463
rect 105046 272399 105098 272405
rect 106486 272457 106538 272463
rect 106486 272399 106538 272405
rect 103894 272235 103946 272241
rect 103894 272177 103946 272183
rect 103606 271791 103658 271797
rect 103606 271733 103658 271739
rect 102646 271421 102698 271427
rect 102646 271363 102698 271369
rect 98038 270755 98090 270761
rect 98038 270697 98090 270703
rect 100726 270755 100778 270761
rect 100726 270697 100778 270703
rect 97174 250553 97226 250559
rect 97174 250495 97226 250501
rect 97186 244713 97214 250495
rect 97846 246039 97898 246045
rect 97846 245981 97898 245987
rect 97858 245897 97886 245981
rect 97846 245891 97898 245897
rect 97846 245833 97898 245839
rect 97174 244707 97226 244713
rect 97174 244649 97226 244655
rect 100738 243825 100766 270697
rect 103618 243899 103646 271733
rect 104374 254919 104426 254925
rect 104374 254861 104426 254867
rect 104386 250115 104414 254861
rect 104374 250109 104426 250115
rect 104374 250051 104426 250057
rect 106498 243973 106526 272399
rect 107458 272167 107486 277870
rect 108720 277856 109406 277884
rect 107446 272161 107498 272167
rect 107446 272103 107498 272109
rect 106582 250109 106634 250115
rect 106582 250051 106634 250057
rect 106594 244861 106622 250051
rect 106582 244855 106634 244861
rect 106582 244797 106634 244803
rect 109378 244047 109406 277856
rect 109858 271131 109886 277870
rect 111106 272389 111134 277870
rect 111094 272383 111146 272389
rect 111094 272325 111146 272331
rect 109846 271125 109898 271131
rect 109846 271067 109898 271073
rect 112258 244121 112286 277870
rect 113506 271353 113534 277870
rect 114658 276723 114686 277870
rect 114644 276714 114700 276723
rect 114644 276649 114700 276658
rect 115220 273162 115276 273171
rect 115220 273097 115276 273106
rect 115234 272431 115262 273097
rect 115316 272570 115372 272579
rect 115316 272505 115372 272514
rect 115220 272422 115276 272431
rect 115220 272357 115276 272366
rect 113494 271347 113546 271353
rect 113494 271289 113546 271295
rect 115330 270803 115358 272505
rect 115316 270794 115372 270803
rect 115810 270761 115838 277870
rect 116962 271279 116990 277870
rect 118114 272463 118142 277870
rect 118102 272457 118154 272463
rect 118102 272399 118154 272405
rect 116950 271273 117002 271279
rect 116950 271215 117002 271221
rect 119362 270761 119390 277870
rect 120514 271205 120542 277870
rect 121762 272537 121790 277870
rect 121750 272531 121802 272537
rect 121750 272473 121802 272479
rect 120982 271717 121034 271723
rect 120788 271682 120844 271691
rect 120788 271617 120790 271626
rect 120842 271617 120844 271626
rect 120980 271682 120982 271691
rect 121034 271682 121036 271691
rect 120980 271617 121036 271626
rect 120790 271585 120842 271591
rect 120502 271199 120554 271205
rect 120502 271141 120554 271147
rect 122914 270761 122942 277870
rect 124162 270761 124190 277870
rect 125314 272759 125342 277870
rect 126576 277856 126686 277884
rect 125302 272753 125354 272759
rect 125302 272695 125354 272701
rect 115316 270729 115372 270738
rect 115798 270755 115850 270761
rect 115798 270697 115850 270703
rect 118006 270755 118058 270761
rect 118006 270697 118058 270703
rect 119350 270755 119402 270761
rect 119350 270697 119402 270703
rect 120886 270755 120938 270761
rect 120886 270697 120938 270703
rect 122902 270755 122954 270761
rect 122902 270697 122954 270703
rect 123766 270755 123818 270761
rect 123766 270697 123818 270703
rect 124150 270755 124202 270761
rect 124150 270697 124202 270703
rect 126550 270755 126602 270761
rect 126550 270697 126602 270703
rect 118018 244195 118046 270697
rect 118102 246187 118154 246193
rect 118102 246129 118154 246135
rect 118114 246045 118142 246129
rect 118102 246039 118154 246045
rect 118102 245981 118154 245987
rect 120898 244269 120926 270697
rect 123778 244343 123806 270697
rect 126562 247377 126590 270697
rect 126550 247371 126602 247377
rect 126550 247313 126602 247319
rect 126658 244417 126686 277856
rect 127714 272611 127742 277870
rect 128962 272685 128990 277870
rect 128950 272679 129002 272685
rect 128950 272621 129002 272627
rect 127702 272605 127754 272611
rect 127702 272547 127754 272553
rect 129526 272605 129578 272611
rect 129526 272547 129578 272553
rect 129538 247303 129566 272547
rect 130114 270835 130142 277870
rect 130102 270829 130154 270835
rect 130102 270771 130154 270777
rect 131266 270761 131294 277870
rect 132514 272759 132542 277870
rect 132502 272753 132554 272759
rect 132502 272695 132554 272701
rect 132406 270829 132458 270835
rect 132406 270771 132458 270777
rect 131254 270755 131306 270761
rect 131254 270697 131306 270703
rect 132310 270755 132362 270761
rect 132310 270697 132362 270703
rect 129526 247297 129578 247303
rect 129526 247239 129578 247245
rect 132322 247155 132350 270697
rect 132310 247149 132362 247155
rect 132310 247091 132362 247097
rect 128086 246187 128138 246193
rect 128086 246129 128138 246135
rect 128098 246045 128126 246129
rect 128086 246039 128138 246045
rect 128086 245981 128138 245987
rect 132418 244491 132446 270771
rect 133570 270761 133598 277870
rect 134832 277856 135230 277884
rect 133558 270755 133610 270761
rect 133558 270697 133610 270703
rect 135202 247229 135230 277856
rect 135284 273162 135340 273171
rect 135284 273097 135340 273106
rect 135298 272431 135326 273097
rect 135970 272833 135998 277870
rect 135958 272827 136010 272833
rect 135958 272769 136010 272775
rect 135284 272422 135340 272431
rect 135284 272357 135340 272366
rect 137218 270761 137246 277870
rect 138370 270761 138398 277870
rect 139618 273129 139646 277870
rect 139606 273123 139658 273129
rect 139606 273065 139658 273071
rect 140770 270817 140798 277870
rect 142018 273055 142046 277870
rect 142006 273049 142058 273055
rect 142006 272991 142058 272997
rect 143170 272981 143198 277870
rect 143926 273049 143978 273055
rect 143926 272991 143978 272997
rect 143158 272975 143210 272981
rect 143158 272917 143210 272923
rect 141046 271717 141098 271723
rect 141044 271682 141046 271691
rect 141334 271717 141386 271723
rect 141098 271682 141100 271691
rect 141044 271617 141100 271626
rect 141332 271682 141334 271691
rect 141386 271682 141388 271691
rect 141332 271617 141388 271626
rect 141142 271569 141194 271575
rect 141140 271534 141142 271543
rect 141622 271569 141674 271575
rect 141194 271534 141196 271543
rect 141140 271469 141196 271478
rect 141620 271534 141622 271543
rect 141674 271534 141676 271543
rect 141620 271469 141676 271478
rect 141140 271386 141196 271395
rect 141140 271321 141196 271330
rect 141620 271386 141676 271395
rect 141620 271321 141676 271330
rect 141154 271261 141182 271321
rect 141634 271261 141662 271321
rect 141154 271233 141662 271261
rect 140770 270789 141086 270817
rect 135286 270755 135338 270761
rect 135286 270697 135338 270703
rect 137206 270755 137258 270761
rect 137206 270697 137258 270703
rect 138166 270755 138218 270761
rect 138166 270697 138218 270703
rect 138358 270755 138410 270761
rect 138358 270697 138410 270703
rect 140950 270755 141002 270761
rect 140950 270697 141002 270703
rect 135190 247223 135242 247229
rect 135190 247165 135242 247171
rect 135298 244565 135326 270697
rect 138178 244639 138206 270697
rect 140962 247081 140990 270697
rect 140950 247075 141002 247081
rect 140950 247017 141002 247023
rect 138166 244633 138218 244639
rect 138166 244575 138218 244581
rect 135286 244559 135338 244565
rect 135286 244501 135338 244507
rect 132406 244485 132458 244491
rect 132406 244427 132458 244433
rect 126646 244411 126698 244417
rect 126646 244353 126698 244359
rect 123766 244337 123818 244343
rect 123766 244279 123818 244285
rect 120886 244263 120938 244269
rect 120886 244205 120938 244211
rect 118006 244189 118058 244195
rect 118006 244131 118058 244137
rect 112246 244115 112298 244121
rect 112246 244057 112298 244063
rect 109366 244041 109418 244047
rect 109366 243983 109418 243989
rect 106486 243967 106538 243973
rect 106486 243909 106538 243915
rect 103606 243893 103658 243899
rect 103606 243835 103658 243841
rect 100726 243819 100778 243825
rect 100726 243761 100778 243767
rect 94966 243745 95018 243751
rect 94966 243687 95018 243693
rect 92086 243671 92138 243677
rect 92086 243613 92138 243619
rect 86326 243597 86378 243603
rect 86326 243539 86378 243545
rect 80566 243523 80618 243529
rect 80566 243465 80618 243471
rect 77686 243449 77738 243455
rect 77686 243391 77738 243397
rect 69046 243375 69098 243381
rect 69046 243317 69098 243323
rect 50326 241969 50378 241975
rect 50326 241911 50378 241917
rect 47542 237899 47594 237905
rect 47542 237841 47594 237847
rect 45142 216513 45194 216519
rect 45142 216455 45194 216461
rect 45046 215773 45098 215779
rect 45046 215715 45098 215721
rect 50338 204457 50366 241911
rect 141058 224659 141086 270789
rect 143938 247007 143966 272991
rect 144418 270835 144446 277870
rect 144406 270829 144458 270835
rect 144406 270771 144458 270777
rect 145570 270761 145598 277870
rect 146722 273129 146750 277870
rect 147970 273203 147998 277870
rect 149136 277856 149630 277884
rect 147958 273197 148010 273203
rect 147958 273139 148010 273145
rect 146710 273123 146762 273129
rect 146710 273065 146762 273071
rect 146902 272753 146954 272759
rect 146902 272695 146954 272701
rect 146914 271797 146942 272695
rect 146902 271791 146954 271797
rect 146902 271733 146954 271739
rect 146806 270829 146858 270835
rect 146806 270771 146858 270777
rect 145558 270755 145610 270761
rect 145558 270697 145610 270703
rect 146710 270755 146762 270761
rect 146710 270697 146762 270703
rect 143926 247001 143978 247007
rect 143926 246943 143978 246949
rect 146722 246933 146750 270697
rect 146710 246927 146762 246933
rect 146710 246869 146762 246875
rect 141142 246039 141194 246045
rect 141142 245981 141194 245987
rect 141154 245897 141182 245981
rect 141142 245891 141194 245897
rect 141142 245833 141194 245839
rect 142486 244707 142538 244713
rect 142486 244649 142538 244655
rect 142498 237651 142526 244649
rect 146132 240602 146188 240611
rect 146132 240537 146188 240546
rect 144116 238678 144172 238687
rect 144116 238613 144172 238622
rect 142484 237642 142540 237651
rect 142484 237577 142540 237586
rect 144020 236310 144076 236319
rect 144130 236277 144158 238613
rect 144020 236245 144076 236254
rect 144118 236271 144170 236277
rect 144034 236203 144062 236245
rect 144118 236213 144170 236219
rect 144022 236197 144074 236203
rect 144022 236139 144074 236145
rect 144020 233646 144076 233655
rect 144020 233581 144076 233590
rect 144034 233317 144062 233581
rect 144022 233311 144074 233317
rect 144022 233253 144074 233259
rect 144116 232166 144172 232175
rect 144116 232101 144172 232110
rect 144020 231426 144076 231435
rect 144020 231361 144076 231370
rect 144034 230579 144062 231361
rect 144022 230573 144074 230579
rect 144022 230515 144074 230521
rect 144130 230505 144158 232101
rect 144118 230499 144170 230505
rect 144118 230441 144170 230447
rect 144212 230242 144268 230251
rect 144212 230177 144268 230186
rect 144116 228466 144172 228475
rect 144116 228401 144172 228410
rect 144020 227874 144076 227883
rect 144020 227809 144076 227818
rect 144034 227767 144062 227809
rect 144022 227761 144074 227767
rect 144022 227703 144074 227709
rect 144130 227693 144158 228401
rect 144118 227687 144170 227693
rect 144118 227629 144170 227635
rect 144226 227619 144254 230177
rect 144214 227613 144266 227619
rect 144214 227555 144266 227561
rect 141046 224653 141098 224659
rect 141046 224595 141098 224601
rect 144404 223730 144460 223739
rect 144404 223665 144460 223674
rect 144418 221847 144446 223665
rect 144406 221841 144458 221847
rect 144406 221783 144458 221789
rect 144404 220178 144460 220187
rect 144404 220113 144460 220122
rect 144418 218961 144446 220113
rect 144406 218955 144458 218961
rect 144406 218897 144458 218903
rect 144212 215294 144268 215303
rect 144212 215229 144268 215238
rect 144226 213189 144254 215229
rect 144214 213183 144266 213189
rect 144214 213125 144266 213131
rect 145364 210558 145420 210567
rect 145364 210493 145420 210502
rect 50326 204451 50378 204457
rect 50326 204393 50378 204399
rect 144980 203306 145036 203315
rect 144980 203241 145036 203250
rect 144994 201645 145022 203241
rect 144982 201639 145034 201645
rect 144982 201581 145034 201587
rect 145076 199014 145132 199023
rect 145076 198949 145132 198958
rect 144596 196646 144652 196655
rect 144596 196581 144652 196590
rect 144404 194870 144460 194879
rect 144404 194805 144460 194814
rect 44758 194535 44810 194541
rect 44758 194477 44810 194483
rect 43126 193499 43178 193505
rect 43126 193441 43178 193447
rect 43030 192241 43082 192247
rect 43030 192183 43082 192189
rect 42934 191501 42986 191507
rect 42934 191443 42986 191449
rect 42932 188358 42988 188367
rect 42932 188293 42988 188302
rect 42166 187727 42218 187733
rect 42166 187669 42218 187675
rect 42838 187727 42890 187733
rect 42838 187669 42890 187675
rect 42178 187442 42206 187669
rect 41780 187174 41836 187183
rect 41780 187109 41836 187118
rect 41794 186776 41822 187109
rect 41780 186434 41836 186443
rect 41780 186369 41836 186378
rect 41794 186184 41822 186369
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42946 125351 42974 188293
rect 144020 181846 144076 181855
rect 144020 181781 144076 181790
rect 144034 181517 144062 181781
rect 144022 181511 144074 181517
rect 144022 181453 144074 181459
rect 144116 176814 144172 176823
rect 144116 176749 144172 176758
rect 144130 175745 144158 176749
rect 144118 175739 144170 175745
rect 144118 175681 144170 175687
rect 144212 163642 144268 163651
rect 144212 163577 144268 163586
rect 144020 159942 144076 159951
rect 144020 159877 144076 159886
rect 144034 127053 144062 159877
rect 144116 158166 144172 158175
rect 144116 158101 144172 158110
rect 144130 127053 144158 158101
rect 144226 127053 144254 163577
rect 144308 155650 144364 155659
rect 144308 155585 144364 155594
rect 144322 144517 144350 155585
rect 144310 144511 144362 144517
rect 144310 144453 144362 144459
rect 144308 144402 144364 144411
rect 144308 144337 144364 144346
rect 144322 144073 144350 144337
rect 144310 144067 144362 144073
rect 144310 144009 144362 144015
rect 144308 142478 144364 142487
rect 144308 142413 144364 142422
rect 144322 141705 144350 142413
rect 144310 141699 144362 141705
rect 144310 141641 144362 141647
rect 144308 141294 144364 141303
rect 144308 141229 144310 141238
rect 144362 141229 144364 141238
rect 144310 141197 144362 141203
rect 144308 139518 144364 139527
rect 144308 139453 144364 139462
rect 144322 138301 144350 139453
rect 144310 138295 144362 138301
rect 144310 138237 144362 138243
rect 144308 137594 144364 137603
rect 144308 137529 144364 137538
rect 144322 135489 144350 137529
rect 144310 135483 144362 135489
rect 144310 135425 144362 135431
rect 144308 134782 144364 134791
rect 144308 134717 144364 134726
rect 144322 132973 144350 134717
rect 144310 132967 144362 132973
rect 144310 132909 144362 132915
rect 144308 132858 144364 132867
rect 144308 132793 144364 132802
rect 144322 132603 144350 132793
rect 144310 132597 144362 132603
rect 144310 132539 144362 132545
rect 144308 130046 144364 130055
rect 144308 129981 144364 129990
rect 144322 129643 144350 129981
rect 144310 129637 144362 129643
rect 144310 129579 144362 129585
rect 144308 129306 144364 129315
rect 144308 129241 144364 129250
rect 144022 127047 144074 127053
rect 144022 126989 144074 126995
rect 144118 127047 144170 127053
rect 144118 126989 144170 126995
rect 144214 127047 144266 127053
rect 144214 126989 144266 126995
rect 144322 126979 144350 129241
rect 144310 126973 144362 126979
rect 144310 126915 144362 126921
rect 144022 126825 144074 126831
rect 144022 126767 144074 126773
rect 144118 126825 144170 126831
rect 144118 126767 144170 126773
rect 144214 126825 144266 126831
rect 144214 126767 144266 126773
rect 144308 126790 144364 126799
rect 143926 126751 143978 126757
rect 143926 126693 143978 126699
rect 143938 126535 143966 126693
rect 143926 126529 143978 126535
rect 143926 126471 143978 126477
rect 39862 125345 39914 125351
rect 39860 125310 39862 125319
rect 42934 125345 42986 125351
rect 39914 125310 39916 125319
rect 42934 125287 42986 125293
rect 39860 125245 39916 125254
rect 143830 106993 143882 106999
rect 143830 106935 143882 106941
rect 141044 104146 141100 104155
rect 141044 104081 141100 104090
rect 141058 103859 141086 104081
rect 141044 103850 141100 103859
rect 141044 103785 141100 103794
rect 143842 103447 143870 106935
rect 143926 106845 143978 106851
rect 143926 106787 143978 106793
rect 143938 106481 143966 106787
rect 143926 106475 143978 106481
rect 143926 106417 143978 106423
rect 143830 103441 143882 103447
rect 143830 103383 143882 103389
rect 144034 94641 144062 126767
rect 144022 94635 144074 94641
rect 144022 94577 144074 94583
rect 144130 92125 144158 126767
rect 144226 94937 144254 126767
rect 144308 126725 144364 126734
rect 144322 124579 144350 126725
rect 144418 125277 144446 194805
rect 144500 183326 144556 183335
rect 144500 183261 144556 183270
rect 144514 181591 144542 183261
rect 144502 181585 144554 181591
rect 144502 181527 144554 181533
rect 144500 151654 144556 151663
rect 144500 151589 144556 151598
rect 144514 146145 144542 151589
rect 144502 146139 144554 146145
rect 144502 146081 144554 146087
rect 144500 146030 144556 146039
rect 144500 145965 144556 145974
rect 144514 144369 144542 145965
rect 144502 144363 144554 144369
rect 144502 144305 144554 144311
rect 144500 143218 144556 143227
rect 144500 143153 144556 143162
rect 144514 141187 144542 143153
rect 144502 141181 144554 141187
rect 144502 141123 144554 141129
rect 144502 140959 144554 140965
rect 144502 140901 144554 140907
rect 144514 135045 144542 140901
rect 144502 135039 144554 135045
rect 144502 134981 144554 134987
rect 144500 134042 144556 134051
rect 144500 133977 144556 133986
rect 144514 132529 144542 133977
rect 144502 132523 144554 132529
rect 144502 132465 144554 132471
rect 144500 131082 144556 131091
rect 144500 131017 144556 131026
rect 144514 129717 144542 131017
rect 144502 129711 144554 129717
rect 144502 129653 144554 129659
rect 144502 129563 144554 129569
rect 144502 129505 144554 129511
rect 144406 125271 144458 125277
rect 144406 125213 144458 125219
rect 144404 125162 144460 125171
rect 144404 125097 144460 125106
rect 144308 124570 144364 124579
rect 144308 124505 144364 124514
rect 144308 124422 144364 124431
rect 144308 124357 144364 124366
rect 144322 124019 144350 124357
rect 144310 124013 144362 124019
rect 144310 123955 144362 123961
rect 144418 123945 144446 125097
rect 144406 123939 144458 123945
rect 144406 123881 144458 123887
rect 144404 122646 144460 122655
rect 144404 122581 144460 122590
rect 144308 121610 144364 121619
rect 144308 121545 144364 121554
rect 144322 121059 144350 121545
rect 144418 121133 144446 122581
rect 144406 121127 144458 121133
rect 144406 121069 144458 121075
rect 144310 121053 144362 121059
rect 144310 120995 144362 121001
rect 144406 120979 144458 120985
rect 144406 120921 144458 120927
rect 144418 119228 144446 120921
rect 144322 119200 144446 119228
rect 144322 118469 144350 119200
rect 144404 119094 144460 119103
rect 144404 119029 144460 119038
rect 144310 118463 144362 118469
rect 144310 118405 144362 118411
rect 144418 118321 144446 119029
rect 144406 118315 144458 118321
rect 144406 118257 144458 118263
rect 144310 118241 144362 118247
rect 144308 118206 144310 118215
rect 144362 118206 144364 118215
rect 144308 118141 144364 118150
rect 144308 116726 144364 116735
rect 144308 116661 144364 116670
rect 144322 116249 144350 116661
rect 144310 116243 144362 116249
rect 144310 116185 144362 116191
rect 144308 115986 144364 115995
rect 144308 115921 144364 115930
rect 144322 115583 144350 115921
rect 144310 115577 144362 115583
rect 144310 115519 144362 115525
rect 144310 115429 144362 115435
rect 144310 115371 144362 115377
rect 144322 113331 144350 115371
rect 144404 114210 144460 114219
rect 144404 114145 144460 114154
rect 144308 113322 144364 113331
rect 144308 113257 144364 113266
rect 144308 113174 144364 113183
rect 144308 113109 144364 113118
rect 144322 112697 144350 113109
rect 144310 112691 144362 112697
rect 144310 112633 144362 112639
rect 144310 112469 144362 112475
rect 144308 112434 144310 112443
rect 144362 112434 144364 112443
rect 144418 112401 144446 114145
rect 144308 112369 144364 112378
rect 144406 112395 144458 112401
rect 144406 112337 144458 112343
rect 144404 111250 144460 111259
rect 144404 111185 144460 111194
rect 144308 109770 144364 109779
rect 144308 109705 144364 109714
rect 144322 109515 144350 109705
rect 144418 109589 144446 111185
rect 144406 109583 144458 109589
rect 144406 109525 144458 109531
rect 144310 109509 144362 109515
rect 144310 109451 144362 109457
rect 144406 109435 144458 109441
rect 144406 109377 144458 109383
rect 144308 107550 144364 107559
rect 144308 107485 144364 107494
rect 144322 106925 144350 107485
rect 144418 106999 144446 109377
rect 144406 106993 144458 106999
rect 144406 106935 144458 106941
rect 144310 106919 144362 106925
rect 144310 106861 144362 106867
rect 144404 106810 144460 106819
rect 144310 106771 144362 106777
rect 144404 106745 144460 106754
rect 144310 106713 144362 106719
rect 144214 94931 144266 94937
rect 144214 94873 144266 94879
rect 144118 92119 144170 92125
rect 144118 92061 144170 92067
rect 144212 87866 144268 87875
rect 144212 87801 144268 87810
rect 144116 87126 144172 87135
rect 144116 87061 144172 87070
rect 144022 75173 144074 75179
rect 144020 75138 144022 75147
rect 144074 75138 144076 75147
rect 144020 75073 144076 75082
rect 144130 75031 144158 87061
rect 144226 75105 144254 87801
rect 144214 75099 144266 75105
rect 144214 75041 144266 75047
rect 144118 75025 144170 75031
rect 144118 74967 144170 74973
rect 144214 74063 144266 74069
rect 144214 74005 144266 74011
rect 144020 69810 144076 69819
rect 144020 69745 144076 69754
rect 144034 69185 144062 69745
rect 144118 69549 144170 69555
rect 144118 69491 144170 69497
rect 144022 69179 144074 69185
rect 144022 69121 144074 69127
rect 144130 56975 144158 69491
rect 144226 64449 144254 74005
rect 144214 64443 144266 64449
rect 144214 64385 144266 64391
rect 144118 56969 144170 56975
rect 144118 56911 144170 56917
rect 144022 56525 144074 56531
rect 144020 56490 144022 56499
rect 144074 56490 144076 56499
rect 144020 56425 144076 56434
rect 144214 54379 144266 54385
rect 144214 54321 144266 54327
rect 144226 52091 144254 54321
rect 144214 52085 144266 52091
rect 144214 52027 144266 52033
rect 144322 50389 144350 106713
rect 144418 100709 144446 106745
rect 144406 100703 144458 100709
rect 144406 100645 144458 100651
rect 144404 77506 144460 77515
rect 144404 77441 144460 77450
rect 144418 74957 144446 77441
rect 144406 74951 144458 74957
rect 144406 74893 144458 74899
rect 144406 74507 144458 74513
rect 144406 74449 144458 74455
rect 144418 72779 144446 74449
rect 144404 72770 144460 72779
rect 144404 72705 144460 72714
rect 144514 64764 144542 129505
rect 144610 125425 144638 196581
rect 144980 174446 145036 174455
rect 144980 174381 145036 174390
rect 144788 173410 144844 173419
rect 144788 173345 144844 173354
rect 144802 172859 144830 173345
rect 144790 172853 144842 172859
rect 144790 172795 144842 172801
rect 144788 168378 144844 168387
rect 144788 168313 144844 168322
rect 144802 167087 144830 168313
rect 144790 167081 144842 167087
rect 144790 167023 144842 167029
rect 144788 166602 144844 166611
rect 144788 166537 144844 166546
rect 144802 164201 144830 166537
rect 144790 164195 144842 164201
rect 144790 164137 144842 164143
rect 144884 162902 144940 162911
rect 144884 162837 144940 162846
rect 144898 161315 144926 162837
rect 144994 162795 145022 174381
rect 144982 162789 145034 162795
rect 144982 162731 145034 162737
rect 144980 161422 145036 161431
rect 144980 161357 145036 161366
rect 144886 161309 144938 161315
rect 144886 161251 144938 161257
rect 144884 159350 144940 159359
rect 144884 159285 144940 159294
rect 144898 158503 144926 159285
rect 144886 158497 144938 158503
rect 144886 158439 144938 158445
rect 144884 156390 144940 156399
rect 144884 156325 144940 156334
rect 144898 155617 144926 156325
rect 144886 155611 144938 155617
rect 144886 155553 144938 155559
rect 144788 154466 144844 154475
rect 144788 154401 144844 154410
rect 144802 152731 144830 154401
rect 144884 152986 144940 152995
rect 144884 152921 144940 152930
rect 144898 152805 144926 152921
rect 144886 152799 144938 152805
rect 144886 152741 144938 152747
rect 144790 152725 144842 152731
rect 144790 152667 144842 152673
rect 144884 150914 144940 150923
rect 144884 150849 144940 150858
rect 144898 149845 144926 150849
rect 144886 149839 144938 149845
rect 144886 149781 144938 149787
rect 144788 149730 144844 149739
rect 144788 149665 144844 149674
rect 144692 146918 144748 146927
rect 144692 146853 144748 146862
rect 144706 136969 144734 146853
rect 144694 136963 144746 136969
rect 144694 136905 144746 136911
rect 144802 136840 144830 149665
rect 144884 147954 144940 147963
rect 144884 147889 144940 147898
rect 144898 146959 144926 147889
rect 144886 146953 144938 146959
rect 144886 146895 144938 146901
rect 144886 146139 144938 146145
rect 144886 146081 144938 146087
rect 144898 137117 144926 146081
rect 144886 137111 144938 137117
rect 144886 137053 144938 137059
rect 144886 136963 144938 136969
rect 144886 136905 144938 136911
rect 144706 136812 144830 136840
rect 144598 125419 144650 125425
rect 144598 125361 144650 125367
rect 144598 125271 144650 125277
rect 144598 125213 144650 125219
rect 144610 120985 144638 125213
rect 144598 120979 144650 120985
rect 144598 120921 144650 120927
rect 144596 120870 144652 120879
rect 144596 120805 144652 120814
rect 144610 118173 144638 120805
rect 144598 118167 144650 118173
rect 144598 118109 144650 118115
rect 144598 118019 144650 118025
rect 144598 117961 144650 117967
rect 144610 109441 144638 117961
rect 144598 109435 144650 109441
rect 144598 109377 144650 109383
rect 144596 108290 144652 108299
rect 144596 108225 144652 108234
rect 144610 106629 144638 108225
rect 144598 106623 144650 106629
rect 144598 106565 144650 106571
rect 144598 106475 144650 106481
rect 144598 106417 144650 106423
rect 144610 100635 144638 106417
rect 144598 100629 144650 100635
rect 144598 100571 144650 100577
rect 144596 80762 144652 80771
rect 144596 80697 144652 80706
rect 144418 64736 144542 64764
rect 144418 50611 144446 64736
rect 144502 64665 144554 64671
rect 144502 64607 144554 64613
rect 144514 54256 144542 64607
rect 144610 54385 144638 80697
rect 144706 64671 144734 136812
rect 144790 136741 144842 136747
rect 144790 136683 144842 136689
rect 144802 64671 144830 136683
rect 144898 129569 144926 136905
rect 144886 129563 144938 129569
rect 144886 129505 144938 129511
rect 144886 129415 144938 129421
rect 144886 129357 144938 129363
rect 144694 64665 144746 64671
rect 144694 64607 144746 64613
rect 144790 64665 144842 64671
rect 144790 64607 144842 64613
rect 144694 64517 144746 64523
rect 144694 64459 144746 64465
rect 144706 54404 144734 64459
rect 144788 54714 144844 54723
rect 144788 54649 144790 54658
rect 144842 54649 144844 54658
rect 144790 54617 144842 54623
rect 144598 54379 144650 54385
rect 144706 54376 144830 54404
rect 144598 54321 144650 54327
rect 144514 54228 144734 54256
rect 144502 54157 144554 54163
rect 144500 54122 144502 54131
rect 144554 54122 144556 54131
rect 144500 54057 144556 54066
rect 144406 50605 144458 50611
rect 144406 50547 144458 50553
rect 144706 50537 144734 54228
rect 144694 50531 144746 50537
rect 144694 50473 144746 50479
rect 144310 50383 144362 50389
rect 144310 50325 144362 50331
rect 144802 50315 144830 54376
rect 144898 50907 144926 129357
rect 144994 51499 145022 161357
rect 145090 126683 145118 198949
rect 145268 179774 145324 179783
rect 145268 179709 145324 179718
rect 145282 178705 145310 179709
rect 145270 178699 145322 178705
rect 145270 178641 145322 178647
rect 145268 172078 145324 172087
rect 145268 172013 145324 172022
rect 145172 164826 145228 164835
rect 145172 164761 145228 164770
rect 145078 126677 145130 126683
rect 145078 126619 145130 126625
rect 145078 126529 145130 126535
rect 145078 126471 145130 126477
rect 145090 106777 145118 126471
rect 145078 106771 145130 106777
rect 145078 106713 145130 106719
rect 145076 106662 145132 106671
rect 145076 106597 145132 106606
rect 145090 103595 145118 106597
rect 145078 103589 145130 103595
rect 145078 103531 145130 103537
rect 145078 103441 145130 103447
rect 145078 103383 145130 103389
rect 145090 100783 145118 103383
rect 145078 100777 145130 100783
rect 145078 100719 145130 100725
rect 145076 84166 145132 84175
rect 145076 84101 145132 84110
rect 145090 52017 145118 84101
rect 145078 52011 145130 52017
rect 145078 51953 145130 51959
rect 144982 51493 145034 51499
rect 144982 51435 145034 51441
rect 145186 51425 145214 164761
rect 145174 51419 145226 51425
rect 145174 51361 145226 51367
rect 144886 50901 144938 50907
rect 144886 50843 144938 50849
rect 145282 50833 145310 172013
rect 145378 51351 145406 210493
rect 145460 208042 145516 208051
rect 145460 207977 145516 207986
rect 145474 69407 145502 207977
rect 145556 205674 145612 205683
rect 145556 205609 145612 205618
rect 145462 69401 145514 69407
rect 145462 69343 145514 69349
rect 145462 69253 145514 69259
rect 145462 69195 145514 69201
rect 145366 51345 145418 51351
rect 145366 51287 145418 51293
rect 145270 50827 145322 50833
rect 145270 50769 145322 50775
rect 144790 50309 144842 50315
rect 144790 50251 144842 50257
rect 145366 49865 145418 49871
rect 145104 49813 145366 49816
rect 145104 49807 145418 49813
rect 145104 49788 145406 49807
rect 145474 49723 145502 69195
rect 145570 64764 145598 205609
rect 145748 205082 145804 205091
rect 145748 205017 145804 205026
rect 145652 201382 145708 201391
rect 145652 201317 145708 201326
rect 145666 69555 145694 201317
rect 145654 69549 145706 69555
rect 145654 69491 145706 69497
rect 145654 69401 145706 69407
rect 145654 69343 145706 69349
rect 145666 64893 145694 69343
rect 145654 64887 145706 64893
rect 145654 64829 145706 64835
rect 145570 64736 145694 64764
rect 145558 64665 145610 64671
rect 145558 64607 145610 64613
rect 145570 50463 145598 64607
rect 145666 51277 145694 64736
rect 145654 51271 145706 51277
rect 145654 51213 145706 51219
rect 145558 50457 145610 50463
rect 145558 50399 145610 50405
rect 145762 50241 145790 205017
rect 145844 193686 145900 193695
rect 145844 193621 145900 193630
rect 145858 69259 145886 193621
rect 145940 190134 145996 190143
rect 145940 190069 145996 190078
rect 145846 69253 145898 69259
rect 145846 69195 145898 69201
rect 145844 69070 145900 69079
rect 145844 69005 145900 69014
rect 145858 66447 145886 69005
rect 145846 66441 145898 66447
rect 145846 66383 145898 66389
rect 145954 64764 145982 190069
rect 146036 189394 146092 189403
rect 146036 189329 146092 189338
rect 145858 64736 145982 64764
rect 145750 50235 145802 50241
rect 145750 50177 145802 50183
rect 145858 50167 145886 64736
rect 145942 64443 145994 64449
rect 145942 64385 145994 64391
rect 145954 50685 145982 64385
rect 146050 51203 146078 189329
rect 146146 144665 146174 240537
rect 146612 239862 146668 239871
rect 146612 239797 146668 239806
rect 146626 239089 146654 239797
rect 146614 239083 146666 239089
rect 146614 239025 146666 239031
rect 146818 237628 146846 270771
rect 149602 245791 149630 277856
rect 149686 273197 149738 273203
rect 149686 273139 149738 273145
rect 149588 245782 149644 245791
rect 149588 245717 149644 245726
rect 149590 244781 149642 244787
rect 149590 244723 149642 244729
rect 149602 239829 149630 244723
rect 149590 239823 149642 239829
rect 149590 239765 149642 239771
rect 146434 237600 146846 237628
rect 148342 237603 148394 237609
rect 146324 236902 146380 236911
rect 146324 236837 146380 236846
rect 146228 185250 146284 185259
rect 146228 185185 146284 185194
rect 146134 144659 146186 144665
rect 146134 144601 146186 144607
rect 146134 144511 146186 144517
rect 146134 144453 146186 144459
rect 146146 129421 146174 144453
rect 146134 129415 146186 129421
rect 146134 129357 146186 129363
rect 146134 128527 146186 128533
rect 146134 128469 146186 128475
rect 146146 124907 146174 128469
rect 146134 124901 146186 124907
rect 146134 124843 146186 124849
rect 146134 124753 146186 124759
rect 146134 124695 146186 124701
rect 146146 115435 146174 124695
rect 146134 115429 146186 115435
rect 146134 115371 146186 115377
rect 146134 115059 146186 115065
rect 146134 115001 146186 115007
rect 146146 103669 146174 115001
rect 146134 103663 146186 103669
rect 146134 103605 146186 103611
rect 146132 99854 146188 99863
rect 146132 99789 146188 99798
rect 146146 97971 146174 99789
rect 146134 97965 146186 97971
rect 146134 97907 146186 97913
rect 146132 89642 146188 89651
rect 146132 89577 146188 89586
rect 146146 89461 146174 89577
rect 146134 89455 146186 89461
rect 146134 89397 146186 89403
rect 146132 83574 146188 83583
rect 146132 83509 146188 83518
rect 146146 75253 146174 83509
rect 146134 75247 146186 75253
rect 146134 75189 146186 75195
rect 146134 75099 146186 75105
rect 146134 75041 146186 75047
rect 146146 51943 146174 75041
rect 146134 51937 146186 51943
rect 146134 51879 146186 51885
rect 146038 51197 146090 51203
rect 146038 51139 146090 51145
rect 146242 51129 146270 185185
rect 146338 144855 146366 236837
rect 146434 224585 146462 237600
rect 148342 237545 148394 237551
rect 146516 235126 146572 235135
rect 146516 235061 146572 235070
rect 146422 224579 146474 224585
rect 146422 224521 146474 224527
rect 146420 186434 146476 186443
rect 146420 186369 146476 186378
rect 146324 144846 146380 144855
rect 146324 144781 146380 144790
rect 146326 144659 146378 144665
rect 146326 144601 146378 144607
rect 146338 140965 146366 144601
rect 146326 140959 146378 140965
rect 146326 140901 146378 140907
rect 146324 138334 146380 138343
rect 146324 138269 146380 138278
rect 146338 126831 146366 138269
rect 146326 126825 146378 126831
rect 146326 126767 146378 126773
rect 146326 126677 146378 126683
rect 146326 126619 146378 126625
rect 146338 125055 146366 126619
rect 146326 125049 146378 125055
rect 146326 124991 146378 124997
rect 146326 124901 146378 124907
rect 146326 124843 146378 124849
rect 146338 104853 146366 124843
rect 146326 104847 146378 104853
rect 146326 104789 146378 104795
rect 146324 104738 146380 104747
rect 146324 104673 146380 104682
rect 146338 103743 146366 104673
rect 146326 103737 146378 103743
rect 146326 103679 146378 103685
rect 146324 102814 146380 102823
rect 146324 102749 146380 102758
rect 146338 100857 146366 102749
rect 146326 100851 146378 100857
rect 146326 100793 146378 100799
rect 146324 99114 146380 99123
rect 146324 99049 146380 99058
rect 146338 98045 146366 99049
rect 146326 98039 146378 98045
rect 146326 97981 146378 97987
rect 146324 96302 146380 96311
rect 146324 96237 146380 96246
rect 146338 95085 146366 96237
rect 146326 95079 146378 95085
rect 146326 95021 146378 95027
rect 146324 94378 146380 94387
rect 146324 94313 146380 94322
rect 146338 92273 146366 94313
rect 146326 92267 146378 92273
rect 146326 92209 146378 92215
rect 146324 91418 146380 91427
rect 146324 91353 146380 91362
rect 146338 89313 146366 91353
rect 146326 89307 146378 89313
rect 146326 89249 146378 89255
rect 146324 79430 146380 79439
rect 146324 79365 146380 79374
rect 146338 77917 146366 79365
rect 146326 77911 146378 77917
rect 146326 77853 146378 77859
rect 146324 75730 146380 75739
rect 146324 75665 146380 75674
rect 146338 75327 146366 75665
rect 146326 75321 146378 75327
rect 146326 75263 146378 75269
rect 146326 75025 146378 75031
rect 146326 74967 146378 74973
rect 146338 52165 146366 74967
rect 146326 52159 146378 52165
rect 146326 52101 146378 52107
rect 146230 51123 146282 51129
rect 146230 51065 146282 51071
rect 146434 51055 146462 186369
rect 146530 128533 146558 235061
rect 146804 226690 146860 226699
rect 146804 226625 146860 226634
rect 146818 225695 146846 226625
rect 146806 225689 146858 225695
rect 146806 225631 146858 225637
rect 146804 225062 146860 225071
rect 146804 224997 146860 225006
rect 146818 224733 146846 224997
rect 146806 224727 146858 224733
rect 146806 224669 146858 224675
rect 146804 222990 146860 222999
rect 146804 222925 146860 222934
rect 146710 221989 146762 221995
rect 146710 221931 146762 221937
rect 146722 221815 146750 221931
rect 146818 221921 146846 222925
rect 146806 221915 146858 221921
rect 146806 221857 146858 221863
rect 146708 221806 146764 221815
rect 146708 221741 146764 221750
rect 146804 218254 146860 218263
rect 146804 218189 146860 218198
rect 146818 216371 146846 218189
rect 146806 216365 146858 216371
rect 146806 216307 146858 216313
rect 146804 213370 146860 213379
rect 146804 213305 146860 213314
rect 146818 213263 146846 213305
rect 146806 213257 146858 213263
rect 146806 213199 146858 213205
rect 146804 211742 146860 211751
rect 146804 211677 146860 211686
rect 146818 210303 146846 211677
rect 146806 210297 146858 210303
rect 146806 210239 146858 210245
rect 148246 210297 148298 210303
rect 148246 210239 148298 210245
rect 146708 209818 146764 209827
rect 146708 209753 146764 209762
rect 146722 207491 146750 209753
rect 146710 207485 146762 207491
rect 146710 207427 146762 207433
rect 146804 207450 146860 207459
rect 146804 207385 146806 207394
rect 146858 207385 146860 207394
rect 146806 207353 146858 207359
rect 146804 202122 146860 202131
rect 146804 202057 146860 202066
rect 146818 201719 146846 202057
rect 146806 201713 146858 201719
rect 146806 201655 146858 201661
rect 146804 199606 146860 199615
rect 146804 199541 146860 199550
rect 146818 198759 146846 199541
rect 146806 198753 146858 198759
rect 146806 198695 146858 198701
rect 146804 197830 146860 197839
rect 146804 197765 146860 197774
rect 146818 195873 146846 197765
rect 146806 195867 146858 195873
rect 146806 195809 146858 195815
rect 146708 192946 146764 192955
rect 146708 192881 146764 192890
rect 146722 190249 146750 192881
rect 146804 191762 146860 191771
rect 146804 191697 146860 191706
rect 146710 190243 146762 190249
rect 146710 190185 146762 190191
rect 146818 190175 146846 191697
rect 146806 190169 146858 190175
rect 146806 190111 146858 190117
rect 146804 188210 146860 188219
rect 146804 188145 146860 188154
rect 146818 187289 146846 188145
rect 146806 187283 146858 187289
rect 146806 187225 146858 187231
rect 146804 184510 146860 184519
rect 146804 184445 146860 184454
rect 146818 184403 146846 184445
rect 146806 184397 146858 184403
rect 146806 184339 146858 184345
rect 146612 180514 146668 180523
rect 146612 180449 146668 180458
rect 146518 128527 146570 128533
rect 146518 128469 146570 128475
rect 146516 127678 146572 127687
rect 146516 127613 146572 127622
rect 146530 126757 146558 127613
rect 146518 126751 146570 126757
rect 146518 126693 146570 126699
rect 146518 125419 146570 125425
rect 146518 125361 146570 125367
rect 146530 106851 146558 125361
rect 146518 106845 146570 106851
rect 146518 106787 146570 106793
rect 146516 106514 146572 106523
rect 146516 106449 146518 106458
rect 146570 106449 146572 106458
rect 146518 106417 146570 106423
rect 146518 104403 146570 104409
rect 146518 104345 146570 104351
rect 146530 104155 146558 104345
rect 146516 104146 146572 104155
rect 146516 104081 146572 104090
rect 146516 101630 146572 101639
rect 146516 101565 146518 101574
rect 146570 101565 146572 101574
rect 146518 101533 146570 101539
rect 146518 98113 146570 98119
rect 146516 98078 146518 98087
rect 146570 98078 146572 98087
rect 146516 98013 146572 98022
rect 146516 95562 146572 95571
rect 146516 95497 146572 95506
rect 146530 95159 146558 95497
rect 146518 95153 146570 95159
rect 146518 95095 146570 95101
rect 146516 92750 146572 92759
rect 146516 92685 146572 92694
rect 146530 92199 146558 92685
rect 146518 92193 146570 92199
rect 146518 92135 146570 92141
rect 146516 90826 146572 90835
rect 146516 90761 146572 90770
rect 146530 89387 146558 90761
rect 146518 89381 146570 89387
rect 146518 89323 146570 89329
rect 146516 85942 146572 85951
rect 146516 85877 146572 85886
rect 146530 85021 146558 85877
rect 146518 85015 146570 85021
rect 146518 84957 146570 84963
rect 146516 82390 146572 82399
rect 146516 82325 146572 82334
rect 146530 82135 146558 82325
rect 146518 82129 146570 82135
rect 146518 82071 146570 82077
rect 146516 78690 146572 78699
rect 146516 78625 146572 78634
rect 146530 77843 146558 78625
rect 146518 77837 146570 77843
rect 146518 77779 146570 77785
rect 146518 75247 146570 75253
rect 146518 75189 146570 75195
rect 146530 52313 146558 75189
rect 146518 52307 146570 52313
rect 146518 52249 146570 52255
rect 146422 51049 146474 51055
rect 146422 50991 146474 50997
rect 146626 50981 146654 180449
rect 146806 178625 146858 178631
rect 146804 178590 146806 178599
rect 146858 178590 146860 178599
rect 146804 178525 146860 178534
rect 146804 176074 146860 176083
rect 146804 176009 146860 176018
rect 146818 175893 146846 176009
rect 146806 175887 146858 175893
rect 146806 175829 146858 175835
rect 146804 171338 146860 171347
rect 146804 171273 146860 171282
rect 146708 170154 146764 170163
rect 146708 170089 146764 170098
rect 146722 162888 146750 170089
rect 146818 169973 146846 171273
rect 146806 169967 146858 169973
rect 146806 169909 146858 169915
rect 146804 167638 146860 167647
rect 146804 167573 146860 167582
rect 146818 167161 146846 167573
rect 146806 167155 146858 167161
rect 146806 167097 146858 167103
rect 146722 162860 146846 162888
rect 146710 162789 146762 162795
rect 146710 162731 146762 162737
rect 146722 74069 146750 162731
rect 146710 74063 146762 74069
rect 146710 74005 146762 74011
rect 146708 73954 146764 73963
rect 146708 73889 146764 73898
rect 146722 72071 146750 73889
rect 146710 72065 146762 72071
rect 146710 72007 146762 72013
rect 146708 70994 146764 71003
rect 146708 70929 146710 70938
rect 146762 70929 146764 70938
rect 146710 70897 146762 70903
rect 146708 67442 146764 67451
rect 146708 67377 146710 67386
rect 146762 67377 146764 67386
rect 146710 67345 146762 67351
rect 146818 66540 146846 162860
rect 146900 136114 146956 136123
rect 146900 136049 146956 136058
rect 146914 136007 146942 136049
rect 146902 136001 146954 136007
rect 146902 135943 146954 135949
rect 146902 135039 146954 135045
rect 146902 134981 146954 134987
rect 146914 115065 146942 134981
rect 146996 126938 147052 126947
rect 146996 126873 146998 126882
rect 147050 126873 147052 126882
rect 146998 126841 147050 126847
rect 148150 115577 148202 115583
rect 148150 115519 148202 115525
rect 146902 115059 146954 115065
rect 146902 115001 146954 115007
rect 147958 112691 148010 112697
rect 147958 112633 148010 112639
rect 147862 109583 147914 109589
rect 147862 109525 147914 109531
rect 147766 106623 147818 106629
rect 147766 106565 147818 106571
rect 146902 104847 146954 104853
rect 146902 104789 146954 104795
rect 146914 103521 146942 104789
rect 146902 103515 146954 103521
rect 146902 103457 146954 103463
rect 146722 66512 146846 66540
rect 146722 65652 146750 66512
rect 146804 66406 146860 66415
rect 146804 66341 146860 66350
rect 146818 66299 146846 66341
rect 146806 66293 146858 66299
rect 146806 66235 146858 66241
rect 146722 65624 146846 65652
rect 146708 65518 146764 65527
rect 146708 65453 146764 65462
rect 146722 64893 146750 65453
rect 146818 64912 146846 65624
rect 146710 64887 146762 64893
rect 146818 64884 146942 64912
rect 146710 64829 146762 64835
rect 146806 64813 146858 64819
rect 146804 64778 146806 64787
rect 146858 64778 146860 64787
rect 146804 64713 146860 64722
rect 146914 64616 146942 64884
rect 146722 64588 146942 64616
rect 146614 50975 146666 50981
rect 146614 50917 146666 50923
rect 146722 50759 146750 64588
rect 146902 63407 146954 63413
rect 146902 63349 146954 63355
rect 146804 62558 146860 62567
rect 146804 62493 146806 62502
rect 146858 62493 146860 62502
rect 146806 62461 146858 62467
rect 146914 62419 146942 63349
rect 146900 62410 146956 62419
rect 146900 62345 146956 62354
rect 146900 60782 146956 60791
rect 146900 60717 146956 60726
rect 146914 60453 146942 60717
rect 146902 60447 146954 60453
rect 146902 60389 146954 60395
rect 146806 59633 146858 59639
rect 146804 59598 146806 59607
rect 146858 59598 146860 59607
rect 146804 59533 146860 59542
rect 146806 59041 146858 59047
rect 146806 58983 146858 58989
rect 146818 58719 146846 58983
rect 146804 58710 146860 58719
rect 146804 58645 146860 58654
rect 146806 57117 146858 57123
rect 146804 57082 146806 57091
rect 146858 57082 146860 57091
rect 146804 57017 146860 57026
rect 146806 56969 146858 56975
rect 146806 56911 146858 56917
rect 146710 50753 146762 50759
rect 146710 50695 146762 50701
rect 145942 50679 145994 50685
rect 145942 50621 145994 50627
rect 145846 50161 145898 50167
rect 145846 50103 145898 50109
rect 146818 49945 146846 56911
rect 146806 49939 146858 49945
rect 146806 49881 146858 49887
rect 145462 49717 145514 49723
rect 145462 49659 145514 49665
rect 145072 48544 145100 49208
rect 145072 48516 145669 48544
rect 142114 46680 142416 46708
rect 142114 40219 142142 46680
rect 145641 45724 145669 48516
rect 147778 47651 147806 106565
rect 147874 47725 147902 109525
rect 147862 47719 147914 47725
rect 147862 47661 147914 47667
rect 147766 47645 147818 47651
rect 147766 47587 147818 47593
rect 147970 47503 147998 112633
rect 148054 112469 148106 112475
rect 148054 112411 148106 112417
rect 148066 47577 148094 112411
rect 148162 48095 148190 115519
rect 148150 48089 148202 48095
rect 148150 48031 148202 48037
rect 148054 47571 148106 47577
rect 148054 47513 148106 47519
rect 147958 47497 148010 47503
rect 147958 47439 148010 47445
rect 148258 47133 148286 210239
rect 148354 74513 148382 237545
rect 149698 224511 149726 273139
rect 150274 272093 150302 277870
rect 151426 273203 151454 277870
rect 152674 273203 152702 277870
rect 153826 273425 153854 277870
rect 155088 277856 155486 277884
rect 153814 273419 153866 273425
rect 153814 273361 153866 273367
rect 151414 273197 151466 273203
rect 151414 273139 151466 273145
rect 152566 273197 152618 273203
rect 152566 273139 152618 273145
rect 152662 273197 152714 273203
rect 152662 273139 152714 273145
rect 155350 273197 155402 273203
rect 155350 273139 155402 273145
rect 150262 272087 150314 272093
rect 150262 272029 150314 272035
rect 151126 246039 151178 246045
rect 151126 245981 151178 245987
rect 151138 245897 151166 245981
rect 151126 245891 151178 245897
rect 151126 245833 151178 245839
rect 151126 230573 151178 230579
rect 151126 230515 151178 230521
rect 149686 224505 149738 224511
rect 149686 224447 149738 224453
rect 148438 190169 148490 190175
rect 148438 190111 148490 190117
rect 148342 74507 148394 74513
rect 148342 74449 148394 74455
rect 148342 60521 148394 60527
rect 148342 60463 148394 60469
rect 148354 54163 148382 60463
rect 148342 54157 148394 54163
rect 148342 54099 148394 54105
rect 148246 47127 148298 47133
rect 148246 47069 148298 47075
rect 148450 46541 148478 190111
rect 148534 181585 148586 181591
rect 148534 181527 148586 181533
rect 148546 47207 148574 181527
rect 148630 178699 148682 178705
rect 148630 178641 148682 178647
rect 148534 47201 148586 47207
rect 148534 47143 148586 47149
rect 148642 46837 148670 178641
rect 148726 175887 148778 175893
rect 148726 175829 148778 175835
rect 148738 46911 148766 175829
rect 148822 167081 148874 167087
rect 148822 167023 148874 167029
rect 148726 46905 148778 46911
rect 148726 46847 148778 46853
rect 148630 46831 148682 46837
rect 148630 46773 148682 46779
rect 148834 46763 148862 167023
rect 148918 164195 148970 164201
rect 148918 164137 148970 164143
rect 148822 46757 148874 46763
rect 148822 46699 148874 46705
rect 148930 46615 148958 164137
rect 149014 161309 149066 161315
rect 149014 161251 149066 161257
rect 149026 46985 149054 161251
rect 149110 158497 149162 158503
rect 149110 158439 149162 158445
rect 149122 47059 149150 158439
rect 149206 141255 149258 141261
rect 149206 141197 149258 141203
rect 149218 48169 149246 141197
rect 149302 136001 149354 136007
rect 149302 135943 149354 135949
rect 149314 48243 149342 135943
rect 149398 126899 149450 126905
rect 149398 126841 149450 126847
rect 149302 48237 149354 48243
rect 149302 48179 149354 48185
rect 149206 48163 149258 48169
rect 149206 48105 149258 48111
rect 149410 48021 149438 126841
rect 149494 121127 149546 121133
rect 149494 121069 149546 121075
rect 149398 48015 149450 48021
rect 149398 47957 149450 47963
rect 149506 47947 149534 121069
rect 149590 121053 149642 121059
rect 149590 120995 149642 121001
rect 149494 47941 149546 47947
rect 149494 47883 149546 47889
rect 149602 47799 149630 120995
rect 149686 116243 149738 116249
rect 149686 116185 149738 116191
rect 149698 47873 149726 116185
rect 151138 100561 151166 230515
rect 152578 224437 152606 273139
rect 155362 245495 155390 273139
rect 155348 245486 155404 245495
rect 155348 245421 155404 245430
rect 152566 224431 152618 224437
rect 152566 224373 152618 224379
rect 155458 221773 155486 277856
rect 156226 273203 156254 277870
rect 157474 273351 157502 277870
rect 157462 273345 157514 273351
rect 157462 273287 157514 273293
rect 156214 273197 156266 273203
rect 158326 273197 158378 273203
rect 156214 273139 156266 273145
rect 156884 273162 156940 273171
rect 158326 273139 158378 273145
rect 156884 273097 156940 273106
rect 156898 272431 156926 273097
rect 156980 272570 157036 272579
rect 156980 272505 157036 272514
rect 156884 272422 156940 272431
rect 156884 272357 156940 272366
rect 156886 271495 156938 271501
rect 156886 271437 156938 271443
rect 156898 271279 156926 271437
rect 156886 271273 156938 271279
rect 156886 271215 156938 271221
rect 156994 270803 157022 272505
rect 156980 270794 157036 270803
rect 156980 270729 157036 270738
rect 158338 245199 158366 273139
rect 158626 270021 158654 277870
rect 158614 270015 158666 270021
rect 158614 269957 158666 269963
rect 159874 263509 159902 277870
rect 161026 273425 161054 277870
rect 160918 273419 160970 273425
rect 160918 273361 160970 273367
rect 161014 273419 161066 273425
rect 161014 273361 161066 273367
rect 161122 273416 161342 273444
rect 160930 273296 160958 273361
rect 161122 273296 161150 273416
rect 160930 273268 161150 273296
rect 161314 273277 161342 273416
rect 161302 273271 161354 273277
rect 161302 273213 161354 273219
rect 162178 273203 162206 277870
rect 163440 277856 164030 277884
rect 162166 273197 162218 273203
rect 162166 273139 162218 273145
rect 160820 271830 160876 271839
rect 161204 271830 161260 271839
rect 160876 271774 161204 271779
rect 160820 271765 161260 271774
rect 160834 271751 161246 271765
rect 161110 271717 161162 271723
rect 161108 271682 161110 271691
rect 161162 271682 161164 271691
rect 161108 271617 161164 271626
rect 161206 270015 161258 270021
rect 161206 269957 161258 269963
rect 159862 263503 159914 263509
rect 159862 263445 159914 263451
rect 161110 263503 161162 263509
rect 161110 263445 161162 263451
rect 158324 245190 158380 245199
rect 158324 245125 158380 245134
rect 161122 245051 161150 263445
rect 161108 245042 161164 245051
rect 161108 244977 161164 244986
rect 157750 239823 157802 239829
rect 157750 239765 157802 239771
rect 157762 237799 157790 239765
rect 157748 237790 157804 237799
rect 157748 237725 157804 237734
rect 156886 225689 156938 225695
rect 156886 225631 156938 225637
rect 155446 221767 155498 221773
rect 155446 221709 155498 221715
rect 154006 216365 154058 216371
rect 154006 216307 154058 216313
rect 151222 190243 151274 190249
rect 151222 190185 151274 190191
rect 151126 100555 151178 100561
rect 151126 100497 151178 100503
rect 151234 94863 151262 190185
rect 151414 129711 151466 129717
rect 151414 129653 151466 129659
rect 151318 100851 151370 100857
rect 151318 100793 151370 100799
rect 151222 94857 151274 94863
rect 151222 94799 151274 94805
rect 151126 89455 151178 89461
rect 151126 89397 151178 89403
rect 151138 71997 151166 89397
rect 151126 71991 151178 71997
rect 151126 71933 151178 71939
rect 149782 70955 149834 70961
rect 149782 70897 149834 70903
rect 149794 69037 149822 70897
rect 149782 69031 149834 69037
rect 149782 68973 149834 68979
rect 149782 62519 149834 62525
rect 149782 62461 149834 62467
rect 149794 60379 149822 62461
rect 151126 60595 151178 60601
rect 151126 60537 151178 60543
rect 149782 60373 149834 60379
rect 149782 60315 149834 60321
rect 151138 54681 151166 60537
rect 151126 54675 151178 54681
rect 151126 54617 151178 54623
rect 151330 52757 151358 100793
rect 151426 83541 151454 129653
rect 154018 97897 154046 216307
rect 154102 144363 154154 144369
rect 154102 144305 154154 144311
rect 154006 97891 154058 97897
rect 154006 97833 154058 97839
rect 154006 92267 154058 92273
rect 154006 92209 154058 92215
rect 151414 83535 151466 83541
rect 151414 83477 151466 83483
rect 154018 74883 154046 92209
rect 154114 86427 154142 144305
rect 156898 97823 156926 225631
rect 161218 221699 161246 269957
rect 164002 247271 164030 277856
rect 164278 273271 164330 273277
rect 164278 273213 164330 273219
rect 164086 273197 164138 273203
rect 164086 273139 164138 273145
rect 163988 247262 164044 247271
rect 163988 247197 164044 247206
rect 161302 237603 161354 237609
rect 161302 237545 161354 237551
rect 161314 237461 161342 237545
rect 161302 237455 161354 237461
rect 161302 237397 161354 237403
rect 161206 221693 161258 221699
rect 161206 221635 161258 221641
rect 164098 221625 164126 273139
rect 164290 272093 164318 273213
rect 164578 272093 164606 277870
rect 164278 272087 164330 272093
rect 164278 272029 164330 272035
rect 164566 272087 164618 272093
rect 164566 272029 164618 272035
rect 165826 271945 165854 277870
rect 165814 271939 165866 271945
rect 165814 271881 165866 271887
rect 166594 271723 166622 278004
rect 182230 277933 182282 277939
rect 168144 277856 168446 277884
rect 169296 277856 169886 277884
rect 182230 277875 182282 277881
rect 166966 272753 167018 272759
rect 166966 272695 167018 272701
rect 166978 272556 167006 272695
rect 166786 272528 167006 272556
rect 166786 271797 166814 272528
rect 166966 271939 167018 271945
rect 166966 271881 167018 271887
rect 166774 271791 166826 271797
rect 166774 271733 166826 271739
rect 166582 271717 166634 271723
rect 166582 271659 166634 271665
rect 166870 271717 166922 271723
rect 166870 271659 166922 271665
rect 166882 244903 166910 271659
rect 166868 244894 166924 244903
rect 166868 244829 166924 244838
rect 165526 233311 165578 233317
rect 165526 233253 165578 233259
rect 164086 221619 164138 221625
rect 164086 221561 164138 221567
rect 159766 201713 159818 201719
rect 159766 201655 159818 201661
rect 156982 167155 157034 167161
rect 156982 167097 157034 167103
rect 156886 97817 156938 97823
rect 156886 97759 156938 97765
rect 156994 89239 157022 167097
rect 157078 101591 157130 101597
rect 157078 101533 157130 101539
rect 156982 89233 157034 89239
rect 156982 89175 157034 89181
rect 154102 86421 154154 86427
rect 154102 86363 154154 86369
rect 157090 77769 157118 101533
rect 159778 100487 159806 201655
rect 162646 201639 162698 201645
rect 162646 201581 162698 201587
rect 159862 169967 159914 169973
rect 159862 169909 159914 169915
rect 159766 100481 159818 100487
rect 159766 100423 159818 100429
rect 159874 89165 159902 169909
rect 159958 106475 160010 106481
rect 159958 106417 160010 106423
rect 159862 89159 159914 89165
rect 159862 89101 159914 89107
rect 157078 77763 157130 77769
rect 157078 77705 157130 77711
rect 156406 75025 156458 75031
rect 156406 74967 156458 74973
rect 154006 74877 154058 74883
rect 154006 74819 154058 74825
rect 153910 72065 153962 72071
rect 153910 72007 153962 72013
rect 153922 68963 153950 72007
rect 153910 68957 153962 68963
rect 153910 68899 153962 68905
rect 156418 68889 156446 74967
rect 156406 68883 156458 68889
rect 156406 68825 156458 68831
rect 152662 67403 152714 67409
rect 152662 67345 152714 67351
rect 152674 66151 152702 67345
rect 158326 66441 158378 66447
rect 158326 66383 158378 66389
rect 152662 66145 152714 66151
rect 152662 66087 152714 66093
rect 158338 66077 158366 66383
rect 158326 66071 158378 66077
rect 158326 66013 158378 66019
rect 156310 60743 156362 60749
rect 156310 60685 156362 60691
rect 152662 60669 152714 60675
rect 152662 60611 152714 60617
rect 152674 56531 152702 60611
rect 156322 57123 156350 60685
rect 156310 57117 156362 57123
rect 156310 57059 156362 57065
rect 152662 56525 152714 56531
rect 152662 56467 152714 56473
rect 159970 52905 159998 106417
rect 160054 104403 160106 104409
rect 160054 104345 160106 104351
rect 160066 77695 160094 104345
rect 160054 77689 160106 77695
rect 160054 77631 160106 77637
rect 160054 75099 160106 75105
rect 160054 75041 160106 75047
rect 160066 68815 160094 75041
rect 161494 74951 161546 74957
rect 161494 74893 161546 74899
rect 161506 71923 161534 74893
rect 161494 71917 161546 71923
rect 161494 71859 161546 71865
rect 160054 68809 160106 68815
rect 160054 68751 160106 68757
rect 160534 60817 160586 60823
rect 160534 60759 160586 60765
rect 160546 59639 160574 60759
rect 160534 59633 160586 59639
rect 160534 59575 160586 59581
rect 159958 52899 160010 52905
rect 159958 52841 160010 52847
rect 151318 52751 151370 52757
rect 151318 52693 151370 52699
rect 162658 48317 162686 201581
rect 162742 172853 162794 172859
rect 162742 172795 162794 172801
rect 162754 89091 162782 172795
rect 162838 106919 162890 106925
rect 162838 106861 162890 106867
rect 162742 89085 162794 89091
rect 162742 89027 162794 89033
rect 162850 77621 162878 106861
rect 162838 77615 162890 77621
rect 162838 77557 162890 77563
rect 162646 48311 162698 48317
rect 162646 48253 162698 48259
rect 165538 48211 165566 233253
rect 166978 221551 167006 271881
rect 168118 271495 168170 271501
rect 168118 271437 168170 271443
rect 168130 271279 168158 271437
rect 168118 271273 168170 271279
rect 168118 271215 168170 271221
rect 168418 270835 168446 277856
rect 168406 270829 168458 270835
rect 168406 270771 168458 270777
rect 168406 236271 168458 236277
rect 168406 236213 168458 236219
rect 166966 221545 167018 221551
rect 166966 221487 167018 221493
rect 165622 207485 165674 207491
rect 165622 207427 165674 207433
rect 165634 94789 165662 207427
rect 165718 132967 165770 132973
rect 165718 132909 165770 132915
rect 165622 94783 165674 94789
rect 165622 94725 165674 94731
rect 165622 89381 165674 89387
rect 165622 89323 165674 89329
rect 165634 71849 165662 89323
rect 165730 83467 165758 132909
rect 165718 83461 165770 83467
rect 165718 83403 165770 83409
rect 165622 71843 165674 71849
rect 165622 71785 165674 71791
rect 168418 48803 168446 236213
rect 169858 221477 169886 277856
rect 170530 271945 170558 277870
rect 170518 271939 170570 271945
rect 170518 271881 170570 271887
rect 171682 271723 171710 277870
rect 172726 271939 172778 271945
rect 172726 271881 172778 271887
rect 171670 271717 171722 271723
rect 171670 271659 171722 271665
rect 172738 246679 172766 271881
rect 172930 269873 172958 277870
rect 172918 269867 172970 269873
rect 172918 269809 172970 269815
rect 174082 269651 174110 277870
rect 175330 271501 175358 277870
rect 176482 271797 176510 277870
rect 177044 273162 177100 273171
rect 177044 273097 177100 273106
rect 177058 272431 177086 273097
rect 177140 272570 177196 272579
rect 177140 272505 177196 272514
rect 177044 272422 177100 272431
rect 177044 272357 177100 272366
rect 176470 271791 176522 271797
rect 176470 271733 176522 271739
rect 175318 271495 175370 271501
rect 175318 271437 175370 271443
rect 175606 270903 175658 270909
rect 175606 270845 175658 270851
rect 175510 270829 175562 270835
rect 175618 270780 175646 270845
rect 177154 270803 177182 272505
rect 177634 271945 177662 277870
rect 177622 271939 177674 271945
rect 177622 271881 177674 271887
rect 178390 271939 178442 271945
rect 178390 271881 178442 271887
rect 175562 270777 175646 270780
rect 175510 270771 175646 270777
rect 175522 270752 175646 270771
rect 177140 270794 177196 270803
rect 177140 270729 177196 270738
rect 175606 269867 175658 269873
rect 175606 269809 175658 269815
rect 174070 269645 174122 269651
rect 174070 269587 174122 269593
rect 175510 269645 175562 269651
rect 175510 269587 175562 269593
rect 175522 247567 175550 269587
rect 175508 247558 175564 247567
rect 175508 247493 175564 247502
rect 172724 246670 172780 246679
rect 172724 246605 172780 246614
rect 170902 246187 170954 246193
rect 170902 246129 170954 246135
rect 170914 246045 170942 246129
rect 170902 246039 170954 246045
rect 170902 245981 170954 245987
rect 174166 239083 174218 239089
rect 174166 239025 174218 239031
rect 171286 237825 171338 237831
rect 171286 237767 171338 237773
rect 171298 237461 171326 237767
rect 171286 237455 171338 237461
rect 171286 237397 171338 237403
rect 171286 236197 171338 236203
rect 171286 236139 171338 236145
rect 169846 221471 169898 221477
rect 169846 221413 169898 221419
rect 168502 213257 168554 213263
rect 168502 213199 168554 213205
rect 168514 94715 168542 213199
rect 168598 138295 168650 138301
rect 168598 138237 168650 138243
rect 168502 94709 168554 94715
rect 168502 94651 168554 94657
rect 168502 89307 168554 89313
rect 168502 89249 168554 89255
rect 168514 71775 168542 89249
rect 168610 83393 168638 138237
rect 168598 83387 168650 83393
rect 168598 83329 168650 83335
rect 168502 71769 168554 71775
rect 168502 71711 168554 71717
rect 168404 48794 168460 48803
rect 168404 48729 168460 48738
rect 171298 48655 171326 236139
rect 171382 213183 171434 213189
rect 171382 213125 171434 213131
rect 171394 97749 171422 213125
rect 171574 141699 171626 141705
rect 171574 141641 171626 141647
rect 171478 118315 171530 118321
rect 171478 118257 171530 118263
rect 171382 97743 171434 97749
rect 171382 97685 171434 97691
rect 171382 92193 171434 92199
rect 171382 92135 171434 92141
rect 171394 71701 171422 92135
rect 171382 71695 171434 71701
rect 171382 71637 171434 71643
rect 171490 52239 171518 118257
rect 171586 83319 171614 141641
rect 171574 83313 171626 83319
rect 171574 83255 171626 83261
rect 171478 52233 171530 52239
rect 171478 52175 171530 52181
rect 171284 48646 171340 48655
rect 171284 48581 171340 48590
rect 174178 48507 174206 239025
rect 174262 218955 174314 218961
rect 174262 218897 174314 218903
rect 174274 97675 174302 218897
rect 175618 218887 175646 269809
rect 178402 243571 178430 271881
rect 178486 271791 178538 271797
rect 178486 271733 178538 271739
rect 178388 243562 178444 243571
rect 178388 243497 178444 243506
rect 177046 221989 177098 221995
rect 177046 221931 177098 221937
rect 175606 218881 175658 218887
rect 175606 218823 175658 218829
rect 174358 146953 174410 146959
rect 174358 146895 174410 146901
rect 174262 97669 174314 97675
rect 174262 97611 174314 97617
rect 174370 86353 174398 146895
rect 174454 95153 174506 95159
rect 174454 95095 174506 95101
rect 174358 86347 174410 86353
rect 174358 86289 174410 86295
rect 174466 74809 174494 95095
rect 174454 74803 174506 74809
rect 174454 74745 174506 74751
rect 174164 48498 174220 48507
rect 174164 48433 174220 48442
rect 165524 48202 165580 48211
rect 165524 48137 165580 48146
rect 149686 47867 149738 47873
rect 149686 47809 149738 47815
rect 149590 47793 149642 47799
rect 149590 47735 149642 47741
rect 177058 47429 177086 221931
rect 178498 218813 178526 271733
rect 178882 271723 178910 277870
rect 180034 271945 180062 277870
rect 180022 271939 180074 271945
rect 180022 271881 180074 271887
rect 178870 271717 178922 271723
rect 178870 271659 178922 271665
rect 181282 247419 181310 277870
rect 181366 271939 181418 271945
rect 181366 271881 181418 271887
rect 181268 247410 181324 247419
rect 181268 247345 181324 247354
rect 179926 221915 179978 221921
rect 179926 221857 179978 221863
rect 178486 218807 178538 218813
rect 178486 218749 178538 218755
rect 177142 149839 177194 149845
rect 177142 149781 177194 149787
rect 177154 86279 177182 149781
rect 177238 95079 177290 95085
rect 177238 95021 177290 95027
rect 177142 86273 177194 86279
rect 177142 86215 177194 86221
rect 177250 74735 177278 95021
rect 177238 74729 177290 74735
rect 177238 74671 177290 74677
rect 177046 47423 177098 47429
rect 177046 47365 177098 47371
rect 179938 47355 179966 221857
rect 181378 218739 181406 271881
rect 182242 262177 182270 277875
rect 182434 271649 182462 277870
rect 183600 277856 184286 277884
rect 182422 271643 182474 271649
rect 182422 271585 182474 271591
rect 182230 262171 182282 262177
rect 182230 262113 182282 262119
rect 181460 247262 181516 247271
rect 181460 247197 181516 247206
rect 181474 246859 181502 247197
rect 181462 246853 181514 246859
rect 181462 246795 181514 246801
rect 181558 246113 181610 246119
rect 181474 246061 181558 246064
rect 181474 246055 181610 246061
rect 181474 246045 181598 246055
rect 181462 246039 181598 246045
rect 181514 246036 181598 246039
rect 181462 245981 181514 245987
rect 181462 237973 181514 237979
rect 181462 237915 181514 237921
rect 181474 237831 181502 237915
rect 181462 237825 181514 237831
rect 181462 237767 181514 237773
rect 182806 221841 182858 221847
rect 182806 221783 182858 221789
rect 181366 218733 181418 218739
rect 181366 218675 181418 218681
rect 180022 152799 180074 152805
rect 180022 152741 180074 152747
rect 180034 86205 180062 152741
rect 180118 98113 180170 98119
rect 180118 98055 180170 98061
rect 180022 86199 180074 86205
rect 180022 86141 180074 86147
rect 180130 74661 180158 98055
rect 182818 97601 182846 221783
rect 184258 218665 184286 277856
rect 184738 271057 184766 277870
rect 185986 271575 186014 277870
rect 187030 271939 187082 271945
rect 186850 271899 187030 271927
rect 186850 271797 186878 271899
rect 187030 271881 187082 271887
rect 186838 271791 186890 271797
rect 186838 271733 186890 271739
rect 187030 271791 187082 271797
rect 187030 271733 187082 271739
rect 185974 271569 186026 271575
rect 187042 271520 187070 271733
rect 185974 271511 186026 271517
rect 186850 271501 187070 271520
rect 186838 271495 187070 271501
rect 186890 271492 187070 271495
rect 186838 271437 186890 271443
rect 184726 271051 184778 271057
rect 184726 270993 184778 270999
rect 187030 271051 187082 271057
rect 187030 270993 187082 270999
rect 187042 246087 187070 270993
rect 187028 246078 187084 246087
rect 187028 246013 187084 246022
rect 184246 218659 184298 218665
rect 184246 218601 184298 218607
rect 187138 216001 187166 277870
rect 188386 271131 188414 277870
rect 188374 271125 188426 271131
rect 188374 271067 188426 271073
rect 189538 270909 189566 277870
rect 190582 273493 190634 273499
rect 190582 273435 190634 273441
rect 190678 273493 190730 273499
rect 190678 273435 190730 273441
rect 190594 271131 190622 273435
rect 190690 272907 190718 273435
rect 190786 272907 190814 277870
rect 190678 272901 190730 272907
rect 190678 272843 190730 272849
rect 190774 272901 190826 272907
rect 190774 272843 190826 272849
rect 190006 271125 190058 271131
rect 190006 271067 190058 271073
rect 190582 271125 190634 271131
rect 190582 271067 190634 271073
rect 189526 270903 189578 270909
rect 189526 270845 189578 270851
rect 190018 247123 190046 271067
rect 191938 270761 191966 277870
rect 192886 272901 192938 272907
rect 192886 272843 192938 272849
rect 191926 270755 191978 270761
rect 191926 270697 191978 270703
rect 190004 247114 190060 247123
rect 190004 247049 190060 247058
rect 187700 246522 187756 246531
rect 187700 246457 187756 246466
rect 187714 245643 187742 246457
rect 187700 245634 187756 245643
rect 187700 245569 187756 245578
rect 188566 227761 188618 227767
rect 188566 227703 188618 227709
rect 187126 215995 187178 216001
rect 187126 215937 187178 215943
rect 185686 195867 185738 195873
rect 185686 195809 185738 195815
rect 182902 152725 182954 152731
rect 182902 152667 182954 152673
rect 182806 97595 182858 97601
rect 182806 97537 182858 97543
rect 182914 86131 182942 152667
rect 182998 98039 183050 98045
rect 182998 97981 183050 97987
rect 182902 86125 182954 86131
rect 182902 86067 182954 86073
rect 180118 74655 180170 74661
rect 180118 74597 180170 74603
rect 183010 74587 183038 97981
rect 182998 74581 183050 74587
rect 182998 74523 183050 74529
rect 185698 48539 185726 195809
rect 185782 175739 185834 175745
rect 185782 175681 185834 175687
rect 185794 89017 185822 175681
rect 185878 109509 185930 109515
rect 185878 109451 185930 109457
rect 185782 89011 185834 89017
rect 185782 88953 185834 88959
rect 185890 77547 185918 109451
rect 185878 77541 185930 77547
rect 185878 77483 185930 77489
rect 188578 48613 188606 227703
rect 192898 215927 192926 272843
rect 193090 270835 193118 277870
rect 193078 270829 193130 270835
rect 193078 270771 193130 270777
rect 194338 270021 194366 277870
rect 195490 270761 195518 277870
rect 196738 275275 196766 277870
rect 196726 275269 196778 275275
rect 196726 275211 196778 275217
rect 198740 273754 198796 273763
rect 198740 273689 198796 273698
rect 198754 273573 198782 273689
rect 198742 273567 198794 273573
rect 198742 273509 198794 273515
rect 197204 273162 197260 273171
rect 197204 273097 197260 273106
rect 197110 272901 197162 272907
rect 197110 272843 197162 272849
rect 197122 272315 197150 272843
rect 197218 272431 197246 273097
rect 197396 272570 197452 272579
rect 197396 272505 197452 272514
rect 197204 272422 197260 272431
rect 197204 272357 197260 272366
rect 197110 272309 197162 272315
rect 197110 272251 197162 272257
rect 197206 272013 197258 272019
rect 197206 271955 197258 271961
rect 197302 272013 197354 272019
rect 197302 271955 197354 271961
rect 195862 271865 195914 271871
rect 195914 271825 195998 271853
rect 195862 271807 195914 271813
rect 195970 271353 195998 271825
rect 195958 271347 196010 271353
rect 195958 271289 196010 271295
rect 197110 271199 197162 271205
rect 195874 271159 196382 271187
rect 195874 271057 195902 271159
rect 195862 271051 195914 271057
rect 195862 270993 195914 270999
rect 196246 271051 196298 271057
rect 196246 270993 196298 270999
rect 195862 270829 195914 270835
rect 196258 270817 196286 270993
rect 196162 270789 196286 270817
rect 196162 270780 196190 270789
rect 195914 270777 196190 270780
rect 195862 270771 196190 270777
rect 195478 270755 195530 270761
rect 195874 270752 196190 270771
rect 195478 270697 195530 270703
rect 196354 270655 196382 271159
rect 197110 271141 197162 271147
rect 196340 270646 196396 270655
rect 196340 270581 196396 270590
rect 194326 270015 194378 270021
rect 194326 269957 194378 269963
rect 192982 262097 193034 262103
rect 192982 262039 193034 262045
rect 192994 253445 193022 262039
rect 197122 257663 197150 271141
rect 197218 267579 197246 271955
rect 197314 271501 197342 271955
rect 197302 271495 197354 271501
rect 197302 271437 197354 271443
rect 197410 270803 197438 272505
rect 197396 270794 197452 270803
rect 197396 270729 197452 270738
rect 197206 267573 197258 267579
rect 197206 267515 197258 267521
rect 199138 266617 199166 277870
rect 200194 275497 200222 277870
rect 200182 275491 200234 275497
rect 200182 275433 200234 275439
rect 199126 266611 199178 266617
rect 199126 266553 199178 266559
rect 201442 265211 201470 277870
rect 202594 271205 202622 277870
rect 202582 271199 202634 271205
rect 202582 271141 202634 271147
rect 203842 270465 203870 277870
rect 204514 271131 204542 278425
rect 265776 278473 266038 278476
rect 265776 278467 266090 278473
rect 265776 278448 266078 278467
rect 263732 278425 263788 278434
rect 223126 278393 223178 278399
rect 204502 271125 204554 271131
rect 204502 271067 204554 271073
rect 203830 270459 203882 270465
rect 203830 270401 203882 270407
rect 204994 267801 205022 277870
rect 205846 271495 205898 271501
rect 205846 271437 205898 271443
rect 205858 270835 205886 271437
rect 205846 270829 205898 270835
rect 205846 270771 205898 270777
rect 206242 270761 206270 277870
rect 207394 274313 207422 277870
rect 208546 276681 208574 277870
rect 208534 276675 208586 276681
rect 208534 276617 208586 276623
rect 207382 274307 207434 274313
rect 207382 274249 207434 274255
rect 209794 272315 209822 277870
rect 209782 272309 209834 272315
rect 209782 272251 209834 272257
rect 207862 272013 207914 272019
rect 207298 271945 207422 271964
rect 207862 271955 207914 271961
rect 207286 271939 207434 271945
rect 207338 271936 207382 271939
rect 207286 271881 207338 271887
rect 207382 271881 207434 271887
rect 207874 271816 207902 271955
rect 210274 271936 210686 271964
rect 210274 271871 210302 271936
rect 208054 271865 208106 271871
rect 207874 271813 208054 271816
rect 207874 271807 208106 271813
rect 210262 271865 210314 271871
rect 210262 271807 210314 271813
rect 210358 271865 210410 271871
rect 210358 271807 210410 271813
rect 207874 271788 208094 271807
rect 206614 271347 206666 271353
rect 206614 271289 206666 271295
rect 206230 270755 206282 270761
rect 206230 270697 206282 270703
rect 204982 267795 205034 267801
rect 204982 267737 205034 267743
rect 201430 265205 201482 265211
rect 201430 265147 201482 265153
rect 197110 257657 197162 257663
rect 197110 257599 197162 257605
rect 192982 253439 193034 253445
rect 192982 253381 193034 253387
rect 198742 253439 198794 253445
rect 198742 253381 198794 253387
rect 198754 247747 198782 253381
rect 205654 249295 205706 249301
rect 205654 249237 205706 249243
rect 198742 247741 198794 247747
rect 196820 247706 196876 247715
rect 198742 247683 198794 247689
rect 196820 247641 196876 247650
rect 196834 242239 196862 247641
rect 197204 247262 197260 247271
rect 197204 247197 197260 247206
rect 197218 246087 197246 247197
rect 197590 246853 197642 246859
rect 197590 246795 197642 246801
rect 197602 246235 197630 246795
rect 205078 246779 205130 246785
rect 205078 246721 205130 246727
rect 204886 246631 204938 246637
rect 204886 246573 204938 246579
rect 204694 246557 204746 246563
rect 204694 246499 204746 246505
rect 197588 246226 197644 246235
rect 197588 246161 197644 246170
rect 197204 246078 197260 246087
rect 197204 246013 197260 246022
rect 204502 244189 204554 244195
rect 204502 244131 204554 244137
rect 196820 242230 196876 242239
rect 196820 242165 196876 242174
rect 201526 237973 201578 237979
rect 201526 237915 201578 237921
rect 201538 237831 201566 237915
rect 201526 237825 201578 237831
rect 201526 237767 201578 237773
rect 202966 230499 203018 230505
rect 202966 230441 203018 230447
rect 194326 227687 194378 227693
rect 194326 227629 194378 227635
rect 192886 215921 192938 215927
rect 192886 215863 192938 215869
rect 191446 198753 191498 198759
rect 191446 198695 191498 198701
rect 188662 181511 188714 181517
rect 188662 181453 188714 181459
rect 188674 91829 188702 181453
rect 188758 118241 188810 118247
rect 188758 118183 188810 118189
rect 188662 91823 188714 91829
rect 188662 91765 188714 91771
rect 188770 80359 188798 118183
rect 188758 80353 188810 80359
rect 188758 80295 188810 80301
rect 190006 77911 190058 77917
rect 190006 77853 190058 77859
rect 190018 77251 190046 77853
rect 190006 77245 190058 77251
rect 190006 77187 190058 77193
rect 188566 48607 188618 48613
rect 188566 48549 188618 48555
rect 185686 48533 185738 48539
rect 185686 48475 185738 48481
rect 179926 47349 179978 47355
rect 179926 47291 179978 47297
rect 149110 47053 149162 47059
rect 149110 46995 149162 47001
rect 149014 46979 149066 46985
rect 149014 46921 149066 46927
rect 148918 46609 148970 46615
rect 148918 46551 148970 46557
rect 148438 46535 148490 46541
rect 148438 46477 148490 46483
rect 191458 46245 191486 198695
rect 191542 178625 191594 178631
rect 191542 178567 191594 178573
rect 191554 88943 191582 178567
rect 191638 112395 191690 112401
rect 191638 112337 191690 112343
rect 191542 88937 191594 88943
rect 191542 88879 191594 88885
rect 191650 77473 191678 112337
rect 191638 77467 191690 77473
rect 191638 77409 191690 77415
rect 193652 66258 193708 66267
rect 193652 66193 193708 66202
rect 193666 66077 193694 66193
rect 193654 66071 193706 66077
rect 193654 66013 193706 66019
rect 194338 48465 194366 227629
rect 197206 227613 197258 227619
rect 197206 227555 197258 227561
rect 196054 221471 196106 221477
rect 196054 221413 196106 221419
rect 196066 219447 196094 221413
rect 196052 219438 196108 219447
rect 196052 219373 196108 219382
rect 194422 184397 194474 184403
rect 194422 184339 194474 184345
rect 194434 90095 194462 184339
rect 194518 118167 194570 118173
rect 194518 118109 194570 118115
rect 194420 90086 194476 90095
rect 194420 90021 194476 90030
rect 194530 78699 194558 118109
rect 194710 100777 194762 100783
rect 194710 100719 194762 100725
rect 194722 98679 194750 100719
rect 194708 98670 194764 98679
rect 194708 98605 194764 98614
rect 195478 94857 195530 94863
rect 195478 94799 195530 94805
rect 194806 94635 194858 94641
rect 194806 94577 194858 94583
rect 194818 92315 194846 94577
rect 195490 93795 195518 94799
rect 195476 93786 195532 93795
rect 195476 93721 195532 93730
rect 194804 92306 194860 92315
rect 194804 92241 194860 92250
rect 196054 86421 196106 86427
rect 196054 86363 196106 86369
rect 196066 83583 196094 86363
rect 196052 83574 196108 83583
rect 196052 83509 196108 83518
rect 194516 78690 194572 78699
rect 194516 78625 194572 78634
rect 196918 77763 196970 77769
rect 196918 77705 196970 77711
rect 196930 75295 196958 77705
rect 196916 75286 196972 75295
rect 196916 75221 196972 75230
rect 195476 68922 195532 68931
rect 195476 68857 195532 68866
rect 196246 68883 196298 68889
rect 195490 68815 195518 68857
rect 196246 68825 196298 68831
rect 195478 68809 195530 68815
rect 195478 68751 195530 68757
rect 196258 68339 196286 68825
rect 196244 68330 196300 68339
rect 196244 68265 196300 68274
rect 195476 63446 195532 63455
rect 195476 63381 195478 63390
rect 195530 63381 195532 63390
rect 195478 63349 195530 63355
rect 195476 60782 195532 60791
rect 195476 60717 195532 60726
rect 195490 60675 195518 60717
rect 195478 60669 195530 60675
rect 195478 60611 195530 60617
rect 194326 48459 194378 48465
rect 194326 48401 194378 48407
rect 197218 48391 197246 227555
rect 200086 224727 200138 224733
rect 200086 224669 200138 224675
rect 199702 224653 199754 224659
rect 199702 224595 199754 224601
rect 199714 224035 199742 224595
rect 199700 224026 199756 224035
rect 199700 223961 199756 223970
rect 198838 221767 198890 221773
rect 198838 221709 198890 221715
rect 198850 221223 198878 221709
rect 198836 221214 198892 221223
rect 198836 221149 198892 221158
rect 197302 187283 197354 187289
rect 197302 187225 197354 187231
rect 197314 90687 197342 187225
rect 197398 124013 197450 124019
rect 197398 123955 197450 123961
rect 197300 90678 197356 90687
rect 197300 90613 197356 90622
rect 197410 79291 197438 123955
rect 198358 100555 198410 100561
rect 198358 100497 198410 100503
rect 198370 100455 198398 100497
rect 198356 100446 198412 100455
rect 198356 100381 198412 100390
rect 197878 89233 197930 89239
rect 197878 89175 197930 89181
rect 197890 86839 197918 89175
rect 197876 86830 197932 86839
rect 197876 86765 197932 86774
rect 198742 86273 198794 86279
rect 198742 86215 198794 86221
rect 197780 85794 197836 85803
rect 197780 85729 197836 85738
rect 197794 85021 197822 85729
rect 197782 85015 197834 85021
rect 197782 84957 197834 84963
rect 198754 84767 198782 86215
rect 198740 84758 198796 84767
rect 198740 84693 198796 84702
rect 197396 79282 197452 79291
rect 197396 79217 197452 79226
rect 198550 66145 198602 66151
rect 198550 66087 198602 66093
rect 198562 65675 198590 66087
rect 198548 65666 198604 65675
rect 198548 65601 198604 65610
rect 198358 60373 198410 60379
rect 198358 60315 198410 60321
rect 198370 59163 198398 60315
rect 198356 59154 198412 59163
rect 198356 59089 198412 59098
rect 197206 48385 197258 48391
rect 197206 48327 197258 48333
rect 200098 47281 200126 224669
rect 201718 224579 201770 224585
rect 201718 224521 201770 224527
rect 201622 224505 201674 224511
rect 201622 224447 201674 224453
rect 201634 222851 201662 224447
rect 201730 223443 201758 224521
rect 201814 224431 201866 224437
rect 201814 224373 201866 224379
rect 201716 223434 201772 223443
rect 201716 223369 201772 223378
rect 201620 222842 201676 222851
rect 201620 222777 201676 222786
rect 201826 221815 201854 224373
rect 201812 221806 201868 221815
rect 201812 221741 201868 221750
rect 201718 221619 201770 221625
rect 201718 221561 201770 221567
rect 201622 221545 201674 221551
rect 201622 221487 201674 221493
rect 201634 219595 201662 221487
rect 201730 220187 201758 221561
rect 201716 220178 201772 220187
rect 201716 220113 201772 220122
rect 201620 219586 201676 219595
rect 201620 219521 201676 219530
rect 200662 218881 200714 218887
rect 200662 218823 200714 218829
rect 200674 218559 200702 218823
rect 201718 218807 201770 218813
rect 201718 218749 201770 218755
rect 201622 218659 201674 218665
rect 201622 218601 201674 218607
rect 200660 218550 200716 218559
rect 200660 218485 200716 218494
rect 201634 216931 201662 218601
rect 201730 217967 201758 218749
rect 201716 217958 201772 217967
rect 201716 217893 201772 217902
rect 201620 216922 201676 216931
rect 201620 216857 201676 216866
rect 201718 215921 201770 215927
rect 201718 215863 201770 215869
rect 201730 215303 201758 215863
rect 201716 215294 201772 215303
rect 201716 215229 201772 215238
rect 200182 155611 200234 155617
rect 200182 155553 200234 155559
rect 200194 91279 200222 155553
rect 200278 123939 200330 123945
rect 200278 123881 200330 123887
rect 200180 91270 200236 91279
rect 200180 91205 200236 91214
rect 200290 80179 200318 123881
rect 201718 100703 201770 100709
rect 201718 100645 201770 100651
rect 201730 99419 201758 100645
rect 201716 99410 201772 99419
rect 201716 99345 201772 99354
rect 200758 97891 200810 97897
rect 200758 97833 200810 97839
rect 200566 97817 200618 97823
rect 200564 97782 200566 97791
rect 200618 97782 200620 97791
rect 200564 97717 200620 97726
rect 200770 96163 200798 97833
rect 201718 97743 201770 97749
rect 201718 97685 201770 97691
rect 201046 97595 201098 97601
rect 201046 97537 201098 97543
rect 201058 97199 201086 97537
rect 201044 97190 201100 97199
rect 201044 97125 201100 97134
rect 200756 96154 200812 96163
rect 200756 96089 200812 96098
rect 201730 95571 201758 97685
rect 201716 95562 201772 95571
rect 201716 95497 201772 95506
rect 201622 94931 201674 94937
rect 201622 94873 201674 94879
rect 201634 92907 201662 94873
rect 201718 94783 201770 94789
rect 201718 94725 201770 94731
rect 201730 94535 201758 94725
rect 201716 94526 201772 94535
rect 201716 94461 201772 94470
rect 201620 92898 201676 92907
rect 201620 92833 201676 92842
rect 201718 91823 201770 91829
rect 201718 91765 201770 91771
rect 201730 89651 201758 91765
rect 201716 89642 201772 89651
rect 201716 89577 201772 89586
rect 201814 89159 201866 89165
rect 201814 89101 201866 89107
rect 201622 89085 201674 89091
rect 201622 89027 201674 89033
rect 201716 89050 201772 89059
rect 201334 89011 201386 89017
rect 201334 88953 201386 88959
rect 201346 88467 201374 88953
rect 201332 88458 201388 88467
rect 201332 88393 201388 88402
rect 201634 88023 201662 89027
rect 201716 88985 201772 88994
rect 201730 88943 201758 88985
rect 201718 88937 201770 88943
rect 201718 88879 201770 88885
rect 201620 88014 201676 88023
rect 201620 87949 201676 87958
rect 201826 87431 201854 89101
rect 201812 87422 201868 87431
rect 201812 87357 201868 87366
rect 201620 86386 201676 86395
rect 201620 86321 201676 86330
rect 201814 86347 201866 86353
rect 201634 86131 201662 86321
rect 201814 86289 201866 86295
rect 201718 86199 201770 86205
rect 201718 86141 201770 86147
rect 201622 86125 201674 86131
rect 201622 86067 201674 86073
rect 201730 85211 201758 86141
rect 201716 85202 201772 85211
rect 201716 85137 201772 85146
rect 201826 84175 201854 86289
rect 201812 84166 201868 84175
rect 201812 84101 201868 84110
rect 201526 83535 201578 83541
rect 201526 83477 201578 83483
rect 201538 80919 201566 83477
rect 201814 83461 201866 83467
rect 201814 83403 201866 83409
rect 201622 83387 201674 83393
rect 201622 83329 201674 83335
rect 201634 82547 201662 83329
rect 201718 83313 201770 83319
rect 201718 83255 201770 83261
rect 201730 83139 201758 83255
rect 201716 83130 201772 83139
rect 201716 83065 201772 83074
rect 201620 82538 201676 82547
rect 201620 82473 201676 82482
rect 201718 82129 201770 82135
rect 201718 82071 201770 82077
rect 201730 81955 201758 82071
rect 201716 81946 201772 81955
rect 201716 81881 201772 81890
rect 201826 81511 201854 83403
rect 201812 81502 201868 81511
rect 201812 81437 201868 81446
rect 201524 80910 201580 80919
rect 201524 80845 201580 80854
rect 200276 80170 200332 80179
rect 200276 80105 200332 80114
rect 201622 77689 201674 77695
rect 201622 77631 201674 77637
rect 201716 77654 201772 77663
rect 200278 77615 200330 77621
rect 200278 77557 200330 77563
rect 200290 76035 200318 77557
rect 200276 76026 200332 76035
rect 200276 75961 200332 75970
rect 201634 75443 201662 77631
rect 201716 77589 201772 77598
rect 201730 77473 201758 77589
rect 201718 77467 201770 77473
rect 201718 77409 201770 77415
rect 201718 77245 201770 77251
rect 201718 77187 201770 77193
rect 201730 77071 201758 77187
rect 201716 77062 201772 77071
rect 201716 76997 201772 77006
rect 201620 75434 201676 75443
rect 201620 75369 201676 75378
rect 201526 74877 201578 74883
rect 201526 74819 201578 74825
rect 201538 72187 201566 74819
rect 201814 74803 201866 74809
rect 201814 74745 201866 74751
rect 201622 74655 201674 74661
rect 201622 74597 201674 74603
rect 201634 73815 201662 74597
rect 201718 74581 201770 74587
rect 201718 74523 201770 74529
rect 201730 74407 201758 74523
rect 201716 74398 201772 74407
rect 201716 74333 201772 74342
rect 201620 73806 201676 73815
rect 201620 73741 201676 73750
rect 201826 72779 201854 74745
rect 201812 72770 201868 72779
rect 201812 72705 201868 72714
rect 201524 72178 201580 72187
rect 201524 72113 201580 72122
rect 200374 71991 200426 71997
rect 200374 71933 200426 71939
rect 200386 69967 200414 71933
rect 201814 71917 201866 71923
rect 201814 71859 201866 71865
rect 201622 71843 201674 71849
rect 201622 71785 201674 71791
rect 201634 70559 201662 71785
rect 201718 71769 201770 71775
rect 201718 71711 201770 71717
rect 201730 71151 201758 71711
rect 201716 71142 201772 71151
rect 201716 71077 201772 71086
rect 201620 70550 201676 70559
rect 201620 70485 201676 70494
rect 200372 69958 200428 69967
rect 200372 69893 200428 69902
rect 201826 69523 201854 71859
rect 201812 69514 201868 69523
rect 201812 69449 201868 69458
rect 201814 69105 201866 69111
rect 201814 69047 201866 69053
rect 201622 69031 201674 69037
rect 201622 68973 201674 68979
rect 201634 67303 201662 68973
rect 201718 68957 201770 68963
rect 201718 68899 201770 68905
rect 201730 67895 201758 68899
rect 201716 67886 201772 67895
rect 201716 67821 201772 67830
rect 201620 67294 201676 67303
rect 201620 67229 201676 67238
rect 201826 66711 201854 69047
rect 201812 66702 201868 66711
rect 201812 66637 201868 66646
rect 201718 66219 201770 66225
rect 201718 66161 201770 66167
rect 201730 65083 201758 66161
rect 201716 65074 201772 65083
rect 201716 65009 201772 65018
rect 201718 64887 201770 64893
rect 201718 64829 201770 64835
rect 201730 64639 201758 64829
rect 201814 64813 201866 64819
rect 201814 64755 201866 64761
rect 201716 64630 201772 64639
rect 201716 64565 201772 64574
rect 201826 64047 201854 64755
rect 201812 64038 201868 64047
rect 201812 63973 201868 63982
rect 201716 63002 201772 63011
rect 201716 62937 201772 62946
rect 201620 62410 201676 62419
rect 201620 62345 201676 62354
rect 201524 61818 201580 61827
rect 201524 61753 201580 61762
rect 201538 60601 201566 61753
rect 201634 60749 201662 62345
rect 201730 60823 201758 62937
rect 201812 61374 201868 61383
rect 201812 61309 201868 61318
rect 201718 60817 201770 60823
rect 201718 60759 201770 60765
rect 201622 60743 201674 60749
rect 201622 60685 201674 60691
rect 201526 60595 201578 60601
rect 201526 60537 201578 60543
rect 201826 60527 201854 61309
rect 201814 60521 201866 60527
rect 201814 60463 201866 60469
rect 201716 60190 201772 60199
rect 201716 60125 201772 60134
rect 201730 59047 201758 60125
rect 201718 59041 201770 59047
rect 201718 58983 201770 58989
rect 202978 48359 203006 230441
rect 204514 227735 204542 244131
rect 204598 243449 204650 243455
rect 204598 243391 204650 243397
rect 204610 228327 204638 243391
rect 204706 232175 204734 246499
rect 204790 246483 204842 246489
rect 204790 246425 204842 246431
rect 204692 232166 204748 232175
rect 204692 232101 204748 232110
rect 204802 231583 204830 246425
rect 204788 231574 204844 231583
rect 204788 231509 204844 231518
rect 204898 230991 204926 246573
rect 204982 244559 205034 244565
rect 204982 244501 205034 244507
rect 204884 230982 204940 230991
rect 204884 230917 204940 230926
rect 204596 228318 204652 228327
rect 204596 228253 204652 228262
rect 204500 227726 204556 227735
rect 204500 227661 204556 227670
rect 204898 227175 204926 230917
rect 204886 227169 204938 227175
rect 204886 227111 204938 227117
rect 204994 225071 205022 244501
rect 205090 232767 205118 246721
rect 205666 244584 205694 249237
rect 205846 246113 205898 246119
rect 205846 246055 205898 246061
rect 205858 245971 205886 246055
rect 205846 245965 205898 245971
rect 205846 245907 205898 245913
rect 205474 244556 205694 244584
rect 205366 244411 205418 244417
rect 205366 244353 205418 244359
rect 205174 244337 205226 244343
rect 205174 244279 205226 244285
rect 205076 232758 205132 232767
rect 205076 232693 205132 232702
rect 205090 232651 205118 232693
rect 205078 232645 205130 232651
rect 205078 232587 205130 232593
rect 205078 232497 205130 232503
rect 205078 232439 205130 232445
rect 204980 225062 205036 225071
rect 204980 224997 205036 225006
rect 205090 224900 205118 232439
rect 205186 226699 205214 244279
rect 205172 226690 205228 226699
rect 205172 226625 205228 226634
rect 205378 226107 205406 244353
rect 205474 230547 205502 244556
rect 205558 244485 205610 244491
rect 205558 244427 205610 244433
rect 205460 230538 205516 230547
rect 205460 230473 205516 230482
rect 205364 226098 205420 226107
rect 205364 226033 205420 226042
rect 205570 225663 205598 244427
rect 205654 244263 205706 244269
rect 205654 244205 205706 244211
rect 205666 227291 205694 244205
rect 206326 244115 206378 244121
rect 206326 244057 206378 244063
rect 205750 243967 205802 243973
rect 205750 243909 205802 243915
rect 205652 227282 205708 227291
rect 205652 227217 205708 227226
rect 205654 227169 205706 227175
rect 205654 227111 205706 227117
rect 205556 225654 205612 225663
rect 205556 225589 205612 225598
rect 204898 224872 205118 224900
rect 203062 207411 203114 207417
rect 203062 207353 203114 207359
rect 203074 93943 203102 207353
rect 203158 126825 203210 126831
rect 203158 126767 203210 126773
rect 203060 93934 203116 93943
rect 203060 93869 203116 93878
rect 203170 80327 203198 126767
rect 204598 103663 204650 103669
rect 204598 103605 204650 103611
rect 204502 103515 204554 103521
rect 204502 103457 204554 103463
rect 204514 101047 204542 103457
rect 204610 102083 204638 103605
rect 204694 103589 204746 103595
rect 204694 103531 204746 103537
rect 204596 102074 204652 102083
rect 204596 102009 204652 102018
rect 204706 101639 204734 103531
rect 204692 101630 204748 101639
rect 204692 101565 204748 101574
rect 204500 101038 204556 101047
rect 204500 100973 204556 100982
rect 204598 100629 204650 100635
rect 204598 100571 204650 100577
rect 204610 98827 204638 100571
rect 204596 98818 204652 98827
rect 204596 98753 204652 98762
rect 203156 80318 203212 80327
rect 203156 80253 203212 80262
rect 204898 53275 204926 224872
rect 205666 54015 205694 227111
rect 205762 223179 205790 243909
rect 206134 243893 206186 243899
rect 206134 243835 206186 243841
rect 205942 243745 205994 243751
rect 205942 243687 205994 243693
rect 205846 241969 205898 241975
rect 205846 241911 205898 241917
rect 205750 223173 205802 223179
rect 205750 223115 205802 223121
rect 205858 222976 205886 241911
rect 205762 222948 205886 222976
rect 205762 202723 205790 222948
rect 205954 214563 205982 243687
rect 206038 243375 206090 243381
rect 206038 243317 206090 243323
rect 206050 229363 206078 243317
rect 206036 229354 206092 229363
rect 206036 229289 206092 229298
rect 206146 223420 206174 243835
rect 206230 243819 206282 243825
rect 206230 243761 206282 243767
rect 206050 223392 206174 223420
rect 206242 223420 206270 243761
rect 206338 230579 206366 244057
rect 206518 244041 206570 244047
rect 206518 243983 206570 243989
rect 206422 243671 206474 243677
rect 206422 243613 206474 243619
rect 206326 230573 206378 230579
rect 206326 230515 206378 230521
rect 206242 223392 206366 223420
rect 205940 214554 205996 214563
rect 205940 214489 205996 214498
rect 206050 213559 206078 223392
rect 206134 223173 206186 223179
rect 206134 223115 206186 223121
rect 206038 213553 206090 213559
rect 206038 213495 206090 213501
rect 206146 212787 206174 223115
rect 206338 213675 206366 223392
rect 206434 214711 206462 243613
rect 206530 233243 206558 243983
rect 206626 243423 206654 271289
rect 210370 271131 210398 271807
rect 210358 271125 210410 271131
rect 210358 271067 210410 271073
rect 210454 271125 210506 271131
rect 210454 271067 210506 271073
rect 210466 270761 210494 271067
rect 210658 270835 210686 271936
rect 210646 270829 210698 270835
rect 210646 270771 210698 270777
rect 210454 270755 210506 270761
rect 210454 270697 210506 270703
rect 210946 268467 210974 277870
rect 212208 277856 212510 277884
rect 212374 273567 212426 273573
rect 212374 273509 212426 273515
rect 211894 271421 211946 271427
rect 211894 271363 211946 271369
rect 211798 271273 211850 271279
rect 211700 271238 211756 271247
rect 211798 271215 211850 271221
rect 211700 271173 211756 271182
rect 211508 268722 211564 268731
rect 211508 268657 211564 268666
rect 210934 268461 210986 268467
rect 210934 268403 210986 268409
rect 211124 268130 211180 268139
rect 211124 268065 211180 268074
rect 211028 267834 211084 267843
rect 211028 267769 211084 267778
rect 210646 264909 210698 264915
rect 210646 264851 210698 264857
rect 207188 261322 207244 261331
rect 207188 261257 207244 261266
rect 206996 249334 207052 249343
rect 206996 249269 207052 249278
rect 206902 249147 206954 249153
rect 206902 249089 206954 249095
rect 206806 244633 206858 244639
rect 206806 244575 206858 244581
rect 206710 243597 206762 243603
rect 206710 243539 206762 243545
rect 206612 243414 206668 243423
rect 206612 243349 206668 243358
rect 206518 233237 206570 233243
rect 206518 233179 206570 233185
rect 206614 233237 206666 233243
rect 206614 233179 206666 233185
rect 206420 214702 206476 214711
rect 206420 214637 206476 214646
rect 206324 213666 206380 213675
rect 206324 213601 206380 213610
rect 206326 213553 206378 213559
rect 206326 213495 206378 213501
rect 206338 213083 206366 213495
rect 206324 213074 206380 213083
rect 206324 213009 206380 213018
rect 206132 212778 206188 212787
rect 206132 212713 206188 212722
rect 206626 212047 206654 233179
rect 206722 216339 206750 243539
rect 206818 224479 206846 244575
rect 206914 230727 206942 249089
rect 207010 243696 207038 249269
rect 207202 243899 207230 261257
rect 209398 247667 209450 247673
rect 209398 247609 209450 247615
rect 207190 243893 207242 243899
rect 207242 243853 207408 243881
rect 207190 243835 207242 243841
rect 207010 243668 207134 243696
rect 206998 243523 207050 243529
rect 206998 243465 207050 243471
rect 206902 230721 206954 230727
rect 206902 230663 206954 230669
rect 206902 230573 206954 230579
rect 206902 230515 206954 230521
rect 206804 224470 206860 224479
rect 206804 224405 206860 224414
rect 206708 216330 206764 216339
rect 206708 216265 206764 216274
rect 206612 212038 206668 212047
rect 206612 211973 206668 211982
rect 206914 211455 206942 230515
rect 207010 222407 207038 243465
rect 207106 237831 207134 243668
rect 207094 237825 207146 237831
rect 207094 237767 207146 237773
rect 207094 230721 207146 230727
rect 207094 230663 207146 230669
rect 207106 229807 207134 230663
rect 207092 229798 207148 229807
rect 207092 229733 207148 229742
rect 206996 222398 207052 222407
rect 206996 222333 207052 222342
rect 207106 222236 207134 229733
rect 207010 222208 207134 222236
rect 206900 211446 206956 211455
rect 206900 211381 206956 211390
rect 207010 202996 207038 222208
rect 206914 202968 207038 202996
rect 205748 202714 205804 202723
rect 205748 202649 205804 202658
rect 206914 192987 206942 202968
rect 206902 192981 206954 192987
rect 206902 192923 206954 192929
rect 206998 192981 207050 192987
rect 206998 192923 207050 192929
rect 207010 169899 207038 192923
rect 206710 169893 206762 169899
rect 206710 169835 206762 169841
rect 206998 169893 207050 169899
rect 206998 169835 207050 169841
rect 206722 142612 206750 169835
rect 206722 142584 207038 142612
rect 207010 126628 207038 142584
rect 207010 126600 207134 126628
rect 207106 120985 207134 126600
rect 207094 120979 207146 120985
rect 207094 120921 207146 120927
rect 207190 120979 207242 120985
rect 207190 120921 207242 120927
rect 207202 97939 207230 120921
rect 207188 97930 207244 97939
rect 207188 97865 207244 97874
rect 206996 57526 207052 57535
rect 206996 57461 207052 57470
rect 206900 55898 206956 55907
rect 206900 55833 206956 55842
rect 205654 54009 205706 54015
rect 205654 53951 205706 53957
rect 204886 53269 204938 53275
rect 204886 53211 204938 53217
rect 203062 52381 203114 52387
rect 203062 52323 203114 52329
rect 203074 52017 203102 52323
rect 203062 52011 203114 52017
rect 203062 51953 203114 51959
rect 202964 48350 203020 48359
rect 202964 48285 203020 48294
rect 200086 47275 200138 47281
rect 200086 47217 200138 47223
rect 191446 46239 191498 46245
rect 191446 46181 191498 46187
rect 145641 45696 206410 45724
rect 206382 42051 206410 45696
rect 206914 42323 206942 55833
rect 207010 46097 207038 57461
rect 206998 46091 207050 46097
rect 206998 46033 207050 46039
rect 206902 42317 206954 42323
rect 206902 42259 206954 42265
rect 207380 42051 207408 243853
rect 209410 239131 209438 247609
rect 209876 247114 209932 247123
rect 209876 247049 209932 247058
rect 209780 246374 209836 246383
rect 209686 246335 209738 246341
rect 209780 246309 209836 246318
rect 209686 246277 209738 246283
rect 209590 246261 209642 246267
rect 209590 246203 209642 246209
rect 209602 245157 209630 246203
rect 209590 245151 209642 245157
rect 209590 245093 209642 245099
rect 209698 244935 209726 246277
rect 209686 244929 209738 244935
rect 209686 244871 209738 244877
rect 209794 243127 209822 246309
rect 209890 246267 209918 247049
rect 209972 246818 210028 246827
rect 209972 246753 210028 246762
rect 210260 246818 210316 246827
rect 210260 246753 210316 246762
rect 209986 246341 210014 246753
rect 210166 246409 210218 246415
rect 210166 246351 210218 246357
rect 209974 246335 210026 246341
rect 209974 246277 210026 246283
rect 209878 246261 209930 246267
rect 209878 246203 209930 246209
rect 209972 245634 210028 245643
rect 209972 245569 210028 245578
rect 209986 243719 210014 245569
rect 210178 245231 210206 246351
rect 210166 245225 210218 245231
rect 210274 245199 210302 246753
rect 210550 245595 210602 245601
rect 210550 245537 210602 245543
rect 210562 245495 210590 245537
rect 210548 245486 210604 245495
rect 210548 245421 210604 245430
rect 210166 245167 210218 245173
rect 210260 245190 210316 245199
rect 210260 245125 210316 245134
rect 210068 245042 210124 245051
rect 210068 244977 210070 244986
rect 210122 244977 210124 244986
rect 210070 244945 210122 244951
rect 210068 244894 210124 244903
rect 210068 244829 210070 244838
rect 210122 244829 210124 244838
rect 210070 244797 210122 244803
rect 209972 243710 210028 243719
rect 209972 243645 210028 243654
rect 210658 243275 210686 264851
rect 210742 249221 210794 249227
rect 210742 249163 210794 249169
rect 210644 243266 210700 243275
rect 210644 243201 210700 243210
rect 209780 243118 209836 243127
rect 209780 243053 209836 243062
rect 209396 239122 209452 239131
rect 209396 239057 209452 239066
rect 209410 238072 209438 239057
rect 209410 238044 209918 238072
rect 209588 237642 209644 237651
rect 209588 237577 209644 237586
rect 208150 233681 208202 233687
rect 208150 233623 208202 233629
rect 207956 232166 208012 232175
rect 207956 232101 208012 232110
rect 207970 53645 207998 232101
rect 208052 97930 208108 97939
rect 208052 97865 208108 97874
rect 207958 53639 208010 53645
rect 207958 53581 208010 53587
rect 208066 53127 208094 97865
rect 208054 53121 208106 53127
rect 208054 53063 208106 53069
rect 208054 50605 208106 50611
rect 208054 50547 208106 50553
rect 208066 50019 208094 50547
rect 208054 50013 208106 50019
rect 208054 49955 208106 49961
rect 208162 48835 208190 233623
rect 209300 231574 209356 231583
rect 209300 231509 209356 231518
rect 209204 202714 209260 202723
rect 209204 202649 209260 202658
rect 208726 144067 208778 144073
rect 208726 144009 208778 144015
rect 208630 129637 208682 129643
rect 208630 129579 208682 129585
rect 208534 126751 208586 126757
rect 208534 126693 208586 126699
rect 208438 103737 208490 103743
rect 208438 103679 208490 103685
rect 208342 97965 208394 97971
rect 208342 97907 208394 97913
rect 208246 77837 208298 77843
rect 208246 77779 208298 77785
rect 208258 50611 208286 77779
rect 208354 53941 208382 97907
rect 208342 53935 208394 53941
rect 208342 53877 208394 53883
rect 208246 50605 208298 50611
rect 208246 50547 208298 50553
rect 208450 50537 208478 103679
rect 208342 50531 208394 50537
rect 208342 50473 208394 50479
rect 208438 50531 208490 50537
rect 208438 50473 208490 50479
rect 208354 49797 208382 50473
rect 208342 49791 208394 49797
rect 208342 49733 208394 49739
rect 208150 48829 208202 48835
rect 208150 48771 208202 48777
rect 208546 48761 208574 126693
rect 208534 48755 208586 48761
rect 208534 48697 208586 48703
rect 208642 48169 208670 129579
rect 208534 48163 208586 48169
rect 208534 48105 208586 48111
rect 208630 48163 208682 48169
rect 208630 48105 208682 48111
rect 208546 46319 208574 48105
rect 208738 46393 208766 144009
rect 208822 141181 208874 141187
rect 208822 141123 208874 141129
rect 208834 46467 208862 141123
rect 208918 135409 208970 135415
rect 208918 135351 208970 135357
rect 208930 48983 208958 135351
rect 209014 132597 209066 132603
rect 209014 132539 209066 132545
rect 208918 48977 208970 48983
rect 208918 48919 208970 48925
rect 209026 48687 209054 132539
rect 209110 132523 209162 132529
rect 209110 132465 209162 132471
rect 209122 50556 209150 132465
rect 209218 50704 209246 202649
rect 209314 54311 209342 231509
rect 209492 230538 209548 230547
rect 209492 230473 209548 230482
rect 209506 62863 209534 230473
rect 209492 62854 209548 62863
rect 209398 62815 209450 62821
rect 209492 62789 209548 62798
rect 209398 62757 209450 62763
rect 209302 54305 209354 54311
rect 209302 54247 209354 54253
rect 209410 53571 209438 62757
rect 209494 62667 209546 62673
rect 209494 62609 209546 62615
rect 209398 53565 209450 53571
rect 209398 53507 209450 53513
rect 209506 53497 209534 62609
rect 209494 53491 209546 53497
rect 209494 53433 209546 53439
rect 209602 51647 209630 237577
rect 209684 236754 209740 236763
rect 209684 236689 209740 236698
rect 209698 54163 209726 236689
rect 209782 233755 209834 233761
rect 209782 233697 209834 233703
rect 209794 71997 209822 233697
rect 209782 71991 209834 71997
rect 209782 71933 209834 71939
rect 209782 71843 209834 71849
rect 209782 71785 209834 71791
rect 209794 54237 209822 71785
rect 209782 54231 209834 54237
rect 209782 54173 209834 54179
rect 209686 54157 209738 54163
rect 209686 54099 209738 54105
rect 209890 51721 209918 238044
rect 210754 236203 210782 249163
rect 211042 247747 211070 267769
rect 211030 247741 211082 247747
rect 211030 247683 211082 247689
rect 210934 246705 210986 246711
rect 210934 246647 210986 246653
rect 210838 245817 210890 245823
rect 210836 245782 210838 245791
rect 210890 245782 210892 245791
rect 210836 245717 210892 245726
rect 210358 236197 210410 236203
rect 210358 236139 210410 236145
rect 210742 236197 210794 236203
rect 210742 236139 210794 236145
rect 210164 234830 210220 234839
rect 210164 234765 210220 234774
rect 210066 233811 210126 233820
rect 210066 233742 210126 233751
rect 209974 233607 210026 233613
rect 209974 233549 210026 233555
rect 209986 71849 210014 233549
rect 209974 71843 210026 71849
rect 209974 71785 210026 71791
rect 209974 71695 210026 71701
rect 209972 71660 209974 71669
rect 210026 71660 210028 71669
rect 209972 71595 210028 71604
rect 209974 60447 210026 60453
rect 209974 60389 210026 60395
rect 209986 59681 210014 60389
rect 209972 59672 210028 59681
rect 209972 59607 210028 59616
rect 209972 56416 210028 56425
rect 209972 56351 210028 56360
rect 209986 53793 210014 56351
rect 209974 53787 210026 53793
rect 209974 53729 210026 53735
rect 209878 51715 209930 51721
rect 209878 51657 209930 51663
rect 209590 51641 209642 51647
rect 209590 51583 209642 51589
rect 209218 50676 209438 50704
rect 209122 50528 209342 50556
rect 209110 50383 209162 50389
rect 209110 50325 209162 50331
rect 209122 50093 209150 50325
rect 209110 50087 209162 50093
rect 209110 50029 209162 50035
rect 209014 48681 209066 48687
rect 209014 48623 209066 48629
rect 209314 48243 209342 50528
rect 209410 50389 209438 50676
rect 209398 50383 209450 50389
rect 209398 50325 209450 50331
rect 210082 48909 210110 233742
rect 210178 228919 210206 234765
rect 210262 233533 210314 233539
rect 210262 233475 210314 233481
rect 210164 228910 210220 228919
rect 210164 228845 210220 228854
rect 210166 221693 210218 221699
rect 210166 221635 210218 221641
rect 210178 220705 210206 221635
rect 210164 220696 210220 220705
rect 210164 220631 210220 220640
rect 210166 218733 210218 218739
rect 210166 218675 210218 218681
rect 210178 217449 210206 218675
rect 210164 217440 210220 217449
rect 210164 217375 210220 217384
rect 210166 215995 210218 216001
rect 210166 215937 210218 215943
rect 210178 215821 210206 215937
rect 210164 215812 210220 215821
rect 210164 215747 210220 215756
rect 210164 205082 210220 205091
rect 210164 205017 210220 205026
rect 210178 164243 210206 205017
rect 210164 164234 210220 164243
rect 210164 164169 210220 164178
rect 210164 125162 210220 125171
rect 210164 125097 210220 125106
rect 210178 121323 210206 125097
rect 210164 121314 210220 121323
rect 210164 121249 210220 121258
rect 210166 100481 210218 100487
rect 210166 100423 210218 100429
rect 210178 99937 210206 100423
rect 210164 99928 210220 99937
rect 210164 99863 210220 99872
rect 210166 97669 210218 97675
rect 210166 97611 210218 97617
rect 210178 96681 210206 97611
rect 210164 96672 210220 96681
rect 210164 96607 210220 96616
rect 210164 95044 210220 95053
rect 210164 94979 210220 94988
rect 210178 94715 210206 94979
rect 210166 94709 210218 94715
rect 210166 94651 210218 94657
rect 210166 92119 210218 92125
rect 210166 92061 210218 92067
rect 210178 91797 210206 92061
rect 210164 91788 210220 91797
rect 210164 91723 210220 91732
rect 210166 80353 210218 80359
rect 210166 80295 210218 80301
rect 210178 78181 210206 80295
rect 210164 78172 210220 78181
rect 210164 78107 210220 78116
rect 210166 77541 210218 77547
rect 210166 77483 210218 77489
rect 210178 76553 210206 77483
rect 210164 76544 210220 76553
rect 210164 76479 210220 76488
rect 210166 74729 210218 74735
rect 210166 74671 210218 74677
rect 210178 73297 210206 74671
rect 210164 73288 210220 73297
rect 210164 73223 210220 73232
rect 210166 71991 210218 71997
rect 210166 71933 210218 71939
rect 210178 62567 210206 71933
rect 210274 62821 210302 233475
rect 210262 62815 210314 62821
rect 210262 62757 210314 62763
rect 210370 62692 210398 236139
rect 210946 233539 210974 246647
rect 211028 246522 211084 246531
rect 211028 246457 211084 246466
rect 211042 243719 211070 246457
rect 211028 243710 211084 243719
rect 211028 243645 211084 243654
rect 211138 241943 211166 268065
rect 211522 267843 211550 268657
rect 211508 267834 211564 267843
rect 211508 267769 211564 267778
rect 211510 267573 211562 267579
rect 211510 267515 211562 267521
rect 211222 264983 211274 264989
rect 211222 264925 211274 264931
rect 211124 241934 211180 241943
rect 211124 241869 211180 241878
rect 211234 238835 211262 264925
rect 211318 247741 211370 247747
rect 211318 247683 211370 247689
rect 211330 238983 211358 247683
rect 211522 243719 211550 267515
rect 211604 247114 211660 247123
rect 211604 247049 211660 247058
rect 211618 246679 211646 247049
rect 211604 246670 211660 246679
rect 211604 246605 211660 246614
rect 211714 246489 211742 271173
rect 211810 246859 211838 271215
rect 211798 246853 211850 246859
rect 211798 246795 211850 246801
rect 211906 246711 211934 271363
rect 212084 271090 212140 271099
rect 212084 271025 212140 271034
rect 212098 257756 212126 271025
rect 212182 270829 212234 270835
rect 212182 270771 212234 270777
rect 212194 257904 212222 270771
rect 212278 267869 212330 267875
rect 212278 267811 212330 267817
rect 212290 264989 212318 267811
rect 212386 265142 212414 273509
rect 212482 265803 212510 277856
rect 213346 272907 213374 277870
rect 214594 274239 214622 277870
rect 215746 276755 215774 277870
rect 215734 276749 215786 276755
rect 215734 276691 215786 276697
rect 214582 274233 214634 274239
rect 214582 274175 214634 274181
rect 213238 272901 213290 272907
rect 213238 272843 213290 272849
rect 213334 272901 213386 272907
rect 213334 272843 213386 272849
rect 216694 272901 216746 272907
rect 216694 272843 216746 272849
rect 212470 265797 212522 265803
rect 212470 265739 212522 265745
rect 213250 265142 213278 272843
rect 216118 272309 216170 272315
rect 216118 272251 216170 272257
rect 215446 271865 215498 271871
rect 215446 271807 215498 271813
rect 214486 270755 214538 270761
rect 214486 270697 214538 270703
rect 213814 270681 213866 270687
rect 213814 270623 213866 270629
rect 213826 265156 213854 270623
rect 213826 265128 214080 265156
rect 214498 265142 214526 270697
rect 214966 266611 215018 266617
rect 214966 266553 215018 266559
rect 214978 265142 215006 266553
rect 215458 265142 215486 271807
rect 215542 271125 215594 271131
rect 215542 271067 215594 271073
rect 215554 265156 215582 271067
rect 216130 265156 216158 272251
rect 215554 265128 215808 265156
rect 216130 265128 216288 265156
rect 216706 265142 216734 272843
rect 216898 265156 216926 277870
rect 217364 273162 217420 273171
rect 217364 273097 217420 273106
rect 217378 272431 217406 273097
rect 217558 272901 217610 272907
rect 217558 272843 217610 272849
rect 217460 272570 217516 272579
rect 217460 272505 217516 272514
rect 217364 272422 217420 272431
rect 217364 272357 217420 272366
rect 217474 270803 217502 272505
rect 217460 270794 217516 270803
rect 217460 270729 217516 270738
rect 216898 265128 217200 265156
rect 217570 265142 217598 272843
rect 218050 268245 218078 277870
rect 219312 277856 219614 277884
rect 218230 272309 218282 272315
rect 218230 272251 218282 272257
rect 218038 268239 218090 268245
rect 218038 268181 218090 268187
rect 218242 265156 218270 272251
rect 219286 271199 219338 271205
rect 219286 271141 219338 271147
rect 218902 271125 218954 271131
rect 218902 271067 218954 271073
rect 218710 270903 218762 270909
rect 218710 270845 218762 270851
rect 218722 265156 218750 270845
rect 218016 265128 218270 265156
rect 218496 265128 218750 265156
rect 218914 265142 218942 271067
rect 219298 265142 219326 271141
rect 219586 267727 219614 277856
rect 220450 272907 220478 277870
rect 220438 272901 220490 272907
rect 220438 272843 220490 272849
rect 221014 272901 221066 272907
rect 221014 272843 221066 272849
rect 220822 271865 220874 271871
rect 220822 271807 220874 271813
rect 220342 271421 220394 271427
rect 220342 271363 220394 271369
rect 219766 271347 219818 271353
rect 219766 271289 219818 271295
rect 219574 267721 219626 267727
rect 219574 267663 219626 267669
rect 219778 265142 219806 271289
rect 220354 265156 220382 271363
rect 220834 265156 220862 271807
rect 220224 265128 220382 265156
rect 220608 265128 220862 265156
rect 221026 265142 221054 272843
rect 221494 269275 221546 269281
rect 221494 269217 221546 269223
rect 221506 265142 221534 269217
rect 221698 265285 221726 277870
rect 223030 274825 223082 274831
rect 223030 274767 223082 274773
rect 221780 271682 221836 271691
rect 221780 271617 221836 271626
rect 221794 271247 221822 271617
rect 221780 271238 221836 271247
rect 221780 271173 221836 271182
rect 221974 270533 222026 270539
rect 221974 270475 222026 270481
rect 221782 267795 221834 267801
rect 221782 267737 221834 267743
rect 221794 267653 221822 267737
rect 221782 267647 221834 267653
rect 221782 267589 221834 267595
rect 221686 265279 221738 265285
rect 221686 265221 221738 265227
rect 221986 265142 222014 270475
rect 222550 268313 222602 268319
rect 222550 268255 222602 268261
rect 222562 265156 222590 268255
rect 223042 265156 223070 274767
rect 224002 272315 224030 277870
rect 225250 277051 225278 277870
rect 225238 277045 225290 277051
rect 225238 276987 225290 276993
rect 226294 274677 226346 274683
rect 226294 274619 226346 274625
rect 225430 274159 225482 274165
rect 225430 274101 225482 274107
rect 225238 274085 225290 274091
rect 225238 274027 225290 274033
rect 224086 273493 224138 273499
rect 224086 273435 224138 273441
rect 223990 272309 224042 272315
rect 223990 272251 224042 272257
rect 223702 272013 223754 272019
rect 223702 271955 223754 271961
rect 223222 268165 223274 268171
rect 223222 268107 223274 268113
rect 222336 265128 222590 265156
rect 222816 265128 223070 265156
rect 223234 265142 223262 268107
rect 223714 265142 223742 271955
rect 224098 265142 224126 273435
rect 224566 272309 224618 272315
rect 224566 272251 224618 272257
rect 224578 265156 224606 272251
rect 225250 265156 225278 274027
rect 224544 265128 224606 265156
rect 225024 265128 225278 265156
rect 225442 265142 225470 274101
rect 225814 268757 225866 268763
rect 225814 268699 225866 268705
rect 225826 265142 225854 268699
rect 226306 265142 226334 274619
rect 226402 265951 226430 277870
rect 227446 275861 227498 275867
rect 227446 275803 227498 275809
rect 226966 269867 227018 269873
rect 226966 269809 227018 269815
rect 226390 265945 226442 265951
rect 226390 265887 226442 265893
rect 226978 265156 227006 269809
rect 227458 265156 227486 275803
rect 227542 273567 227594 273573
rect 227542 273509 227594 273515
rect 227554 272759 227582 273509
rect 227542 272753 227594 272759
rect 227542 272695 227594 272701
rect 227650 270909 227678 277870
rect 228022 275195 228074 275201
rect 228022 275137 228074 275143
rect 227638 270903 227690 270909
rect 227638 270845 227690 270851
rect 227542 269497 227594 269503
rect 227542 269439 227594 269445
rect 226752 265128 227006 265156
rect 227232 265128 227486 265156
rect 227554 265142 227582 269439
rect 228034 265142 228062 275137
rect 228502 269349 228554 269355
rect 228502 269291 228554 269297
rect 228514 265142 228542 269291
rect 228802 268393 228830 277870
rect 229078 275047 229130 275053
rect 229078 274989 229130 274995
rect 228790 268387 228842 268393
rect 228790 268329 228842 268335
rect 229090 265156 229118 274989
rect 229750 273789 229802 273795
rect 229750 273731 229802 273737
rect 229558 268905 229610 268911
rect 229558 268847 229610 268853
rect 229570 265156 229598 268847
rect 228864 265128 229118 265156
rect 229344 265128 229598 265156
rect 229762 265142 229790 273731
rect 230050 266247 230078 277870
rect 230614 273863 230666 273869
rect 230614 273805 230666 273811
rect 230230 268979 230282 268985
rect 230230 268921 230282 268927
rect 230038 266241 230090 266247
rect 230038 266183 230090 266189
rect 230242 265142 230270 268921
rect 230626 265142 230654 273805
rect 231202 271131 231230 277870
rect 231958 276379 232010 276385
rect 231958 276321 232010 276327
rect 231766 273715 231818 273721
rect 231766 273657 231818 273663
rect 231190 271125 231242 271131
rect 231190 271067 231242 271073
rect 231286 270607 231338 270613
rect 231286 270549 231338 270555
rect 231298 265156 231326 270549
rect 231778 265156 231806 273657
rect 231072 265128 231326 265156
rect 231552 265128 231806 265156
rect 231970 265142 231998 276321
rect 232342 276305 232394 276311
rect 232342 276247 232394 276253
rect 232354 265142 232382 276247
rect 232450 273943 232478 277870
rect 233506 277125 233534 277870
rect 233494 277119 233546 277125
rect 233494 277061 233546 277067
rect 233494 276009 233546 276015
rect 233494 275951 233546 275957
rect 232438 273937 232490 273943
rect 232438 273879 232490 273885
rect 232822 270311 232874 270317
rect 232822 270253 232874 270259
rect 232834 265142 232862 270253
rect 233506 265156 233534 275951
rect 234070 275713 234122 275719
rect 234070 275655 234122 275661
rect 233974 270237 234026 270243
rect 233974 270179 234026 270185
rect 233986 265156 234014 270179
rect 233280 265128 233534 265156
rect 233760 265128 234014 265156
rect 234082 265142 234110 275655
rect 234658 271205 234686 277870
rect 235030 275417 235082 275423
rect 235030 275359 235082 275365
rect 234646 271199 234698 271205
rect 234646 271141 234698 271147
rect 234550 270089 234602 270095
rect 234550 270031 234602 270037
rect 234562 265142 234590 270031
rect 235042 265142 235070 275359
rect 235702 269719 235754 269725
rect 235702 269661 235754 269667
rect 235714 265156 235742 269661
rect 235906 268097 235934 277870
rect 237168 277856 237470 277884
rect 235990 275343 236042 275349
rect 235990 275285 236042 275291
rect 235894 268091 235946 268097
rect 235894 268033 235946 268039
rect 236002 265156 236030 275285
rect 236758 275121 236810 275127
rect 236758 275063 236810 275069
rect 236278 273641 236330 273647
rect 236278 273583 236330 273589
rect 236182 271865 236234 271871
rect 236290 271853 236318 273583
rect 236234 271825 236318 271853
rect 236182 271807 236234 271813
rect 236278 269571 236330 269577
rect 236278 269513 236330 269519
rect 235488 265128 235742 265156
rect 235872 265128 236030 265156
rect 236290 265142 236318 269513
rect 236770 265142 236798 275063
rect 237142 268535 237194 268541
rect 237142 268477 237194 268483
rect 237154 265142 237182 268477
rect 237442 266543 237470 277856
rect 237814 274381 237866 274387
rect 237814 274323 237866 274329
rect 237430 266537 237482 266543
rect 237430 266479 237482 266485
rect 237826 265156 237854 274323
rect 238306 271353 238334 277870
rect 239350 274529 239402 274535
rect 239350 274471 239402 274477
rect 238486 274455 238538 274461
rect 238486 274397 238538 274403
rect 238294 271347 238346 271353
rect 238294 271289 238346 271295
rect 238294 268609 238346 268615
rect 238294 268551 238346 268557
rect 238306 265156 238334 268551
rect 237600 265128 237854 265156
rect 238080 265128 238334 265156
rect 238498 265142 238526 274397
rect 238870 268683 238922 268689
rect 238870 268625 238922 268631
rect 238882 265142 238910 268625
rect 239362 265142 239390 274471
rect 239458 274017 239486 277870
rect 240706 277273 240734 277870
rect 240694 277267 240746 277273
rect 240694 277209 240746 277215
rect 240502 274603 240554 274609
rect 240502 274545 240554 274551
rect 239446 274011 239498 274017
rect 239446 273953 239498 273959
rect 240022 268831 240074 268837
rect 240022 268773 240074 268779
rect 240034 265156 240062 268773
rect 240514 265156 240542 274545
rect 241556 271534 241612 271543
rect 241556 271469 241612 271478
rect 241570 271353 241598 271469
rect 241858 271427 241886 277870
rect 242998 274899 243050 274905
rect 242998 274841 243050 274847
rect 242230 274751 242282 274757
rect 242230 274693 242282 274699
rect 242036 271534 242092 271543
rect 242036 271469 242092 271478
rect 241846 271421 241898 271427
rect 241652 271386 241708 271395
rect 241558 271347 241610 271353
rect 241846 271363 241898 271369
rect 241940 271386 241996 271395
rect 241708 271330 241940 271335
rect 242050 271353 242078 271469
rect 241652 271321 241996 271330
rect 242038 271347 242090 271353
rect 241666 271307 241982 271321
rect 241558 271289 241610 271295
rect 242038 271289 242090 271295
rect 241846 270977 241898 270983
rect 241846 270919 241898 270925
rect 241942 270977 241994 270983
rect 241942 270919 241994 270925
rect 241858 270817 241886 270919
rect 241954 270817 241982 270919
rect 241858 270789 241982 270817
rect 241558 269127 241610 269133
rect 241558 269069 241610 269075
rect 240886 269053 240938 269059
rect 240886 268995 240938 269001
rect 240898 265156 240926 268995
rect 241078 267869 241130 267875
rect 241078 267811 241130 267817
rect 239808 265128 240062 265156
rect 240288 265128 240542 265156
rect 240672 265128 240926 265156
rect 241090 265142 241118 267811
rect 241570 265142 241598 269069
rect 241846 267573 241898 267579
rect 241846 267515 241898 267521
rect 241858 267431 241886 267515
rect 241846 267425 241898 267431
rect 241846 267367 241898 267373
rect 242242 265156 242270 274693
rect 242614 269201 242666 269207
rect 242614 269143 242666 269149
rect 242626 265156 242654 269143
rect 243010 265156 243038 274841
rect 243106 267949 243134 277870
rect 243766 276453 243818 276459
rect 243766 276395 243818 276401
rect 243286 270681 243338 270687
rect 243286 270623 243338 270629
rect 243094 267943 243146 267949
rect 243094 267885 243146 267891
rect 242016 265128 242270 265156
rect 242400 265128 242654 265156
rect 242880 265128 243038 265156
rect 243298 265142 243326 270623
rect 243778 265142 243806 276395
rect 244258 266617 244286 277870
rect 244726 276231 244778 276237
rect 244726 276173 244778 276179
rect 244246 266611 244298 266617
rect 244246 266553 244298 266559
rect 244150 266463 244202 266469
rect 244150 266405 244202 266411
rect 244162 265142 244190 266405
rect 244738 265156 244766 276173
rect 245398 276157 245450 276163
rect 245398 276099 245450 276105
rect 245302 270385 245354 270391
rect 245302 270327 245354 270333
rect 245314 265156 245342 270327
rect 244608 265128 244766 265156
rect 245088 265128 245342 265156
rect 245410 265142 245438 276099
rect 245506 273647 245534 277870
rect 246358 276083 246410 276089
rect 246358 276025 246410 276031
rect 245494 273641 245546 273647
rect 245494 273583 245546 273589
rect 246164 271682 246220 271691
rect 246164 271617 246220 271626
rect 246178 271247 246206 271617
rect 246164 271238 246220 271247
rect 246164 271173 246220 271182
rect 245878 270163 245930 270169
rect 245878 270105 245930 270111
rect 245890 265142 245918 270105
rect 246370 265142 246398 276025
rect 246658 271427 246686 277870
rect 247906 277421 247934 277870
rect 247894 277415 247946 277421
rect 247894 277357 247946 277363
rect 247414 275935 247466 275941
rect 247414 275877 247466 275883
rect 246646 271421 246698 271427
rect 246646 271363 246698 271369
rect 247030 269941 247082 269947
rect 247030 269883 247082 269889
rect 247042 265156 247070 269883
rect 247426 265156 247454 275877
rect 248086 275787 248138 275793
rect 248086 275729 248138 275735
rect 247606 273567 247658 273573
rect 247606 273509 247658 273515
rect 247618 272759 247646 273509
rect 247606 272753 247658 272759
rect 247606 272695 247658 272701
rect 247606 269793 247658 269799
rect 247606 269735 247658 269741
rect 246816 265128 247070 265156
rect 247200 265128 247454 265156
rect 247618 265142 247646 269735
rect 248098 265142 248126 275729
rect 249058 272907 249086 277870
rect 249142 275639 249194 275645
rect 249142 275581 249194 275587
rect 249046 272901 249098 272907
rect 249046 272843 249098 272849
rect 248566 269645 248618 269651
rect 248566 269587 248618 269593
rect 248578 265142 248606 269587
rect 249154 265156 249182 275581
rect 249814 275565 249866 275571
rect 249814 275507 249866 275513
rect 249622 269423 249674 269429
rect 249622 269365 249674 269371
rect 249634 265156 249662 269365
rect 248928 265128 249182 265156
rect 249408 265128 249662 265156
rect 249826 265142 249854 275507
rect 250210 271871 250238 277870
rect 251376 277856 251678 277884
rect 250676 274198 250732 274207
rect 250676 274133 250732 274142
rect 250198 271865 250250 271871
rect 250198 271807 250250 271813
rect 250292 268574 250348 268583
rect 250292 268509 250348 268518
rect 250306 265142 250334 268509
rect 250690 265142 250718 274133
rect 251254 270755 251306 270761
rect 251254 270697 251306 270703
rect 251266 269281 251294 270697
rect 251254 269275 251306 269281
rect 251254 269217 251306 269223
rect 251350 269275 251402 269281
rect 251350 269217 251402 269223
rect 251362 265156 251390 269217
rect 251650 266913 251678 277856
rect 252226 277856 252528 277884
rect 251828 274346 251884 274355
rect 251828 274281 251884 274290
rect 251638 266907 251690 266913
rect 251638 266849 251690 266855
rect 251842 265156 251870 274281
rect 252226 270761 252254 277856
rect 252404 274494 252460 274503
rect 252404 274429 252460 274438
rect 252214 270755 252266 270761
rect 252214 270697 252266 270703
rect 252020 268870 252076 268879
rect 252020 268805 252076 268814
rect 251926 267795 251978 267801
rect 251926 267737 251978 267743
rect 251938 267653 251966 267737
rect 251926 267647 251978 267653
rect 251926 267589 251978 267595
rect 251136 265128 251390 265156
rect 251616 265128 251870 265156
rect 252034 265142 252062 268805
rect 252418 265142 252446 274429
rect 253762 271353 253790 277870
rect 254914 276829 254942 277870
rect 254902 276823 254954 276829
rect 254902 276765 254954 276771
rect 254132 274790 254188 274799
rect 254132 274725 254188 274734
rect 253940 274642 253996 274651
rect 253940 274577 253996 274586
rect 253750 271347 253802 271353
rect 253750 271289 253802 271295
rect 253364 270498 253420 270507
rect 253364 270433 253420 270442
rect 252884 269018 252940 269027
rect 252884 268953 252940 268962
rect 252898 265142 252926 268953
rect 253378 265156 253406 270433
rect 253954 265156 253982 274577
rect 253344 265128 253406 265156
rect 253728 265128 253982 265156
rect 254146 265142 254174 274725
rect 256162 270539 256190 277870
rect 256820 273902 256876 273911
rect 256820 273837 256876 273846
rect 256150 270533 256202 270539
rect 256150 270475 256202 270481
rect 254612 267982 254668 267991
rect 254612 267917 254668 267926
rect 254626 265142 254654 267917
rect 256150 267499 256202 267505
rect 256150 267441 256202 267447
rect 255094 266093 255146 266099
rect 255094 266035 255146 266041
rect 255106 265142 255134 266035
rect 256162 265156 256190 267441
rect 255456 265137 255710 265156
rect 255456 265131 255722 265137
rect 255456 265128 255670 265131
rect 255936 265128 256190 265156
rect 256834 265142 256862 273837
rect 257314 270835 257342 277870
rect 258562 274979 258590 277870
rect 258550 274973 258602 274979
rect 258550 274915 258602 274921
rect 259604 273162 259660 273171
rect 259604 273097 259660 273106
rect 258358 272901 258410 272907
rect 258358 272843 258410 272849
rect 257686 271421 257738 271427
rect 257686 271363 257738 271369
rect 257698 270983 257726 271363
rect 257686 270977 257738 270983
rect 257686 270919 257738 270925
rect 257302 270829 257354 270835
rect 257302 270771 257354 270777
rect 257396 268722 257452 268731
rect 257396 268657 257452 268666
rect 257300 268130 257356 268139
rect 257300 268065 257356 268074
rect 257314 265156 257342 268065
rect 257232 265128 257342 265156
rect 257410 265156 257438 268657
rect 258370 265156 258398 272843
rect 259318 271791 259370 271797
rect 259318 271733 259370 271739
rect 259330 271099 259358 271733
rect 259316 271090 259372 271099
rect 259316 271025 259372 271034
rect 258932 268426 258988 268435
rect 258932 268361 258988 268370
rect 258550 267869 258602 267875
rect 258550 267811 258602 267817
rect 257410 265128 257664 265156
rect 258144 265128 258398 265156
rect 258562 265142 258590 267811
rect 258646 267795 258698 267801
rect 258646 267737 258698 267743
rect 258658 266099 258686 267737
rect 258646 266093 258698 266099
rect 258646 266035 258698 266041
rect 258946 265142 258974 268361
rect 259618 265156 259646 273097
rect 259714 268319 259742 277870
rect 260962 271131 260990 277870
rect 261620 275678 261676 275687
rect 261620 275613 261676 275622
rect 260950 271125 261002 271131
rect 260950 271067 261002 271073
rect 260660 270794 260716 270803
rect 260660 270729 260716 270738
rect 260564 269166 260620 269175
rect 260564 269101 260620 269110
rect 259702 268313 259754 268319
rect 259702 268255 259754 268261
rect 260086 268313 260138 268319
rect 260086 268255 260138 268261
rect 260098 265156 260126 268255
rect 260578 265156 260606 269101
rect 259440 265128 259646 265156
rect 259872 265128 260126 265156
rect 260352 265128 260606 265156
rect 260674 265142 260702 270729
rect 261332 268574 261388 268583
rect 261332 268509 261388 268518
rect 261346 268287 261374 268509
rect 261140 268278 261196 268287
rect 261140 268213 261196 268222
rect 261332 268278 261388 268287
rect 261332 268213 261388 268222
rect 261154 265142 261182 268213
rect 261634 265142 261662 275613
rect 262006 268017 262058 268023
rect 261922 267977 262006 268005
rect 261814 267647 261866 267653
rect 261814 267589 261866 267595
rect 261826 267431 261854 267589
rect 261814 267425 261866 267431
rect 261814 267367 261866 267373
rect 261922 266469 261950 267977
rect 262006 267959 262058 267965
rect 262004 267834 262060 267843
rect 262004 267769 262060 267778
rect 261910 266463 261962 266469
rect 261910 266405 261962 266411
rect 262018 265156 262046 267769
rect 262114 267135 262142 277870
rect 262868 274938 262924 274947
rect 262868 274873 262924 274882
rect 262678 273641 262730 273647
rect 262678 273583 262730 273589
rect 262390 273567 262442 273573
rect 262390 273509 262442 273515
rect 262402 272019 262430 273509
rect 262390 272013 262442 272019
rect 262390 271955 262442 271961
rect 262196 271682 262252 271691
rect 262196 271617 262252 271626
rect 262210 271279 262238 271617
rect 262198 271273 262250 271279
rect 262198 271215 262250 271221
rect 262102 267129 262154 267135
rect 262102 267071 262154 267077
rect 261984 265128 262046 265156
rect 262102 265205 262154 265211
rect 262690 265156 262718 273583
rect 262102 265147 262154 265153
rect 255670 265073 255722 265079
rect 262114 265063 262142 265147
rect 262464 265128 262718 265156
rect 262882 265142 262910 274873
rect 263362 274831 263390 277870
rect 263350 274825 263402 274831
rect 263350 274767 263402 274773
rect 263348 274050 263404 274059
rect 263348 273985 263404 273994
rect 263362 265142 263390 273985
rect 263746 265142 263774 278425
rect 293782 278377 293834 278383
rect 293782 278319 293834 278325
rect 292054 278303 292106 278309
rect 292054 278245 292106 278251
rect 290806 278007 290858 278013
rect 290806 277949 290858 277955
rect 264404 275530 264460 275539
rect 264404 275465 264460 275474
rect 264418 265156 264446 275465
rect 264514 271353 264542 277870
rect 265940 275382 265996 275391
rect 265940 275317 265996 275326
rect 264502 271347 264554 271353
rect 264502 271289 264554 271295
rect 265460 271238 265516 271247
rect 265460 271173 265516 271182
rect 264884 269758 264940 269767
rect 264884 269693 264940 269702
rect 264898 265156 264926 269693
rect 265076 268722 265132 268731
rect 265076 268657 265132 268666
rect 264192 265128 264446 265156
rect 264672 265128 264926 265156
rect 265090 265142 265118 268657
rect 265474 265142 265502 271173
rect 265954 265142 265982 275317
rect 266612 269610 266668 269619
rect 266612 269545 266668 269554
rect 266626 265156 266654 269545
rect 266818 268171 266846 277870
rect 267092 275234 267148 275243
rect 267092 275169 267148 275178
rect 266806 268165 266858 268171
rect 266806 268107 266858 268113
rect 267106 265156 267134 275169
rect 267188 275086 267244 275095
rect 267188 275021 267244 275030
rect 266400 265128 266654 265156
rect 266880 265128 267134 265156
rect 267202 265142 267230 275021
rect 268066 272019 268094 277870
rect 269218 274831 269246 277870
rect 269206 274825 269258 274831
rect 269206 274767 269258 274773
rect 270370 273573 270398 277870
rect 270742 275491 270794 275497
rect 270742 275433 270794 275439
rect 270550 275269 270602 275275
rect 270550 275211 270602 275217
rect 270358 273567 270410 273573
rect 270358 273509 270410 273515
rect 270454 273567 270506 273573
rect 270454 273509 270506 273515
rect 268054 272013 268106 272019
rect 268054 271955 268106 271961
rect 270466 271205 270494 273509
rect 269398 271199 269450 271205
rect 269398 271141 269450 271147
rect 270454 271199 270506 271205
rect 270454 271141 270506 271147
rect 268726 270755 268778 270761
rect 268726 270697 268778 270703
rect 267668 269462 267724 269471
rect 267668 269397 267724 269406
rect 267382 268165 267434 268171
rect 267382 268107 267434 268113
rect 267394 267843 267422 268107
rect 267380 267834 267436 267843
rect 267380 267769 267436 267778
rect 267478 267795 267530 267801
rect 267478 267737 267530 267743
rect 267490 267653 267518 267737
rect 267478 267647 267530 267653
rect 267478 267589 267530 267595
rect 267682 265142 267710 269397
rect 268148 269314 268204 269323
rect 268148 269249 268204 269258
rect 268054 268165 268106 268171
rect 268054 268107 268106 268113
rect 268066 267843 268094 268107
rect 267764 267834 267820 267843
rect 267764 267769 267820 267778
rect 268052 267834 268108 267843
rect 268052 267769 268108 267778
rect 267778 267653 267806 267769
rect 267766 267647 267818 267653
rect 267766 267589 267818 267595
rect 268162 265142 268190 269249
rect 268244 267834 268300 267843
rect 268244 267769 268300 267778
rect 267574 265131 267626 265137
rect 267574 265073 267626 265079
rect 262102 265057 262154 265063
rect 256368 264989 256670 265008
rect 262102 264999 262154 265005
rect 212278 264983 212330 264989
rect 256368 264983 256682 264989
rect 256368 264980 256630 264983
rect 212278 264925 212330 264931
rect 267586 264931 267614 265073
rect 268258 264989 268286 267769
rect 268738 265156 268766 270697
rect 269204 269906 269260 269915
rect 269204 269841 269260 269850
rect 269014 267499 269066 267505
rect 269014 267441 269066 267447
rect 269026 265507 269054 267441
rect 269014 265501 269066 265507
rect 269014 265443 269066 265449
rect 269218 265156 269246 269841
rect 269302 267795 269354 267801
rect 269302 267737 269354 267743
rect 269314 267431 269342 267737
rect 269302 267425 269354 267431
rect 269302 267367 269354 267373
rect 268512 265128 268766 265156
rect 268992 265128 269246 265156
rect 269410 265142 269438 271141
rect 269878 271051 269930 271057
rect 269878 270993 269930 270999
rect 269890 265142 269918 270993
rect 270562 265156 270590 275211
rect 270754 265156 270782 275433
rect 271318 274307 271370 274313
rect 271318 274249 271370 274255
rect 271414 274307 271466 274313
rect 271414 274249 271466 274255
rect 270934 270459 270986 270465
rect 270934 270401 270986 270407
rect 270288 265128 270590 265156
rect 270720 265128 270782 265156
rect 270946 265156 270974 270401
rect 271330 265156 271358 274249
rect 271426 273573 271454 274249
rect 271618 273573 271646 277870
rect 272470 274233 272522 274239
rect 272470 274175 272522 274181
rect 271414 273567 271466 273573
rect 271414 273509 271466 273515
rect 271606 273567 271658 273573
rect 271606 273509 271658 273515
rect 271990 268461 272042 268467
rect 271990 268403 272042 268409
rect 270946 265128 271200 265156
rect 271330 265128 271632 265156
rect 272002 265142 272030 268403
rect 272482 265142 272510 274175
rect 272770 268467 272798 277870
rect 273622 277045 273674 277051
rect 273622 276987 273674 276993
rect 273526 271791 273578 271797
rect 273526 271733 273578 271739
rect 273538 271099 273566 271733
rect 273524 271090 273580 271099
rect 273524 271025 273580 271034
rect 272758 268461 272810 268467
rect 272758 268403 272810 268409
rect 272662 268239 272714 268245
rect 272662 268181 272714 268187
rect 272674 265156 272702 268181
rect 273142 265279 273194 265285
rect 273142 265221 273194 265227
rect 273154 265156 273182 265221
rect 273634 265156 273662 276987
rect 274018 273499 274046 277870
rect 274678 273937 274730 273943
rect 274678 273879 274730 273885
rect 274006 273493 274058 273499
rect 274006 273435 274058 273441
rect 274198 268387 274250 268393
rect 274198 268329 274250 268335
rect 272674 265128 272928 265156
rect 273154 265128 273408 265156
rect 273634 265128 273792 265156
rect 274210 265142 274238 268329
rect 274690 265142 274718 273879
rect 275170 273499 275198 277870
rect 276418 274313 276446 277870
rect 276406 274307 276458 274313
rect 276406 274249 276458 274255
rect 275254 274011 275306 274017
rect 275254 273953 275306 273959
rect 275158 273493 275210 273499
rect 275158 273435 275210 273441
rect 274870 268091 274922 268097
rect 274870 268033 274922 268039
rect 274882 265156 274910 268033
rect 275266 265156 275294 273953
rect 277570 272315 277598 277870
rect 278818 272315 278846 277870
rect 279478 273567 279530 273573
rect 279478 273509 279530 273515
rect 277558 272309 277610 272315
rect 277558 272251 277610 272257
rect 278806 272309 278858 272315
rect 278806 272251 278858 272257
rect 278998 272013 279050 272019
rect 278998 271955 279050 271961
rect 276790 271865 276842 271871
rect 276790 271807 276842 271813
rect 276214 270977 276266 270983
rect 276214 270919 276266 270925
rect 275734 267943 275786 267949
rect 275734 267885 275786 267891
rect 275746 265156 275774 267885
rect 276226 265156 276254 270919
rect 274882 265128 275136 265156
rect 275266 265128 275520 265156
rect 275746 265128 276000 265156
rect 276226 265128 276432 265156
rect 276802 265142 276830 271807
rect 277270 271421 277322 271427
rect 277270 271363 277322 271369
rect 277282 265142 277310 271363
rect 278518 271347 278570 271353
rect 278518 271289 278570 271295
rect 278134 271125 278186 271131
rect 278134 271067 278186 271073
rect 277462 270829 277514 270835
rect 277462 270771 277514 270777
rect 277474 265156 277502 270771
rect 277844 268722 277900 268731
rect 277844 268657 277900 268666
rect 277654 268239 277706 268245
rect 277654 268181 277706 268187
rect 277666 268139 277694 268181
rect 277858 268139 277886 268657
rect 277652 268130 277708 268139
rect 277652 268065 277708 268074
rect 277844 268130 277900 268139
rect 277844 268065 277900 268074
rect 278146 265156 278174 271067
rect 277474 265128 277728 265156
rect 278146 265128 278208 265156
rect 278530 265142 278558 271289
rect 279010 265142 279038 271955
rect 279490 265142 279518 273509
rect 279670 273493 279722 273499
rect 279670 273435 279722 273441
rect 279682 265156 279710 273435
rect 279970 267579 279998 277870
rect 281122 274091 281150 277870
rect 281110 274085 281162 274091
rect 281110 274027 281162 274033
rect 281206 273493 281258 273499
rect 281206 273435 281258 273441
rect 280054 272309 280106 272315
rect 280054 272251 280106 272257
rect 280726 272309 280778 272315
rect 280726 272251 280778 272257
rect 279958 267573 280010 267579
rect 279958 267515 280010 267521
rect 280066 265156 280094 272251
rect 279682 265128 279936 265156
rect 280066 265128 280320 265156
rect 280738 265142 280766 272251
rect 280820 269166 280876 269175
rect 280820 269101 280876 269110
rect 280834 268731 280862 269101
rect 280820 268722 280876 268731
rect 280820 268657 280876 268666
rect 281218 265142 281246 273435
rect 282370 272315 282398 277870
rect 282358 272309 282410 272315
rect 282358 272251 282410 272257
rect 283414 271865 283466 271871
rect 283414 271807 283466 271813
rect 282164 271682 282220 271691
rect 282164 271617 282220 271626
rect 282178 271279 282206 271617
rect 282934 271347 282986 271353
rect 282934 271289 282986 271295
rect 282166 271273 282218 271279
rect 282166 271215 282218 271221
rect 282742 271199 282794 271205
rect 282742 271141 282794 271147
rect 282166 271125 282218 271131
rect 282166 271067 282218 271073
rect 281686 271051 281738 271057
rect 281686 270993 281738 270999
rect 281698 265142 281726 270993
rect 282178 265156 282206 271067
rect 282260 269018 282316 269027
rect 282260 268953 282316 268962
rect 282274 268245 282302 268953
rect 282262 268239 282314 268245
rect 282262 268181 282314 268187
rect 282048 265128 282206 265156
rect 282262 265205 282314 265211
rect 282754 265156 282782 271141
rect 282262 265147 282314 265153
rect 282274 265063 282302 265147
rect 282528 265128 282782 265156
rect 282946 265142 282974 271289
rect 283426 265142 283454 271807
rect 283522 268245 283550 277870
rect 284674 274165 284702 277870
rect 284950 275269 285002 275275
rect 284950 275211 285002 275217
rect 284662 274159 284714 274165
rect 284662 274101 284714 274107
rect 284470 273567 284522 273573
rect 284470 273509 284522 273515
rect 283798 272013 283850 272019
rect 283798 271955 283850 271961
rect 283510 268239 283562 268245
rect 283510 268181 283562 268187
rect 283810 265142 283838 271955
rect 284482 265156 284510 273509
rect 284962 265156 284990 275211
rect 285826 273499 285854 277870
rect 287074 274239 287102 277870
rect 287254 277859 287306 277865
rect 287254 277801 287306 277807
rect 287062 274233 287114 274239
rect 287062 274175 287114 274181
rect 286774 274159 286826 274165
rect 286774 274101 286826 274107
rect 285814 273493 285866 273499
rect 285814 273435 285866 273441
rect 285526 272309 285578 272315
rect 285526 272251 285578 272257
rect 285046 267943 285098 267949
rect 285046 267885 285098 267891
rect 284256 265128 284510 265156
rect 284736 265128 284990 265156
rect 285058 265142 285086 267885
rect 285538 265142 285566 272251
rect 286006 268091 286058 268097
rect 286006 268033 286058 268039
rect 286018 265142 286046 268033
rect 286786 266044 286814 274101
rect 287062 268387 287114 268393
rect 287062 268329 287114 268335
rect 286498 266016 286814 266044
rect 286498 265156 286526 266016
rect 287074 265156 287102 268329
rect 286464 265128 286526 265156
rect 286848 265128 287102 265156
rect 287266 265142 287294 277801
rect 288020 270054 288076 270063
rect 288020 269989 288076 269998
rect 288034 268435 288062 269989
rect 288226 268763 288254 277870
rect 289270 276897 289322 276903
rect 289270 276839 289322 276845
rect 288406 276527 288458 276533
rect 288406 276469 288458 276475
rect 288214 268757 288266 268763
rect 288214 268699 288266 268705
rect 288308 268722 288364 268731
rect 288308 268657 288364 268666
rect 288322 268435 288350 268657
rect 288020 268426 288076 268435
rect 288020 268361 288076 268370
rect 288308 268426 288364 268435
rect 288308 268361 288364 268370
rect 287540 267834 287596 267843
rect 287540 267769 287596 267778
rect 282262 265057 282314 265063
rect 282262 264999 282314 265005
rect 287554 264989 287582 267769
rect 287734 267647 287786 267653
rect 287734 267589 287786 267595
rect 287746 265142 287774 267589
rect 288418 265156 288446 276469
rect 288500 267834 288556 267843
rect 288500 267769 288556 267778
rect 288514 265507 288542 267769
rect 288790 266759 288842 266765
rect 288790 266701 288842 266707
rect 288502 265501 288554 265507
rect 288502 265443 288554 265449
rect 288802 265156 288830 266701
rect 289282 265156 289310 276839
rect 289474 271057 289502 277870
rect 289942 277785 289994 277791
rect 289942 277727 289994 277733
rect 289462 271051 289514 271057
rect 289462 270993 289514 270999
rect 289462 267277 289514 267283
rect 289462 267219 289514 267225
rect 288240 265128 288446 265156
rect 288576 265128 288830 265156
rect 289056 265128 289310 265156
rect 289474 265142 289502 267219
rect 289954 265142 289982 277727
rect 290626 268763 290654 277870
rect 290818 277273 290846 277949
rect 291478 277711 291530 277717
rect 291478 277653 291530 277659
rect 290806 277267 290858 277273
rect 290806 277209 290858 277215
rect 290806 277045 290858 277051
rect 290806 276987 290858 276993
rect 290614 268757 290666 268763
rect 290614 268699 290666 268705
rect 290326 267425 290378 267431
rect 290326 267367 290378 267373
rect 290338 265142 290366 267367
rect 290818 265156 290846 276987
rect 290902 273567 290954 273573
rect 290902 273509 290954 273515
rect 290914 271131 290942 273509
rect 290902 271125 290954 271131
rect 290902 271067 290954 271073
rect 291490 265156 291518 277653
rect 291874 274683 291902 277870
rect 291862 274677 291914 274683
rect 291862 274619 291914 274625
rect 291860 268722 291916 268731
rect 291860 268657 291916 268666
rect 291874 268139 291902 268657
rect 291860 268130 291916 268139
rect 291860 268065 291916 268074
rect 291670 267351 291722 267357
rect 291670 267293 291722 267299
rect 290784 265128 290846 265156
rect 291264 265128 291518 265156
rect 291682 265142 291710 267293
rect 292066 265142 292094 278245
rect 292246 277415 292298 277421
rect 292246 277357 292298 277363
rect 292258 276607 292286 277357
rect 292246 276601 292298 276607
rect 292246 276543 292298 276549
rect 293026 273573 293054 277870
rect 293206 277563 293258 277569
rect 293206 277505 293258 277511
rect 293014 273567 293066 273573
rect 293014 273509 293066 273515
rect 292534 271199 292586 271205
rect 292534 271141 292586 271147
rect 292150 270533 292202 270539
rect 292150 270475 292202 270481
rect 292162 268319 292190 270475
rect 292150 268313 292202 268319
rect 292150 268255 292202 268261
rect 292546 265142 292574 271141
rect 293218 265156 293246 277505
rect 293590 267203 293642 267209
rect 293590 267145 293642 267151
rect 293602 265156 293630 267145
rect 292992 265128 293246 265156
rect 293376 265128 293630 265156
rect 293794 265142 293822 278319
rect 294288 277856 294590 277884
rect 294262 271051 294314 271057
rect 294262 270993 294314 270999
rect 294274 265142 294302 270993
rect 294562 268171 294590 277856
rect 294742 273567 294794 273573
rect 294742 273509 294794 273515
rect 294550 268165 294602 268171
rect 294550 268107 294602 268113
rect 294754 265142 294782 273509
rect 295426 269873 295454 277870
rect 295414 269867 295466 269873
rect 295414 269809 295466 269815
rect 295318 267055 295370 267061
rect 295318 266997 295370 267003
rect 295330 265156 295358 266997
rect 295810 265156 295838 278541
rect 303380 278342 303436 278351
rect 303380 278277 303436 278286
rect 301846 278229 301898 278235
rect 301846 278171 301898 278177
rect 297526 278081 297578 278087
rect 297526 278023 297578 278029
rect 296470 277637 296522 277643
rect 296470 277579 296522 277585
rect 295990 266981 296042 266987
rect 295990 266923 296042 266929
rect 295104 265128 295358 265156
rect 295584 265128 295838 265156
rect 296002 265142 296030 266923
rect 296482 265142 296510 277579
rect 296674 274091 296702 277870
rect 296662 274085 296714 274091
rect 296662 274027 296714 274033
rect 297142 274085 297194 274091
rect 297142 274027 297194 274033
rect 296854 271939 296906 271945
rect 296854 271881 296906 271887
rect 296950 271939 297002 271945
rect 296950 271881 297002 271887
rect 296866 271853 296894 271881
rect 296962 271853 296990 271881
rect 296866 271825 296990 271853
rect 296662 271791 296714 271797
rect 296662 271733 296714 271739
rect 296674 271668 296702 271733
rect 296674 271640 296798 271668
rect 296866 271649 297086 271668
rect 296770 271099 296798 271640
rect 296854 271643 297098 271649
rect 296906 271640 297046 271643
rect 296854 271585 296906 271591
rect 297046 271585 297098 271591
rect 297154 271131 297182 274027
rect 297142 271125 297194 271131
rect 296756 271090 296812 271099
rect 297142 271067 297194 271073
rect 296756 271025 296812 271034
rect 296660 269166 296716 269175
rect 296660 269101 296716 269110
rect 296674 268319 296702 269101
rect 296662 268313 296714 268319
rect 296662 268255 296714 268261
rect 297142 267425 297194 267431
rect 297142 267367 297194 267373
rect 296854 266833 296906 266839
rect 296854 266775 296906 266781
rect 296866 265142 296894 266775
rect 297154 266765 297182 267367
rect 297142 266759 297194 266765
rect 297142 266701 297194 266707
rect 297538 265156 297566 278023
rect 301558 277933 301610 277939
rect 301296 277881 301558 277884
rect 301296 277875 301610 277881
rect 297826 274683 297854 277870
rect 298198 277415 298250 277421
rect 298198 277357 298250 277363
rect 297814 274677 297866 274683
rect 297814 274619 297866 274625
rect 298006 266759 298058 266765
rect 298006 266701 298058 266707
rect 298018 265156 298046 266701
rect 297312 265128 297566 265156
rect 297792 265128 298046 265156
rect 298210 265142 298238 277357
rect 298978 275867 299006 277870
rect 299062 277267 299114 277273
rect 299062 277209 299114 277215
rect 298966 275861 299018 275867
rect 298966 275803 299018 275809
rect 298582 266685 298634 266691
rect 298582 266627 298634 266633
rect 298594 265142 298622 266627
rect 299074 265142 299102 277209
rect 300130 271353 300158 277870
rect 301296 277856 301598 277875
rect 300214 277193 300266 277199
rect 300214 277135 300266 277141
rect 300118 271347 300170 271353
rect 300118 271289 300170 271295
rect 299734 266463 299786 266469
rect 299734 266405 299786 266411
rect 299746 265156 299774 266405
rect 300226 265156 300254 277135
rect 300790 276971 300842 276977
rect 300790 276913 300842 276919
rect 300310 266389 300362 266395
rect 300310 266331 300362 266337
rect 299520 265128 299774 265156
rect 300000 265128 300254 265156
rect 300322 265142 300350 266331
rect 300802 265142 300830 276913
rect 301270 266315 301322 266321
rect 301270 266257 301322 266263
rect 301282 265142 301310 266257
rect 301858 265156 301886 278171
rect 302530 269503 302558 277870
rect 302806 271125 302858 271131
rect 302806 271067 302858 271073
rect 302518 269497 302570 269503
rect 302518 269439 302570 269445
rect 302326 266167 302378 266173
rect 302326 266109 302378 266115
rect 302338 265156 302366 266109
rect 302818 265156 302846 271067
rect 302998 266093 303050 266099
rect 302998 266035 303050 266041
rect 301632 265128 301886 265156
rect 302112 265128 302366 265156
rect 302544 265128 302846 265156
rect 303010 265142 303038 266035
rect 303394 265142 303422 278277
rect 304532 278194 304588 278203
rect 304532 278129 304588 278138
rect 303682 271871 303710 277870
rect 303670 271865 303722 271871
rect 303670 271807 303722 271813
rect 304054 266019 304106 266025
rect 304054 265961 304106 265967
rect 304066 265156 304094 265961
rect 304546 265156 304574 278129
rect 305204 277898 305260 277907
rect 304930 274091 304958 277870
rect 305204 277833 305260 277842
rect 304918 274085 304970 274091
rect 304918 274027 304970 274033
rect 304918 270533 304970 270539
rect 304918 270475 304970 270481
rect 304930 270211 304958 270475
rect 304916 270202 304972 270211
rect 304916 270137 304972 270146
rect 304726 265871 304778 265877
rect 304726 265813 304778 265819
rect 303840 265128 304094 265156
rect 304320 265128 304574 265156
rect 304738 265142 304766 265813
rect 305218 265156 305246 277833
rect 306082 275201 306110 277870
rect 307124 277750 307180 277759
rect 307124 277685 307180 277694
rect 306070 275195 306122 275201
rect 306070 275137 306122 275143
rect 306262 271273 306314 271279
rect 306262 271215 306314 271221
rect 305590 265723 305642 265729
rect 305590 265665 305642 265671
rect 305136 265128 305246 265156
rect 305602 265142 305630 265665
rect 306274 265156 306302 271215
rect 306742 265649 306794 265655
rect 306742 265591 306794 265597
rect 306754 265156 306782 265591
rect 307138 265156 307166 277685
rect 307330 272019 307358 277870
rect 308372 277602 308428 277611
rect 308372 277537 308428 277546
rect 307990 277489 308042 277495
rect 307990 277431 308042 277437
rect 308002 276607 308030 277431
rect 307990 276601 308042 276607
rect 307990 276543 308042 276549
rect 307318 272013 307370 272019
rect 307318 271955 307370 271961
rect 307798 270459 307850 270465
rect 307798 270401 307850 270407
rect 307318 265575 307370 265581
rect 307318 265517 307370 265523
rect 306048 265128 306302 265156
rect 306528 265128 306782 265156
rect 306912 265128 307166 265156
rect 307330 265142 307358 265517
rect 307810 265142 307838 270401
rect 308084 270054 308140 270063
rect 308084 269989 308140 269998
rect 308098 268435 308126 269989
rect 308084 268426 308140 268435
rect 308084 268361 308140 268370
rect 308386 265156 308414 277537
rect 308482 272019 308510 277870
rect 308854 273937 308906 273943
rect 308854 273879 308906 273885
rect 308470 272013 308522 272019
rect 308470 271955 308522 271961
rect 308866 265156 308894 273879
rect 309058 273573 309086 278541
rect 317108 278046 317164 278055
rect 309430 278007 309482 278013
rect 309430 277949 309482 277955
rect 311830 278007 311882 278013
rect 311830 277949 311882 277955
rect 316930 278004 317108 278032
rect 309442 277019 309470 277949
rect 309524 277454 309580 277463
rect 309524 277389 309580 277398
rect 309428 277010 309484 277019
rect 309428 276945 309484 276954
rect 309046 273567 309098 273573
rect 309046 273509 309098 273515
rect 309430 267129 309482 267135
rect 309430 267071 309482 267077
rect 309334 265501 309386 265507
rect 309334 265443 309386 265449
rect 309346 265156 309374 265443
rect 308256 265128 308414 265156
rect 308640 265128 308894 265156
rect 309120 265128 309374 265156
rect 309442 265063 309470 267071
rect 309538 265142 309566 277389
rect 309620 276862 309676 276871
rect 309620 276797 309676 276806
rect 309634 276681 309662 276797
rect 309622 276675 309674 276681
rect 309622 276617 309674 276623
rect 309730 269355 309758 277870
rect 310882 273499 310910 277870
rect 310964 277306 311020 277315
rect 310964 277241 311020 277250
rect 310870 273493 310922 273499
rect 310870 273435 310922 273441
rect 310390 269867 310442 269873
rect 310390 269809 310442 269815
rect 309718 269349 309770 269355
rect 309718 269291 309770 269297
rect 309622 267869 309674 267875
rect 309622 267811 309674 267817
rect 309634 267135 309662 267811
rect 309622 267129 309674 267135
rect 309622 267071 309674 267077
rect 309910 265427 309962 265433
rect 309910 265369 309962 265375
rect 309922 265142 309950 265369
rect 310402 265142 310430 269809
rect 310978 265156 311006 277241
rect 311842 276755 311870 277949
rect 311926 277933 311978 277939
rect 312406 277933 312458 277939
rect 311926 277875 311978 277881
rect 312144 277881 312406 277884
rect 312144 277875 312458 277881
rect 311938 276755 311966 277875
rect 312144 277856 312446 277875
rect 312404 277158 312460 277167
rect 312404 277093 312460 277102
rect 311830 276749 311882 276755
rect 311830 276691 311882 276697
rect 311926 276749 311978 276755
rect 311926 276691 311978 276697
rect 311542 275861 311594 275867
rect 311542 275803 311594 275809
rect 311554 265156 311582 275803
rect 312116 267834 312172 267843
rect 312022 267795 312074 267801
rect 312116 267769 312118 267778
rect 312022 267737 312074 267743
rect 312170 267769 312172 267778
rect 312118 267737 312170 267743
rect 311638 265353 311690 265359
rect 311638 265295 311690 265301
rect 310848 265128 311006 265156
rect 311328 265128 311582 265156
rect 311650 265142 311678 265295
rect 312034 265211 312062 267737
rect 312022 265205 312074 265211
rect 312418 265156 312446 277093
rect 313282 275053 313310 277870
rect 314434 275275 314462 277870
rect 315092 276566 315148 276575
rect 315092 276501 315148 276510
rect 314422 275269 314474 275275
rect 314422 275211 314474 275217
rect 313270 275047 313322 275053
rect 313270 274989 313322 274995
rect 313654 271865 313706 271871
rect 313654 271807 313706 271813
rect 312598 269497 312650 269503
rect 312598 269439 312650 269445
rect 312022 265147 312074 265153
rect 312144 265128 312446 265156
rect 312610 265142 312638 269439
rect 312694 268313 312746 268319
rect 312694 268255 312746 268261
rect 312706 268139 312734 268255
rect 312692 268130 312748 268139
rect 312692 268065 312748 268074
rect 313270 265279 313322 265285
rect 313270 265221 313322 265227
rect 313282 265156 313310 265221
rect 313666 265156 313694 271807
rect 314326 271421 314378 271427
rect 314326 271363 314378 271369
rect 313846 269349 313898 269355
rect 313846 269291 313898 269297
rect 313056 265128 313310 265156
rect 313440 265128 313694 265156
rect 313858 265142 313886 269291
rect 314338 265142 314366 271363
rect 315106 270951 315134 276501
rect 315298 271381 315518 271409
rect 315190 271273 315242 271279
rect 315190 271215 315242 271221
rect 315092 270942 315148 270951
rect 315202 270909 315230 271215
rect 315298 271205 315326 271381
rect 315382 271347 315434 271353
rect 315382 271289 315434 271295
rect 315286 271199 315338 271205
rect 315286 271141 315338 271147
rect 315092 270877 315148 270886
rect 315190 270903 315242 270909
rect 315190 270845 315242 270851
rect 314806 270829 314858 270835
rect 314806 270771 314858 270777
rect 314818 265142 314846 270771
rect 315394 265156 315422 271289
rect 315490 271205 315518 271381
rect 315682 271279 315710 277870
rect 316354 277856 316752 277884
rect 316054 275269 316106 275275
rect 316054 275211 316106 275217
rect 315670 271273 315722 271279
rect 315670 271215 315722 271221
rect 315478 271199 315530 271205
rect 315478 271141 315530 271147
rect 315572 270350 315628 270359
rect 315572 270285 315628 270294
rect 315586 268731 315614 270285
rect 315572 268722 315628 268731
rect 315572 268657 315628 268666
rect 315764 268722 315820 268731
rect 315764 268657 315820 268666
rect 315778 265156 315806 268657
rect 315168 265128 315422 265156
rect 315648 265128 315806 265156
rect 316066 265142 316094 275211
rect 316354 268911 316382 277856
rect 316726 271791 316778 271797
rect 316726 271733 316778 271739
rect 316738 271520 316766 271733
rect 316642 271492 316766 271520
rect 316532 271386 316588 271395
rect 316532 271321 316588 271330
rect 316546 270063 316574 271321
rect 316642 271099 316670 271492
rect 316724 271386 316780 271395
rect 316724 271321 316780 271330
rect 316628 271090 316684 271099
rect 316628 271025 316684 271034
rect 316738 270761 316766 271321
rect 316930 270909 316958 278004
rect 317108 277981 317164 277990
rect 317026 277856 318000 277884
rect 316918 270903 316970 270909
rect 316918 270845 316970 270851
rect 316726 270755 316778 270761
rect 316726 270697 316778 270703
rect 316726 270533 316778 270539
rect 316726 270475 316778 270481
rect 316532 270054 316588 270063
rect 316532 269989 316588 269998
rect 316738 269915 316766 270475
rect 316724 269906 316780 269915
rect 316724 269841 316780 269850
rect 317026 269152 317054 277856
rect 318070 277489 318122 277495
rect 318070 277431 318122 277437
rect 318082 276607 318110 277431
rect 318178 276681 318206 278615
rect 370486 278599 370538 278605
rect 370966 278599 371018 278605
rect 370538 278559 370966 278587
rect 370486 278541 370538 278547
rect 373172 278573 373228 278582
rect 373364 278638 373420 278647
rect 379042 278633 379358 278661
rect 379042 278605 379070 278633
rect 373364 278573 373420 278582
rect 379030 278599 379082 278605
rect 370966 278541 371018 278547
rect 373186 278531 373214 278573
rect 334390 278525 334442 278531
rect 334390 278467 334442 278473
rect 338326 278525 338378 278531
rect 338326 278467 338378 278473
rect 358582 278525 358634 278531
rect 358582 278467 358634 278473
rect 373174 278525 373226 278531
rect 373174 278467 373226 278473
rect 329110 278451 329162 278457
rect 329110 278393 329162 278399
rect 325270 278155 325322 278161
rect 325270 278097 325322 278103
rect 326614 278155 326666 278161
rect 326614 278097 326666 278103
rect 319152 277856 319358 277884
rect 318358 277489 318410 277495
rect 318358 277431 318410 277437
rect 318370 277019 318398 277431
rect 318454 277341 318506 277347
rect 318454 277283 318506 277289
rect 318356 277010 318412 277019
rect 318356 276945 318412 276954
rect 318466 276871 318494 277283
rect 318452 276862 318508 276871
rect 318452 276797 318508 276806
rect 318166 276675 318218 276681
rect 318166 276617 318218 276623
rect 318070 276601 318122 276607
rect 318070 276543 318122 276549
rect 318644 276418 318700 276427
rect 318644 276353 318700 276362
rect 317302 275195 317354 275201
rect 317302 275137 317354 275143
rect 317110 270755 317162 270761
rect 317110 270697 317162 270703
rect 317122 270655 317150 270697
rect 317108 270646 317164 270655
rect 317108 270581 317164 270590
rect 317108 270202 317164 270211
rect 317108 270137 317164 270146
rect 316450 269124 317054 269152
rect 316342 268905 316394 268911
rect 316342 268847 316394 268853
rect 316450 268708 316478 269124
rect 316162 268680 316478 268708
rect 316162 267949 316190 268680
rect 316918 268461 316970 268467
rect 316918 268403 316970 268409
rect 316534 268239 316586 268245
rect 316930 268227 316958 268403
rect 317122 268319 317150 270137
rect 317110 268313 317162 268319
rect 317110 268255 317162 268261
rect 316586 268199 316958 268227
rect 316534 268181 316586 268187
rect 316246 268091 316298 268097
rect 316246 268033 316298 268039
rect 317110 268091 317162 268097
rect 317110 268033 317162 268039
rect 316258 267949 316286 268033
rect 316150 267943 316202 267949
rect 316150 267885 316202 267891
rect 316246 267943 316298 267949
rect 316246 267885 316298 267891
rect 317122 267579 317150 268033
rect 317110 267573 317162 267579
rect 317110 267515 317162 267521
rect 317206 267573 317258 267579
rect 317206 267515 317258 267521
rect 317218 267228 317246 267515
rect 316642 267200 317246 267228
rect 316642 265211 316670 267200
rect 317314 265304 317342 275137
rect 318070 275047 318122 275053
rect 318070 274989 318122 274995
rect 317492 270942 317548 270951
rect 317492 270877 317548 270886
rect 317218 265276 317342 265304
rect 316630 265205 316682 265211
rect 316464 265137 316574 265156
rect 317218 265156 317246 265276
rect 317506 265156 317534 270877
rect 317972 270646 318028 270655
rect 317972 270581 318028 270590
rect 317986 270359 318014 270581
rect 317972 270350 318028 270359
rect 317972 270285 318028 270294
rect 317588 269018 317644 269027
rect 317780 269018 317836 269027
rect 317588 268953 317644 268962
rect 317698 268976 317780 269004
rect 317602 268139 317630 268953
rect 317588 268130 317644 268139
rect 317588 268065 317644 268074
rect 317698 265211 317726 268976
rect 317780 268953 317836 268962
rect 317974 268979 318026 268985
rect 317974 268921 318026 268927
rect 317986 268763 318014 268921
rect 317974 268757 318026 268763
rect 317974 268699 318026 268705
rect 317878 267869 317930 267875
rect 317878 267811 317930 267817
rect 317890 267135 317918 267811
rect 317878 267129 317930 267135
rect 317878 267071 317930 267077
rect 316630 265147 316682 265153
rect 316464 265131 316586 265137
rect 316464 265128 316534 265131
rect 316944 265128 317246 265156
rect 317376 265128 317534 265156
rect 317686 265205 317738 265211
rect 318082 265156 318110 274989
rect 318164 270350 318220 270359
rect 318164 270285 318220 270294
rect 317686 265147 317738 265153
rect 317856 265128 318110 265156
rect 318178 265142 318206 270285
rect 318274 270160 318590 270188
rect 318274 268911 318302 270160
rect 318562 270021 318590 270160
rect 318454 270015 318506 270021
rect 318454 269957 318506 269963
rect 318550 270015 318602 270021
rect 318550 269957 318602 269963
rect 318262 268905 318314 268911
rect 318262 268847 318314 268853
rect 318358 268905 318410 268911
rect 318358 268847 318410 268853
rect 318262 268757 318314 268763
rect 318262 268699 318314 268705
rect 318274 268393 318302 268699
rect 318262 268387 318314 268393
rect 318262 268329 318314 268335
rect 318370 268171 318398 268847
rect 318466 268171 318494 269957
rect 318550 268387 318602 268393
rect 318550 268329 318602 268335
rect 318358 268165 318410 268171
rect 318358 268107 318410 268113
rect 318454 268165 318506 268171
rect 318454 268107 318506 268113
rect 318562 267949 318590 268329
rect 318550 267943 318602 267949
rect 318550 267885 318602 267891
rect 318658 267783 318686 276353
rect 319330 271131 319358 277856
rect 320098 277856 320400 277884
rect 319604 276270 319660 276279
rect 319604 276205 319660 276214
rect 319318 271125 319370 271131
rect 319318 271067 319370 271073
rect 319508 271090 319564 271099
rect 319030 271051 319082 271057
rect 319508 271025 319564 271034
rect 319030 270993 319082 270999
rect 319042 270928 319070 270993
rect 319042 270900 319262 270928
rect 318370 267755 318686 267783
rect 318262 267721 318314 267727
rect 318262 267663 318314 267669
rect 318274 267135 318302 267663
rect 318262 267129 318314 267135
rect 318262 267071 318314 267077
rect 318370 266044 318398 267755
rect 319234 267653 319262 270900
rect 319412 270202 319468 270211
rect 319412 270137 319468 270146
rect 318454 267647 318506 267653
rect 318454 267589 318506 267595
rect 319222 267647 319274 267653
rect 319222 267589 319274 267595
rect 318274 266016 318398 266044
rect 316534 265073 316586 265079
rect 309430 265057 309482 265063
rect 309430 264999 309482 265005
rect 318274 265008 318302 266016
rect 318466 265951 318494 267589
rect 318658 266016 319358 266044
rect 318358 265945 318410 265951
rect 318358 265887 318410 265893
rect 318454 265945 318506 265951
rect 318454 265887 318506 265893
rect 318370 265859 318398 265887
rect 318658 265859 318686 266016
rect 318370 265831 318686 265859
rect 318754 265905 319070 265933
rect 318754 265655 318782 265905
rect 318850 265831 318974 265859
rect 318850 265803 318878 265831
rect 318946 265803 318974 265831
rect 318838 265797 318890 265803
rect 318838 265739 318890 265745
rect 318934 265797 318986 265803
rect 318934 265739 318986 265745
rect 319042 265655 319070 265905
rect 318742 265649 318794 265655
rect 318742 265591 318794 265597
rect 319030 265649 319082 265655
rect 319030 265591 319082 265597
rect 318550 265427 318602 265433
rect 319222 265427 319274 265433
rect 318550 265369 318602 265375
rect 318850 265387 319222 265415
rect 318562 265137 318590 265369
rect 318850 265285 318878 265387
rect 319222 265369 319274 265375
rect 318934 265353 318986 265359
rect 318986 265313 319262 265341
rect 318934 265295 318986 265301
rect 318838 265279 318890 265285
rect 318838 265221 318890 265227
rect 318742 265205 318794 265211
rect 318742 265147 318794 265153
rect 318550 265131 318602 265137
rect 318550 265073 318602 265079
rect 268246 264983 268298 264989
rect 256630 264925 256682 264931
rect 267570 264922 267630 264931
rect 268246 264925 268298 264931
rect 287542 264983 287594 264989
rect 318274 264980 318672 265008
rect 318754 264989 318782 265147
rect 319234 265137 319262 265313
rect 319330 265211 319358 266016
rect 319318 265205 319370 265211
rect 319318 265147 319370 265153
rect 318934 265131 318986 265137
rect 318934 265073 318986 265079
rect 319222 265131 319274 265137
rect 319222 265073 319274 265079
rect 318946 264989 318974 265073
rect 319426 265008 319454 270137
rect 319522 270063 319550 271025
rect 319508 270054 319564 270063
rect 319508 269989 319564 269998
rect 319618 265156 319646 276205
rect 319702 273863 319754 273869
rect 319702 273805 319754 273811
rect 319714 273499 319742 273805
rect 320098 273795 320126 277856
rect 321428 277010 321484 277019
rect 321428 276945 321484 276954
rect 320852 276122 320908 276131
rect 320852 276057 320908 276066
rect 320086 273789 320138 273795
rect 320086 273731 320138 273737
rect 319798 273567 319850 273573
rect 319798 273509 319850 273515
rect 319702 273493 319754 273499
rect 319702 273435 319754 273441
rect 319810 272315 319838 273509
rect 319798 272309 319850 272315
rect 319798 272251 319850 272257
rect 320374 272309 320426 272315
rect 320374 272251 320426 272257
rect 319702 270829 319754 270835
rect 319702 270771 319754 270777
rect 319714 270063 319742 270771
rect 319700 270054 319756 270063
rect 319700 269989 319756 269998
rect 320180 269906 320236 269915
rect 320180 269841 320236 269850
rect 319702 265427 319754 265433
rect 319702 265369 319754 265375
rect 319714 265285 319742 265369
rect 319702 265279 319754 265285
rect 319702 265221 319754 265227
rect 320194 265156 320222 269841
rect 319584 265128 319646 265156
rect 319968 265128 320222 265156
rect 320386 265142 320414 272251
rect 320866 265142 320894 276057
rect 321334 267943 321386 267949
rect 321334 267885 321386 267891
rect 321046 265427 321098 265433
rect 321046 265369 321098 265375
rect 318742 264983 318794 264989
rect 287542 264925 287594 264931
rect 318742 264925 318794 264931
rect 318934 264983 318986 264989
rect 319152 264980 319454 265008
rect 321058 264989 321086 265369
rect 321346 265142 321374 267885
rect 321442 265156 321470 276945
rect 321538 273573 321566 277870
rect 322100 276714 322156 276723
rect 322100 276649 322156 276658
rect 321526 273567 321578 273573
rect 321526 273509 321578 273515
rect 322114 271279 322142 276649
rect 322786 273943 322814 277870
rect 323554 277856 323952 277884
rect 324898 277856 325200 277884
rect 323254 275491 323306 275497
rect 323254 275433 323306 275439
rect 322774 273937 322826 273943
rect 322774 273879 322826 273885
rect 322594 272824 323006 272852
rect 322594 272611 322622 272824
rect 322978 272611 323006 272824
rect 322582 272605 322634 272611
rect 322582 272547 322634 272553
rect 322966 272605 323018 272611
rect 322966 272547 323018 272553
rect 322582 272457 322634 272463
rect 322582 272399 322634 272405
rect 322774 272457 322826 272463
rect 322774 272399 322826 272405
rect 322594 272260 322622 272399
rect 322786 272260 322814 272399
rect 322594 272232 322814 272260
rect 322582 271939 322634 271945
rect 322582 271881 322634 271887
rect 323062 271939 323114 271945
rect 323062 271881 323114 271887
rect 322594 271816 322622 271881
rect 323074 271816 323102 271881
rect 322594 271788 323102 271816
rect 323266 271409 323294 275433
rect 322690 271381 323294 271409
rect 322690 271353 322718 271381
rect 322678 271347 322730 271353
rect 322678 271289 322730 271295
rect 322774 271347 322826 271353
rect 322774 271289 322826 271295
rect 322006 271273 322058 271279
rect 322006 271215 322058 271221
rect 322102 271273 322154 271279
rect 322786 271261 322814 271289
rect 322102 271215 322154 271221
rect 322306 271233 322814 271261
rect 322018 270909 322046 271215
rect 322306 271057 322334 271233
rect 322498 271159 322814 271187
rect 322388 271090 322444 271099
rect 322294 271051 322346 271057
rect 322498 271076 322526 271159
rect 322786 271131 322814 271159
rect 322774 271125 322826 271131
rect 322444 271048 322526 271076
rect 322580 271090 322636 271099
rect 322388 271025 322444 271034
rect 322774 271067 322826 271073
rect 322580 271025 322636 271034
rect 322294 270993 322346 270999
rect 322006 270903 322058 270909
rect 322006 270845 322058 270851
rect 322594 268245 322622 271025
rect 322966 270829 323018 270835
rect 322966 270771 323018 270777
rect 322978 268393 323006 270771
rect 323554 270188 323582 277856
rect 323924 275974 323980 275983
rect 323924 275909 323980 275918
rect 323362 270160 323582 270188
rect 323362 270021 323390 270160
rect 323350 270015 323402 270021
rect 323350 269957 323402 269963
rect 323446 270015 323498 270021
rect 323446 269957 323498 269963
rect 322966 268387 323018 268393
rect 322966 268329 323018 268335
rect 323062 268387 323114 268393
rect 323062 268329 323114 268335
rect 322582 268239 322634 268245
rect 322582 268181 322634 268187
rect 322870 268239 322922 268245
rect 322870 268181 322922 268187
rect 322486 267573 322538 267579
rect 322486 267515 322538 267521
rect 322498 265156 322526 267515
rect 322882 265156 322910 268181
rect 321442 265128 321696 265156
rect 322176 265128 322526 265156
rect 322608 265128 322910 265156
rect 323074 265142 323102 268329
rect 323458 265142 323486 269957
rect 323938 268245 323966 275909
rect 324898 270835 324926 277856
rect 325076 276862 325132 276871
rect 325076 276797 325132 276806
rect 324886 270829 324938 270835
rect 324886 270771 324938 270777
rect 324982 270829 325034 270835
rect 324982 270771 325034 270777
rect 324994 268449 325022 270771
rect 324514 268421 325022 268449
rect 324514 268245 324542 268421
rect 325090 268375 325118 276797
rect 325282 273869 325310 278097
rect 325556 276714 325612 276723
rect 325556 276649 325612 276658
rect 325270 273863 325322 273869
rect 325270 273805 325322 273811
rect 325462 273715 325514 273721
rect 325462 273657 325514 273663
rect 325474 273573 325502 273657
rect 325462 273567 325514 273573
rect 325462 273509 325514 273515
rect 324994 268347 325118 268375
rect 323926 268239 323978 268245
rect 323926 268181 323978 268187
rect 324022 268239 324074 268245
rect 324022 268181 324074 268187
rect 324502 268239 324554 268245
rect 324502 268181 324554 268187
rect 324598 268239 324650 268245
rect 324598 268181 324650 268187
rect 324034 268023 324062 268181
rect 324022 268017 324074 268023
rect 324022 267959 324074 267965
rect 324118 268017 324170 268023
rect 324118 267959 324170 267965
rect 324130 265156 324158 267959
rect 324610 265156 324638 268181
rect 324994 265156 325022 268347
rect 323904 265128 324158 265156
rect 324384 265128 324638 265156
rect 324720 265128 325022 265156
rect 325570 265008 325598 276649
rect 325942 273863 325994 273869
rect 325942 273805 325994 273811
rect 325654 273715 325706 273721
rect 325654 273657 325706 273663
rect 325666 271353 325694 273657
rect 325654 271347 325706 271353
rect 325654 271289 325706 271295
rect 325654 268165 325706 268171
rect 325654 268107 325706 268113
rect 325666 265142 325694 268107
rect 325954 265156 325982 273805
rect 326338 271279 326366 277870
rect 326326 271273 326378 271279
rect 326326 271215 326378 271221
rect 326626 268023 326654 278097
rect 328150 278007 328202 278013
rect 328150 277949 328202 277955
rect 327382 277341 327434 277347
rect 327382 277283 327434 277289
rect 327094 271199 327146 271205
rect 327094 271141 327146 271147
rect 326710 268313 326762 268319
rect 326710 268255 326762 268261
rect 326806 268313 326858 268319
rect 326806 268255 326858 268261
rect 326722 268023 326750 268255
rect 326614 268017 326666 268023
rect 326614 267959 326666 267965
rect 326710 268017 326762 268023
rect 326710 267959 326762 267965
rect 326818 267653 326846 268255
rect 326998 268091 327050 268097
rect 326998 268033 327050 268039
rect 327010 267727 327038 268033
rect 326902 267721 326954 267727
rect 326902 267663 326954 267669
rect 326998 267721 327050 267727
rect 326998 267663 327050 267669
rect 326806 267647 326858 267653
rect 326806 267589 326858 267595
rect 326470 265353 326522 265359
rect 326470 265295 326522 265301
rect 326614 265353 326666 265359
rect 326614 265295 326666 265301
rect 325954 265128 326112 265156
rect 326482 265142 326510 265295
rect 326626 265137 326654 265295
rect 326914 265142 326942 267663
rect 327106 267653 327134 271141
rect 327094 267647 327146 267653
rect 327094 267589 327146 267595
rect 327394 265142 327422 277283
rect 327490 273499 327518 277870
rect 327670 277341 327722 277347
rect 327670 277283 327722 277289
rect 327682 273721 327710 277283
rect 327670 273715 327722 273721
rect 327670 273657 327722 273663
rect 327478 273493 327530 273499
rect 327478 273435 327530 273441
rect 327574 273493 327626 273499
rect 327574 273435 327626 273441
rect 327586 271427 327614 273435
rect 327574 271421 327626 271427
rect 327574 271363 327626 271369
rect 327478 271347 327530 271353
rect 327478 271289 327530 271295
rect 327490 271057 327518 271289
rect 327958 271199 328010 271205
rect 327958 271141 328010 271147
rect 327478 271051 327530 271057
rect 327478 270993 327530 270999
rect 327766 268091 327818 268097
rect 327766 268033 327818 268039
rect 327778 267801 327806 268033
rect 327860 267834 327916 267843
rect 327766 267795 327818 267801
rect 327860 267769 327862 267778
rect 327766 267737 327818 267743
rect 327914 267769 327916 267778
rect 327862 267737 327914 267743
rect 327970 265803 327998 271141
rect 328162 267783 328190 277949
rect 328532 275826 328588 275835
rect 328532 275761 328588 275770
rect 328546 271395 328574 275761
rect 328738 274165 328766 277870
rect 328726 274159 328778 274165
rect 328726 274101 328778 274107
rect 328532 271386 328588 271395
rect 328532 271321 328588 271330
rect 328628 270942 328684 270951
rect 328628 270877 328684 270886
rect 328246 270829 328298 270835
rect 328246 270771 328298 270777
rect 328342 270829 328394 270835
rect 328342 270771 328394 270777
rect 328258 270188 328286 270771
rect 328354 270317 328382 270771
rect 328438 270607 328490 270613
rect 328438 270549 328490 270555
rect 328450 270317 328478 270549
rect 328342 270311 328394 270317
rect 328342 270253 328394 270259
rect 328438 270311 328490 270317
rect 328438 270253 328490 270259
rect 328258 270160 328382 270188
rect 328354 268023 328382 270160
rect 328642 270063 328670 270877
rect 328436 270054 328492 270063
rect 328436 269989 328492 269998
rect 328628 270054 328684 270063
rect 328628 269989 328684 269998
rect 328450 268171 328478 269989
rect 328438 268165 328490 268171
rect 328438 268107 328490 268113
rect 328246 268017 328298 268023
rect 328246 267959 328298 267965
rect 328342 268017 328394 268023
rect 328342 267959 328394 267965
rect 328258 267931 328286 267959
rect 328258 267903 328670 267931
rect 328162 267755 328382 267783
rect 327862 265797 327914 265803
rect 327862 265739 327914 265745
rect 327958 265797 328010 265803
rect 327958 265739 328010 265745
rect 327874 265142 327902 265739
rect 328354 265304 328382 267755
rect 328642 267135 328670 267903
rect 328534 267129 328586 267135
rect 328534 267071 328586 267077
rect 328630 267129 328682 267135
rect 328630 267071 328682 267077
rect 328258 265276 328382 265304
rect 328258 265156 328286 265276
rect 326614 265131 326666 265137
rect 328224 265128 328286 265156
rect 328546 265156 328574 267071
rect 328546 265128 328704 265156
rect 329122 265142 329150 278393
rect 329986 271353 330014 277870
rect 330166 277119 330218 277125
rect 330166 277061 330218 277067
rect 329974 271347 330026 271353
rect 329974 271289 330026 271295
rect 329974 266241 330026 266247
rect 329974 266183 330026 266189
rect 329302 265205 329354 265211
rect 329354 265153 329616 265156
rect 329302 265147 329616 265153
rect 329314 265128 329616 265147
rect 329986 265142 330014 266183
rect 330178 265156 330206 277061
rect 331138 270317 331166 277870
rect 331318 277489 331370 277495
rect 331318 277431 331370 277437
rect 331222 270829 331274 270835
rect 331222 270771 331274 270777
rect 331234 270317 331262 270771
rect 331126 270311 331178 270317
rect 331126 270253 331178 270259
rect 331222 270311 331274 270317
rect 331222 270253 331274 270259
rect 330646 266537 330698 266543
rect 330646 266479 330698 266485
rect 330658 265156 330686 266479
rect 330178 265128 330432 265156
rect 330658 265128 330912 265156
rect 331330 265142 331358 277431
rect 332182 276601 332234 276607
rect 332182 276543 332234 276549
rect 331414 272013 331466 272019
rect 331414 271955 331466 271961
rect 331426 266543 331454 271955
rect 331702 266611 331754 266617
rect 331702 266553 331754 266559
rect 331414 266537 331466 266543
rect 331414 266479 331466 266485
rect 331714 265142 331742 266553
rect 332194 265142 332222 276543
rect 332290 271099 332318 277870
rect 332758 276823 332810 276829
rect 332758 276765 332810 276771
rect 332276 271090 332332 271099
rect 332276 271025 332332 271034
rect 332278 268313 332330 268319
rect 332278 268255 332330 268261
rect 332566 268313 332618 268319
rect 332566 268255 332618 268261
rect 332290 265211 332318 268255
rect 332578 267875 332606 268255
rect 332566 267869 332618 267875
rect 332566 267811 332618 267817
rect 332374 266907 332426 266913
rect 332374 266849 332426 266855
rect 332278 265205 332330 265211
rect 332278 265147 332330 265153
rect 332386 265156 332414 266849
rect 332770 265156 332798 276765
rect 333142 274973 333194 274979
rect 333142 274915 333194 274921
rect 333154 265156 333182 274915
rect 333442 271427 333470 277870
rect 334102 271791 334154 271797
rect 334102 271733 334154 271739
rect 333430 271421 333482 271427
rect 334114 271395 334142 271733
rect 333430 271363 333482 271369
rect 334100 271386 334156 271395
rect 334100 271321 334156 271330
rect 334100 269166 334156 269175
rect 334100 269101 334156 269110
rect 334114 267875 334142 269101
rect 334102 267869 334154 267875
rect 334102 267811 334154 267817
rect 332386 265128 332640 265156
rect 332770 265128 333024 265156
rect 333154 265128 333456 265156
rect 334402 265142 334430 278467
rect 334486 274825 334538 274831
rect 334486 274767 334538 274773
rect 334498 265156 334526 274767
rect 334594 273573 334622 277870
rect 335554 277865 335856 277884
rect 335542 277859 335856 277865
rect 335594 277856 335856 277859
rect 335542 277801 335594 277807
rect 335638 274307 335690 274313
rect 335638 274249 335690 274255
rect 334582 273567 334634 273573
rect 334582 273509 334634 273515
rect 334966 268757 335018 268763
rect 334966 268699 335018 268705
rect 335062 268757 335114 268763
rect 335062 268699 335114 268705
rect 334978 265156 335006 268699
rect 335074 267875 335102 268699
rect 335062 267869 335114 267875
rect 335062 267811 335114 267817
rect 334498 265128 334752 265156
rect 334978 265128 335232 265156
rect 335650 265142 335678 274249
rect 336994 272019 337022 277870
rect 338242 276385 338270 277870
rect 338338 276681 338366 278467
rect 350326 278451 350378 278457
rect 350326 278393 350378 278399
rect 339958 277933 340010 277939
rect 339106 277856 339408 277884
rect 339958 277875 340010 277881
rect 338710 276749 338762 276755
rect 338710 276691 338762 276697
rect 338326 276675 338378 276681
rect 338326 276617 338378 276623
rect 338230 276379 338282 276385
rect 338230 276321 338282 276327
rect 337942 274677 337994 274683
rect 337942 274619 337994 274625
rect 337558 274233 337610 274239
rect 337558 274175 337610 274181
rect 336982 272013 337034 272019
rect 336982 271955 337034 271961
rect 337270 268979 337322 268985
rect 337270 268921 337322 268927
rect 336502 268461 336554 268467
rect 336502 268403 336554 268409
rect 336598 268461 336650 268467
rect 336598 268403 336650 268409
rect 336212 268130 336268 268139
rect 336212 268065 336268 268074
rect 336404 268130 336460 268139
rect 336404 268065 336406 268074
rect 336226 267727 336254 268065
rect 336458 268065 336460 268074
rect 336406 268033 336458 268039
rect 336118 267721 336170 267727
rect 336118 267663 336170 267669
rect 336214 267721 336266 267727
rect 336214 267663 336266 267669
rect 336130 265142 336158 267663
rect 336514 265142 336542 268403
rect 336610 267949 336638 268403
rect 336982 268165 337034 268171
rect 336980 268130 336982 268139
rect 337034 268130 337036 268139
rect 336980 268065 337036 268074
rect 336598 267943 336650 267949
rect 336598 267885 336650 267891
rect 337282 265156 337310 268921
rect 337366 268461 337418 268467
rect 337366 268403 337418 268409
rect 337378 268097 337406 268403
rect 337462 268313 337514 268319
rect 337462 268255 337514 268261
rect 337366 268091 337418 268097
rect 337366 268033 337418 268039
rect 337474 267875 337502 268255
rect 337462 267869 337514 267875
rect 337462 267811 337514 267817
rect 336960 265137 337118 265156
rect 336960 265131 337130 265137
rect 336960 265128 337078 265131
rect 326614 265073 326666 265079
rect 337282 265128 337440 265156
rect 337570 265137 337598 274175
rect 337846 268905 337898 268911
rect 337846 268847 337898 268853
rect 337750 268461 337802 268467
rect 337750 268403 337802 268409
rect 337762 267801 337790 268403
rect 337750 267795 337802 267801
rect 337750 267737 337802 267743
rect 337858 265142 337886 268847
rect 337954 265156 337982 274619
rect 338516 270350 338572 270359
rect 338050 270308 338516 270336
rect 338050 270063 338078 270308
rect 338516 270285 338572 270294
rect 338036 270054 338092 270063
rect 338036 269989 338092 269998
rect 338326 268387 338378 268393
rect 338326 268329 338378 268335
rect 338338 267949 338366 268329
rect 338326 267943 338378 267949
rect 338326 267885 338378 267891
rect 338038 267795 338090 267801
rect 338038 267737 338090 267743
rect 338050 267579 338078 267737
rect 338038 267573 338090 267579
rect 338038 267515 338090 267521
rect 338326 267499 338378 267505
rect 338326 267441 338378 267447
rect 338338 266617 338366 267441
rect 338326 266611 338378 266617
rect 338326 266553 338378 266559
rect 337558 265131 337610 265137
rect 337078 265073 337130 265079
rect 337954 265128 338256 265156
rect 338722 265142 338750 276691
rect 338902 274085 338954 274091
rect 338902 274027 338954 274033
rect 338914 265156 338942 274027
rect 339106 265951 339134 277856
rect 339862 270829 339914 270835
rect 339862 270771 339914 270777
rect 339874 270317 339902 270771
rect 339862 270311 339914 270317
rect 339862 270253 339914 270259
rect 339382 266537 339434 266543
rect 339382 266479 339434 266485
rect 339094 265945 339146 265951
rect 339094 265887 339146 265893
rect 339394 265156 339422 266479
rect 339970 265156 339998 277875
rect 340642 273573 340670 277870
rect 341794 276311 341822 277870
rect 342946 276533 342974 277870
rect 342934 276527 342986 276533
rect 342934 276469 342986 276475
rect 341782 276305 341834 276311
rect 341782 276247 341834 276253
rect 341302 273937 341354 273943
rect 341302 273879 341354 273885
rect 340630 273567 340682 273573
rect 340630 273509 340682 273515
rect 340918 271125 340970 271131
rect 340918 271067 340970 271073
rect 340438 270903 340490 270909
rect 340438 270845 340490 270851
rect 338914 265128 339168 265156
rect 339394 265128 339648 265156
rect 339970 265128 340032 265156
rect 340450 265142 340478 270845
rect 340930 265142 340958 271067
rect 341314 265142 341342 273879
rect 343510 273567 343562 273573
rect 343510 273509 343562 273515
rect 343030 272013 343082 272019
rect 343030 271955 343082 271961
rect 342646 271421 342698 271427
rect 342646 271363 342698 271369
rect 341974 271347 342026 271353
rect 341974 271289 342026 271295
rect 341494 271273 341546 271279
rect 341494 271215 341546 271221
rect 341506 265156 341534 271215
rect 341986 265156 342014 271289
rect 341506 265128 341760 265156
rect 341986 265128 342240 265156
rect 342658 265142 342686 271363
rect 343042 265142 343070 271955
rect 343522 265142 343550 273509
rect 344194 265156 344222 277870
rect 344662 273567 344714 273573
rect 344662 273509 344714 273515
rect 344674 265156 344702 273509
rect 345238 271125 345290 271131
rect 345238 271067 345290 271073
rect 344758 270903 344810 270909
rect 344758 270845 344810 270851
rect 343968 265128 344222 265156
rect 344448 265128 344702 265156
rect 344770 265142 344798 270845
rect 344854 267647 344906 267653
rect 344854 267589 344906 267595
rect 344866 265137 344894 267589
rect 345250 265142 345278 271067
rect 345346 270835 345374 277870
rect 345718 271273 345770 271279
rect 345718 271215 345770 271221
rect 345334 270829 345386 270835
rect 345334 270771 345386 270777
rect 345730 265142 345758 271215
rect 346390 271199 346442 271205
rect 346390 271141 346442 271147
rect 346402 265156 346430 271141
rect 346594 267431 346622 277870
rect 346774 276379 346826 276385
rect 346774 276321 346826 276327
rect 346582 267425 346634 267431
rect 346582 267367 346634 267373
rect 346786 265156 346814 276321
rect 347746 273573 347774 277870
rect 348886 276823 348938 276829
rect 348886 276765 348938 276771
rect 348406 276305 348458 276311
rect 348406 276247 348458 276253
rect 347734 273567 347786 273573
rect 347734 273509 347786 273515
rect 347926 272013 347978 272019
rect 347926 271955 347978 271961
rect 347446 271421 347498 271427
rect 347446 271363 347498 271369
rect 347252 269166 347308 269175
rect 347252 269101 347308 269110
rect 347266 267431 347294 269101
rect 347254 267425 347306 267431
rect 347254 267367 347306 267373
rect 347254 266241 347306 266247
rect 347254 266183 347306 266189
rect 347266 265156 347294 266183
rect 344854 265131 344906 265137
rect 337558 265073 337610 265079
rect 346176 265128 346430 265156
rect 346560 265128 346814 265156
rect 346992 265128 347294 265156
rect 347458 265142 347486 271363
rect 347830 270829 347882 270835
rect 347830 270771 347882 270777
rect 347540 269166 347596 269175
rect 347540 269101 347596 269110
rect 347554 268245 347582 269101
rect 347542 268239 347594 268245
rect 347542 268181 347594 268187
rect 347842 266247 347870 270771
rect 347830 266241 347882 266247
rect 347830 266183 347882 266189
rect 347938 265142 347966 271955
rect 348020 269166 348076 269175
rect 348020 269101 348076 269110
rect 348034 268763 348062 269101
rect 348022 268757 348074 268763
rect 348022 268699 348074 268705
rect 348418 265156 348446 276247
rect 348596 268426 348652 268435
rect 348596 268361 348652 268370
rect 348502 268313 348554 268319
rect 348502 268255 348554 268261
rect 348514 267135 348542 268255
rect 348610 268097 348638 268361
rect 348598 268091 348650 268097
rect 348598 268033 348650 268039
rect 348502 267129 348554 267135
rect 348502 267071 348554 267077
rect 348598 267129 348650 267135
rect 348598 267071 348650 267077
rect 348502 265797 348554 265803
rect 348502 265739 348554 265745
rect 348288 265128 348446 265156
rect 344854 265073 344906 265079
rect 321046 264983 321098 264989
rect 318934 264925 318986 264931
rect 325200 264980 325598 265008
rect 333622 265057 333674 265063
rect 333674 265005 333936 265008
rect 333622 264999 333936 265005
rect 333634 264980 333936 264999
rect 321046 264925 321098 264931
rect 212470 264909 212522 264915
rect 348514 264915 348542 265739
rect 348610 264989 348638 267071
rect 348898 265156 348926 276765
rect 348994 276015 349022 277870
rect 349078 277119 349130 277125
rect 349078 277061 349130 277067
rect 348982 276009 349034 276015
rect 348982 275951 349034 275957
rect 349090 272260 349118 277061
rect 350050 276903 350078 277870
rect 350038 276897 350090 276903
rect 350038 276839 350090 276845
rect 349172 272570 349228 272579
rect 349172 272505 349228 272514
rect 349186 272408 349214 272505
rect 349460 272422 349516 272431
rect 349186 272380 349460 272408
rect 349460 272357 349516 272366
rect 349090 272232 349214 272260
rect 349078 268979 349130 268985
rect 349078 268921 349130 268927
rect 349090 267875 349118 268921
rect 349078 267869 349130 267875
rect 349078 267811 349130 267817
rect 348768 265128 348926 265156
rect 349186 265142 349214 272232
rect 349558 266907 349610 266913
rect 349558 266849 349610 266855
rect 349570 265142 349598 266849
rect 350338 265156 350366 278393
rect 353494 278007 353546 278013
rect 353494 277949 353546 277955
rect 357430 278007 357482 278013
rect 357430 277949 357482 277955
rect 351094 276527 351146 276533
rect 351094 276469 351146 276475
rect 350710 265797 350762 265803
rect 350710 265739 350762 265745
rect 350722 265156 350750 265739
rect 351106 265156 351134 276469
rect 351298 270909 351326 277870
rect 352246 274233 352298 274239
rect 352246 274175 352298 274181
rect 351286 270903 351338 270909
rect 351286 270845 351338 270851
rect 351766 268905 351818 268911
rect 351766 268847 351818 268853
rect 351286 267647 351338 267653
rect 351286 267589 351338 267595
rect 350064 265128 350366 265156
rect 350496 265128 350750 265156
rect 350976 265128 351134 265156
rect 351298 265142 351326 267589
rect 351778 265142 351806 268847
rect 352258 265142 352286 274175
rect 352450 270243 352478 277870
rect 352918 277489 352970 277495
rect 352918 277431 352970 277437
rect 352438 270237 352490 270243
rect 352438 270179 352490 270185
rect 352930 265156 352958 277431
rect 353302 267573 353354 267579
rect 353302 267515 353354 267521
rect 353314 265156 353342 267515
rect 352704 265128 352958 265156
rect 353088 265128 353342 265156
rect 353506 265142 353534 277949
rect 355510 277933 355562 277939
rect 355510 277875 355562 277881
rect 353698 267283 353726 277870
rect 354454 273715 354506 273721
rect 354454 273657 354506 273663
rect 353974 268091 354026 268097
rect 353974 268033 354026 268039
rect 353686 267277 353738 267283
rect 353686 267219 353738 267225
rect 353986 265142 354014 268033
rect 354466 265142 354494 273657
rect 354850 271131 354878 277870
rect 354838 271125 354890 271131
rect 354838 271067 354890 271073
rect 355030 267499 355082 267505
rect 355030 267441 355082 267447
rect 355042 265156 355070 267441
rect 355522 265156 355550 277875
rect 356098 275719 356126 277870
rect 356854 277859 356906 277865
rect 356854 277801 356906 277807
rect 357058 277856 357264 277884
rect 356086 275713 356138 275719
rect 356086 275655 356138 275661
rect 356182 273863 356234 273869
rect 356182 273805 356234 273811
rect 355702 268165 355754 268171
rect 355702 268107 355754 268113
rect 354816 265128 355070 265156
rect 355296 265128 355550 265156
rect 355714 265142 355742 268107
rect 356194 265142 356222 273805
rect 356866 272852 356894 277801
rect 357058 277791 357086 277856
rect 357046 277785 357098 277791
rect 357046 277727 357098 277733
rect 356950 277711 357002 277717
rect 356950 277653 357002 277659
rect 356962 273573 356990 277653
rect 357442 277495 357470 277949
rect 358114 277856 358416 277884
rect 357430 277489 357482 277495
rect 357430 277431 357482 277437
rect 356950 273567 357002 273573
rect 356950 273509 357002 273515
rect 356866 272824 356990 272852
rect 356566 267277 356618 267283
rect 356566 267219 356618 267225
rect 356578 265142 356606 267219
rect 356962 265452 356990 272824
rect 357046 271791 357098 271797
rect 357046 271733 357098 271739
rect 357058 271395 357086 271733
rect 357044 271386 357100 271395
rect 357044 271321 357100 271330
rect 357334 271347 357386 271353
rect 357334 271289 357386 271295
rect 357346 267727 357374 271289
rect 358114 271279 358142 277856
rect 358594 276607 358622 278467
rect 358870 277711 358922 277717
rect 358870 277653 358922 277659
rect 358582 276601 358634 276607
rect 358582 276543 358634 276549
rect 358774 274307 358826 274313
rect 358774 274249 358826 274255
rect 358306 272528 358622 272556
rect 358306 272431 358334 272528
rect 358292 272422 358348 272431
rect 358292 272357 358348 272366
rect 358484 272422 358540 272431
rect 358484 272357 358540 272366
rect 358498 272135 358526 272357
rect 358484 272126 358540 272135
rect 358594 272112 358622 272528
rect 358676 272126 358732 272135
rect 358594 272084 358676 272112
rect 358484 272061 358540 272070
rect 358676 272061 358732 272070
rect 358102 271273 358154 271279
rect 358102 271215 358154 271221
rect 357718 271125 357770 271131
rect 357718 271067 357770 271073
rect 357622 270311 357674 270317
rect 357622 270253 357674 270259
rect 357634 269725 357662 270253
rect 357622 269719 357674 269725
rect 357622 269661 357674 269667
rect 357334 267721 357386 267727
rect 357334 267663 357386 267669
rect 357430 267721 357482 267727
rect 357430 267663 357482 267669
rect 357442 266913 357470 267663
rect 357430 266907 357482 266913
rect 357430 266849 357482 266855
rect 356962 265424 357038 265452
rect 357010 265142 357038 265424
rect 357730 265156 357758 271067
rect 358486 270237 358538 270243
rect 358486 270179 358538 270185
rect 358498 269577 358526 270179
rect 358786 269744 358814 274249
rect 358582 269719 358634 269725
rect 358582 269661 358634 269667
rect 358690 269716 358814 269744
rect 358486 269571 358538 269577
rect 358486 269513 358538 269519
rect 358594 268541 358622 269661
rect 358582 268535 358634 268541
rect 358582 268477 358634 268483
rect 358690 268412 358718 269716
rect 358594 268384 358718 268412
rect 357814 266241 357866 266247
rect 357814 266183 357866 266189
rect 357504 265128 357758 265156
rect 357826 265142 357854 266183
rect 358594 265156 358622 268384
rect 358882 268264 358910 277653
rect 359650 270095 359678 277870
rect 360502 274085 360554 274091
rect 360502 274027 360554 274033
rect 360022 273937 360074 273943
rect 360022 273879 360074 273885
rect 359638 270089 359690 270095
rect 359638 270031 359690 270037
rect 358320 265128 358622 265156
rect 358786 268236 358910 268264
rect 359446 268239 359498 268245
rect 358786 265142 358814 268236
rect 359446 268181 359498 268187
rect 359458 265156 359486 268181
rect 359830 266907 359882 266913
rect 359830 266849 359882 266855
rect 359842 265156 359870 266849
rect 359232 265128 359486 265156
rect 359616 265128 359870 265156
rect 360034 265142 360062 273879
rect 360514 265142 360542 274027
rect 360802 266617 360830 277870
rect 361558 277489 361610 277495
rect 361558 277431 361610 277437
rect 360982 268387 361034 268393
rect 360982 268329 361034 268335
rect 360790 266611 360842 266617
rect 360790 266553 360842 266559
rect 360994 265142 361022 268329
rect 361570 265156 361598 277431
rect 362050 271205 362078 277870
rect 363202 275423 363230 277870
rect 364450 277051 364478 277870
rect 364438 277045 364490 277051
rect 364438 276987 364490 276993
rect 364822 277045 364874 277051
rect 364822 276987 364874 276993
rect 363766 276675 363818 276681
rect 363766 276617 363818 276623
rect 363190 275417 363242 275423
rect 363190 275359 363242 275365
rect 362038 271199 362090 271205
rect 362038 271141 362090 271147
rect 362038 270829 362090 270835
rect 362038 270771 362090 270777
rect 362050 265156 362078 270771
rect 363094 270089 363146 270095
rect 363094 270031 363146 270037
rect 362230 266611 362282 266617
rect 362230 266553 362282 266559
rect 361344 265128 361598 265156
rect 361824 265128 362078 265156
rect 362242 265142 362270 266553
rect 362710 266537 362762 266543
rect 362710 266479 362762 266485
rect 362722 265142 362750 266479
rect 363106 265142 363134 270031
rect 363778 265156 363806 276617
rect 364246 275713 364298 275719
rect 364246 275655 364298 275661
rect 364258 265156 364286 275655
rect 364342 274159 364394 274165
rect 364342 274101 364394 274107
rect 363552 265128 363806 265156
rect 364032 265128 364286 265156
rect 364354 265142 364382 274101
rect 364834 265142 364862 276987
rect 365302 276897 365354 276903
rect 365302 276839 365354 276845
rect 365206 267425 365258 267431
rect 365206 267367 365258 267373
rect 365218 264989 365246 267367
rect 365314 265142 365342 276839
rect 365602 276385 365630 277870
rect 365590 276379 365642 276385
rect 365590 276321 365642 276327
rect 366454 271347 366506 271353
rect 366454 271289 366506 271295
rect 366466 268467 366494 271289
rect 366754 270317 366782 277870
rect 367906 273573 367934 277870
rect 368578 276681 368798 276700
rect 368566 276675 368810 276681
rect 368618 276672 368758 276675
rect 368566 276617 368618 276623
rect 368758 276617 368810 276623
rect 368086 274973 368138 274979
rect 368086 274915 368138 274921
rect 367894 273567 367946 273573
rect 367894 273509 367946 273515
rect 367126 271273 367178 271279
rect 367124 271238 367126 271247
rect 367178 271238 367180 271247
rect 367124 271173 367180 271182
rect 367124 271090 367180 271099
rect 367124 271025 367180 271034
rect 366742 270311 366794 270317
rect 366742 270253 366794 270259
rect 367030 270311 367082 270317
rect 367030 270253 367082 270259
rect 366646 270015 366698 270021
rect 366646 269957 366698 269963
rect 366742 270015 366794 270021
rect 366742 269957 366794 269963
rect 366550 268535 366602 268541
rect 366550 268477 366602 268483
rect 366454 268461 366506 268467
rect 366454 268403 366506 268409
rect 366358 267869 366410 267875
rect 366358 267811 366410 267817
rect 366370 265156 366398 267811
rect 366144 265128 366398 265156
rect 366562 265142 366590 268477
rect 366658 268467 366686 269957
rect 366754 268615 366782 269957
rect 366742 268609 366794 268615
rect 366742 268551 366794 268557
rect 366646 268461 366698 268467
rect 366646 268403 366698 268409
rect 367042 267357 367070 270253
rect 367138 269175 367166 271025
rect 367124 269166 367180 269175
rect 367124 269101 367180 269110
rect 367510 268757 367562 268763
rect 367510 268699 367562 268705
rect 367030 267351 367082 267357
rect 367030 267293 367082 267299
rect 367126 267351 367178 267357
rect 367126 267293 367178 267299
rect 367138 267209 367166 267293
rect 367126 267203 367178 267209
rect 367126 267145 367178 267151
rect 367318 267129 367370 267135
rect 367318 267071 367370 267077
rect 367030 265945 367082 265951
rect 367030 265887 367082 265893
rect 367042 265142 367070 265887
rect 367330 265211 367358 267071
rect 367318 265205 367370 265211
rect 367318 265147 367370 265153
rect 367522 265142 367550 268699
rect 367798 267721 367850 267727
rect 367798 267663 367850 267669
rect 367810 267505 367838 267663
rect 367798 267499 367850 267505
rect 367798 267441 367850 267447
rect 368098 265156 368126 274915
rect 368660 271386 368716 271395
rect 368660 271321 368716 271330
rect 368564 270942 368620 270951
rect 368564 270877 368620 270886
rect 368578 270780 368606 270877
rect 368674 270780 368702 271321
rect 369154 270909 369182 277870
rect 370306 275349 370334 277870
rect 371568 277856 371678 277884
rect 370966 276897 371018 276903
rect 370966 276839 371018 276845
rect 370978 276755 371006 276839
rect 370966 276749 371018 276755
rect 370966 276691 371018 276697
rect 370966 276379 371018 276385
rect 370966 276321 371018 276327
rect 370390 276009 370442 276015
rect 370390 275951 370442 275957
rect 370294 275343 370346 275349
rect 370294 275285 370346 275291
rect 369236 274938 369292 274947
rect 369236 274873 369292 274882
rect 369250 270909 369278 274873
rect 369526 274677 369578 274683
rect 369526 274619 369578 274625
rect 369142 270903 369194 270909
rect 369142 270845 369194 270851
rect 369238 270903 369290 270909
rect 369238 270845 369290 270851
rect 368578 270752 368702 270780
rect 369430 270829 369482 270835
rect 369430 270771 369482 270777
rect 369442 270655 369470 270771
rect 368468 270646 368524 270655
rect 369428 270646 369484 270655
rect 368468 270581 368470 270590
rect 368522 270581 368524 270590
rect 368758 270607 368810 270613
rect 368470 270549 368522 270555
rect 369428 270581 369484 270590
rect 368758 270549 368810 270555
rect 368470 269571 368522 269577
rect 368470 269513 368522 269519
rect 368482 265156 368510 269513
rect 368770 269175 368798 270549
rect 368756 269166 368812 269175
rect 368756 269101 368812 269110
rect 368566 267721 368618 267727
rect 368566 267663 368618 267669
rect 368578 265803 368606 267663
rect 369058 267607 369374 267635
rect 368758 267499 368810 267505
rect 368758 267441 368810 267447
rect 368770 265803 368798 267441
rect 369058 267283 369086 267607
rect 369142 267499 369194 267505
rect 369142 267441 369194 267447
rect 369046 267277 369098 267283
rect 369046 267219 369098 267225
rect 368566 265797 368618 265803
rect 368566 265739 368618 265745
rect 368758 265797 368810 265803
rect 368758 265739 368810 265745
rect 369154 265156 369182 267441
rect 369346 267283 369374 267607
rect 369334 267277 369386 267283
rect 369334 267219 369386 267225
rect 367872 265128 368126 265156
rect 368352 265128 368510 265156
rect 368784 265128 369182 265156
rect 365974 265057 366026 265063
rect 365760 265005 365974 265008
rect 369538 265008 369566 274619
rect 369910 270829 369962 270835
rect 369910 270771 369962 270777
rect 369812 270646 369868 270655
rect 369812 270581 369868 270590
rect 369826 268985 369854 270581
rect 369814 268979 369866 268985
rect 369814 268921 369866 268927
rect 369922 265156 369950 270771
rect 370004 270646 370060 270655
rect 370004 270581 370060 270590
rect 370018 270539 370046 270581
rect 370006 270533 370058 270539
rect 370006 270475 370058 270481
rect 370402 265156 370430 275951
rect 370774 268609 370826 268615
rect 370774 268551 370826 268557
rect 370786 265156 370814 268551
rect 369648 265128 369950 265156
rect 370080 265128 370430 265156
rect 370560 265128 370814 265156
rect 370978 265142 371006 276321
rect 371542 273271 371594 273277
rect 371542 273213 371594 273219
rect 371554 271131 371582 273213
rect 371446 271125 371498 271131
rect 371446 271067 371498 271073
rect 371542 271125 371594 271131
rect 371542 271067 371594 271073
rect 371458 270539 371486 271067
rect 371446 270533 371498 270539
rect 371446 270475 371498 270481
rect 371650 270317 371678 277856
rect 371830 275417 371882 275423
rect 371830 275359 371882 275365
rect 371638 270311 371690 270317
rect 371638 270253 371690 270259
rect 371350 268979 371402 268985
rect 371350 268921 371402 268927
rect 371362 265142 371390 268921
rect 371842 265142 371870 275359
rect 372310 274825 372362 274831
rect 372310 274767 372362 274773
rect 372322 274387 372350 274767
rect 372310 274381 372362 274387
rect 372310 274323 372362 274329
rect 372406 274233 372458 274239
rect 372406 274175 372458 274181
rect 372418 273647 372446 274175
rect 372406 273641 372458 273647
rect 372406 273583 372458 273589
rect 372706 271427 372734 277870
rect 373378 276575 373406 278573
rect 379030 278541 379082 278547
rect 379126 278599 379178 278605
rect 379126 278541 379178 278547
rect 374818 278309 375120 278328
rect 374806 278303 375120 278309
rect 374858 278300 375120 278303
rect 375478 278303 375530 278309
rect 374806 278245 374858 278251
rect 375478 278245 375530 278251
rect 373474 277856 373872 277884
rect 373364 276566 373420 276575
rect 373364 276501 373420 276510
rect 372886 275343 372938 275349
rect 372886 275285 372938 275291
rect 372694 271421 372746 271427
rect 372694 271363 372746 271369
rect 372502 270607 372554 270613
rect 372502 270549 372554 270555
rect 372514 265156 372542 270549
rect 372898 265156 372926 275285
rect 372982 271273 373034 271279
rect 372982 271215 373034 271221
rect 372994 269577 373022 271215
rect 373366 270311 373418 270317
rect 373366 270253 373418 270259
rect 372982 269571 373034 269577
rect 372982 269513 373034 269519
rect 373378 265156 373406 270253
rect 373474 270243 373502 277856
rect 373940 276566 373996 276575
rect 373940 276501 373996 276510
rect 373954 273444 373982 276501
rect 375490 276385 375518 278245
rect 375478 276379 375530 276385
rect 375478 276321 375530 276327
rect 375574 276379 375626 276385
rect 375574 276321 375626 276327
rect 374134 274233 374186 274239
rect 374134 274175 374186 274181
rect 374146 273467 374174 274175
rect 374326 274159 374378 274165
rect 374326 274101 374378 274107
rect 374338 273615 374366 274101
rect 374324 273606 374380 273615
rect 374324 273541 374380 273550
rect 373762 273416 373982 273444
rect 374132 273458 374188 273467
rect 373462 270237 373514 270243
rect 373462 270179 373514 270185
rect 373558 270237 373610 270243
rect 373558 270179 373610 270185
rect 372288 265128 372542 265156
rect 372672 265128 372926 265156
rect 373152 265128 373406 265156
rect 373570 265142 373598 270179
rect 373762 270021 373790 273416
rect 374132 273393 374188 273402
rect 374708 273310 374764 273319
rect 374326 273271 374378 273277
rect 373858 273231 374326 273259
rect 373858 273129 373886 273231
rect 374708 273245 374764 273254
rect 374326 273213 374378 273219
rect 373846 273123 373898 273129
rect 373846 273065 373898 273071
rect 374614 273123 374666 273129
rect 374614 273065 374666 273071
rect 374626 273000 374654 273065
rect 374434 272981 374654 273000
rect 374422 272975 374654 272981
rect 374474 272972 374654 272975
rect 374422 272917 374474 272923
rect 374326 272901 374378 272907
rect 374614 272901 374666 272907
rect 374378 272849 374614 272852
rect 374326 272843 374666 272849
rect 374338 272824 374654 272843
rect 374722 272727 374750 273245
rect 374806 272827 374858 272833
rect 374806 272769 374858 272775
rect 374708 272718 374764 272727
rect 374708 272653 374764 272662
rect 374818 272112 374846 272769
rect 375188 272126 375244 272135
rect 374530 272084 374846 272112
rect 374914 272084 375188 272112
rect 374530 272019 374558 272084
rect 374518 272013 374570 272019
rect 374518 271955 374570 271961
rect 374710 272013 374762 272019
rect 374914 271987 374942 272084
rect 375188 272061 375244 272070
rect 374710 271955 374762 271961
rect 374900 271978 374956 271987
rect 374324 270942 374380 270951
rect 374324 270877 374380 270886
rect 373750 270015 373802 270021
rect 373750 269957 373802 269963
rect 374038 270015 374090 270021
rect 374038 269957 374090 269963
rect 374050 265142 374078 269957
rect 374338 268319 374366 270877
rect 374422 270829 374474 270835
rect 374422 270771 374474 270777
rect 374518 270829 374570 270835
rect 374518 270771 374570 270777
rect 374434 269577 374462 270771
rect 374530 270021 374558 270771
rect 374518 270015 374570 270021
rect 374518 269957 374570 269963
rect 374422 269571 374474 269577
rect 374422 269513 374474 269519
rect 374326 268313 374378 268319
rect 374326 268255 374378 268261
rect 374422 268313 374474 268319
rect 374422 268255 374474 268261
rect 374434 266044 374462 268255
rect 374242 266016 374462 266044
rect 374242 265137 374270 266016
rect 374722 265156 374750 271955
rect 374900 271913 374956 271922
rect 374902 270015 374954 270021
rect 374902 269957 374954 269963
rect 374806 267499 374858 267505
rect 374806 267441 374858 267447
rect 374818 265433 374846 267441
rect 374806 265427 374858 265433
rect 374806 265369 374858 265375
rect 374914 265304 374942 269957
rect 375010 267681 375422 267709
rect 375010 267579 375038 267681
rect 375190 267647 375242 267653
rect 375190 267589 375242 267595
rect 374998 267573 375050 267579
rect 374998 267515 375050 267521
rect 375202 267135 375230 267589
rect 375394 267579 375422 267681
rect 375382 267573 375434 267579
rect 375382 267515 375434 267521
rect 375190 267129 375242 267135
rect 375190 267071 375242 267077
rect 374230 265131 374282 265137
rect 374448 265128 374750 265156
rect 374866 265276 374942 265304
rect 374866 265142 374894 265276
rect 375586 265156 375614 276321
rect 376258 272833 376286 277870
rect 376546 277412 377054 277440
rect 376546 276589 376574 277412
rect 376642 277264 376958 277292
rect 376642 276977 376670 277264
rect 376930 276977 376958 277264
rect 377026 277051 377054 277412
rect 377014 277045 377066 277051
rect 377014 276987 377066 276993
rect 376630 276971 376682 276977
rect 376630 276913 376682 276919
rect 376918 276971 376970 276977
rect 376918 276913 376970 276919
rect 376546 276561 376670 276589
rect 376532 273014 376588 273023
rect 376532 272949 376588 272958
rect 376246 272827 376298 272833
rect 376246 272769 376298 272775
rect 376342 272827 376394 272833
rect 376342 272769 376394 272775
rect 375668 272570 375724 272579
rect 375668 272505 375724 272514
rect 375682 269725 375710 272505
rect 375670 269719 375722 269725
rect 375670 269661 375722 269667
rect 375766 269719 375818 269725
rect 375766 269661 375818 269667
rect 375360 265128 375614 265156
rect 375778 265142 375806 269661
rect 376354 268319 376382 272769
rect 376546 272283 376574 272949
rect 376532 272274 376588 272283
rect 376532 272209 376588 272218
rect 376342 268313 376394 268319
rect 376342 268255 376394 268261
rect 375958 267129 376010 267135
rect 375958 267071 376010 267077
rect 375970 266247 375998 267071
rect 375958 266241 376010 266247
rect 375958 266183 376010 266189
rect 376438 265427 376490 265433
rect 376438 265369 376490 265375
rect 376450 265156 376478 265369
rect 376176 265128 376478 265156
rect 376642 265142 376670 276561
rect 377506 275127 377534 277870
rect 377698 277856 378672 277884
rect 377590 275343 377642 275349
rect 377590 275285 377642 275291
rect 377602 275127 377630 275285
rect 377494 275121 377546 275127
rect 377494 275063 377546 275069
rect 377590 275121 377642 275127
rect 377590 275063 377642 275069
rect 377492 274938 377548 274947
rect 377492 274873 377548 274882
rect 377506 273795 377534 274873
rect 377494 273789 377546 273795
rect 377494 273731 377546 273737
rect 377590 273789 377642 273795
rect 377590 273731 377642 273737
rect 377300 273458 377356 273467
rect 377492 273458 377548 273467
rect 377300 273393 377356 273402
rect 377410 273416 377492 273444
rect 377314 273023 377342 273393
rect 377300 273014 377356 273023
rect 377300 272949 377356 272958
rect 377410 272833 377438 273416
rect 377492 273393 377548 273402
rect 377398 272827 377450 272833
rect 377398 272769 377450 272775
rect 377494 272827 377546 272833
rect 377494 272769 377546 272775
rect 377506 271797 377534 272769
rect 377494 271791 377546 271797
rect 377494 271733 377546 271739
rect 377300 271238 377356 271247
rect 377110 271199 377162 271205
rect 377206 271199 377258 271205
rect 377162 271159 377206 271187
rect 377110 271141 377162 271147
rect 377300 271173 377356 271182
rect 377206 271141 377258 271147
rect 377026 271057 377150 271076
rect 377014 271051 377162 271057
rect 377066 271048 377110 271051
rect 377014 270993 377066 270999
rect 377110 270993 377162 270999
rect 376834 269272 377054 269300
rect 376834 268615 376862 269272
rect 376916 269166 376972 269175
rect 377026 269152 377054 269272
rect 377108 269166 377164 269175
rect 377026 269124 377108 269152
rect 376916 269101 376972 269110
rect 377108 269101 377164 269110
rect 376822 268609 376874 268615
rect 376822 268551 376874 268557
rect 376822 268313 376874 268319
rect 376822 268255 376874 268261
rect 376834 267843 376862 268255
rect 376820 267834 376876 267843
rect 376820 267769 376876 267778
rect 376930 267653 376958 269101
rect 377014 268609 377066 268615
rect 377014 268551 377066 268557
rect 377026 267949 377054 268551
rect 377204 267982 377260 267991
rect 377014 267943 377066 267949
rect 377314 267968 377342 271173
rect 377602 268116 377630 273731
rect 377698 273467 377726 277856
rect 378550 277045 378602 277051
rect 378550 276987 378602 276993
rect 378646 277045 378698 277051
rect 378646 276987 378698 276993
rect 378562 276552 378590 276987
rect 378658 276681 378686 276987
rect 378646 276675 378698 276681
rect 378646 276617 378698 276623
rect 378742 276675 378794 276681
rect 378742 276617 378794 276623
rect 378754 276552 378782 276617
rect 379138 276607 379166 278541
rect 379330 278365 379358 278633
rect 384020 278638 384076 278647
rect 379702 278599 379754 278605
rect 396226 278605 396528 278624
rect 403330 278605 403632 278624
rect 384020 278573 384076 278582
rect 396214 278599 396528 278605
rect 379702 278541 379754 278547
rect 379714 278365 379742 278541
rect 379330 278337 379742 278365
rect 379522 278004 379920 278032
rect 378562 276524 378782 276552
rect 379126 276601 379178 276607
rect 379126 276543 379178 276549
rect 379522 276311 379550 278004
rect 380002 277856 381072 277884
rect 380002 276811 380030 277856
rect 382306 277569 382334 277870
rect 382294 277563 382346 277569
rect 382294 277505 382346 277511
rect 383362 276829 383390 277870
rect 379618 276783 380030 276811
rect 383350 276823 383402 276829
rect 379510 276305 379562 276311
rect 379510 276247 379562 276253
rect 377878 275417 377930 275423
rect 377878 275359 377930 275365
rect 377684 273458 377740 273467
rect 377684 273393 377740 273402
rect 377782 271791 377834 271797
rect 377782 271733 377834 271739
rect 377260 267940 377342 267968
rect 377506 268088 377630 268116
rect 377204 267917 377260 267926
rect 377014 267885 377066 267891
rect 377012 267834 377068 267843
rect 377012 267769 377068 267778
rect 376822 267647 376874 267653
rect 376822 267589 376874 267595
rect 376918 267647 376970 267653
rect 376918 267589 376970 267595
rect 376834 267524 376862 267589
rect 376834 267496 376958 267524
rect 376930 267117 376958 267496
rect 377026 267209 377054 267769
rect 377506 267376 377534 268088
rect 377122 267348 377534 267376
rect 377014 267203 377066 267209
rect 377014 267145 377066 267151
rect 377122 267117 377150 267348
rect 377206 267203 377258 267209
rect 377206 267145 377258 267151
rect 376930 267089 377150 267117
rect 376918 266241 376970 266247
rect 376918 266183 376970 266189
rect 376930 265600 376958 266183
rect 376738 265572 376958 265600
rect 374230 265073 374282 265079
rect 376738 265063 376766 265572
rect 377218 265433 377246 267145
rect 377206 265427 377258 265433
rect 377206 265369 377258 265375
rect 377794 265156 377822 271733
rect 377890 270188 377918 275359
rect 379414 275343 379466 275349
rect 379414 275285 379466 275291
rect 379510 275343 379562 275349
rect 379510 275285 379562 275291
rect 378562 275044 378782 275072
rect 378562 274683 378590 275044
rect 378754 274979 378782 275044
rect 378646 274973 378698 274979
rect 378646 274915 378698 274921
rect 378742 274973 378794 274979
rect 379426 274947 379454 275285
rect 378742 274915 378794 274921
rect 379028 274938 379084 274947
rect 378658 274683 378686 274915
rect 379028 274873 379084 274882
rect 379412 274938 379468 274947
rect 379412 274873 379468 274882
rect 378550 274677 378602 274683
rect 378550 274619 378602 274625
rect 378646 274677 378698 274683
rect 378646 274619 378698 274625
rect 378466 274452 378878 274480
rect 378466 274239 378494 274452
rect 378850 274387 378878 274452
rect 378742 274381 378794 274387
rect 378742 274323 378794 274329
rect 378838 274381 378890 274387
rect 378838 274323 378890 274329
rect 378454 274233 378506 274239
rect 378454 274175 378506 274181
rect 378550 274233 378602 274239
rect 378550 274175 378602 274181
rect 378562 274017 378590 274175
rect 378646 274085 378698 274091
rect 378646 274027 378698 274033
rect 378550 274011 378602 274017
rect 378550 273953 378602 273959
rect 378260 273902 378316 273911
rect 378260 273837 378316 273846
rect 378452 273902 378508 273911
rect 378452 273837 378508 273846
rect 378274 273467 378302 273837
rect 378260 273458 378316 273467
rect 378260 273393 378316 273402
rect 378466 272907 378494 273837
rect 378658 273777 378686 274027
rect 378754 273943 378782 274323
rect 378838 274159 378890 274165
rect 378838 274101 378890 274107
rect 378742 273937 378794 273943
rect 378742 273879 378794 273885
rect 378850 273777 378878 274101
rect 378658 273749 378878 273777
rect 378454 272901 378506 272907
rect 378082 272861 378398 272889
rect 378082 272389 378110 272861
rect 378166 272827 378218 272833
rect 378166 272769 378218 272775
rect 378070 272383 378122 272389
rect 378178 272371 378206 272769
rect 378370 272593 378398 272861
rect 378454 272843 378506 272849
rect 378562 272824 378878 272852
rect 378454 272753 378506 272759
rect 378562 272704 378590 272824
rect 378850 272759 378878 272824
rect 378506 272701 378590 272704
rect 378454 272695 378590 272701
rect 378838 272753 378890 272759
rect 378838 272695 378890 272701
rect 378466 272676 378590 272695
rect 378742 272679 378794 272685
rect 378742 272621 378794 272627
rect 378754 272593 378782 272621
rect 378370 272565 378782 272593
rect 378742 272531 378794 272537
rect 378370 272491 378686 272519
rect 378178 272343 378302 272371
rect 378070 272325 378122 272331
rect 378164 272126 378220 272135
rect 378164 272061 378220 272070
rect 378274 272075 378302 272343
rect 378370 272167 378398 272491
rect 378454 272457 378506 272463
rect 378658 272445 378686 272491
rect 378794 272491 378974 272519
rect 378742 272473 378794 272479
rect 378838 272457 378890 272463
rect 378658 272417 378838 272445
rect 378454 272399 378506 272405
rect 378838 272399 378890 272405
rect 378358 272161 378410 272167
rect 378466 272149 378494 272399
rect 378946 272389 378974 272491
rect 378934 272383 378986 272389
rect 378934 272325 378986 272331
rect 379042 272241 379070 274873
rect 379222 272531 379274 272537
rect 379222 272473 379274 272479
rect 379126 272457 379178 272463
rect 379126 272399 379178 272405
rect 379030 272235 379082 272241
rect 379030 272177 379082 272183
rect 378466 272121 378878 272149
rect 378358 272103 378410 272109
rect 378178 271247 378206 272061
rect 378274 272047 378686 272075
rect 378658 272019 378686 272047
rect 378550 272013 378602 272019
rect 378550 271955 378602 271961
rect 378646 272013 378698 272019
rect 378646 271955 378698 271961
rect 378164 271238 378220 271247
rect 378164 271173 378220 271182
rect 378562 270965 378590 271955
rect 378742 271791 378794 271797
rect 378742 271733 378794 271739
rect 378754 271631 378782 271733
rect 378850 271705 378878 272121
rect 379028 272126 379084 272135
rect 379028 272061 379084 272070
rect 379042 271797 379070 272061
rect 379030 271791 379082 271797
rect 379030 271733 379082 271739
rect 379138 271705 379166 272399
rect 378850 271677 379166 271705
rect 379234 271631 379262 272473
rect 378754 271603 379262 271631
rect 378658 271159 379358 271187
rect 378658 271057 378686 271159
rect 378646 271051 378698 271057
rect 378646 270993 378698 270999
rect 378742 271051 378794 271057
rect 378742 270993 378794 270999
rect 378754 270965 378782 270993
rect 378562 270937 378782 270965
rect 377890 270160 378014 270188
rect 377878 268461 377930 268467
rect 377986 268449 378014 270160
rect 379126 270015 379178 270021
rect 379126 269957 379178 269963
rect 379222 270015 379274 270021
rect 379222 269957 379274 269963
rect 379138 269725 379166 269957
rect 379030 269719 379082 269725
rect 379030 269661 379082 269667
rect 379126 269719 379178 269725
rect 379126 269661 379178 269667
rect 379042 269577 379070 269661
rect 378934 269571 378986 269577
rect 378934 269513 378986 269519
rect 379030 269571 379082 269577
rect 379030 269513 379082 269519
rect 378454 268979 378506 268985
rect 378506 268939 378782 268967
rect 378454 268921 378506 268927
rect 378646 268905 378698 268911
rect 378646 268847 378698 268853
rect 378754 268856 378782 268939
rect 378550 268831 378602 268837
rect 378550 268773 378602 268779
rect 378358 268683 378410 268689
rect 378358 268625 378410 268631
rect 378370 268597 378398 268625
rect 378562 268615 378590 268773
rect 378550 268609 378602 268615
rect 378370 268569 378494 268597
rect 377986 268421 378110 268449
rect 377878 268403 377930 268409
rect 377890 267949 377918 268403
rect 377878 267943 377930 267949
rect 377878 267885 377930 267891
rect 377974 267869 378026 267875
rect 377972 267834 377974 267843
rect 378026 267834 378028 267843
rect 377972 267769 378028 267778
rect 378082 265156 378110 268421
rect 378164 268426 378220 268435
rect 378164 268361 378220 268370
rect 377568 265128 377822 265156
rect 377904 265128 378110 265156
rect 378178 265156 378206 268361
rect 378262 267943 378314 267949
rect 378262 267885 378314 267891
rect 378274 265785 378302 267885
rect 378358 267869 378410 267875
rect 378358 267811 378410 267817
rect 378370 267653 378398 267811
rect 378358 267647 378410 267653
rect 378358 267589 378410 267595
rect 378466 267357 378494 268569
rect 378550 268551 378602 268557
rect 378658 268541 378686 268847
rect 378754 268828 378878 268856
rect 378742 268757 378794 268763
rect 378742 268699 378794 268705
rect 378646 268535 378698 268541
rect 378646 268477 378698 268483
rect 378550 267943 378602 267949
rect 378550 267885 378602 267891
rect 378358 267351 378410 267357
rect 378358 267293 378410 267299
rect 378454 267351 378506 267357
rect 378454 267293 378506 267299
rect 378370 267228 378398 267293
rect 378562 267228 378590 267885
rect 378754 267843 378782 268699
rect 378850 268541 378878 268828
rect 378838 268535 378890 268541
rect 378838 268477 378890 268483
rect 378946 268467 378974 269513
rect 379234 269175 379262 269957
rect 379220 269166 379276 269175
rect 379220 269101 379276 269110
rect 378934 268461 378986 268467
rect 378934 268403 378986 268409
rect 379330 267843 379358 271159
rect 378740 267834 378796 267843
rect 378740 267769 378796 267778
rect 379316 267834 379372 267843
rect 379316 267769 379372 267778
rect 378838 267721 378890 267727
rect 378838 267663 378890 267669
rect 378370 267200 378590 267228
rect 378850 267061 378878 267663
rect 378838 267055 378890 267061
rect 378838 266997 378890 267003
rect 378934 267055 378986 267061
rect 378934 266997 378986 267003
rect 378946 266044 378974 266997
rect 378370 266016 378974 266044
rect 378370 265951 378398 266016
rect 378358 265945 378410 265951
rect 378358 265887 378410 265893
rect 378454 265945 378506 265951
rect 378454 265887 378506 265893
rect 378466 265785 378494 265887
rect 378274 265757 378494 265785
rect 378742 265797 378794 265803
rect 378742 265739 378794 265745
rect 378838 265797 378890 265803
rect 378838 265739 378890 265745
rect 378754 265359 378782 265739
rect 378742 265353 378794 265359
rect 378742 265295 378794 265301
rect 378178 265128 378384 265156
rect 378850 265142 378878 265739
rect 379126 265501 379178 265507
rect 378946 265449 379126 265452
rect 378946 265443 379178 265449
rect 378946 265433 379166 265443
rect 378934 265427 379166 265433
rect 378986 265424 379166 265427
rect 378934 265369 378986 265375
rect 379522 265156 379550 275285
rect 379618 272579 379646 276783
rect 383350 276765 383402 276771
rect 383734 276823 383786 276829
rect 383734 276765 383786 276771
rect 379798 276601 379850 276607
rect 379798 276543 379850 276549
rect 379604 272570 379660 272579
rect 379604 272505 379660 272514
rect 379810 265156 379838 276543
rect 380470 276379 380522 276385
rect 380470 276321 380522 276327
rect 380566 276379 380618 276385
rect 380566 276321 380618 276327
rect 379990 276305 380042 276311
rect 379990 276247 380042 276253
rect 380002 275127 380030 276247
rect 380482 275719 380510 276321
rect 380278 275713 380330 275719
rect 380278 275655 380330 275661
rect 380470 275713 380522 275719
rect 380470 275655 380522 275661
rect 379990 275121 380042 275127
rect 379990 275063 380042 275069
rect 380086 275121 380138 275127
rect 380086 275063 380138 275069
rect 379988 274938 380044 274947
rect 380098 274924 380126 275063
rect 380044 274896 380126 274924
rect 380180 274938 380236 274947
rect 379988 274873 380044 274882
rect 380180 274873 380236 274882
rect 380194 274239 380222 274873
rect 380290 274239 380318 275655
rect 380578 275127 380606 276321
rect 380566 275121 380618 275127
rect 380566 275063 380618 275069
rect 381430 275121 381482 275127
rect 381430 275063 381482 275069
rect 380182 274233 380234 274239
rect 380182 274175 380234 274181
rect 380278 274233 380330 274239
rect 380278 274175 380330 274181
rect 380278 273567 380330 273573
rect 380278 273509 380330 273515
rect 380374 273567 380426 273573
rect 380374 273509 380426 273515
rect 380290 273023 380318 273509
rect 380084 273014 380140 273023
rect 380084 272949 380140 272958
rect 380276 273014 380332 273023
rect 380276 272949 380332 272958
rect 380098 272704 380126 272949
rect 380386 272907 380414 273509
rect 380482 272972 381278 273000
rect 380374 272901 380426 272907
rect 380374 272843 380426 272849
rect 380482 272704 380510 272972
rect 380566 272901 380618 272907
rect 380566 272843 380618 272849
rect 381140 272866 381196 272875
rect 380098 272676 380510 272704
rect 380180 272570 380236 272579
rect 380180 272505 380236 272514
rect 380194 271427 380222 272505
rect 380276 272126 380332 272135
rect 380276 272061 380332 272070
rect 380182 271421 380234 271427
rect 380182 271363 380234 271369
rect 380290 270909 380318 272061
rect 380374 271421 380426 271427
rect 380374 271363 380426 271369
rect 380278 270903 380330 270909
rect 380278 270845 380330 270851
rect 380386 270835 380414 271363
rect 380374 270829 380426 270835
rect 380374 270771 380426 270777
rect 380084 269166 380140 269175
rect 380084 269101 380140 269110
rect 379296 265128 379550 265156
rect 379680 265128 379838 265156
rect 380098 265142 380126 269101
rect 380578 265142 380606 272843
rect 381250 272852 381278 272972
rect 381332 272866 381388 272875
rect 381250 272824 381332 272852
rect 381140 272801 381196 272810
rect 381332 272801 381388 272810
rect 380950 270903 381002 270909
rect 380950 270845 381002 270851
rect 380962 265142 380990 270845
rect 381154 265156 381182 272801
rect 381442 270909 381470 275063
rect 382964 274050 383020 274059
rect 383156 274050 383212 274059
rect 383074 274017 383156 274036
rect 382964 273985 383020 273994
rect 383062 274011 383156 274017
rect 382978 273615 383006 273985
rect 383114 274008 383156 274011
rect 383156 273985 383212 273994
rect 383062 273953 383114 273959
rect 382772 273606 382828 273615
rect 382772 273541 382828 273550
rect 382964 273606 383020 273615
rect 382964 273541 383020 273550
rect 382786 273444 382814 273541
rect 382786 273416 383102 273444
rect 383074 272875 383102 273416
rect 383060 272866 383116 272875
rect 383060 272801 383116 272810
rect 382292 272718 382348 272727
rect 382292 272653 382348 272662
rect 381812 272274 381868 272283
rect 381812 272209 381868 272218
rect 381826 271987 381854 272209
rect 381620 271978 381676 271987
rect 381620 271913 381676 271922
rect 381812 271978 381868 271987
rect 381812 271913 381868 271922
rect 381430 270903 381482 270909
rect 381430 270845 381482 270851
rect 381634 265156 381662 271913
rect 381154 265128 381408 265156
rect 381634 265128 381888 265156
rect 382306 265142 382334 272653
rect 383060 272274 383116 272283
rect 383060 272209 383116 272218
rect 383074 272167 383102 272209
rect 383062 272161 383114 272167
rect 383254 272161 383306 272167
rect 383062 272103 383114 272109
rect 383170 272121 383254 272149
rect 382966 272087 383018 272093
rect 383170 272075 383198 272121
rect 383254 272103 383306 272109
rect 383350 272087 383402 272093
rect 383018 272047 383198 272075
rect 383266 272047 383350 272075
rect 382966 272029 383018 272035
rect 383266 271945 383294 272047
rect 383350 272029 383402 272035
rect 383254 271939 383306 271945
rect 383446 271939 383498 271945
rect 383254 271881 383306 271887
rect 383362 271899 383446 271927
rect 383362 271871 383390 271899
rect 383446 271881 383498 271887
rect 383350 271865 383402 271871
rect 383350 271807 383402 271813
rect 383746 271797 383774 276765
rect 383828 273310 383884 273319
rect 383828 273245 383884 273254
rect 383734 271791 383786 271797
rect 383734 271733 383786 271739
rect 382966 271717 383018 271723
rect 383254 271717 383306 271723
rect 383018 271677 383254 271705
rect 382966 271659 383018 271665
rect 383254 271659 383306 271665
rect 383062 271643 383114 271649
rect 383062 271585 383114 271591
rect 383074 270909 383102 271585
rect 383446 271421 383498 271427
rect 383446 271363 383498 271369
rect 383158 271347 383210 271353
rect 383158 271289 383210 271295
rect 383062 270903 383114 270909
rect 383062 270845 383114 270851
rect 383170 270835 383198 271289
rect 383458 271224 383486 271363
rect 383362 271196 383486 271224
rect 383158 270829 383210 270835
rect 383158 270771 383210 270777
rect 383362 265156 383390 271196
rect 383444 267834 383500 267843
rect 383444 267769 383500 267778
rect 383184 265128 383390 265156
rect 365760 264999 366026 265005
rect 348598 264983 348650 264989
rect 348598 264925 348650 264931
rect 365206 264983 365258 264989
rect 365760 264980 366014 264999
rect 369264 264980 369566 265008
rect 376726 265057 376778 265063
rect 377206 265057 377258 265063
rect 376726 264999 376778 265005
rect 377088 265005 377206 265008
rect 377088 264999 377258 265005
rect 377088 264980 377246 264999
rect 382402 264980 382704 265008
rect 365206 264925 365258 264931
rect 382402 264915 382430 264980
rect 383458 264915 383486 267769
rect 383842 265156 383870 273245
rect 383616 265128 383870 265156
rect 384034 265156 384062 278573
rect 396266 278596 396528 278599
rect 403318 278599 403632 278605
rect 396214 278541 396266 278547
rect 403370 278596 403632 278599
rect 403318 278541 403370 278547
rect 387766 278525 387818 278531
rect 387766 278467 387818 278473
rect 388342 278525 388394 278531
rect 490198 278525 490250 278531
rect 388342 278467 388394 278473
rect 385078 278303 385130 278309
rect 385078 278245 385130 278251
rect 384610 274831 384638 277870
rect 385090 276385 385118 278245
rect 385474 277856 385776 277884
rect 385078 276379 385130 276385
rect 385078 276321 385130 276327
rect 384886 276305 384938 276311
rect 384886 276247 384938 276253
rect 384898 276015 384926 276247
rect 384790 276009 384842 276015
rect 384790 275951 384842 275957
rect 384886 276009 384938 276015
rect 384886 275951 384938 275957
rect 384802 274979 384830 275951
rect 384694 274973 384746 274979
rect 384694 274915 384746 274921
rect 384790 274973 384842 274979
rect 384790 274915 384842 274921
rect 384706 274831 384734 274915
rect 384598 274825 384650 274831
rect 384598 274767 384650 274773
rect 384694 274825 384746 274831
rect 384694 274767 384746 274773
rect 384884 272866 384940 272875
rect 384884 272801 384940 272810
rect 384116 272422 384172 272431
rect 384116 272357 384172 272366
rect 384130 271427 384158 272357
rect 384404 271978 384460 271987
rect 384404 271913 384460 271922
rect 384118 271421 384170 271427
rect 384118 271363 384170 271369
rect 384214 271421 384266 271427
rect 384214 271363 384266 271369
rect 384226 271057 384254 271363
rect 384214 271051 384266 271057
rect 384214 270993 384266 270999
rect 384034 265128 384096 265156
rect 384418 265142 384446 271913
rect 384898 265142 384926 272801
rect 385364 272718 385420 272727
rect 385364 272653 385420 272662
rect 385270 272235 385322 272241
rect 385270 272177 385322 272183
rect 385282 271945 385310 272177
rect 385270 271939 385322 271945
rect 385270 271881 385322 271887
rect 385378 265142 385406 272653
rect 385474 267949 385502 277856
rect 387010 277125 387038 277870
rect 386998 277119 387050 277125
rect 386998 277061 387050 277067
rect 387778 276256 387806 278467
rect 387874 277856 388176 277884
rect 387874 276575 387902 277856
rect 387860 276566 387916 276575
rect 387860 276501 387916 276510
rect 387778 276228 387902 276256
rect 385558 274381 385610 274387
rect 385558 274323 385610 274329
rect 385846 274381 385898 274387
rect 385846 274323 385898 274329
rect 385570 272241 385598 274323
rect 385750 274085 385802 274091
rect 385750 274027 385802 274033
rect 385558 272235 385610 272241
rect 385558 272177 385610 272183
rect 385654 271051 385706 271057
rect 385654 270993 385706 270999
rect 385558 268979 385610 268985
rect 385558 268921 385610 268927
rect 385570 267949 385598 268921
rect 385462 267943 385514 267949
rect 385462 267885 385514 267891
rect 385558 267943 385610 267949
rect 385558 267885 385610 267891
rect 385666 264989 385694 270993
rect 385762 265304 385790 274027
rect 385858 267357 385886 274323
rect 385940 272866 385996 272875
rect 385940 272801 385996 272810
rect 386612 272866 386668 272875
rect 386612 272801 386668 272810
rect 385846 267351 385898 267357
rect 385846 267293 385898 267299
rect 385762 265276 385886 265304
rect 385858 265156 385886 265276
rect 385824 265128 385886 265156
rect 385954 265156 385982 272801
rect 386324 271978 386380 271987
rect 386324 271913 386380 271922
rect 386338 270835 386366 271913
rect 386326 270829 386378 270835
rect 386326 270771 386378 270777
rect 385954 265128 386208 265156
rect 386626 265142 386654 272801
rect 386806 272235 386858 272241
rect 386806 272177 386858 272183
rect 386818 265156 386846 272177
rect 387478 271939 387530 271945
rect 387478 271881 387530 271887
rect 387490 270835 387518 271881
rect 387764 271238 387820 271247
rect 387764 271173 387820 271182
rect 387478 270829 387530 270835
rect 386914 270752 387422 270780
rect 387478 270771 387530 270777
rect 386914 270021 386942 270752
rect 387394 270613 387422 270752
rect 387286 270607 387338 270613
rect 387286 270549 387338 270555
rect 387382 270607 387434 270613
rect 387382 270549 387434 270555
rect 387190 270311 387242 270317
rect 387190 270253 387242 270259
rect 387094 270237 387146 270243
rect 387094 270179 387146 270185
rect 386998 270089 387050 270095
rect 386998 270031 387050 270037
rect 386902 270015 386954 270021
rect 386902 269957 386954 269963
rect 387010 268985 387038 270031
rect 387106 270021 387134 270179
rect 387202 270095 387230 270253
rect 387298 270243 387326 270549
rect 387382 270311 387434 270317
rect 387382 270253 387434 270259
rect 387286 270237 387338 270243
rect 387286 270179 387338 270185
rect 387190 270089 387242 270095
rect 387190 270031 387242 270037
rect 387094 270015 387146 270021
rect 387094 269957 387146 269963
rect 386998 268979 387050 268985
rect 386998 268921 387050 268927
rect 387394 268597 387422 270253
rect 387298 268569 387422 268597
rect 387298 268541 387326 268569
rect 387286 268535 387338 268541
rect 387286 268477 387338 268483
rect 387478 267351 387530 267357
rect 387478 267293 387530 267299
rect 387490 267209 387518 267293
rect 387478 267203 387530 267209
rect 387478 267145 387530 267151
rect 387574 267203 387626 267209
rect 387574 267145 387626 267151
rect 387190 265501 387242 265507
rect 387190 265443 387242 265449
rect 387202 265415 387230 265443
rect 387586 265415 387614 267145
rect 387202 265387 387614 265415
rect 387778 265156 387806 271173
rect 387874 265452 387902 276228
rect 388354 273319 388382 278467
rect 393826 278457 394128 278476
rect 598484 278490 598540 278499
rect 490250 278473 490512 278476
rect 490198 278467 490512 278473
rect 393814 278451 394128 278457
rect 393866 278448 394128 278451
rect 490210 278448 490512 278467
rect 598540 278448 598800 278476
rect 598484 278425 598540 278434
rect 393814 278393 393866 278399
rect 389014 278377 389066 278383
rect 467540 278342 467596 278351
rect 389066 278325 389328 278328
rect 389014 278319 389328 278325
rect 389026 278300 389328 278319
rect 467596 278300 467856 278328
rect 467540 278277 467596 278286
rect 453238 278229 453290 278235
rect 474740 278194 474796 278203
rect 453290 278177 453552 278180
rect 453238 278171 453552 278177
rect 453250 278152 453552 278171
rect 474796 278152 475056 278180
rect 635266 278161 635568 278180
rect 635254 278155 635568 278161
rect 474740 278129 474796 278138
rect 635306 278152 635568 278155
rect 635254 278097 635306 278103
rect 417622 278081 417674 278087
rect 415330 278013 415632 278032
rect 488948 278046 489004 278055
rect 417674 278029 417936 278032
rect 417622 278023 417936 278029
rect 415318 278007 415632 278013
rect 415370 278004 415632 278007
rect 417634 278004 417936 278023
rect 489004 278004 489264 278032
rect 488948 277981 489004 277990
rect 415318 277949 415370 277955
rect 422326 277933 422378 277939
rect 388438 277119 388490 277125
rect 388438 277061 388490 277067
rect 388340 273310 388396 273319
rect 388340 273245 388396 273254
rect 388148 271830 388204 271839
rect 388148 271765 388204 271774
rect 387874 265424 387950 265452
rect 386818 265128 387120 265156
rect 387600 265128 387806 265156
rect 387922 265142 387950 265424
rect 388162 265156 388190 271765
rect 388450 268615 388478 277061
rect 388918 274085 388970 274091
rect 388642 274059 388918 274073
rect 388628 274050 388918 274059
rect 388684 274045 388918 274050
rect 388918 274027 388970 274033
rect 388628 273985 388684 273994
rect 389494 272383 389546 272389
rect 389494 272325 389546 272331
rect 389590 272383 389642 272389
rect 389590 272325 389642 272331
rect 389108 271830 389164 271839
rect 389108 271765 389164 271774
rect 388534 268979 388586 268985
rect 388534 268921 388586 268927
rect 388726 268979 388778 268985
rect 388822 268979 388874 268985
rect 388778 268939 388822 268967
rect 388726 268921 388778 268927
rect 388822 268921 388874 268927
rect 388438 268609 388490 268615
rect 388438 268551 388490 268557
rect 388546 268541 388574 268921
rect 388918 268609 388970 268615
rect 388642 268569 388918 268597
rect 388534 268535 388586 268541
rect 388534 268477 388586 268483
rect 388438 268461 388490 268467
rect 388642 268435 388670 268569
rect 388918 268551 388970 268557
rect 388438 268403 388490 268409
rect 388628 268426 388684 268435
rect 388450 268116 388478 268403
rect 388820 268426 388876 268435
rect 388628 268361 388684 268370
rect 388738 268384 388820 268412
rect 388738 268319 388766 268384
rect 388820 268361 388876 268370
rect 388726 268313 388778 268319
rect 388726 268255 388778 268261
rect 388822 268313 388874 268319
rect 388822 268255 388874 268261
rect 388834 268116 388862 268255
rect 388450 268088 388862 268116
rect 389122 265156 389150 271765
rect 389300 271682 389356 271691
rect 389300 271617 389356 271626
rect 389206 268683 389258 268689
rect 389206 268625 389258 268631
rect 389218 268435 389246 268625
rect 389204 268426 389260 268435
rect 389204 268361 389260 268370
rect 389314 265156 389342 271617
rect 389506 268615 389534 272325
rect 389602 272019 389630 272325
rect 389590 272013 389642 272019
rect 389590 271955 389642 271961
rect 389684 271682 389740 271691
rect 389684 271617 389740 271626
rect 389398 268609 389450 268615
rect 389398 268551 389450 268557
rect 389494 268609 389546 268615
rect 389494 268551 389546 268557
rect 389410 268435 389438 268551
rect 389396 268426 389452 268435
rect 389396 268361 389452 268370
rect 388162 265128 388416 265156
rect 388848 265128 389150 265156
rect 389232 265128 389342 265156
rect 389698 265142 389726 271617
rect 389876 271534 389932 271543
rect 389876 271469 389932 271478
rect 389890 265156 389918 271469
rect 390562 265359 390590 277870
rect 391714 274461 391742 277870
rect 391702 274455 391754 274461
rect 391702 274397 391754 274403
rect 392962 273795 392990 277870
rect 395362 274387 395390 277870
rect 397474 277856 397776 277884
rect 395350 274381 395402 274387
rect 395350 274323 395402 274329
rect 392950 273789 393002 273795
rect 391412 273754 391468 273763
rect 392950 273731 393002 273737
rect 391412 273689 391468 273698
rect 390836 273310 390892 273319
rect 390836 273245 390892 273254
rect 390550 265353 390602 265359
rect 390550 265295 390602 265301
rect 390850 265156 390878 273245
rect 390932 272422 390988 272431
rect 390932 272357 390988 272366
rect 389890 265128 390144 265156
rect 390624 265128 390878 265156
rect 390946 265142 390974 272357
rect 391426 265142 391454 273689
rect 397364 273606 397420 273615
rect 396214 273567 396266 273573
rect 396214 273509 396266 273515
rect 396310 273567 396362 273573
rect 397364 273541 397420 273550
rect 396310 273509 396362 273515
rect 392852 273458 392908 273467
rect 392852 273393 392908 273402
rect 393140 273458 393196 273467
rect 393140 273393 393196 273402
rect 392470 272679 392522 272685
rect 392470 272621 392522 272627
rect 392566 272679 392618 272685
rect 392566 272621 392618 272627
rect 391702 272605 391754 272611
rect 391702 272547 391754 272553
rect 391606 272013 391658 272019
rect 391606 271955 391658 271961
rect 391618 270951 391646 271955
rect 391604 270942 391660 270951
rect 391604 270877 391660 270886
rect 391714 265156 391742 272547
rect 392086 270755 392138 270761
rect 392086 270697 392138 270703
rect 392098 265156 392126 270697
rect 392482 265156 392510 272621
rect 392578 272093 392606 272621
rect 392566 272087 392618 272093
rect 392566 272029 392618 272035
rect 392758 271643 392810 271649
rect 392758 271585 392810 271591
rect 392770 270909 392798 271585
rect 392866 270909 392894 273393
rect 392948 270942 393004 270951
rect 392758 270903 392810 270909
rect 392758 270845 392810 270851
rect 392854 270903 392906 270909
rect 392948 270877 393004 270886
rect 392854 270845 392906 270851
rect 392854 265353 392906 265359
rect 392854 265295 392906 265301
rect 391714 265128 391920 265156
rect 392098 265128 392352 265156
rect 392482 265128 392736 265156
rect 392866 264989 392894 265295
rect 385654 264983 385706 264989
rect 385654 264925 385706 264931
rect 392854 264983 392906 264989
rect 392854 264925 392906 264931
rect 212522 264857 212784 264860
rect 212470 264851 212784 264857
rect 267570 264853 267630 264862
rect 348502 264909 348554 264915
rect 348502 264851 348554 264857
rect 382390 264909 382442 264915
rect 382390 264851 382442 264857
rect 383446 264909 383498 264915
rect 388979 264913 389039 264922
rect 392962 264921 392990 270877
rect 393154 265142 393182 273393
rect 394484 273014 394540 273023
rect 394484 272949 394540 272958
rect 395636 273014 395692 273023
rect 395636 272949 395692 272958
rect 394292 272570 394348 272579
rect 394498 272556 394526 272949
rect 395650 272727 395678 272949
rect 395636 272718 395692 272727
rect 395636 272653 395692 272662
rect 395828 272718 395884 272727
rect 395828 272653 395884 272662
rect 394498 272537 394622 272556
rect 394498 272531 394634 272537
rect 394498 272528 394582 272531
rect 394292 272505 394348 272514
rect 394198 272457 394250 272463
rect 394004 272422 394060 272431
rect 394198 272399 394250 272405
rect 394004 272357 394060 272366
rect 393622 265353 393674 265359
rect 393622 265295 393674 265301
rect 393634 265142 393662 265295
rect 394018 265156 394046 272357
rect 394102 271791 394154 271797
rect 394102 271733 394154 271739
rect 394114 270983 394142 271733
rect 394102 270977 394154 270983
rect 394102 270919 394154 270925
rect 394210 265156 394238 272399
rect 394306 270983 394334 272505
rect 394582 272473 394634 272479
rect 394486 272457 394538 272463
rect 394486 272399 394538 272405
rect 394498 272135 394526 272399
rect 394484 272126 394540 272135
rect 394484 272061 394540 272070
rect 394390 271939 394442 271945
rect 394390 271881 394442 271887
rect 394294 270977 394346 270983
rect 394294 270919 394346 270925
rect 394402 270803 394430 271881
rect 395156 271534 395212 271543
rect 395156 271469 395212 271478
rect 394484 271090 394540 271099
rect 394484 271025 394540 271034
rect 394388 270794 394444 270803
rect 394498 270761 394526 271025
rect 394388 270729 394444 270738
rect 394486 270755 394538 270761
rect 394486 270697 394538 270703
rect 395170 265156 395198 271469
rect 395350 268609 395402 268615
rect 395350 268551 395402 268557
rect 395446 268609 395498 268615
rect 395446 268551 395498 268557
rect 393334 265131 393386 265137
rect 394018 265128 394128 265156
rect 394210 265128 394464 265156
rect 394944 265128 395198 265156
rect 395362 265142 395390 268551
rect 395458 267991 395486 268551
rect 395444 267982 395500 267991
rect 395444 267917 395500 267926
rect 395842 265142 395870 272653
rect 396226 265142 396254 273509
rect 396322 271987 396350 273509
rect 396982 272975 397034 272981
rect 396982 272917 397034 272923
rect 396790 272605 396842 272611
rect 396790 272547 396842 272553
rect 396406 272161 396458 272167
rect 396406 272103 396458 272109
rect 396308 271978 396364 271987
rect 396308 271913 396364 271922
rect 396418 271927 396446 272103
rect 396802 272019 396830 272547
rect 396790 272013 396842 272019
rect 396790 271955 396842 271961
rect 396694 271939 396746 271945
rect 396418 271899 396694 271927
rect 396694 271881 396746 271887
rect 396884 271238 396940 271247
rect 396884 271173 396940 271182
rect 396898 265156 396926 271173
rect 396672 265128 396926 265156
rect 393334 265073 393386 265079
rect 393346 264989 393374 265073
rect 396994 264989 397022 272917
rect 397078 272827 397130 272833
rect 397078 272769 397130 272775
rect 397090 265156 397118 272769
rect 397378 272611 397406 273541
rect 397366 272605 397418 272611
rect 397366 272547 397418 272553
rect 397270 267869 397322 267875
rect 397270 267811 397322 267817
rect 397282 266987 397310 267811
rect 397474 267653 397502 277856
rect 398914 274535 398942 277870
rect 398902 274529 398954 274535
rect 398902 274471 398954 274477
rect 399670 273049 399722 273055
rect 399670 272991 399722 272997
rect 398326 272753 398378 272759
rect 398326 272695 398378 272701
rect 397748 271090 397804 271099
rect 397748 271025 397804 271034
rect 397556 267982 397612 267991
rect 397556 267917 397558 267926
rect 397610 267917 397612 267926
rect 397558 267885 397610 267891
rect 397462 267647 397514 267653
rect 397462 267589 397514 267595
rect 397558 267647 397610 267653
rect 397558 267589 397610 267595
rect 397570 267505 397598 267589
rect 397558 267499 397610 267505
rect 397558 267441 397610 267447
rect 397654 267499 397706 267505
rect 397654 267441 397706 267447
rect 397666 267228 397694 267441
rect 397378 267200 397694 267228
rect 397174 266981 397226 266987
rect 397174 266923 397226 266929
rect 397270 266981 397322 266987
rect 397270 266923 397322 266929
rect 397186 266784 397214 266923
rect 397378 266784 397406 267200
rect 397186 266756 397406 266784
rect 397762 265156 397790 271025
rect 397844 267834 397900 267843
rect 397844 267769 397900 267778
rect 397858 265951 397886 267769
rect 398230 267055 398282 267061
rect 398230 266997 398282 267003
rect 398242 265951 398270 266997
rect 397846 265945 397898 265951
rect 397846 265887 397898 265893
rect 398230 265945 398282 265951
rect 398230 265887 398282 265893
rect 398338 265156 398366 272695
rect 398420 272422 398476 272431
rect 398420 272357 398476 272366
rect 397090 265128 397152 265156
rect 397488 265128 397790 265156
rect 397968 265128 398366 265156
rect 398434 265142 398462 272357
rect 398998 271125 399050 271131
rect 398818 271073 398998 271076
rect 398818 271067 399050 271073
rect 398818 271057 399038 271067
rect 398806 271051 399038 271057
rect 398858 271048 399038 271051
rect 398806 270993 398858 270999
rect 399476 270942 399532 270951
rect 399476 270877 399532 270886
rect 399286 268535 399338 268541
rect 399286 268477 399338 268483
rect 398818 267644 399134 267672
rect 398818 267505 398846 267644
rect 398806 267499 398858 267505
rect 398806 267441 398858 267447
rect 398902 267499 398954 267505
rect 398902 267441 398954 267447
rect 398518 267203 398570 267209
rect 398518 267145 398570 267151
rect 398806 267203 398858 267209
rect 398806 267145 398858 267151
rect 398530 266987 398558 267145
rect 398518 266981 398570 266987
rect 398518 266923 398570 266929
rect 398818 266765 398846 267145
rect 398914 266839 398942 267441
rect 399106 266839 399134 267644
rect 399190 266981 399242 266987
rect 399190 266923 399242 266929
rect 398902 266833 398954 266839
rect 398902 266775 398954 266781
rect 399094 266833 399146 266839
rect 399094 266775 399146 266781
rect 398806 266759 398858 266765
rect 398806 266701 398858 266707
rect 399202 265803 399230 266923
rect 399298 266765 399326 268477
rect 399286 266759 399338 266765
rect 399286 266701 399338 266707
rect 399094 265797 399146 265803
rect 399094 265739 399146 265745
rect 399190 265797 399242 265803
rect 399190 265739 399242 265745
rect 398710 265353 398762 265359
rect 398530 265313 398710 265341
rect 398530 265211 398558 265313
rect 398710 265295 398762 265301
rect 398998 265279 399050 265285
rect 398998 265221 399050 265227
rect 398518 265205 398570 265211
rect 398518 265147 398570 265153
rect 399010 265063 399038 265221
rect 399106 265063 399134 265739
rect 399490 265156 399518 270877
rect 399574 268609 399626 268615
rect 399574 268551 399626 268557
rect 399264 265128 399518 265156
rect 398998 265057 399050 265063
rect 398626 264989 398880 265008
rect 398998 264999 399050 265005
rect 399094 265057 399146 265063
rect 399094 264999 399146 265005
rect 399586 264989 399614 268551
rect 399682 265142 399710 272991
rect 400066 267727 400094 277870
rect 401218 276533 401246 277870
rect 402466 277125 402494 277870
rect 404674 277856 404784 277884
rect 402454 277119 402506 277125
rect 402454 277061 402506 277067
rect 401206 276527 401258 276533
rect 401206 276469 401258 276475
rect 404086 273345 404138 273351
rect 404086 273287 404138 273293
rect 401302 273271 401354 273277
rect 401302 273213 401354 273219
rect 400630 273123 400682 273129
rect 400630 273065 400682 273071
rect 400148 272274 400204 272283
rect 400148 272209 400204 272218
rect 400054 267721 400106 267727
rect 400054 267663 400106 267669
rect 399862 265427 399914 265433
rect 399862 265369 399914 265375
rect 399874 265211 399902 265369
rect 399862 265205 399914 265211
rect 399862 265147 399914 265153
rect 400162 265142 400190 272209
rect 400642 265142 400670 273065
rect 401204 270794 401260 270803
rect 401204 270729 401260 270738
rect 401218 265156 401246 270729
rect 400992 265128 401246 265156
rect 401314 265156 401342 273213
rect 403222 273197 403274 273203
rect 403222 273139 403274 273145
rect 402740 272126 402796 272135
rect 402740 272061 402796 272070
rect 401876 271978 401932 271987
rect 401876 271913 401932 271922
rect 401684 267982 401740 267991
rect 401684 267917 401740 267926
rect 401698 267727 401726 267917
rect 401686 267721 401738 267727
rect 401686 267663 401738 267669
rect 401314 265128 401472 265156
rect 401890 265142 401918 271913
rect 402358 271051 402410 271057
rect 402358 270993 402410 270999
rect 402370 265142 402398 270993
rect 402754 265142 402782 272061
rect 402838 270977 402890 270983
rect 402934 270977 402986 270983
rect 402890 270937 402934 270965
rect 402838 270919 402890 270925
rect 402934 270919 402986 270925
rect 403234 265156 403262 273139
rect 403702 268535 403754 268541
rect 403702 268477 403754 268483
rect 403714 268435 403742 268477
rect 403700 268426 403756 268435
rect 403700 268361 403756 268370
rect 403892 268426 403948 268435
rect 403892 268361 403948 268370
rect 403906 265156 403934 268361
rect 403200 265128 403262 265156
rect 403680 265128 403934 265156
rect 404098 265142 404126 273287
rect 404674 267653 404702 277856
rect 406018 274609 406046 277870
rect 406006 274603 406058 274609
rect 406006 274545 406058 274551
rect 404950 273419 405002 273425
rect 404950 273361 405002 273367
rect 404756 267982 404812 267991
rect 404756 267917 404812 267926
rect 404662 267647 404714 267653
rect 404662 267589 404714 267595
rect 404770 265156 404798 267917
rect 404496 265128 404798 265156
rect 404962 265142 404990 273361
rect 406676 271978 406732 271987
rect 405718 271939 405770 271945
rect 406676 271913 406732 271922
rect 405718 271881 405770 271887
rect 405620 267982 405676 267991
rect 405620 267917 405676 267926
rect 405634 265156 405662 267917
rect 405730 265452 405758 271881
rect 406582 271791 406634 271797
rect 406582 271733 406634 271739
rect 406102 268535 406154 268541
rect 406102 268477 406154 268483
rect 406114 268435 406142 268477
rect 406100 268426 406156 268435
rect 406100 268361 406156 268370
rect 405730 265424 405806 265452
rect 405408 265128 405662 265156
rect 405778 265142 405806 265424
rect 406486 265205 406538 265211
rect 406272 265153 406486 265156
rect 406272 265147 406538 265153
rect 406594 265156 406622 271733
rect 406690 271247 406718 271913
rect 406676 271238 406732 271247
rect 406676 271173 406732 271182
rect 407170 266839 407198 277870
rect 407254 272679 407306 272685
rect 407254 272621 407306 272627
rect 407158 266833 407210 266839
rect 407158 266775 407210 266781
rect 407266 265156 407294 272621
rect 408130 272537 408350 272556
rect 408118 272531 408350 272537
rect 408170 272528 408350 272531
rect 408118 272473 408170 272479
rect 408322 272389 408350 272528
rect 408214 272383 408266 272389
rect 408214 272325 408266 272331
rect 408310 272383 408362 272389
rect 408310 272325 408362 272331
rect 408118 265205 408170 265211
rect 406272 265128 406526 265147
rect 406594 265128 406704 265156
rect 407266 265128 407568 265156
rect 408118 265147 408170 265153
rect 408226 265156 408254 272325
rect 408418 267875 408446 277870
rect 409270 271717 409322 271723
rect 409270 271659 409322 271665
rect 408980 270794 409036 270803
rect 408980 270729 409036 270738
rect 408994 270063 409022 270729
rect 408980 270054 409036 270063
rect 408980 269989 409036 269998
rect 408596 267982 408652 267991
rect 408596 267917 408652 267926
rect 408788 267982 408844 267991
rect 408788 267917 408790 267926
rect 408406 267869 408458 267875
rect 408406 267811 408458 267817
rect 408610 265156 408638 267917
rect 408842 267917 408844 267926
rect 408790 267885 408842 267891
rect 408788 267834 408844 267843
rect 408788 267769 408844 267778
rect 408802 266765 408830 267769
rect 408790 266759 408842 266765
rect 408790 266701 408842 266707
rect 393334 264983 393386 264989
rect 393334 264925 393386 264931
rect 396982 264983 397034 264989
rect 396982 264925 397034 264931
rect 398614 264983 398880 264989
rect 398666 264980 398880 264983
rect 399574 264983 399626 264989
rect 398614 264925 398666 264931
rect 408130 264942 408158 265147
rect 408226 265128 408480 265156
rect 408610 265128 408912 265156
rect 409282 265142 409310 271659
rect 409570 269059 409598 277870
rect 410818 277643 410846 277870
rect 410806 277637 410858 277643
rect 410806 277579 410858 277585
rect 411970 273647 411998 277870
rect 412258 277856 413232 277884
rect 481844 277898 481900 277907
rect 422378 277881 422640 277884
rect 422326 277875 422640 277881
rect 411958 273641 412010 273647
rect 411958 273583 412010 273589
rect 409942 271643 409994 271649
rect 409942 271585 409994 271591
rect 409558 269053 409610 269059
rect 409558 268995 409610 269001
rect 409954 265156 409982 271585
rect 410998 271569 411050 271575
rect 410998 271511 411050 271517
rect 409954 265128 410208 265156
rect 411010 265142 411038 271511
rect 411958 271495 412010 271501
rect 411958 271437 412010 271443
rect 411766 265205 411818 265211
rect 411504 265153 411766 265156
rect 411504 265147 411818 265153
rect 411504 265128 411806 265147
rect 411970 265142 411998 271437
rect 412054 265205 412106 265211
rect 412054 265147 412106 265153
rect 399574 264925 399626 264931
rect 388977 264857 388979 264909
rect 389039 264857 389041 264909
rect 392962 264899 393023 264921
rect 383446 264851 383498 264857
rect 392962 264855 393014 264899
rect 212482 264832 212784 264851
rect 388979 264844 389039 264853
rect 393005 264839 393014 264855
rect 393074 264839 393083 264899
rect 407094 264880 407103 264940
rect 407163 264938 407172 264940
rect 407163 264882 407202 264938
rect 407697 264918 407706 264934
rect 407694 264890 407706 264918
rect 407163 264880 407172 264882
rect 407697 264874 407706 264890
rect 407766 264918 407775 264934
rect 408114 264933 408174 264942
rect 409948 264937 410009 264939
rect 407766 264890 408013 264918
rect 407766 264874 407775 264890
rect 409739 264921 410009 264937
rect 409739 264909 409996 264921
rect 409948 264877 409996 264909
rect 408114 264864 408174 264873
rect 409987 264861 409996 264877
rect 410056 264861 410065 264921
rect 410524 264881 410533 264941
rect 410593 264927 410602 264941
rect 410593 264895 410697 264927
rect 410593 264881 410602 264895
rect 412066 264587 412094 265147
rect 412052 264578 412108 264587
rect 412052 264513 412108 264522
rect 212194 257876 212318 257904
rect 212098 257728 212222 257756
rect 212086 257657 212138 257663
rect 212086 257599 212138 257605
rect 211988 255402 212044 255411
rect 211988 255337 212044 255346
rect 211894 246705 211946 246711
rect 211894 246647 211946 246653
rect 211702 246483 211754 246489
rect 211702 246425 211754 246431
rect 212002 246193 212030 255337
rect 212098 246415 212126 257599
rect 212194 246563 212222 257728
rect 212290 246785 212318 257876
rect 216444 253065 216472 255902
rect 412148 247558 412204 247567
rect 412258 247544 412286 277856
rect 412916 267834 412972 267843
rect 412916 267769 412972 267778
rect 412822 267721 412874 267727
rect 412822 267663 412874 267669
rect 412834 265327 412862 267663
rect 412930 265475 412958 267769
rect 414370 267505 414398 277870
rect 416674 269133 416702 277870
rect 418964 270350 419020 270359
rect 418964 270285 419020 270294
rect 416662 269127 416714 269133
rect 416662 269069 416714 269075
rect 416278 269053 416330 269059
rect 416278 268995 416330 269001
rect 416290 268837 416318 268995
rect 416278 268831 416330 268837
rect 416278 268773 416330 268779
rect 415126 268683 415178 268689
rect 415126 268625 415178 268631
rect 415138 267695 415166 268625
rect 418978 267991 419006 270285
rect 418964 267982 419020 267991
rect 418964 267917 419020 267926
rect 414932 267686 414988 267695
rect 414932 267621 414988 267630
rect 415124 267686 415180 267695
rect 415124 267621 415180 267630
rect 414358 267499 414410 267505
rect 414358 267441 414410 267447
rect 413686 266981 413738 266987
rect 413686 266923 413738 266929
rect 413698 266215 413726 266923
rect 413684 266206 413740 266215
rect 413684 266141 413740 266150
rect 414946 265919 414974 267621
rect 419074 267579 419102 277870
rect 420226 274757 420254 277870
rect 420214 274751 420266 274757
rect 420214 274693 420266 274699
rect 419156 270794 419212 270803
rect 419156 270729 419212 270738
rect 419170 270359 419198 270729
rect 419156 270350 419212 270359
rect 419156 270285 419212 270294
rect 419062 267573 419114 267579
rect 419062 267515 419114 267521
rect 421474 267209 421502 277870
rect 422338 277856 422640 277875
rect 421846 271495 421898 271501
rect 421846 271437 421898 271443
rect 421858 271279 421886 271437
rect 421846 271273 421898 271279
rect 421846 271215 421898 271221
rect 423874 269207 423902 277870
rect 425026 277421 425054 277870
rect 425014 277415 425066 277421
rect 425014 277357 425066 277363
rect 423862 269201 423914 269207
rect 423862 269143 423914 269149
rect 426274 268097 426302 277870
rect 427426 274905 427454 277870
rect 427414 274899 427466 274905
rect 427414 274841 427466 274847
rect 428182 271051 428234 271057
rect 428182 270993 428234 270999
rect 428194 270951 428222 270993
rect 428180 270942 428236 270951
rect 428180 270877 428236 270886
rect 426262 268091 426314 268097
rect 426262 268033 426314 268039
rect 421462 267203 421514 267209
rect 421462 267145 421514 267151
rect 428674 266691 428702 277870
rect 429826 273721 429854 277870
rect 429814 273715 429866 273721
rect 429814 273657 429866 273663
rect 428962 270752 429278 270780
rect 428962 270211 428990 270752
rect 429250 270211 429278 270752
rect 431074 270687 431102 277870
rect 432226 277273 432254 277870
rect 432214 277267 432266 277273
rect 432214 277209 432266 277215
rect 431926 271495 431978 271501
rect 431926 271437 431978 271443
rect 431938 271279 431966 271437
rect 431926 271273 431978 271279
rect 431926 271215 431978 271221
rect 431638 271199 431690 271205
rect 431638 271141 431690 271147
rect 431830 271199 431882 271205
rect 431830 271141 431882 271147
rect 431650 270965 431678 271141
rect 431842 270965 431870 271141
rect 431650 270937 431870 270965
rect 431062 270681 431114 270687
rect 431062 270623 431114 270629
rect 428948 270202 429004 270211
rect 428948 270137 429004 270146
rect 429236 270202 429292 270211
rect 429236 270137 429292 270146
rect 433378 267431 433406 277870
rect 434530 276459 434558 277870
rect 434518 276453 434570 276459
rect 434518 276395 434570 276401
rect 433366 267425 433418 267431
rect 433366 267367 433418 267373
rect 428662 266685 428714 266691
rect 428662 266627 428714 266633
rect 435682 266469 435710 277870
rect 436642 277865 436944 277884
rect 436630 277859 436944 277865
rect 436682 277856 436944 277859
rect 436630 277801 436682 277807
rect 438082 268023 438110 277870
rect 439330 277199 439358 277870
rect 439318 277193 439370 277199
rect 439318 277135 439370 277141
rect 438932 270350 438988 270359
rect 438932 270285 438988 270294
rect 438070 268017 438122 268023
rect 438070 267959 438122 267965
rect 438946 267820 438974 270285
rect 440482 268171 440510 277870
rect 441730 276237 441758 277870
rect 441718 276231 441770 276237
rect 441718 276173 441770 276179
rect 440470 268165 440522 268171
rect 440470 268107 440522 268113
rect 439126 268017 439178 268023
rect 439124 267982 439126 267991
rect 439178 267982 439180 267991
rect 439124 267917 439180 267926
rect 439316 267982 439372 267991
rect 439316 267917 439372 267926
rect 439330 267820 439358 267917
rect 438946 267792 439358 267820
rect 435670 266463 435722 266469
rect 435670 266405 435722 266411
rect 442882 266395 442910 277870
rect 444130 273869 444158 277870
rect 444118 273863 444170 273869
rect 444118 273805 444170 273811
rect 445282 270391 445310 277870
rect 446530 276977 446558 277870
rect 446518 276971 446570 276977
rect 446518 276913 446570 276919
rect 446326 271051 446378 271057
rect 446326 270993 446378 270999
rect 446338 270951 446366 270993
rect 446324 270942 446380 270951
rect 446324 270877 446380 270886
rect 445270 270385 445322 270391
rect 445270 270327 445322 270333
rect 447682 267283 447710 277870
rect 448834 276163 448862 277870
rect 448822 276157 448874 276163
rect 448822 276099 448874 276105
rect 449300 271238 449356 271247
rect 449300 271173 449356 271182
rect 449588 271238 449644 271247
rect 449588 271173 449644 271182
rect 449314 271131 449342 271173
rect 449602 271131 449630 271173
rect 449302 271125 449354 271131
rect 449302 271067 449354 271073
rect 449590 271125 449642 271131
rect 449590 271067 449642 271073
rect 449204 270350 449260 270359
rect 449122 270308 449204 270336
rect 449122 268023 449150 270308
rect 449204 270285 449260 270294
rect 449204 270054 449260 270063
rect 449204 269989 449260 269998
rect 449110 268017 449162 268023
rect 449218 267991 449246 269989
rect 449110 267959 449162 267965
rect 449204 267982 449260 267991
rect 449204 267917 449260 267926
rect 447670 267277 447722 267283
rect 447670 267219 447722 267225
rect 442870 266389 442922 266395
rect 442870 266331 442922 266337
rect 449986 266321 450014 277870
rect 450850 277856 451152 277884
rect 450850 277791 450878 277856
rect 450838 277785 450890 277791
rect 450838 277727 450890 277733
rect 452180 271090 452236 271099
rect 452180 271025 452182 271034
rect 452234 271025 452236 271034
rect 452182 270993 452234 270999
rect 452180 270942 452236 270951
rect 452180 270877 452182 270886
rect 452234 270877 452236 270886
rect 452182 270845 452234 270851
rect 452180 270794 452236 270803
rect 452180 270729 452182 270738
rect 452234 270729 452236 270738
rect 452182 270697 452234 270703
rect 452386 270169 452414 277870
rect 452468 270942 452524 270951
rect 452468 270877 452470 270886
rect 452522 270877 452524 270886
rect 452470 270845 452522 270851
rect 452660 270794 452716 270803
rect 452660 270729 452662 270738
rect 452714 270729 452716 270738
rect 452662 270697 452714 270703
rect 454786 270539 454814 277870
rect 455938 276089 455966 277870
rect 455926 276083 455978 276089
rect 455926 276025 455978 276031
rect 454774 270533 454826 270539
rect 454774 270475 454826 270481
rect 452374 270163 452426 270169
rect 452374 270105 452426 270111
rect 449974 266315 450026 266321
rect 449974 266257 450026 266263
rect 457186 266173 457214 277870
rect 458338 267135 458366 277870
rect 459586 269947 459614 277870
rect 460738 277347 460766 277870
rect 460726 277341 460778 277347
rect 460726 277283 460778 277289
rect 461986 273943 462014 277870
rect 463138 275941 463166 277870
rect 463126 275935 463178 275941
rect 463126 275877 463178 275883
rect 461974 273937 462026 273943
rect 461974 273879 462026 273885
rect 459574 269941 459626 269947
rect 459574 269883 459626 269889
rect 458326 267129 458378 267135
rect 458326 267071 458378 267077
rect 457174 266167 457226 266173
rect 457174 266109 457226 266115
rect 464290 266099 464318 277870
rect 465538 277717 465566 277870
rect 465526 277711 465578 277717
rect 465526 277653 465578 277659
rect 466594 269799 466622 277870
rect 466582 269793 466634 269799
rect 466582 269735 466634 269741
rect 468994 268245 469022 277870
rect 470242 275793 470270 277870
rect 470230 275787 470282 275793
rect 470230 275729 470282 275735
rect 469460 271090 469516 271099
rect 469460 271025 469462 271034
rect 469514 271025 469516 271034
rect 469462 270993 469514 270999
rect 469460 270350 469516 270359
rect 469460 270285 469516 270294
rect 468982 268239 469034 268245
rect 468982 268181 469034 268187
rect 469474 267991 469502 270285
rect 469460 267982 469516 267991
rect 469460 267917 469516 267926
rect 464278 266093 464330 266099
rect 464278 266035 464330 266041
rect 471394 266025 471422 277870
rect 472642 266913 472670 277870
rect 473794 269651 473822 277870
rect 476194 274091 476222 277870
rect 477442 275645 477470 277870
rect 477430 275639 477482 275645
rect 477430 275581 477482 275587
rect 476182 274085 476234 274091
rect 476182 274027 476234 274033
rect 473782 269645 473834 269651
rect 473782 269587 473834 269593
rect 472630 266907 472682 266913
rect 472630 266849 472682 266855
rect 471382 266019 471434 266025
rect 471382 265961 471434 265967
rect 414932 265910 414988 265919
rect 478594 265877 478622 277870
rect 479746 274165 479774 277870
rect 481008 277856 481406 277884
rect 479734 274159 479786 274165
rect 479734 274101 479786 274107
rect 480982 271273 481034 271279
rect 480980 271238 480982 271247
rect 481034 271238 481036 271247
rect 480980 271173 481036 271182
rect 481078 271125 481130 271131
rect 481174 271125 481226 271131
rect 481130 271073 481174 271076
rect 481078 271067 481226 271073
rect 481090 271048 481214 271067
rect 481378 269429 481406 277856
rect 481900 277856 482160 277884
rect 481844 277833 481900 277842
rect 481366 269423 481418 269429
rect 481366 269365 481418 269371
rect 483298 268393 483326 277870
rect 484450 275571 484478 277870
rect 484438 275565 484490 275571
rect 484438 275507 484490 275513
rect 483286 268387 483338 268393
rect 483286 268329 483338 268335
rect 414932 265845 414988 265854
rect 478582 265871 478634 265877
rect 478582 265813 478634 265819
rect 485698 265729 485726 277870
rect 486850 277495 486878 277870
rect 486838 277489 486890 277495
rect 486838 277431 486890 277437
rect 486646 269201 486698 269207
rect 486646 269143 486698 269149
rect 486658 269059 486686 269143
rect 486646 269053 486698 269059
rect 486646 268995 486698 269001
rect 488098 268287 488126 277870
rect 491650 274207 491678 277870
rect 491636 274198 491692 274207
rect 491636 274133 491692 274142
rect 489538 271057 489662 271076
rect 489526 271051 489662 271057
rect 489578 271048 489662 271051
rect 489526 270993 489578 270999
rect 489634 270983 489662 271048
rect 489622 270977 489674 270983
rect 489622 270919 489674 270925
rect 489524 270350 489580 270359
rect 489524 270285 489580 270294
rect 488084 268278 488140 268287
rect 488084 268213 488140 268222
rect 489538 267991 489566 270285
rect 489622 268979 489674 268985
rect 489718 268979 489770 268985
rect 489674 268939 489718 268967
rect 489622 268921 489674 268927
rect 489718 268921 489770 268927
rect 489524 267982 489580 267991
rect 489524 267917 489580 267926
rect 485686 265723 485738 265729
rect 485686 265665 485738 265671
rect 492898 265655 492926 277870
rect 494050 266617 494078 277870
rect 495202 269281 495230 277870
rect 496162 277856 496464 277884
rect 496162 277759 496190 277856
rect 496148 277750 496204 277759
rect 496148 277685 496204 277694
rect 495190 269275 495242 269281
rect 495190 269217 495242 269223
rect 494038 266611 494090 266617
rect 494038 266553 494090 266559
rect 497602 266543 497630 277870
rect 498850 274355 498878 277870
rect 498836 274346 498892 274355
rect 498836 274281 498892 274290
rect 497590 266537 497642 266543
rect 497590 266479 497642 266485
rect 492886 265649 492938 265655
rect 492886 265591 492938 265597
rect 499906 265581 499934 277870
rect 501046 271273 501098 271279
rect 501044 271238 501046 271247
rect 501098 271238 501100 271247
rect 501044 271173 501100 271182
rect 501154 268467 501182 277870
rect 502306 268583 502334 277870
rect 503554 270465 503582 277870
rect 504706 277051 504734 277870
rect 504694 277045 504746 277051
rect 504694 276987 504746 276993
rect 505954 274503 505982 277870
rect 507106 277611 507134 277870
rect 507092 277602 507148 277611
rect 507092 277537 507148 277546
rect 505940 274494 505996 274503
rect 505940 274429 505996 274438
rect 508354 274239 508382 277870
rect 508342 274233 508394 274239
rect 508342 274175 508394 274181
rect 503542 270459 503594 270465
rect 503542 270401 503594 270407
rect 509506 268879 509534 277870
rect 510658 270835 510686 277870
rect 511906 274313 511934 277870
rect 511894 274307 511946 274313
rect 511894 274249 511946 274255
rect 510646 270829 510698 270835
rect 510646 270771 510698 270777
rect 513058 270507 513086 277870
rect 513044 270498 513100 270507
rect 513044 270433 513100 270442
rect 509492 268870 509548 268879
rect 509492 268805 509548 268814
rect 502292 268574 502348 268583
rect 502292 268509 502348 268518
rect 501142 268461 501194 268467
rect 501142 268403 501194 268409
rect 499894 265575 499946 265581
rect 499894 265517 499946 265523
rect 514306 265507 514334 277870
rect 515458 276903 515486 277870
rect 515446 276897 515498 276903
rect 515446 276839 515498 276845
rect 516610 274651 516638 277870
rect 517762 277463 517790 277870
rect 517748 277454 517804 277463
rect 517748 277389 517804 277398
rect 519010 276755 519038 277870
rect 518998 276749 519050 276755
rect 518998 276691 519050 276697
rect 520162 274799 520190 277870
rect 520148 274790 520204 274799
rect 520148 274725 520204 274734
rect 516596 274642 516652 274651
rect 516596 274577 516652 274586
rect 518434 271057 518558 271076
rect 518422 271051 518570 271057
rect 518474 271048 518518 271051
rect 518422 270993 518474 270999
rect 518518 270993 518570 270999
rect 518326 269053 518378 269059
rect 518378 269001 518462 269004
rect 518326 268995 518462 269001
rect 518338 268985 518462 268995
rect 518338 268979 518474 268985
rect 518338 268976 518422 268979
rect 518422 268921 518474 268927
rect 514294 265501 514346 265507
rect 412916 265466 412972 265475
rect 514294 265443 514346 265449
rect 521410 265433 521438 277870
rect 522562 266247 522590 277870
rect 523810 276829 523838 277870
rect 523798 276823 523850 276829
rect 523798 276765 523850 276771
rect 524962 269873 524990 277870
rect 524950 269867 525002 269873
rect 524950 269809 525002 269815
rect 526114 268763 526142 277870
rect 526102 268757 526154 268763
rect 526102 268699 526154 268705
rect 522550 266241 522602 266247
rect 522550 266183 522602 266189
rect 412916 265401 412972 265410
rect 521398 265427 521450 265433
rect 521398 265369 521450 265375
rect 527362 265327 527390 277870
rect 528514 277315 528542 277870
rect 528500 277306 528556 277315
rect 528500 277241 528556 277250
rect 529762 268911 529790 277870
rect 529750 268905 529802 268911
rect 529750 268847 529802 268853
rect 412820 265318 412876 265327
rect 412820 265253 412876 265262
rect 527348 265318 527404 265327
rect 527348 265253 527404 265262
rect 530914 265179 530942 277870
rect 532162 275867 532190 277870
rect 532150 275861 532202 275867
rect 532150 275803 532202 275809
rect 533218 265951 533246 277870
rect 534466 271131 534494 277870
rect 534454 271125 534506 271131
rect 534454 271067 534506 271073
rect 533206 265945 533258 265951
rect 533206 265887 533258 265893
rect 535618 265359 535646 277870
rect 536866 269059 536894 277870
rect 536854 269053 536906 269059
rect 536854 268995 536906 269001
rect 535606 265353 535658 265359
rect 535606 265295 535658 265301
rect 412724 265170 412780 265179
rect 412724 265105 412780 265114
rect 530900 265170 530956 265179
rect 530900 265105 530956 265114
rect 412628 265022 412684 265031
rect 412628 264957 412630 264966
rect 412682 264957 412684 264966
rect 412630 264925 412682 264931
rect 412738 264915 412766 265105
rect 538018 265031 538046 277870
rect 539266 277167 539294 277870
rect 539252 277158 539308 277167
rect 539252 277093 539308 277102
rect 540418 274683 540446 277870
rect 540406 274677 540458 274683
rect 540406 274619 540458 274625
rect 541570 270909 541598 277870
rect 541558 270903 541610 270909
rect 541558 270845 541610 270851
rect 539924 270202 539980 270211
rect 539924 270137 539980 270146
rect 539938 268879 539966 270137
rect 540020 270054 540076 270063
rect 540020 269989 540076 269998
rect 539924 268870 539980 268879
rect 539924 268805 539980 268814
rect 540034 268583 540062 269989
rect 542818 269503 542846 277870
rect 543970 271279 543998 277870
rect 543958 271273 544010 271279
rect 543958 271215 544010 271221
rect 545218 271205 545246 277870
rect 545206 271199 545258 271205
rect 545206 271141 545258 271147
rect 542806 269497 542858 269503
rect 542806 269439 542858 269445
rect 540020 268574 540076 268583
rect 540020 268509 540076 268518
rect 546370 265285 546398 277870
rect 547618 265803 547646 277870
rect 547714 277856 548784 277884
rect 547606 265797 547658 265803
rect 547606 265739 547658 265745
rect 546358 265279 546410 265285
rect 546358 265221 546410 265227
rect 538004 265022 538060 265031
rect 538004 264957 538060 264966
rect 412726 264909 412778 264915
rect 412726 264851 412778 264857
rect 489524 264874 489580 264883
rect 489524 264809 489580 264818
rect 489538 264767 489566 264809
rect 449398 264761 449450 264767
rect 449396 264726 449398 264735
rect 469366 264761 469418 264767
rect 449450 264726 449452 264735
rect 449396 264661 449452 264670
rect 469364 264726 469366 264735
rect 475798 264761 475850 264767
rect 469418 264726 469420 264735
rect 469364 264661 469420 264670
rect 475796 264726 475798 264735
rect 489526 264761 489578 264767
rect 475850 264726 475852 264735
rect 489526 264703 489578 264709
rect 475796 264661 475852 264670
rect 547714 257756 547742 277856
rect 549922 271871 549950 277870
rect 551074 274831 551102 277870
rect 551062 274825 551114 274831
rect 551062 274767 551114 274773
rect 552322 274059 552350 277870
rect 552308 274050 552364 274059
rect 552308 273985 552364 273994
rect 549910 271865 549962 271871
rect 549910 271807 549962 271813
rect 548566 271051 548618 271057
rect 548566 270993 548618 270999
rect 548578 270909 548606 270993
rect 548566 270903 548618 270909
rect 548566 270845 548618 270851
rect 548566 270533 548618 270539
rect 548564 270498 548566 270507
rect 548618 270498 548620 270507
rect 548564 270433 548620 270442
rect 553474 269355 553502 277870
rect 553462 269349 553514 269355
rect 553462 269291 553514 269297
rect 554722 268319 554750 277870
rect 554710 268313 554762 268319
rect 554710 268255 554762 268261
rect 555874 264587 555902 277870
rect 557026 273499 557054 277870
rect 558274 274979 558302 277870
rect 558262 274973 558314 274979
rect 558262 274915 558314 274921
rect 557014 273493 557066 273499
rect 557014 273435 557066 273441
rect 559426 271395 559454 277870
rect 559412 271386 559468 271395
rect 559412 271321 559468 271330
rect 558646 271051 558698 271057
rect 558646 270993 558698 270999
rect 558658 270909 558686 270993
rect 558646 270903 558698 270909
rect 558646 270845 558698 270851
rect 560180 270202 560236 270211
rect 560180 270137 560236 270146
rect 560084 270054 560140 270063
rect 560084 269989 560140 269998
rect 560098 268583 560126 269989
rect 560194 268879 560222 270137
rect 560180 268870 560236 268879
rect 560180 268805 560236 268814
rect 560084 268574 560140 268583
rect 560084 268509 560140 268518
rect 560674 268139 560702 277870
rect 561826 270613 561854 277870
rect 563074 273171 563102 277870
rect 564226 275497 564254 277870
rect 565474 276385 565502 277870
rect 565462 276379 565514 276385
rect 565462 276321 565514 276327
rect 564214 275491 564266 275497
rect 564214 275433 564266 275439
rect 563060 273162 563116 273171
rect 563060 273097 563116 273106
rect 566530 272241 566558 277870
rect 566518 272235 566570 272241
rect 566518 272177 566570 272183
rect 564500 271090 564556 271099
rect 564500 271025 564502 271034
rect 564554 271025 564556 271034
rect 564502 270993 564554 270999
rect 561814 270607 561866 270613
rect 561814 270549 561866 270555
rect 567778 268731 567806 277870
rect 568930 270317 568958 277870
rect 570178 270761 570206 277870
rect 571330 275275 571358 277870
rect 572482 276311 572510 277870
rect 572470 276305 572522 276311
rect 572470 276247 572522 276253
rect 571318 275269 571370 275275
rect 571318 275211 571370 275217
rect 573730 272167 573758 277870
rect 573718 272161 573770 272167
rect 573718 272103 573770 272109
rect 570166 270755 570218 270761
rect 570166 270697 570218 270703
rect 568918 270311 568970 270317
rect 568918 270253 568970 270259
rect 574882 269027 574910 277870
rect 575830 270533 575882 270539
rect 575830 270475 575882 270481
rect 575924 270498 575980 270507
rect 575842 270336 575870 270475
rect 575924 270433 575980 270442
rect 575938 270336 575966 270433
rect 575842 270308 575966 270336
rect 576130 270243 576158 277870
rect 576226 277856 577296 277884
rect 576118 270237 576170 270243
rect 576118 270179 576170 270185
rect 574868 269018 574924 269027
rect 574868 268953 574924 268962
rect 567764 268722 567820 268731
rect 567764 268657 567820 268666
rect 560660 268130 560716 268139
rect 560660 268065 560716 268074
rect 555860 264578 555916 264587
rect 555860 264513 555916 264522
rect 547522 257728 547742 257756
rect 412258 247516 412670 247544
rect 412148 247493 412204 247502
rect 412052 247262 412108 247271
rect 412052 247197 412108 247206
rect 406496 246834 406612 246840
rect 226388 246818 226444 246827
rect 212278 246779 212330 246785
rect 227348 246818 227404 246827
rect 226388 246753 226444 246762
rect 227062 246779 227114 246785
rect 212278 246721 212330 246727
rect 212182 246557 212234 246563
rect 212182 246499 212234 246505
rect 212086 246409 212138 246415
rect 212086 246351 212138 246357
rect 211990 246187 212042 246193
rect 211990 246129 212042 246135
rect 211508 243710 211564 243719
rect 211508 243645 211564 243654
rect 211316 238974 211372 238983
rect 211316 238909 211372 238918
rect 211220 238826 211276 238835
rect 211220 238761 211276 238770
rect 212180 236754 212236 236763
rect 212180 236689 212236 236698
rect 211303 233811 211363 233820
rect 212194 233761 212222 236689
rect 212386 235135 212414 246494
rect 212770 240643 212798 246494
rect 213142 244929 213194 244935
rect 213142 244871 213194 244877
rect 212758 240637 212810 240643
rect 212758 240579 212810 240585
rect 213046 236197 213098 236203
rect 213046 236139 213098 236145
rect 212372 235126 212428 235135
rect 212372 235061 212428 235070
rect 212564 233942 212620 233951
rect 212564 233877 212620 233886
rect 212276 233794 212332 233803
rect 211303 233742 211363 233751
rect 212182 233755 212234 233761
rect 210934 233533 210986 233539
rect 211319 233532 211347 233742
rect 212276 233729 212332 233738
rect 212182 233697 212234 233703
rect 212084 233646 212140 233655
rect 212084 233581 212140 233590
rect 211299 233526 211374 233532
rect 210986 233481 211200 233484
rect 210934 233475 211200 233481
rect 210946 233456 211200 233475
rect 211299 233474 211307 233526
rect 211359 233474 211374 233526
rect 211700 233498 211756 233507
rect 211299 233465 211374 233474
rect 211584 233456 211700 233484
rect 212098 233484 212126 233581
rect 211968 233456 212126 233484
rect 212290 233470 212318 233729
rect 212578 233655 212606 233877
rect 212564 233646 212620 233655
rect 212564 233581 212620 233590
rect 212578 233484 212606 233581
rect 212578 233456 212688 233484
rect 213058 233470 213086 236139
rect 213154 233613 213182 244871
rect 213250 242979 213278 246494
rect 213696 246480 213950 246508
rect 214080 246480 214238 246508
rect 213526 245151 213578 245157
rect 213526 245093 213578 245099
rect 213236 242970 213292 242979
rect 213236 242905 213292 242914
rect 213538 233687 213566 245093
rect 213922 241605 213950 246480
rect 214006 245225 214058 245231
rect 214006 245167 214058 245173
rect 213910 241599 213962 241605
rect 213910 241541 213962 241547
rect 213526 233681 213578 233687
rect 213526 233623 213578 233629
rect 213142 233607 213194 233613
rect 213142 233549 213194 233555
rect 213154 233484 213182 233549
rect 213538 233484 213566 233623
rect 213910 233533 213962 233539
rect 213154 233456 213408 233484
rect 213538 233456 213792 233484
rect 214018 233484 214046 245167
rect 214210 234987 214238 246480
rect 214294 245077 214346 245083
rect 214294 245019 214346 245025
rect 214196 234978 214252 234987
rect 214196 234913 214252 234922
rect 214306 233507 214334 245019
rect 214498 239755 214526 246494
rect 214978 243127 215006 246494
rect 214964 243118 215020 243127
rect 214964 243053 215020 243062
rect 215458 241827 215486 246494
rect 215808 246480 215966 246508
rect 216288 246480 216542 246508
rect 215446 241821 215498 241827
rect 215446 241763 215498 241769
rect 214486 239749 214538 239755
rect 214486 239691 214538 239697
rect 215938 239681 215966 246480
rect 216022 246113 216074 246119
rect 216022 246055 216074 246061
rect 216034 245675 216062 246055
rect 216022 245669 216074 245675
rect 216022 245611 216074 245617
rect 216514 244935 216542 246480
rect 216598 245225 216650 245231
rect 216598 245167 216650 245173
rect 216502 244929 216554 244935
rect 216502 244871 216554 244877
rect 215926 239675 215978 239681
rect 215926 239617 215978 239623
rect 215828 238234 215884 238243
rect 215828 238169 215884 238178
rect 215252 238086 215308 238095
rect 215252 238021 215308 238030
rect 214868 237938 214924 237947
rect 214868 237873 214924 237882
rect 214772 237642 214828 237651
rect 214772 237577 214828 237586
rect 214786 236615 214814 237577
rect 214772 236606 214828 236615
rect 214772 236541 214828 236550
rect 214292 233498 214348 233507
rect 213962 233481 214176 233484
rect 213910 233475 214176 233481
rect 213922 233456 214176 233475
rect 211700 233433 211756 233442
rect 214348 233456 214512 233484
rect 214882 233470 214910 237873
rect 215266 233470 215294 238021
rect 215842 233484 215870 238169
rect 216212 237642 216268 237651
rect 216212 237577 216268 237586
rect 216226 233484 216254 237577
rect 216610 233484 216638 245167
rect 216706 240939 216734 246494
rect 217186 242091 217214 246494
rect 217172 242082 217228 242091
rect 217172 242017 217228 242026
rect 216694 240933 216746 240939
rect 216694 240875 216746 240881
rect 217570 240199 217598 246494
rect 218016 246480 218270 246508
rect 218496 246480 218750 246508
rect 217558 240193 217610 240199
rect 217558 240135 217610 240141
rect 218038 238343 218090 238349
rect 218038 238285 218090 238291
rect 216692 237790 216748 237799
rect 216692 237725 216748 237734
rect 215616 233456 215870 233484
rect 216000 233456 216254 233484
rect 216384 233456 216638 233484
rect 216706 233470 216734 237725
rect 217078 237307 217130 237313
rect 217078 237249 217130 237255
rect 217090 233470 217118 237249
rect 217462 236197 217514 236203
rect 217462 236139 217514 236145
rect 217474 233470 217502 236139
rect 218050 233484 218078 238285
rect 218242 235283 218270 246480
rect 218722 241901 218750 246480
rect 218914 242831 218942 246494
rect 218900 242822 218956 242831
rect 218900 242757 218956 242766
rect 218710 241895 218762 241901
rect 218710 241837 218762 241843
rect 219298 241753 219326 246494
rect 219286 241747 219338 241753
rect 219286 241689 219338 241695
rect 219286 240859 219338 240865
rect 219286 240801 219338 240807
rect 218806 240711 218858 240717
rect 218806 240653 218858 240659
rect 218422 240341 218474 240347
rect 218422 240283 218474 240289
rect 218228 235274 218284 235283
rect 218228 235209 218284 235218
rect 218434 233484 218462 240283
rect 218818 233484 218846 240653
rect 218902 239675 218954 239681
rect 218902 239617 218954 239623
rect 217824 233456 218078 233484
rect 218208 233456 218462 233484
rect 218592 233456 218846 233484
rect 218914 233470 218942 239617
rect 219298 233470 219326 240801
rect 219670 240415 219722 240421
rect 219670 240357 219722 240363
rect 219682 233470 219710 240357
rect 219778 235727 219806 246494
rect 220224 246480 220478 246508
rect 220608 246480 220862 246508
rect 221040 246480 221342 246508
rect 220450 241013 220478 246480
rect 220834 242683 220862 246480
rect 221206 243523 221258 243529
rect 221206 243465 221258 243471
rect 221218 243275 221246 243465
rect 221204 243266 221260 243275
rect 221204 243201 221260 243210
rect 220820 242674 220876 242683
rect 220820 242609 220876 242618
rect 220438 241007 220490 241013
rect 220438 240949 220490 240955
rect 220246 240489 220298 240495
rect 220246 240431 220298 240437
rect 219764 235718 219820 235727
rect 219764 235653 219820 235662
rect 220258 233484 220286 240431
rect 220630 240045 220682 240051
rect 220630 239987 220682 239993
rect 220642 233484 220670 239987
rect 221110 238417 221162 238423
rect 221110 238359 221162 238365
rect 221014 237751 221066 237757
rect 221014 237693 221066 237699
rect 221026 233484 221054 237693
rect 220032 233456 220286 233484
rect 220416 233456 220670 233484
rect 220800 233456 221054 233484
rect 221122 233470 221150 238359
rect 221314 235875 221342 246480
rect 221396 243266 221452 243275
rect 221396 243201 221452 243210
rect 221410 241827 221438 243201
rect 221398 241821 221450 241827
rect 221398 241763 221450 241769
rect 221506 241679 221534 246494
rect 221782 246409 221834 246415
rect 221878 246409 221930 246415
rect 221834 246369 221878 246397
rect 221782 246351 221834 246357
rect 221878 246351 221930 246357
rect 221986 242419 222014 246494
rect 222336 246480 222590 246508
rect 222816 246480 223070 246508
rect 221974 242413 222026 242419
rect 221974 242355 222026 242361
rect 221494 241673 221546 241679
rect 221494 241615 221546 241621
rect 221782 240563 221834 240569
rect 221782 240505 221834 240511
rect 221494 237381 221546 237387
rect 221494 237323 221546 237329
rect 221300 235866 221356 235875
rect 221300 235801 221356 235810
rect 221506 233470 221534 237323
rect 221794 236203 221822 240505
rect 222562 240125 222590 246480
rect 222550 240119 222602 240125
rect 222550 240061 222602 240067
rect 221878 238269 221930 238275
rect 221878 238211 221930 238217
rect 221782 236197 221834 236203
rect 221782 236139 221834 236145
rect 221890 233470 221918 238211
rect 222838 238195 222890 238201
rect 222838 238137 222890 238143
rect 221974 237825 222026 237831
rect 221974 237767 222026 237773
rect 221986 233484 222014 237767
rect 222850 233484 222878 238137
rect 223042 235579 223070 246480
rect 223234 241531 223262 246494
rect 223714 242239 223742 246494
rect 223700 242230 223756 242239
rect 223700 242165 223756 242174
rect 223222 241525 223274 241531
rect 223222 241467 223274 241473
rect 224098 239311 224126 246494
rect 224530 246212 224558 246494
rect 225024 246480 225278 246508
rect 224482 246184 224558 246212
rect 224086 239305 224138 239311
rect 224086 239247 224138 239253
rect 223222 238121 223274 238127
rect 223222 238063 223274 238069
rect 223028 235570 223084 235579
rect 223028 235505 223084 235514
rect 223234 233484 223262 238063
rect 223318 237973 223370 237979
rect 223318 237915 223370 237921
rect 221986 233456 222240 233484
rect 222624 233456 222878 233484
rect 223008 233456 223262 233484
rect 223330 233470 223358 237915
rect 224086 237899 224138 237905
rect 224086 237841 224138 237847
rect 223702 236937 223754 236943
rect 223702 236879 223754 236885
rect 223714 233470 223742 236879
rect 224098 233470 224126 237841
rect 224482 235431 224510 246184
rect 225250 241087 225278 246480
rect 225442 241235 225470 246494
rect 225430 241229 225482 241235
rect 225430 241171 225482 241177
rect 225238 241081 225290 241087
rect 225238 241023 225290 241029
rect 225142 239749 225194 239755
rect 225142 239691 225194 239697
rect 225046 237825 225098 237831
rect 225046 237767 225098 237773
rect 224566 237011 224618 237017
rect 224566 236953 224618 236959
rect 224468 235422 224524 235431
rect 224468 235357 224524 235366
rect 224578 233484 224606 236953
rect 225058 233484 225086 237767
rect 224448 233456 224606 233484
rect 224832 233456 225086 233484
rect 225154 233484 225182 239691
rect 225526 236419 225578 236425
rect 225526 236361 225578 236367
rect 225154 233456 225216 233484
rect 225538 233470 225566 236361
rect 225826 236171 225854 246494
rect 226004 243710 226060 243719
rect 226004 243645 226060 243654
rect 226018 243233 226046 243645
rect 226006 243227 226058 243233
rect 226006 243169 226058 243175
rect 226306 241309 226334 246494
rect 226402 245157 226430 246753
rect 227348 246753 227404 246762
rect 237044 246818 237100 246827
rect 237716 246818 237772 246827
rect 237044 246753 237100 246762
rect 237250 246776 237600 246804
rect 227062 246721 227114 246727
rect 226752 246480 226814 246508
rect 226390 245151 226442 245157
rect 226390 245093 226442 245099
rect 226786 243455 226814 246480
rect 226966 246483 227018 246489
rect 226966 246425 227018 246431
rect 226978 245749 227006 246425
rect 227074 246045 227102 246721
rect 227218 246212 227246 246494
rect 227218 246184 227294 246212
rect 227062 246039 227114 246045
rect 227062 245981 227114 245987
rect 226966 245743 227018 245749
rect 226966 245685 227018 245691
rect 226774 243449 226826 243455
rect 226774 243391 226826 243397
rect 226294 241303 226346 241309
rect 226294 241245 226346 241251
rect 227266 239607 227294 246184
rect 227362 245823 227390 246753
rect 232150 246557 232202 246563
rect 227568 246480 227870 246508
rect 227350 245817 227402 245823
rect 227350 245759 227402 245765
rect 227444 243710 227500 243719
rect 227444 243645 227500 243654
rect 227458 243529 227486 243645
rect 227446 243523 227498 243529
rect 227446 243465 227498 243471
rect 227732 242378 227788 242387
rect 227732 242313 227788 242322
rect 227746 242271 227774 242313
rect 227350 242265 227402 242271
rect 227350 242207 227402 242213
rect 227734 242265 227786 242271
rect 227734 242207 227786 242213
rect 227362 242091 227390 242207
rect 227348 242082 227404 242091
rect 227348 242017 227404 242026
rect 227254 239601 227306 239607
rect 227254 239543 227306 239549
rect 227254 238787 227306 238793
rect 227254 238729 227306 238735
rect 226294 238713 226346 238719
rect 226294 238655 226346 238661
rect 225910 237085 225962 237091
rect 225910 237027 225962 237033
rect 225812 236162 225868 236171
rect 225812 236097 225868 236106
rect 225922 233470 225950 237027
rect 226306 233470 226334 238655
rect 226870 236715 226922 236721
rect 226870 236657 226922 236663
rect 226882 233484 226910 236657
rect 227266 233484 227294 238729
rect 227734 238565 227786 238571
rect 227734 238507 227786 238513
rect 227350 237455 227402 237461
rect 227350 237397 227402 237403
rect 226656 233456 226910 233484
rect 227040 233456 227294 233484
rect 214292 233433 214348 233442
rect 227362 233336 227390 237397
rect 227444 236754 227500 236763
rect 227636 236754 227692 236763
rect 227500 236712 227636 236740
rect 227444 236689 227500 236698
rect 227636 236689 227692 236698
rect 227746 233470 227774 238507
rect 227842 234723 227870 246480
rect 228034 239755 228062 246494
rect 228514 243381 228542 246494
rect 228864 246480 229214 246508
rect 229344 246480 229598 246508
rect 228502 243375 228554 243381
rect 228502 243317 228554 243323
rect 228212 243266 228268 243275
rect 228212 243201 228268 243210
rect 228226 242091 228254 243201
rect 228212 242082 228268 242091
rect 228212 242017 228268 242026
rect 229186 241772 229214 246480
rect 229186 241744 229406 241772
rect 229174 241599 229226 241605
rect 229174 241541 229226 241547
rect 228022 239749 228074 239755
rect 228022 239691 228074 239697
rect 229078 239675 229130 239681
rect 229078 239617 229130 239623
rect 228502 239009 228554 239015
rect 228502 238951 228554 238957
rect 228118 238935 228170 238941
rect 228118 238877 228170 238883
rect 227830 234717 227882 234723
rect 227830 234659 227882 234665
rect 228130 233470 228158 238877
rect 228514 233470 228542 238951
rect 229090 233484 229118 239617
rect 229186 233780 229214 241541
rect 229186 233752 229262 233780
rect 228864 233456 229118 233484
rect 229234 233470 229262 233752
rect 229378 233484 229406 241744
rect 229570 236023 229598 246480
rect 229762 243529 229790 246494
rect 229750 243523 229802 243529
rect 229750 243465 229802 243471
rect 229942 239749 229994 239755
rect 229942 239691 229994 239697
rect 229556 236014 229612 236023
rect 229556 235949 229612 235958
rect 229378 233456 229632 233484
rect 229954 233470 229982 239691
rect 230242 239681 230270 246494
rect 230230 239675 230282 239681
rect 230230 239617 230282 239623
rect 230326 239601 230378 239607
rect 230326 239543 230378 239549
rect 230338 233470 230366 239543
rect 230626 234797 230654 246494
rect 230818 246480 231072 246508
rect 231552 246480 231806 246508
rect 232150 246499 232202 246505
rect 230710 241303 230762 241309
rect 230710 241245 230762 241251
rect 230614 234791 230666 234797
rect 230614 234733 230666 234739
rect 230722 233470 230750 241245
rect 230818 239015 230846 246480
rect 231778 243677 231806 246480
rect 231862 246409 231914 246415
rect 231862 246351 231914 246357
rect 231874 246045 231902 246351
rect 231862 246039 231914 246045
rect 231862 245981 231914 245987
rect 231766 243671 231818 243677
rect 231766 243613 231818 243619
rect 230902 241229 230954 241235
rect 230902 241171 230954 241177
rect 230806 239009 230858 239015
rect 230806 238951 230858 238957
rect 230914 233484 230942 241171
rect 231190 241081 231242 241087
rect 231190 241023 231242 241029
rect 231202 233484 231230 241023
rect 231574 239305 231626 239311
rect 231574 239247 231626 239253
rect 231586 233484 231614 239247
rect 231970 238941 231998 246494
rect 232162 245749 232190 246499
rect 232150 245743 232202 245749
rect 232150 245685 232202 245691
rect 232150 241525 232202 241531
rect 232150 241467 232202 241473
rect 231958 238935 232010 238941
rect 231958 238877 232010 238883
rect 230914 233456 231072 233484
rect 231202 233456 231456 233484
rect 231586 233456 231840 233484
rect 232162 233470 232190 241467
rect 232354 240791 232382 246494
rect 232342 240785 232394 240791
rect 232342 240727 232394 240733
rect 232534 240119 232586 240125
rect 232534 240061 232586 240067
rect 232546 233470 232574 240061
rect 232834 238571 232862 246494
rect 233280 246480 233534 246508
rect 233506 241827 233534 246480
rect 233602 246480 233760 246508
rect 233494 241821 233546 241827
rect 233494 241763 233546 241769
rect 232918 241673 232970 241679
rect 232918 241615 232970 241621
rect 232822 238565 232874 238571
rect 232822 238507 232874 238513
rect 232930 233470 232958 241615
rect 233398 241007 233450 241013
rect 233398 240949 233450 240955
rect 233302 240637 233354 240643
rect 233302 240579 233354 240585
rect 233314 233484 233342 240579
rect 233280 233456 233342 233484
rect 233410 233484 233438 240949
rect 233602 237461 233630 246480
rect 233782 241747 233834 241753
rect 233782 241689 233834 241695
rect 233590 237455 233642 237461
rect 233590 237397 233642 237403
rect 233794 233484 233822 241689
rect 234082 238793 234110 246494
rect 234562 241901 234590 246494
rect 234358 241895 234410 241901
rect 234358 241837 234410 241843
rect 234550 241895 234602 241901
rect 234550 241837 234602 241843
rect 234070 238787 234122 238793
rect 234070 238729 234122 238735
rect 233410 233456 233664 233484
rect 233794 233456 234048 233484
rect 234370 233470 234398 241837
rect 234742 240193 234794 240199
rect 234742 240135 234794 240141
rect 234754 233470 234782 240135
rect 235042 236721 235070 246494
rect 235488 246480 235550 246508
rect 235126 244263 235178 244269
rect 235126 244205 235178 244211
rect 235030 236715 235082 236721
rect 235030 236657 235082 236663
rect 235138 233470 235166 244205
rect 235522 239237 235550 246480
rect 235618 246480 235872 246508
rect 235510 239231 235562 239237
rect 235510 239173 235562 239179
rect 235618 238719 235646 246480
rect 236086 245965 236138 245971
rect 236086 245907 236138 245913
rect 236098 245675 236126 245907
rect 236086 245669 236138 245675
rect 236086 245611 236138 245617
rect 236290 243603 236318 246494
rect 236278 243597 236330 243603
rect 236278 243539 236330 243545
rect 236182 243227 236234 243233
rect 236182 243169 236234 243175
rect 236194 243085 236222 243169
rect 236182 243079 236234 243085
rect 236182 243021 236234 243027
rect 236470 241673 236522 241679
rect 236470 241615 236522 241621
rect 236182 240933 236234 240939
rect 236182 240875 236234 240881
rect 236194 239089 236222 240875
rect 236182 239083 236234 239089
rect 236182 239025 236234 239031
rect 235606 238713 235658 238719
rect 235606 238655 235658 238661
rect 235702 235901 235754 235907
rect 235702 235843 235754 235849
rect 235714 233484 235742 235843
rect 236086 235457 236138 235463
rect 236086 235399 236138 235405
rect 236098 233484 236126 235399
rect 236482 233484 236510 241615
rect 236566 239971 236618 239977
rect 236566 239913 236618 239919
rect 235488 233456 235742 233484
rect 235872 233456 236126 233484
rect 236256 233456 236510 233484
rect 236578 233470 236606 239913
rect 236770 237091 236798 246494
rect 237058 245897 237086 246753
rect 237046 245891 237098 245897
rect 237046 245833 237098 245839
rect 236950 240193 237002 240199
rect 236950 240135 237002 240141
rect 236758 237085 236810 237091
rect 236758 237027 236810 237033
rect 236962 233470 236990 240135
rect 237154 239163 237182 246494
rect 237142 239157 237194 239163
rect 237142 239099 237194 239105
rect 237250 236425 237278 246776
rect 237716 246753 237772 246762
rect 240020 246818 240076 246827
rect 240020 246753 240076 246762
rect 240500 246818 240556 246827
rect 240500 246753 240556 246762
rect 241748 246818 241804 246827
rect 241748 246753 241804 246762
rect 242516 246818 242572 246827
rect 242516 246753 242572 246762
rect 252500 246818 252556 246827
rect 252500 246753 252556 246762
rect 252692 246818 252748 246827
rect 252692 246753 252748 246762
rect 266708 246818 266764 246827
rect 266708 246753 266764 246762
rect 268628 246818 268684 246827
rect 286100 246818 286156 246827
rect 278544 246776 278942 246804
rect 268628 246753 268684 246762
rect 237730 246119 237758 246753
rect 237814 246705 237866 246711
rect 237814 246647 237866 246653
rect 237826 246267 237854 246647
rect 238080 246480 238334 246508
rect 237814 246261 237866 246267
rect 237814 246203 237866 246209
rect 237718 246113 237770 246119
rect 237718 246055 237770 246061
rect 237716 242822 237772 242831
rect 237442 242780 237716 242808
rect 237442 242683 237470 242780
rect 237716 242757 237772 242766
rect 237428 242674 237484 242683
rect 237428 242609 237484 242618
rect 238306 242197 238334 246480
rect 238294 242191 238346 242197
rect 238294 242133 238346 242139
rect 237526 241081 237578 241087
rect 237526 241023 237578 241029
rect 237430 240933 237482 240939
rect 237430 240875 237482 240881
rect 237334 240119 237386 240125
rect 237334 240061 237386 240067
rect 237238 236419 237290 236425
rect 237238 236361 237290 236367
rect 237346 233470 237374 240061
rect 237442 240051 237470 240875
rect 237538 240569 237566 241023
rect 237622 241007 237674 241013
rect 237622 240949 237674 240955
rect 237526 240563 237578 240569
rect 237526 240505 237578 240511
rect 237634 240347 237662 240949
rect 237622 240341 237674 240347
rect 237622 240283 237674 240289
rect 237910 240267 237962 240273
rect 237910 240209 237962 240215
rect 237430 240045 237482 240051
rect 237430 239987 237482 239993
rect 237922 233484 237950 240209
rect 238498 239089 238526 246494
rect 238678 240785 238730 240791
rect 238678 240727 238730 240733
rect 238198 239083 238250 239089
rect 238198 239025 238250 239031
rect 238486 239083 238538 239089
rect 238486 239025 238538 239031
rect 238054 233755 238106 233761
rect 238054 233697 238106 233703
rect 237696 233456 237950 233484
rect 238066 233470 238094 233697
rect 238210 233484 238238 239025
rect 238690 234395 238718 240727
rect 238882 237831 238910 246494
rect 239362 243751 239390 246494
rect 239650 246480 239808 246508
rect 239350 243745 239402 243751
rect 239350 243687 239402 243693
rect 238966 241969 239018 241975
rect 238966 241911 239018 241917
rect 238978 241827 239006 241911
rect 238966 241821 239018 241827
rect 238966 241763 239018 241769
rect 239062 241821 239114 241827
rect 239062 241763 239114 241769
rect 238966 239231 239018 239237
rect 238966 239173 239018 239179
rect 238870 237825 238922 237831
rect 238870 237767 238922 237773
rect 238774 237455 238826 237461
rect 238774 237397 238826 237403
rect 238676 234386 238732 234395
rect 238676 234321 238732 234330
rect 238210 233456 238464 233484
rect 238786 233470 238814 237397
rect 238978 234543 239006 239173
rect 238964 234534 239020 234543
rect 238964 234469 239020 234478
rect 239074 233761 239102 241763
rect 239158 241525 239210 241531
rect 239158 241467 239210 241473
rect 239062 233755 239114 233761
rect 239062 233697 239114 233703
rect 239170 233470 239198 241467
rect 239542 238935 239594 238941
rect 239542 238877 239594 238883
rect 239554 233470 239582 238877
rect 239650 237017 239678 246480
rect 240034 246045 240062 246753
rect 240274 246212 240302 246494
rect 240514 246267 240542 246753
rect 240610 246480 240672 246508
rect 241104 246480 241502 246508
rect 240502 246261 240554 246267
rect 240274 246184 240350 246212
rect 240502 246203 240554 246209
rect 240022 246039 240074 246045
rect 240022 245981 240074 245987
rect 240322 239385 240350 246184
rect 240310 239379 240362 239385
rect 240310 239321 240362 239327
rect 240502 239009 240554 239015
rect 240502 238951 240554 238957
rect 240118 238861 240170 238867
rect 240118 238803 240170 238809
rect 239638 237011 239690 237017
rect 239638 236953 239690 236959
rect 240130 233484 240158 238803
rect 240514 233484 240542 238951
rect 240610 237905 240638 246480
rect 241474 242049 241502 246480
rect 241462 242043 241514 242049
rect 241462 241985 241514 241991
rect 240980 240454 241036 240463
rect 240980 240389 241036 240398
rect 240886 240341 240938 240347
rect 240886 240283 240938 240289
rect 240598 237899 240650 237905
rect 240598 237841 240650 237847
rect 240898 233484 240926 240283
rect 239904 233456 240158 233484
rect 240288 233456 240542 233484
rect 240672 233456 240926 233484
rect 240994 233470 241022 240389
rect 241364 238530 241420 238539
rect 241364 238465 241420 238474
rect 241378 233470 241406 238465
rect 241570 236943 241598 246494
rect 241762 246045 241790 246753
rect 242146 246628 242400 246656
rect 242016 246480 242078 246508
rect 241750 246039 241802 246045
rect 241750 245981 241802 245987
rect 241748 240602 241804 240611
rect 241748 240537 241804 240546
rect 241654 239157 241706 239163
rect 241654 239099 241706 239105
rect 241558 236937 241610 236943
rect 241558 236879 241610 236885
rect 241666 235241 241694 239099
rect 241654 235235 241706 235241
rect 241654 235177 241706 235183
rect 241762 233470 241790 240537
rect 241846 239083 241898 239089
rect 241846 239025 241898 239031
rect 241858 235093 241886 239025
rect 242050 235167 242078 246480
rect 242146 237979 242174 246628
rect 242530 246119 242558 246753
rect 242626 246480 242880 246508
rect 242518 246113 242570 246119
rect 242518 246055 242570 246061
rect 242324 238530 242380 238539
rect 242324 238465 242380 238474
rect 242134 237973 242186 237979
rect 242134 237915 242186 237921
rect 242038 235161 242090 235167
rect 242038 235103 242090 235109
rect 241846 235087 241898 235093
rect 241846 235029 241898 235035
rect 242338 233484 242366 238465
rect 242626 238127 242654 246480
rect 243188 241046 243244 241055
rect 243188 240981 243244 240990
rect 242708 240750 242764 240759
rect 242708 240685 242764 240694
rect 242614 238121 242666 238127
rect 242614 238063 242666 238069
rect 242722 233484 242750 240685
rect 243092 237346 243148 237355
rect 243092 237281 243148 237290
rect 243106 233484 243134 237281
rect 242112 233456 242366 233484
rect 242496 233456 242750 233484
rect 242880 233456 243134 233484
rect 243202 233470 243230 240981
rect 243298 234945 243326 246494
rect 243572 238678 243628 238687
rect 243572 238613 243628 238622
rect 243286 234939 243338 234945
rect 243286 234881 243338 234887
rect 243586 233470 243614 238613
rect 243778 238201 243806 246494
rect 244162 242271 244190 246494
rect 244594 246212 244622 246494
rect 244834 246480 245088 246508
rect 244594 246184 244670 246212
rect 244150 242265 244202 242271
rect 244150 242207 244202 242213
rect 244532 241342 244588 241351
rect 244532 241277 244588 241286
rect 244150 239379 244202 239385
rect 244150 239321 244202 239327
rect 243766 238195 243818 238201
rect 243766 238137 243818 238143
rect 243956 237494 244012 237503
rect 243956 237429 244012 237438
rect 243970 233470 243998 237429
rect 244162 234871 244190 239321
rect 244150 234865 244202 234871
rect 244150 234807 244202 234813
rect 244546 233484 244574 241277
rect 244642 239163 244670 246184
rect 244726 241155 244778 241161
rect 244726 241097 244778 241103
rect 244630 239157 244682 239163
rect 244630 239099 244682 239105
rect 244738 233780 244766 241097
rect 244834 238275 244862 246480
rect 245410 243825 245438 246494
rect 245398 243819 245450 243825
rect 245398 243761 245450 243767
rect 245396 241786 245452 241795
rect 245396 241721 245452 241730
rect 244822 238269 244874 238275
rect 244822 238211 244874 238217
rect 245300 237198 245356 237207
rect 245300 237133 245356 237142
rect 244320 233456 244574 233484
rect 244690 233752 244766 233780
rect 244690 233470 244718 233752
rect 245314 233484 245342 237133
rect 245088 233456 245342 233484
rect 245410 233470 245438 241721
rect 245782 237677 245834 237683
rect 245782 237619 245834 237625
rect 245794 233470 245822 237619
rect 245890 237387 245918 246494
rect 246384 246480 246494 246508
rect 246262 239157 246314 239163
rect 246262 239099 246314 239105
rect 246166 237603 246218 237609
rect 246166 237545 246218 237551
rect 245878 237381 245930 237387
rect 245878 237323 245930 237329
rect 246178 233470 246206 237545
rect 246274 235389 246302 239099
rect 246262 235383 246314 235389
rect 246262 235325 246314 235331
rect 246466 235019 246494 246480
rect 246562 246480 246816 246508
rect 246946 246480 247200 246508
rect 246562 238423 246590 246480
rect 246740 241638 246796 241647
rect 246740 241573 246796 241582
rect 246550 238417 246602 238423
rect 246550 238359 246602 238365
rect 246454 235013 246506 235019
rect 246454 234955 246506 234961
rect 246754 233484 246782 241573
rect 246946 237757 246974 246480
rect 247222 246335 247274 246341
rect 247222 246277 247274 246283
rect 247234 246045 247262 246277
rect 247222 246039 247274 246045
rect 247222 245981 247274 245987
rect 247618 244177 247646 246494
rect 247426 244149 247646 244177
rect 247426 241383 247454 244149
rect 247508 242526 247564 242535
rect 247700 242526 247756 242535
rect 247508 242461 247510 242470
rect 247562 242461 247564 242470
rect 247618 242484 247700 242512
rect 247510 242429 247562 242435
rect 247618 242419 247646 242484
rect 247700 242461 247756 242470
rect 247606 242413 247658 242419
rect 247606 242355 247658 242361
rect 247414 241377 247466 241383
rect 247414 241319 247466 241325
rect 248098 240939 248126 246494
rect 248578 241901 248606 246494
rect 248674 246480 248928 246508
rect 249408 246480 249662 246508
rect 248566 241895 248618 241901
rect 248566 241837 248618 241843
rect 248086 240933 248138 240939
rect 248086 240875 248138 240881
rect 248674 240495 248702 246480
rect 249634 245379 249662 246480
rect 249622 245373 249674 245379
rect 249622 245315 249674 245321
rect 248662 240489 248714 240495
rect 248662 240431 248714 240437
rect 249718 240489 249770 240495
rect 249718 240431 249770 240437
rect 247700 240158 247756 240167
rect 247700 240093 247756 240102
rect 247714 238220 247742 240093
rect 247988 240010 248044 240019
rect 247988 239945 248044 239954
rect 247522 238192 247742 238220
rect 247126 237825 247178 237831
rect 247126 237767 247178 237773
rect 246934 237751 246986 237757
rect 246934 237693 246986 237699
rect 247138 233484 247166 237767
rect 247522 233484 247550 238192
rect 247606 237751 247658 237757
rect 247606 237693 247658 237699
rect 246528 233456 246782 233484
rect 246912 233456 247166 233484
rect 247296 233456 247550 233484
rect 247618 233470 247646 237693
rect 248002 233470 248030 239945
rect 248374 239823 248426 239829
rect 248374 239765 248426 239771
rect 248386 233470 248414 239765
rect 248950 238639 249002 238645
rect 248950 238581 249002 238587
rect 248962 233484 248990 238581
rect 249334 237899 249386 237905
rect 249334 237841 249386 237847
rect 249346 233484 249374 237841
rect 249730 233484 249758 240431
rect 249826 240421 249854 246494
rect 250306 245527 250334 246494
rect 250294 245521 250346 245527
rect 250294 245463 250346 245469
rect 250390 241377 250442 241383
rect 250390 241319 250442 241325
rect 250198 240563 250250 240569
rect 250198 240505 250250 240511
rect 249814 240415 249866 240421
rect 249814 240357 249866 240363
rect 249814 237973 249866 237979
rect 249814 237915 249866 237921
rect 248736 233456 248990 233484
rect 249120 233456 249374 233484
rect 249504 233456 249758 233484
rect 249826 233470 249854 237915
rect 250210 233470 250238 240505
rect 250402 235315 250430 241319
rect 250690 240865 250718 246494
rect 251136 246480 251390 246508
rect 251616 246480 251870 246508
rect 251362 245823 251390 246480
rect 251350 245817 251402 245823
rect 251350 245759 251402 245765
rect 250678 240859 250730 240865
rect 250678 240801 250730 240807
rect 251542 240859 251594 240865
rect 251542 240801 251594 240807
rect 250582 240637 250634 240643
rect 250582 240579 250634 240585
rect 250390 235309 250442 235315
rect 250390 235251 250442 235257
rect 250594 233470 250622 240579
rect 251158 238121 251210 238127
rect 251158 238063 251210 238069
rect 251170 233484 251198 238063
rect 251554 233484 251582 240801
rect 251842 240791 251870 246480
rect 251926 245151 251978 245157
rect 251926 245093 251978 245099
rect 251938 244861 251966 245093
rect 251926 244855 251978 244861
rect 251926 244797 251978 244803
rect 251830 240785 251882 240791
rect 251830 240727 251882 240733
rect 252034 240717 252062 246494
rect 252418 245305 252446 246494
rect 252514 246045 252542 246753
rect 252502 246039 252554 246045
rect 252502 245981 252554 245987
rect 252706 245897 252734 246753
rect 266722 246563 266750 246753
rect 268642 246711 268670 246753
rect 267478 246705 267530 246711
rect 267478 246647 267530 246653
rect 267574 246705 267626 246711
rect 267574 246647 267626 246653
rect 268630 246705 268682 246711
rect 268630 246647 268682 246653
rect 276694 246705 276746 246711
rect 276694 246647 276746 246653
rect 278806 246705 278858 246711
rect 278806 246647 278858 246653
rect 266614 246557 266666 246563
rect 252694 245891 252746 245897
rect 252694 245833 252746 245839
rect 252406 245299 252458 245305
rect 252406 245241 252458 245247
rect 252118 245003 252170 245009
rect 252118 244945 252170 244951
rect 252130 244787 252158 244945
rect 252118 244781 252170 244787
rect 252118 244723 252170 244729
rect 252790 241599 252842 241605
rect 252790 241541 252842 241547
rect 252310 240933 252362 240939
rect 252310 240875 252362 240881
rect 252022 240711 252074 240717
rect 252022 240653 252074 240659
rect 251926 238047 251978 238053
rect 251926 237989 251978 237995
rect 251938 233484 251966 237989
rect 252322 233484 252350 240875
rect 252406 238269 252458 238275
rect 252406 238211 252458 238217
rect 250944 233456 251198 233484
rect 251328 233456 251582 233484
rect 251712 233456 251966 233484
rect 252048 233456 252350 233484
rect 252418 233470 252446 238211
rect 252802 233470 252830 241541
rect 252898 241013 252926 246494
rect 253344 246480 253406 246508
rect 253378 245453 253406 246480
rect 253474 246480 253728 246508
rect 253366 245447 253418 245453
rect 253366 245389 253418 245395
rect 253366 243227 253418 243233
rect 253366 243169 253418 243175
rect 253378 243085 253406 243169
rect 253366 243079 253418 243085
rect 253366 243021 253418 243027
rect 252886 241007 252938 241013
rect 252886 240949 252938 240955
rect 253474 238349 253502 246480
rect 254146 245749 254174 246494
rect 254134 245743 254186 245749
rect 254134 245685 254186 245691
rect 254230 241303 254282 241309
rect 254230 241245 254282 241251
rect 253750 241229 253802 241235
rect 253750 241171 253802 241177
rect 253462 238343 253514 238349
rect 253462 238285 253514 238291
rect 253366 238195 253418 238201
rect 253366 238137 253418 238143
rect 253378 233484 253406 238137
rect 253762 233484 253790 241171
rect 254134 238417 254186 238423
rect 254134 238359 254186 238365
rect 254146 233484 254174 238359
rect 253152 233456 253406 233484
rect 253536 233456 253790 233484
rect 253920 233456 254174 233484
rect 254242 233470 254270 241245
rect 254626 241087 254654 246494
rect 255106 245897 255134 246494
rect 255202 246480 255456 246508
rect 255682 246480 255936 246508
rect 255094 245891 255146 245897
rect 255094 245833 255146 245839
rect 254998 241377 255050 241383
rect 254998 241319 255050 241325
rect 254614 241081 254666 241087
rect 254614 241023 254666 241029
rect 254614 238491 254666 238497
rect 254614 238433 254666 238439
rect 254626 233470 254654 238433
rect 255010 233470 255038 241319
rect 255094 241007 255146 241013
rect 255094 240949 255146 240955
rect 255106 240347 255134 240949
rect 255094 240341 255146 240347
rect 255094 240283 255146 240289
rect 255202 237313 255230 246480
rect 255682 239015 255710 246480
rect 256354 244121 256382 246494
rect 256534 244337 256586 244343
rect 256534 244279 256586 244285
rect 256342 244115 256394 244121
rect 256342 244057 256394 244063
rect 256066 243520 256286 243548
rect 256066 243423 256094 243520
rect 256258 243423 256286 243520
rect 256052 243414 256108 243423
rect 256052 243349 256108 243358
rect 256244 243414 256300 243423
rect 256244 243349 256300 243358
rect 256546 243275 256574 244279
rect 256244 243266 256300 243275
rect 256244 243201 256246 243210
rect 256298 243201 256300 243210
rect 256532 243266 256588 243275
rect 256532 243201 256588 243210
rect 256246 243169 256298 243175
rect 256340 243118 256396 243127
rect 256724 243118 256780 243127
rect 256546 243076 256724 243104
rect 256546 243067 256574 243076
rect 256396 243062 256574 243067
rect 256340 243053 256574 243062
rect 256724 243053 256780 243062
rect 256354 243039 256574 243053
rect 255958 241451 256010 241457
rect 255958 241393 256010 241399
rect 255670 239009 255722 239015
rect 255670 238951 255722 238957
rect 255574 238565 255626 238571
rect 255574 238507 255626 238513
rect 255190 237307 255242 237313
rect 255190 237249 255242 237255
rect 255586 233484 255614 238507
rect 255970 233484 255998 241393
rect 256438 239897 256490 239903
rect 256438 239839 256490 239845
rect 256246 238713 256298 238719
rect 256246 238655 256298 238661
rect 256258 233484 256286 238655
rect 255360 233456 255614 233484
rect 255744 233456 255998 233484
rect 256128 233456 256286 233484
rect 256450 233470 256478 239839
rect 256834 238867 256862 246494
rect 257232 246480 257342 246508
rect 257206 239675 257258 239681
rect 257206 239617 257258 239623
rect 256822 238861 256874 238867
rect 256822 238803 256874 238809
rect 257110 238861 257162 238867
rect 257110 238803 257162 238809
rect 257122 233484 257150 238803
rect 256848 233456 257150 233484
rect 257218 233470 257246 239617
rect 257314 235611 257342 246480
rect 257410 246480 257664 246508
rect 258144 246480 258398 246508
rect 257410 238941 257438 246480
rect 258370 244047 258398 246480
rect 258358 244041 258410 244047
rect 258358 243983 258410 243989
rect 258562 241531 258590 246494
rect 258550 241525 258602 241531
rect 258550 241467 258602 241473
rect 257878 240637 257930 240643
rect 257698 240585 257878 240588
rect 257698 240579 257930 240585
rect 257698 240560 257918 240579
rect 257698 240495 257726 240560
rect 257686 240489 257738 240495
rect 257686 240431 257738 240437
rect 257878 240489 257930 240495
rect 257878 240431 257930 240437
rect 257890 239829 257918 240431
rect 257878 239823 257930 239829
rect 257878 239765 257930 239771
rect 257398 238935 257450 238941
rect 257398 238877 257450 238883
rect 257782 238787 257834 238793
rect 257782 238729 257834 238735
rect 257302 235605 257354 235611
rect 257302 235547 257354 235553
rect 257794 233484 257822 238729
rect 258644 238382 258700 238391
rect 258550 238343 258602 238349
rect 258644 238317 258700 238326
rect 258550 238285 258602 238291
rect 258166 236641 258218 236647
rect 258166 236583 258218 236589
rect 258178 233484 258206 236583
rect 258562 233484 258590 238285
rect 257568 233456 257822 233484
rect 257952 233456 258206 233484
rect 258336 233456 258590 233484
rect 258658 233470 258686 238317
rect 258946 235759 258974 246494
rect 259028 240898 259084 240907
rect 259028 240833 259084 240842
rect 258934 235753 258986 235759
rect 258934 235695 258986 235701
rect 259042 233470 259070 240833
rect 259426 237461 259454 246494
rect 259872 246480 260126 246508
rect 260352 246480 260606 246508
rect 260098 244195 260126 246480
rect 260086 244189 260138 244195
rect 260086 244131 260138 244137
rect 259604 241194 259660 241203
rect 259604 241129 259660 241138
rect 259414 237455 259466 237461
rect 259414 237397 259466 237403
rect 259124 236754 259180 236763
rect 259124 236689 259180 236698
rect 259138 236319 259166 236689
rect 259124 236310 259180 236319
rect 259124 236245 259180 236254
rect 259618 233484 259646 241129
rect 260374 239009 260426 239015
rect 260374 238951 260426 238957
rect 259990 238935 260042 238941
rect 259990 238877 260042 238883
rect 260002 233484 260030 238877
rect 260386 233484 260414 238951
rect 260578 235537 260606 246480
rect 260674 241827 260702 246494
rect 260854 245077 260906 245083
rect 260854 245019 260906 245025
rect 260758 245003 260810 245009
rect 260758 244945 260810 244951
rect 260662 241821 260714 241827
rect 260662 241763 260714 241769
rect 260566 235531 260618 235537
rect 260566 235473 260618 235479
rect 260770 233484 260798 244945
rect 259440 233456 259646 233484
rect 259776 233456 260030 233484
rect 260160 233456 260414 233484
rect 260544 233456 260798 233484
rect 260866 233470 260894 245019
rect 261154 243973 261182 246494
rect 261142 243967 261194 243973
rect 261142 243909 261194 243915
rect 261236 241490 261292 241499
rect 261236 241425 261292 241434
rect 261250 233470 261278 241425
rect 261634 240273 261662 246494
rect 261970 246212 261998 246494
rect 261922 246184 261998 246212
rect 262210 246480 262464 246508
rect 261814 245151 261866 245157
rect 261814 245093 261866 245099
rect 261622 240267 261674 240273
rect 261622 240209 261674 240215
rect 261826 233484 261854 245093
rect 261922 235685 261950 246184
rect 262006 241747 262058 241753
rect 262006 241689 262058 241695
rect 261910 235679 261962 235685
rect 261910 235621 261962 235627
rect 262018 233484 262046 241689
rect 262102 240341 262154 240347
rect 262102 240283 262154 240289
rect 262114 236647 262142 240283
rect 262210 240125 262238 246480
rect 262582 246039 262634 246045
rect 262582 245981 262634 245987
rect 262198 240119 262250 240125
rect 262198 240061 262250 240067
rect 262102 236641 262154 236647
rect 262102 236583 262154 236589
rect 262594 233484 262622 245981
rect 262882 243159 262910 246494
rect 263062 245669 263114 245675
rect 263062 245611 263114 245617
rect 262870 243153 262922 243159
rect 262870 243095 262922 243101
rect 262964 240306 263020 240315
rect 262964 240241 263020 240250
rect 262978 233484 263006 240241
rect 261648 233456 261854 233484
rect 261984 233456 262046 233484
rect 262368 233456 262622 233484
rect 262752 233456 263006 233484
rect 263074 233470 263102 245611
rect 263362 240199 263390 246494
rect 263446 244485 263498 244491
rect 263446 244427 263498 244433
rect 263350 240193 263402 240199
rect 263350 240135 263402 240141
rect 263458 233470 263486 244427
rect 263746 235833 263774 246494
rect 263938 246480 264192 246508
rect 264418 246480 264672 246508
rect 263830 245965 263882 245971
rect 263830 245907 263882 245913
rect 263734 235827 263786 235833
rect 263734 235769 263786 235775
rect 263842 233470 263870 245907
rect 263938 240051 263966 246480
rect 264310 241747 264362 241753
rect 264310 241689 264362 241695
rect 263926 240045 263978 240051
rect 263926 239987 263978 239993
rect 264322 233484 264350 241689
rect 264418 241679 264446 246480
rect 264790 244411 264842 244417
rect 264790 244353 264842 244359
rect 264406 241673 264458 241679
rect 264406 241615 264458 241621
rect 264802 233484 264830 244353
rect 264886 236049 264938 236055
rect 264886 235991 264938 235997
rect 264192 233456 264350 233484
rect 264576 233456 264830 233484
rect 264898 233484 264926 235991
rect 265090 235981 265118 246494
rect 265270 242635 265322 242641
rect 265270 242577 265322 242583
rect 265078 235975 265130 235981
rect 265078 235917 265130 235923
rect 264898 233456 264960 233484
rect 265282 233470 265310 242577
rect 265474 235463 265502 246494
rect 265954 243307 265982 246494
rect 266146 246480 266400 246508
rect 266614 246499 266666 246505
rect 266710 246557 266762 246563
rect 266710 246499 266762 246505
rect 265942 243301 265994 243307
rect 265942 243243 265994 243249
rect 266038 243005 266090 243011
rect 266038 242947 266090 242953
rect 265654 236123 265706 236129
rect 265654 236065 265706 236071
rect 265462 235457 265514 235463
rect 265462 235399 265514 235405
rect 265666 233470 265694 236065
rect 266050 233470 266078 242947
rect 266146 235907 266174 246480
rect 266626 246119 266654 246499
rect 266880 246480 267134 246508
rect 266518 246113 266570 246119
rect 266518 246055 266570 246061
rect 266614 246113 266666 246119
rect 266614 246055 266666 246061
rect 266530 244639 266558 246055
rect 266518 244633 266570 244639
rect 266518 244575 266570 244581
rect 266614 242857 266666 242863
rect 266614 242799 266666 242805
rect 266134 235901 266186 235907
rect 266134 235843 266186 235849
rect 266626 233484 266654 242799
rect 267106 235907 267134 246480
rect 267202 244269 267230 246494
rect 267490 246397 267518 246647
rect 267586 246563 267614 246647
rect 269302 246631 269354 246637
rect 269302 246573 269354 246579
rect 267574 246557 267626 246563
rect 267958 246557 268010 246563
rect 267574 246499 267626 246505
rect 267696 246505 267958 246508
rect 267696 246499 268010 246505
rect 267696 246480 267998 246499
rect 268176 246480 268382 246508
rect 268512 246480 268766 246508
rect 268992 246480 269150 246508
rect 267490 246369 267902 246397
rect 267766 246335 267818 246341
rect 267766 246277 267818 246283
rect 267778 246193 267806 246277
rect 267874 246193 267902 246369
rect 267766 246187 267818 246193
rect 267766 246129 267818 246135
rect 267862 246187 267914 246193
rect 267862 246129 267914 246135
rect 268246 244707 268298 244713
rect 268246 244649 268298 244655
rect 267190 244263 267242 244269
rect 267190 244205 267242 244211
rect 268258 243899 268286 244649
rect 268150 243893 268202 243899
rect 268150 243835 268202 243841
rect 268246 243893 268298 243899
rect 268246 243835 268298 243841
rect 267382 243227 267434 243233
rect 267382 243169 267434 243175
rect 267094 235901 267146 235907
rect 267094 235843 267146 235849
rect 266998 234569 267050 234575
rect 266998 234511 267050 234517
rect 267010 233484 267038 234511
rect 267394 233484 267422 243169
rect 268162 242937 268190 243835
rect 268150 242931 268202 242937
rect 268150 242873 268202 242879
rect 267862 242487 267914 242493
rect 267862 242429 267914 242435
rect 267478 234421 267530 234427
rect 267478 234363 267530 234369
rect 266400 233456 266654 233484
rect 266784 233456 267038 233484
rect 267168 233456 267422 233484
rect 267490 233470 267518 234363
rect 267874 233470 267902 242429
rect 268246 239749 268298 239755
rect 268246 239691 268298 239697
rect 268258 233470 268286 239691
rect 268354 236351 268382 246480
rect 268738 239903 268766 246480
rect 268726 239897 268778 239903
rect 268726 239839 268778 239845
rect 268342 236345 268394 236351
rect 268342 236287 268394 236293
rect 268822 234125 268874 234131
rect 268822 234067 268874 234073
rect 268834 233484 268862 234067
rect 269122 233613 269150 246480
rect 269314 246193 269342 246573
rect 276706 246563 276734 246647
rect 276886 246631 276938 246637
rect 276886 246573 276938 246579
rect 277366 246631 277418 246637
rect 277366 246573 277418 246579
rect 278614 246631 278666 246637
rect 278818 246619 278846 246647
rect 278666 246591 278846 246619
rect 278614 246573 278666 246579
rect 276598 246557 276650 246563
rect 269302 246187 269354 246193
rect 269302 246129 269354 246135
rect 269206 242783 269258 242789
rect 269206 242725 269258 242731
rect 269110 233607 269162 233613
rect 269110 233549 269162 233555
rect 269218 233484 269246 242725
rect 269302 241599 269354 241605
rect 269302 241541 269354 241547
rect 269314 240273 269342 241541
rect 269302 240267 269354 240273
rect 269302 240209 269354 240215
rect 269300 239862 269356 239871
rect 269300 239797 269356 239806
rect 269314 239681 269342 239797
rect 269302 239675 269354 239681
rect 269302 239617 269354 239623
rect 269410 239607 269438 246494
rect 269686 242709 269738 242715
rect 269686 242651 269738 242657
rect 269398 239601 269450 239607
rect 269398 239543 269450 239549
rect 269590 234051 269642 234057
rect 269590 233993 269642 233999
rect 269602 233484 269630 233993
rect 268608 233456 268862 233484
rect 268992 233456 269246 233484
rect 269376 233456 269630 233484
rect 269698 233470 269726 242651
rect 269890 242567 269918 246494
rect 269878 242561 269930 242567
rect 269878 242503 269930 242509
rect 270274 239681 270302 246494
rect 270720 246480 270878 246508
rect 270850 243085 270878 246480
rect 270946 246480 271200 246508
rect 270838 243079 270890 243085
rect 270838 243021 270890 243027
rect 270946 239755 270974 246480
rect 271508 241342 271564 241351
rect 271508 241277 271564 241286
rect 271522 241055 271550 241277
rect 271316 241046 271372 241055
rect 271316 240981 271372 240990
rect 271508 241046 271564 241055
rect 271508 240981 271564 240990
rect 271330 240463 271358 240981
rect 271124 240454 271180 240463
rect 271124 240389 271180 240398
rect 271316 240454 271372 240463
rect 271316 240389 271372 240398
rect 270934 239749 270986 239755
rect 271138 239723 271166 240389
rect 270934 239691 270986 239697
rect 271124 239714 271180 239723
rect 270262 239675 270314 239681
rect 271124 239649 271180 239658
rect 270262 239617 270314 239623
rect 271030 239453 271082 239459
rect 271030 239395 271082 239401
rect 270070 233755 270122 233761
rect 270070 233697 270122 233703
rect 270082 233470 270110 233697
rect 270646 233681 270698 233687
rect 270646 233623 270698 233629
rect 270658 233484 270686 233623
rect 271042 233484 271070 239395
rect 271414 236271 271466 236277
rect 271414 236213 271466 236219
rect 271426 233484 271454 236213
rect 271618 234353 271646 246494
rect 272002 241753 272030 246494
rect 271990 241747 272042 241753
rect 271990 241689 272042 241695
rect 272482 240125 272510 246494
rect 272928 246480 273182 246508
rect 272854 246187 272906 246193
rect 272854 246129 272906 246135
rect 272866 244491 272894 246129
rect 272854 244485 272906 244491
rect 272854 244427 272906 244433
rect 273154 241087 273182 246480
rect 273394 246212 273422 246494
rect 273792 246480 274046 246508
rect 273394 246184 273470 246212
rect 273142 241081 273194 241087
rect 273142 241023 273194 241029
rect 272470 240119 272522 240125
rect 272470 240061 272522 240067
rect 272278 239675 272330 239681
rect 272278 239617 272330 239623
rect 271798 239231 271850 239237
rect 271798 239173 271850 239179
rect 271606 234347 271658 234353
rect 271606 234289 271658 234295
rect 271810 233484 271838 239173
rect 271894 236641 271946 236647
rect 271894 236583 271946 236589
rect 270480 233456 270686 233484
rect 270816 233456 271070 233484
rect 271200 233456 271454 233484
rect 271584 233456 271838 233484
rect 271906 233470 271934 236583
rect 272290 233470 272318 239617
rect 272662 239157 272714 239163
rect 272662 239099 272714 239105
rect 272674 233470 272702 239099
rect 273238 237307 273290 237313
rect 273238 237249 273290 237255
rect 273250 233484 273278 237249
rect 273442 236425 273470 246184
rect 273526 242413 273578 242419
rect 273526 242355 273578 242361
rect 273538 241901 273566 242355
rect 274018 241901 274046 246480
rect 273526 241895 273578 241901
rect 273526 241837 273578 241843
rect 274006 241895 274058 241901
rect 274006 241837 274058 241843
rect 274210 239829 274238 246494
rect 274390 240785 274442 240791
rect 274390 240727 274442 240733
rect 274486 240785 274538 240791
rect 274486 240727 274538 240733
rect 274198 239823 274250 239829
rect 274198 239765 274250 239771
rect 273526 239675 273578 239681
rect 273526 239617 273578 239623
rect 273430 236419 273482 236425
rect 273430 236361 273482 236367
rect 273538 233484 273566 239617
rect 274006 237233 274058 237239
rect 274006 237175 274058 237181
rect 274018 233484 274046 237175
rect 274102 236715 274154 236721
rect 274102 236657 274154 236663
rect 273024 233456 273278 233484
rect 273408 233456 273566 233484
rect 273792 233456 274046 233484
rect 274114 233470 274142 236657
rect 274402 235463 274430 240727
rect 274390 235457 274442 235463
rect 274390 235399 274442 235405
rect 274498 233470 274526 240727
rect 274690 240421 274718 246494
rect 275136 246480 275390 246508
rect 275520 246480 275774 246508
rect 274678 240415 274730 240421
rect 274678 240357 274730 240363
rect 275362 237535 275390 246480
rect 275746 240199 275774 246480
rect 275842 246480 276000 246508
rect 276598 246499 276650 246505
rect 276694 246557 276746 246563
rect 276694 246499 276746 246505
rect 275734 240193 275786 240199
rect 275734 240135 275786 240141
rect 275446 240045 275498 240051
rect 275446 239987 275498 239993
rect 275350 237529 275402 237535
rect 275350 237471 275402 237477
rect 274870 233903 274922 233909
rect 274870 233845 274922 233851
rect 274882 233470 274910 233845
rect 275458 233484 275486 239987
rect 275842 239755 275870 246480
rect 276310 244337 276362 244343
rect 276310 244279 276362 244285
rect 275926 244263 275978 244269
rect 275926 244205 275978 244211
rect 275830 239749 275882 239755
rect 275830 239691 275882 239697
rect 275830 237455 275882 237461
rect 275830 237397 275882 237403
rect 275842 233484 275870 237397
rect 275938 236499 275966 244205
rect 276322 243252 276350 244279
rect 276418 244269 276446 246494
rect 276610 244269 276638 246499
rect 276406 244263 276458 244269
rect 276406 244205 276458 244211
rect 276598 244263 276650 244269
rect 276598 244205 276650 244211
rect 276404 243266 276460 243275
rect 276322 243224 276404 243252
rect 276404 243201 276460 243210
rect 276310 239601 276362 239607
rect 276310 239543 276362 239549
rect 276214 239305 276266 239311
rect 276214 239247 276266 239253
rect 275926 236493 275978 236499
rect 275926 236435 275978 236441
rect 276226 233484 276254 239247
rect 275232 233456 275486 233484
rect 275616 233456 275870 233484
rect 276000 233456 276254 233484
rect 276322 233470 276350 239543
rect 276694 239379 276746 239385
rect 276694 239321 276746 239327
rect 276706 233470 276734 239321
rect 276802 237017 276830 246494
rect 276898 246489 276926 246573
rect 276886 246483 276938 246489
rect 276886 246425 276938 246431
rect 277078 239527 277130 239533
rect 277078 239469 277130 239475
rect 276790 237011 276842 237017
rect 276790 236953 276842 236959
rect 277090 233470 277118 239469
rect 277282 236869 277310 246494
rect 277378 246267 277406 246573
rect 278710 246557 278762 246563
rect 278626 246517 278710 246545
rect 277474 246480 277728 246508
rect 277858 246480 278208 246508
rect 277366 246261 277418 246267
rect 277366 246203 277418 246209
rect 277366 244559 277418 244565
rect 277366 244501 277418 244507
rect 277378 242641 277406 244501
rect 277366 242635 277418 242641
rect 277366 242577 277418 242583
rect 277474 240273 277502 246480
rect 277858 246101 277886 246480
rect 278038 246187 278090 246193
rect 278038 246129 278090 246135
rect 278134 246187 278186 246193
rect 278134 246129 278186 246135
rect 277666 246073 277886 246101
rect 277666 242919 277694 246073
rect 277750 246039 277802 246045
rect 277750 245981 277802 245987
rect 277762 245916 277790 245981
rect 278050 245971 278078 246129
rect 278038 245965 278090 245971
rect 277762 245888 277982 245916
rect 278038 245907 278090 245913
rect 277954 245675 277982 245888
rect 277942 245669 277994 245675
rect 278146 245620 278174 246129
rect 278626 246119 278654 246517
rect 278710 246499 278762 246505
rect 278614 246113 278666 246119
rect 278614 246055 278666 246061
rect 278710 246113 278762 246119
rect 278710 246055 278762 246061
rect 277942 245611 277994 245617
rect 277750 245595 277802 245601
rect 278050 245592 278174 245620
rect 278050 245583 278078 245592
rect 277802 245555 278078 245583
rect 277750 245537 277802 245543
rect 278722 245176 278750 246055
rect 278050 245148 278750 245176
rect 278050 244880 278078 245148
rect 277954 244852 278078 244880
rect 277954 244713 277982 244852
rect 277942 244707 277994 244713
rect 277942 244649 277994 244655
rect 278038 244707 278090 244713
rect 278038 244649 278090 244655
rect 277750 244633 277802 244639
rect 277750 244575 277802 244581
rect 277762 243011 277790 244575
rect 277846 244411 277898 244417
rect 277846 244353 277898 244359
rect 277858 243307 277886 244353
rect 277942 244337 277994 244343
rect 277942 244279 277994 244285
rect 277846 243301 277898 243307
rect 277846 243243 277898 243249
rect 277954 243159 277982 244279
rect 277942 243153 277994 243159
rect 277942 243095 277994 243101
rect 277750 243005 277802 243011
rect 277750 242947 277802 242953
rect 277846 243005 277898 243011
rect 277846 242947 277898 242953
rect 277858 242919 277886 242947
rect 277666 242891 277886 242919
rect 278050 242863 278078 244649
rect 278038 242857 278090 242863
rect 278038 242799 278090 242805
rect 278914 242771 278942 246776
rect 286100 246753 286156 246762
rect 286292 246818 286348 246827
rect 286292 246753 286348 246762
rect 288884 246818 288940 246827
rect 288884 246753 288940 246762
rect 291956 246818 292012 246827
rect 291956 246753 292012 246762
rect 292244 246818 292300 246827
rect 292244 246753 292300 246762
rect 292628 246818 292684 246827
rect 387380 246818 387436 246827
rect 292628 246753 292684 246762
rect 307906 246776 308256 246804
rect 362736 246776 362942 246804
rect 278818 242743 278942 242771
rect 277558 242561 277610 242567
rect 277846 242561 277898 242567
rect 277610 242509 277846 242512
rect 277558 242503 277898 242509
rect 277570 242484 277886 242503
rect 277748 241786 277804 241795
rect 277748 241721 277804 241730
rect 278134 241747 278186 241753
rect 277762 241351 277790 241721
rect 278134 241689 278186 241695
rect 277748 241342 277804 241351
rect 277748 241277 277804 241286
rect 278036 240750 278092 240759
rect 277570 240708 278036 240736
rect 277570 240463 277598 240708
rect 278036 240685 278092 240694
rect 277556 240454 277612 240463
rect 277556 240389 277612 240398
rect 278146 240347 278174 241689
rect 278230 241525 278282 241531
rect 278230 241467 278282 241473
rect 278134 240341 278186 240347
rect 278134 240283 278186 240289
rect 277462 240267 277514 240273
rect 277462 240209 277514 240215
rect 278242 239871 278270 241467
rect 278326 240341 278378 240347
rect 278326 240283 278378 240289
rect 278228 239862 278284 239871
rect 278228 239797 278284 239806
rect 278338 239681 278366 240283
rect 278326 239675 278378 239681
rect 278326 239617 278378 239623
rect 277654 239601 277706 239607
rect 277654 239543 277706 239549
rect 277940 239566 277996 239575
rect 277270 236863 277322 236869
rect 277270 236805 277322 236811
rect 277666 233484 277694 239543
rect 277940 239501 277996 239510
rect 277954 239459 277982 239501
rect 277942 239453 277994 239459
rect 277942 239395 277994 239401
rect 278038 239453 278090 239459
rect 278038 239395 278090 239401
rect 277846 238935 277898 238941
rect 277846 238877 277898 238883
rect 277858 237387 277886 238877
rect 277846 237381 277898 237387
rect 277846 237323 277898 237329
rect 278050 233484 278078 239395
rect 278518 238935 278570 238941
rect 278518 238877 278570 238883
rect 278422 236567 278474 236573
rect 278422 236509 278474 236515
rect 278434 233484 278462 236509
rect 277440 233456 277694 233484
rect 277824 233456 278078 233484
rect 278208 233456 278462 233484
rect 278530 233470 278558 238877
rect 278818 237091 278846 242743
rect 278902 239675 278954 239681
rect 278902 239617 278954 239623
rect 278806 237085 278858 237091
rect 278806 237027 278858 237033
rect 278914 233470 278942 239617
rect 279010 233484 279038 246494
rect 279382 243005 279434 243011
rect 279382 242947 279434 242953
rect 279394 233484 279422 242947
rect 279490 239977 279518 246494
rect 279682 246480 279936 246508
rect 280320 246480 280574 246508
rect 279478 239971 279530 239977
rect 279478 239913 279530 239919
rect 279682 239681 279710 246480
rect 280546 241087 280574 246480
rect 280438 241081 280490 241087
rect 280438 241023 280490 241029
rect 280534 241081 280586 241087
rect 280534 241023 280586 241029
rect 280450 239903 280478 241023
rect 280150 239897 280202 239903
rect 280150 239839 280202 239845
rect 280438 239897 280490 239903
rect 280438 239839 280490 239845
rect 279670 239675 279722 239681
rect 279670 239617 279722 239623
rect 279766 239675 279818 239681
rect 279766 239617 279818 239623
rect 279778 239575 279806 239617
rect 279764 239566 279820 239575
rect 279764 239501 279820 239510
rect 279766 236863 279818 236869
rect 279766 236805 279818 236811
rect 279778 233484 279806 236805
rect 280162 233484 280190 239839
rect 280534 239749 280586 239755
rect 280534 239691 280586 239697
rect 280546 233484 280574 239691
rect 280738 238941 280766 246494
rect 280918 239009 280970 239015
rect 280918 238951 280970 238957
rect 280726 238935 280778 238941
rect 280726 238877 280778 238883
rect 280930 238349 280958 238951
rect 280918 238343 280970 238349
rect 280918 238285 280970 238291
rect 281110 237529 281162 237535
rect 281110 237471 281162 237477
rect 279010 233456 279312 233484
rect 279394 233456 279648 233484
rect 279778 233456 280032 233484
rect 280162 233456 280416 233484
rect 280546 233456 280752 233484
rect 281122 233470 281150 237471
rect 281218 236573 281246 246494
rect 281602 246480 281712 246508
rect 281794 246480 282048 246508
rect 282528 246480 282782 246508
rect 281494 239823 281546 239829
rect 281494 239765 281546 239771
rect 281206 236567 281258 236573
rect 281206 236509 281258 236515
rect 281506 233470 281534 239765
rect 281602 236592 281630 246480
rect 281686 240193 281738 240199
rect 281686 240135 281738 240141
rect 281698 239681 281726 240135
rect 281686 239675 281738 239681
rect 281686 239617 281738 239623
rect 281794 239459 281822 246480
rect 282454 244633 282506 244639
rect 282274 244593 282454 244621
rect 282274 244565 282302 244593
rect 282454 244575 282506 244581
rect 282262 244559 282314 244565
rect 282262 244501 282314 244507
rect 281974 241895 282026 241901
rect 281974 241837 282026 241843
rect 281878 240785 281930 240791
rect 281878 240727 281930 240733
rect 281890 240199 281918 240727
rect 281878 240193 281930 240199
rect 281878 240135 281930 240141
rect 281986 239459 282014 241837
rect 282262 240785 282314 240791
rect 282262 240727 282314 240733
rect 282166 239971 282218 239977
rect 282166 239913 282218 239919
rect 282178 239755 282206 239913
rect 282166 239749 282218 239755
rect 282166 239691 282218 239697
rect 281782 239453 281834 239459
rect 281782 239395 281834 239401
rect 281974 239453 282026 239459
rect 281974 239395 282026 239401
rect 282274 238941 282302 240727
rect 282262 238935 282314 238941
rect 282262 238877 282314 238883
rect 281602 236564 281726 236592
rect 281590 236419 281642 236425
rect 281590 236361 281642 236367
rect 281602 233484 281630 236361
rect 281698 236203 281726 236564
rect 282754 236351 282782 246480
rect 282946 239607 282974 246494
rect 283222 243005 283274 243011
rect 283222 242947 283274 242953
rect 283030 239897 283082 239903
rect 283030 239839 283082 239845
rect 283042 239607 283070 239839
rect 282934 239601 282986 239607
rect 282934 239543 282986 239549
rect 283030 239601 283082 239607
rect 283030 239543 283082 239549
rect 282742 236345 282794 236351
rect 282742 236287 282794 236293
rect 281686 236197 281738 236203
rect 281686 236139 281738 236145
rect 282454 234643 282506 234649
rect 282454 234585 282506 234591
rect 282466 233484 282494 234585
rect 282838 234495 282890 234501
rect 282838 234437 282890 234443
rect 282850 233484 282878 234437
rect 283234 233484 283262 242947
rect 283426 239089 283454 246494
rect 283702 243301 283754 243307
rect 283702 243243 283754 243249
rect 283414 239083 283466 239089
rect 283414 239025 283466 239031
rect 283318 238343 283370 238349
rect 283318 238285 283370 238291
rect 281602 233456 281856 233484
rect 282240 233456 282494 233484
rect 282624 233456 282878 233484
rect 282960 233456 283262 233484
rect 283330 233470 283358 238285
rect 283714 233470 283742 243243
rect 283810 239533 283838 246494
rect 284256 246480 284414 246508
rect 283894 240415 283946 240421
rect 283894 240357 283946 240363
rect 284086 240415 284138 240421
rect 284086 240357 284138 240363
rect 283906 239533 283934 240357
rect 283990 240341 284042 240347
rect 283990 240283 284042 240289
rect 284002 239903 284030 240283
rect 283990 239897 284042 239903
rect 283990 239839 284042 239845
rect 284098 239829 284126 240357
rect 284086 239823 284138 239829
rect 284086 239765 284138 239771
rect 283798 239527 283850 239533
rect 283798 239469 283850 239475
rect 283894 239527 283946 239533
rect 283894 239469 283946 239475
rect 284386 238941 284414 246480
rect 284482 246480 284736 246508
rect 284482 239385 284510 246480
rect 284950 243153 285002 243159
rect 284950 243095 285002 243101
rect 284854 239971 284906 239977
rect 284854 239913 284906 239919
rect 284470 239379 284522 239385
rect 284470 239321 284522 239327
rect 284374 238935 284426 238941
rect 284374 238877 284426 238883
rect 284866 238349 284894 239913
rect 284854 238343 284906 238349
rect 284854 238285 284906 238291
rect 284662 234273 284714 234279
rect 284662 234215 284714 234221
rect 284278 234199 284330 234205
rect 284278 234141 284330 234147
rect 284290 233484 284318 234141
rect 284674 233484 284702 234215
rect 284962 233484 284990 243095
rect 285058 239385 285086 246494
rect 285552 246480 285854 246508
rect 285718 244781 285770 244787
rect 285718 244723 285770 244729
rect 285730 242715 285758 244723
rect 285526 242709 285578 242715
rect 285526 242651 285578 242657
rect 285718 242709 285770 242715
rect 285718 242651 285770 242657
rect 285538 242493 285566 242651
rect 285526 242487 285578 242493
rect 285526 242429 285578 242435
rect 285526 240119 285578 240125
rect 285526 240061 285578 240067
rect 285046 239379 285098 239385
rect 285046 239321 285098 239327
rect 285142 233977 285194 233983
rect 285142 233919 285194 233925
rect 284064 233456 284318 233484
rect 284448 233456 284702 233484
rect 284832 233456 284990 233484
rect 285154 233470 285182 233919
rect 285538 233470 285566 240061
rect 285826 238349 285854 246480
rect 285910 246113 285962 246119
rect 285910 246055 285962 246061
rect 285922 244787 285950 246055
rect 285910 244781 285962 244787
rect 285910 244723 285962 244729
rect 285910 242857 285962 242863
rect 285910 242799 285962 242805
rect 285814 238343 285866 238349
rect 285814 238285 285866 238291
rect 285922 233470 285950 242799
rect 286018 239311 286046 246494
rect 286114 246119 286142 246753
rect 286102 246113 286154 246119
rect 286102 246055 286154 246061
rect 286306 242493 286334 246753
rect 288022 246705 288074 246711
rect 288074 246665 288158 246693
rect 288022 246647 288074 246653
rect 286450 246212 286478 246494
rect 286402 246184 286478 246212
rect 286594 246480 286848 246508
rect 287280 246480 287390 246508
rect 286294 242487 286346 242493
rect 286294 242429 286346 242435
rect 286006 239305 286058 239311
rect 286006 239247 286058 239253
rect 286402 236943 286430 246184
rect 286486 242487 286538 242493
rect 286486 242429 286538 242435
rect 286390 236937 286442 236943
rect 286390 236879 286442 236885
rect 286498 233484 286526 242429
rect 286594 237461 286622 246480
rect 286870 241895 286922 241901
rect 286870 241837 286922 241843
rect 286582 237455 286634 237461
rect 286582 237397 286634 237403
rect 286882 233484 286910 241837
rect 287254 240341 287306 240347
rect 287254 240283 287306 240289
rect 287266 233484 287294 240283
rect 287362 239237 287390 246480
rect 287458 246480 287760 246508
rect 287458 240051 287486 246480
rect 287638 246261 287690 246267
rect 287638 246203 287690 246209
rect 287542 242931 287594 242937
rect 287542 242873 287594 242879
rect 287446 240045 287498 240051
rect 287446 239987 287498 239993
rect 287350 239231 287402 239237
rect 287350 239173 287402 239179
rect 287350 236567 287402 236573
rect 287350 236509 287402 236515
rect 286272 233456 286526 233484
rect 286656 233456 286910 233484
rect 287040 233456 287294 233484
rect 287362 233470 287390 236509
rect 287554 233484 287582 242873
rect 287650 239575 287678 246203
rect 288130 246193 288158 246665
rect 288898 246637 288926 246753
rect 288886 246631 288938 246637
rect 288886 246573 288938 246579
rect 288240 246480 288446 246508
rect 288576 246480 288638 246508
rect 289056 246480 289406 246508
rect 288118 246187 288170 246193
rect 288118 246129 288170 246135
rect 288214 244707 288266 244713
rect 287938 244667 288214 244695
rect 287938 243899 287966 244667
rect 288214 244649 288266 244655
rect 288022 244633 288074 244639
rect 288022 244575 288074 244581
rect 288034 243899 288062 244575
rect 287926 243893 287978 243899
rect 287926 243835 287978 243841
rect 288022 243893 288074 243899
rect 288022 243835 288074 243841
rect 287926 242413 287978 242419
rect 287842 242373 287926 242401
rect 287734 242339 287786 242345
rect 287734 242281 287786 242287
rect 287746 241943 287774 242281
rect 287732 241934 287788 241943
rect 287732 241869 287788 241878
rect 287842 239977 287870 242373
rect 287926 242355 287978 242361
rect 287830 239971 287882 239977
rect 287830 239913 287882 239919
rect 287636 239566 287692 239575
rect 287636 239501 287692 239510
rect 288418 238941 288446 246480
rect 288310 238935 288362 238941
rect 288310 238877 288362 238883
rect 288406 238935 288458 238941
rect 288406 238877 288458 238883
rect 288118 237529 288170 237535
rect 288118 237471 288170 237477
rect 288022 237455 288074 237461
rect 288022 237397 288074 237403
rect 287926 237381 287978 237387
rect 288034 237369 288062 237397
rect 287978 237341 288062 237369
rect 287926 237323 287978 237329
rect 287830 237307 287882 237313
rect 288130 237295 288158 237471
rect 287882 237267 288158 237295
rect 287830 237249 287882 237255
rect 288322 237165 288350 238877
rect 288310 237159 288362 237165
rect 288310 237101 288362 237107
rect 288214 236863 288266 236869
rect 288214 236805 288266 236811
rect 288226 236721 288254 236805
rect 288214 236715 288266 236721
rect 288214 236657 288266 236663
rect 288118 236419 288170 236425
rect 288118 236361 288170 236367
rect 287554 233456 287760 233484
rect 288130 233470 288158 236361
rect 288610 233909 288638 246480
rect 288694 240045 288746 240051
rect 288694 239987 288746 239993
rect 288598 233903 288650 233909
rect 288598 233845 288650 233851
rect 288706 233484 288734 239987
rect 289378 237387 289406 246480
rect 289474 240199 289502 246494
rect 289652 241342 289708 241351
rect 289652 241277 289708 241286
rect 289844 241342 289900 241351
rect 289844 241277 289900 241286
rect 289462 240193 289514 240199
rect 289462 240135 289514 240141
rect 289558 240119 289610 240125
rect 289558 240061 289610 240067
rect 289462 239823 289514 239829
rect 289462 239765 289514 239771
rect 289366 237381 289418 237387
rect 289366 237323 289418 237329
rect 288980 236310 289036 236319
rect 288980 236245 288982 236254
rect 289034 236245 289036 236254
rect 289078 236271 289130 236277
rect 288982 236213 289034 236219
rect 289078 236213 289130 236219
rect 289090 233484 289118 236213
rect 289474 233484 289502 239765
rect 288480 233456 288734 233484
rect 288864 233456 289118 233484
rect 289248 233456 289502 233484
rect 289570 233470 289598 240061
rect 289666 239871 289694 241277
rect 289858 240759 289886 241277
rect 289844 240750 289900 240759
rect 289844 240685 289900 240694
rect 289652 239862 289708 239871
rect 289652 239797 289708 239806
rect 289954 236869 289982 246494
rect 290146 246480 290352 246508
rect 290434 246480 290784 246508
rect 291264 246480 291518 246508
rect 290146 237313 290174 246480
rect 290434 240144 290462 246480
rect 291382 242931 291434 242937
rect 291382 242873 291434 242879
rect 291394 242715 291422 242873
rect 291382 242709 291434 242715
rect 291382 242651 291434 242657
rect 290614 241081 290666 241087
rect 290614 241023 290666 241029
rect 290242 240116 290462 240144
rect 290134 237307 290186 237313
rect 290134 237249 290186 237255
rect 290242 237239 290270 240116
rect 290422 239971 290474 239977
rect 290422 239913 290474 239919
rect 290434 239311 290462 239913
rect 290422 239305 290474 239311
rect 290422 239247 290474 239253
rect 290518 239305 290570 239311
rect 290518 239247 290570 239253
rect 290230 237233 290282 237239
rect 290230 237175 290282 237181
rect 290422 237159 290474 237165
rect 290422 237101 290474 237107
rect 289942 236863 289994 236869
rect 289942 236805 289994 236811
rect 290434 236721 290462 237101
rect 290422 236715 290474 236721
rect 290422 236657 290474 236663
rect 289942 236419 289994 236425
rect 289942 236361 289994 236367
rect 289954 233470 289982 236361
rect 290530 233484 290558 239247
rect 290626 237165 290654 241023
rect 291094 240193 291146 240199
rect 291094 240135 291146 240141
rect 290722 239524 291038 239552
rect 290614 237159 290666 237165
rect 290614 237101 290666 237107
rect 290722 236277 290750 239524
rect 291010 239459 291038 239524
rect 290806 239453 290858 239459
rect 290806 239395 290858 239401
rect 290998 239453 291050 239459
rect 290998 239395 291050 239401
rect 290818 236277 290846 239395
rect 291106 239163 291134 240135
rect 291490 239237 291518 246480
rect 291574 243079 291626 243085
rect 291574 243021 291626 243027
rect 291586 242715 291614 243021
rect 291574 242709 291626 242715
rect 291574 242651 291626 242657
rect 291682 239903 291710 246494
rect 291970 244565 291998 246753
rect 292080 246480 292190 246508
rect 292162 246175 292190 246480
rect 292258 246267 292286 246753
rect 292450 246480 292560 246508
rect 292246 246261 292298 246267
rect 292246 246203 292298 246209
rect 292342 246261 292394 246267
rect 292342 246203 292394 246209
rect 292354 246175 292382 246203
rect 292162 246147 292382 246175
rect 292450 245028 292478 246480
rect 292642 246119 292670 246753
rect 297922 246665 298142 246693
rect 296880 246628 297182 246656
rect 297922 246637 297950 246665
rect 292992 246480 293246 246508
rect 292630 246113 292682 246119
rect 292630 246055 292682 246061
rect 292726 246113 292778 246119
rect 292726 246055 292778 246061
rect 292066 245000 292478 245028
rect 291862 244559 291914 244565
rect 291862 244501 291914 244507
rect 291958 244559 292010 244565
rect 292066 244547 292094 245000
rect 292738 244787 292766 246055
rect 292726 244781 292778 244787
rect 292726 244723 292778 244729
rect 292822 244781 292874 244787
rect 292822 244723 292874 244729
rect 292066 244519 292382 244547
rect 291958 244501 292010 244507
rect 291874 244140 291902 244501
rect 291874 244112 292286 244140
rect 292258 243899 292286 244112
rect 292150 243893 292202 243899
rect 292150 243835 292202 243841
rect 292246 243893 292298 243899
rect 292246 243835 292298 243841
rect 291766 243079 291818 243085
rect 291766 243021 291818 243027
rect 291778 242567 291806 243021
rect 291766 242561 291818 242567
rect 291766 242503 291818 242509
rect 292162 242493 292190 243835
rect 292150 242487 292202 242493
rect 292150 242429 292202 242435
rect 291958 241081 292010 241087
rect 291958 241023 292010 241029
rect 291862 240045 291914 240051
rect 291862 239987 291914 239993
rect 291670 239897 291722 239903
rect 291670 239839 291722 239845
rect 291874 239829 291902 239987
rect 291862 239823 291914 239829
rect 291862 239765 291914 239771
rect 291478 239231 291530 239237
rect 291478 239173 291530 239179
rect 291094 239157 291146 239163
rect 291094 239099 291146 239105
rect 291970 237461 291998 241023
rect 292150 239601 292202 239607
rect 292150 239543 292202 239549
rect 291958 237455 292010 237461
rect 291958 237397 292010 237403
rect 291670 237233 291722 237239
rect 291670 237175 291722 237181
rect 291286 236789 291338 236795
rect 291286 236731 291338 236737
rect 290710 236271 290762 236277
rect 290710 236213 290762 236219
rect 290806 236271 290858 236277
rect 290806 236213 290858 236219
rect 290900 233498 290956 233507
rect 290352 233456 290558 233484
rect 290688 233456 290900 233484
rect 291298 233484 291326 236731
rect 291682 233484 291710 237175
rect 291766 236863 291818 236869
rect 291766 236805 291818 236811
rect 291072 233456 291326 233484
rect 291456 233456 291710 233484
rect 291778 233470 291806 236805
rect 292054 236641 292106 236647
rect 292054 236583 292106 236589
rect 291862 236567 291914 236573
rect 292066 236555 292094 236583
rect 291914 236527 292094 236555
rect 291862 236509 291914 236515
rect 292162 233470 292190 239543
rect 292354 237535 292382 244519
rect 292834 242937 292862 244723
rect 292822 242931 292874 242937
rect 292822 242873 292874 242879
rect 292918 242931 292970 242937
rect 292918 242873 292970 242879
rect 292930 242493 292958 242873
rect 292918 242487 292970 242493
rect 292918 242429 292970 242435
rect 293218 239681 293246 246480
rect 293314 246480 293376 246508
rect 293808 246480 294110 246508
rect 293314 240199 293342 246480
rect 293398 242709 293450 242715
rect 293398 242651 293450 242657
rect 293494 242709 293546 242715
rect 293494 242651 293546 242657
rect 293302 240193 293354 240199
rect 293302 240135 293354 240141
rect 293206 239675 293258 239681
rect 293206 239617 293258 239623
rect 293410 239427 293438 242651
rect 293396 239418 293452 239427
rect 293396 239353 293452 239362
rect 292342 237529 292394 237535
rect 292342 237471 292394 237477
rect 292534 233903 292586 233909
rect 292534 233845 292586 233851
rect 292546 233470 292574 233845
rect 293110 233829 293162 233835
rect 293110 233771 293162 233777
rect 293122 233484 293150 233771
rect 293506 233484 293534 242651
rect 293590 242487 293642 242493
rect 293590 242429 293642 242435
rect 292896 233456 293150 233484
rect 293280 233456 293534 233484
rect 293602 233484 293630 242429
rect 293782 240193 293834 240199
rect 293782 240135 293834 240141
rect 293794 239829 293822 240135
rect 293782 239823 293834 239829
rect 293782 239765 293834 239771
rect 293780 239566 293836 239575
rect 293780 239501 293836 239510
rect 293794 237535 293822 239501
rect 293972 239270 294028 239279
rect 293972 239205 294028 239214
rect 293986 239015 294014 239205
rect 294082 239015 294110 246480
rect 294166 246261 294218 246267
rect 294166 246203 294218 246209
rect 293974 239009 294026 239015
rect 293974 238951 294026 238957
rect 294070 239009 294122 239015
rect 294070 238951 294122 238957
rect 293782 237529 293834 237535
rect 293782 237471 293834 237477
rect 294178 237461 294206 246203
rect 294274 239829 294302 246494
rect 294466 246480 294768 246508
rect 295104 246480 295262 246508
rect 294262 239823 294314 239829
rect 294262 239765 294314 239771
rect 294358 239527 294410 239533
rect 294358 239469 294410 239475
rect 294166 237455 294218 237461
rect 294166 237397 294218 237403
rect 294068 236310 294124 236319
rect 293974 236271 294026 236277
rect 294068 236245 294070 236254
rect 293974 236213 294026 236219
rect 294122 236245 294124 236254
rect 294070 236213 294122 236219
rect 293602 233456 293664 233484
rect 293986 233470 294014 236213
rect 294370 233470 294398 239469
rect 294466 236573 294494 246480
rect 294550 246261 294602 246267
rect 294550 246203 294602 246209
rect 294562 242789 294590 246203
rect 294742 243079 294794 243085
rect 294742 243021 294794 243027
rect 294754 242956 294782 243021
rect 294754 242928 295166 242956
rect 295138 242863 295166 242928
rect 295126 242857 295178 242863
rect 294658 242789 295070 242808
rect 295126 242799 295178 242805
rect 294550 242783 294602 242789
rect 294550 242725 294602 242731
rect 294658 242783 295082 242789
rect 294658 242780 295030 242783
rect 294658 242715 294686 242780
rect 295030 242725 295082 242731
rect 294646 242709 294698 242715
rect 294646 242651 294698 242657
rect 295234 240144 295262 246480
rect 295426 246480 295584 246508
rect 295318 243079 295370 243085
rect 295318 243021 295370 243027
rect 295330 242641 295358 243021
rect 295318 242635 295370 242641
rect 295318 242577 295370 242583
rect 295138 240116 295262 240144
rect 294742 239601 294794 239607
rect 294742 239543 294794 239549
rect 294454 236567 294506 236573
rect 294454 236509 294506 236515
rect 294754 233470 294782 239543
rect 295138 238072 295166 240116
rect 295222 239971 295274 239977
rect 295426 239959 295454 246480
rect 295606 240267 295658 240273
rect 295606 240209 295658 240215
rect 295274 239931 295454 239959
rect 295222 239913 295274 239919
rect 295138 238044 295262 238072
rect 295030 237085 295082 237091
rect 295030 237027 295082 237033
rect 295042 236499 295070 237027
rect 295234 237017 295262 238044
rect 295126 237011 295178 237017
rect 295126 236953 295178 236959
rect 295222 237011 295274 237017
rect 295222 236953 295274 236959
rect 294838 236493 294890 236499
rect 294838 236435 294890 236441
rect 295030 236493 295082 236499
rect 295030 236435 295082 236441
rect 294850 233484 294878 236435
rect 295138 233780 295166 236953
rect 295138 233752 295262 233780
rect 295234 233484 295262 233752
rect 295618 233484 295646 240209
rect 296002 239607 296030 246494
rect 296278 240045 296330 240051
rect 296278 239987 296330 239993
rect 295990 239601 296042 239607
rect 295990 239543 296042 239549
rect 296290 239279 296318 239987
rect 296276 239270 296332 239279
rect 296276 239205 296332 239214
rect 296182 236493 296234 236499
rect 296182 236435 296234 236441
rect 294850 233456 295104 233484
rect 295234 233456 295488 233484
rect 295618 233456 295872 233484
rect 296194 233470 296222 236435
rect 296482 236277 296510 246494
rect 297154 240199 297182 246628
rect 297910 246631 297962 246637
rect 297910 246573 297962 246579
rect 298006 246631 298058 246637
rect 298006 246573 298058 246579
rect 297312 246480 297374 246508
rect 297346 240421 297374 246480
rect 297730 246480 297792 246508
rect 297622 242857 297674 242863
rect 297622 242799 297674 242805
rect 297334 240415 297386 240421
rect 297334 240357 297386 240363
rect 297142 240193 297194 240199
rect 297142 240135 297194 240141
rect 297634 239755 297662 242799
rect 297730 242549 297758 246480
rect 298018 246415 298046 246573
rect 298114 246415 298142 246665
rect 302422 246631 302474 246637
rect 302422 246573 302474 246579
rect 298224 246480 298526 246508
rect 298006 246409 298058 246415
rect 298006 246351 298058 246357
rect 298102 246409 298154 246415
rect 298102 246351 298154 246357
rect 298102 243301 298154 243307
rect 298102 243243 298154 243249
rect 298294 243301 298346 243307
rect 298294 243243 298346 243249
rect 298006 243153 298058 243159
rect 298006 243095 298058 243101
rect 298018 242863 298046 243095
rect 298006 242857 298058 242863
rect 298006 242799 298058 242805
rect 298114 242789 298142 243243
rect 297814 242783 297866 242789
rect 297814 242725 297866 242731
rect 298102 242783 298154 242789
rect 298102 242725 298154 242731
rect 297826 242660 297854 242725
rect 298306 242660 298334 243243
rect 297826 242632 298334 242660
rect 297730 242521 297854 242549
rect 297826 241901 297854 242521
rect 297718 241895 297770 241901
rect 297718 241837 297770 241843
rect 297814 241895 297866 241901
rect 297814 241837 297866 241843
rect 297730 240421 297758 241837
rect 297826 241448 298142 241476
rect 297826 241351 297854 241448
rect 297812 241342 297868 241351
rect 297812 241277 297868 241286
rect 298004 241342 298060 241351
rect 298004 241277 298060 241286
rect 298018 241055 298046 241277
rect 298004 241046 298060 241055
rect 298114 241032 298142 241448
rect 298196 241046 298252 241055
rect 298114 241004 298196 241032
rect 298004 240981 298060 240990
rect 298196 240981 298252 240990
rect 298004 240454 298060 240463
rect 297718 240415 297770 240421
rect 298004 240389 298060 240398
rect 297718 240357 297770 240363
rect 296566 239749 296618 239755
rect 296566 239691 296618 239697
rect 297622 239749 297674 239755
rect 298018 239723 298046 240389
rect 297622 239691 297674 239697
rect 298004 239714 298060 239723
rect 296470 236271 296522 236277
rect 296470 236213 296522 236219
rect 296578 233470 296606 239691
rect 298004 239649 298060 239658
rect 298390 239083 298442 239089
rect 298390 239025 298442 239031
rect 296950 237085 297002 237091
rect 296950 237027 297002 237033
rect 296962 233470 296990 237027
rect 297814 236345 297866 236351
rect 297814 236287 297866 236293
rect 297430 236197 297482 236203
rect 297430 236139 297482 236145
rect 297046 233607 297098 233613
rect 297046 233549 297098 233555
rect 297058 233484 297086 233549
rect 297442 233484 297470 236139
rect 297826 233484 297854 236287
rect 298198 233607 298250 233613
rect 298198 233549 298250 233555
rect 298210 233507 298238 233549
rect 298196 233498 298252 233507
rect 297058 233456 297312 233484
rect 297442 233456 297696 233484
rect 297826 233456 298080 233484
rect 290900 233433 290956 233442
rect 298402 233470 298430 239025
rect 298498 233687 298526 246480
rect 298594 233761 298622 246494
rect 298870 239379 298922 239385
rect 298870 239321 298922 239327
rect 298774 236715 298826 236721
rect 298774 236657 298826 236663
rect 298582 233755 298634 233761
rect 298582 233697 298634 233703
rect 298486 233681 298538 233687
rect 298486 233623 298538 233629
rect 298786 233470 298814 236657
rect 298882 233484 298910 239321
rect 299074 238349 299102 246494
rect 299266 246480 299520 246508
rect 300000 246480 300254 246508
rect 299266 246415 299294 246480
rect 299254 246409 299306 246415
rect 299254 246351 299306 246357
rect 299638 243301 299690 243307
rect 299638 243243 299690 243249
rect 299650 242641 299678 243243
rect 299638 242635 299690 242641
rect 299638 242577 299690 242583
rect 300022 239157 300074 239163
rect 300022 239099 300074 239105
rect 298966 238343 299018 238349
rect 298966 238285 299018 238291
rect 299062 238343 299114 238349
rect 299062 238285 299114 238291
rect 298978 238220 299006 238285
rect 298978 238192 299582 238220
rect 299554 233484 299582 238192
rect 299638 236937 299690 236943
rect 299638 236879 299690 236885
rect 298882 233456 299184 233484
rect 299520 233456 299582 233484
rect 299650 233484 299678 236879
rect 300034 233484 300062 239099
rect 300226 236573 300254 246480
rect 300214 236567 300266 236573
rect 300214 236509 300266 236515
rect 300322 234057 300350 246494
rect 300802 238941 300830 246494
rect 301282 246267 301310 246494
rect 301632 246480 301886 246508
rect 301270 246261 301322 246267
rect 301270 246203 301322 246209
rect 301366 246261 301418 246267
rect 301366 246203 301418 246209
rect 301378 244565 301406 246203
rect 301366 244559 301418 244565
rect 301366 244501 301418 244507
rect 301858 239755 301886 246480
rect 301954 246480 302112 246508
rect 301078 239749 301130 239755
rect 301078 239691 301130 239697
rect 301846 239749 301898 239755
rect 301846 239691 301898 239697
rect 300598 238935 300650 238941
rect 300598 238877 300650 238883
rect 300790 238935 300842 238941
rect 300790 238877 300842 238883
rect 300310 234051 300362 234057
rect 300310 233993 300362 233999
rect 299650 233456 299904 233484
rect 300034 233456 300288 233484
rect 300610 233470 300638 238877
rect 300982 237381 301034 237387
rect 300982 237323 301034 237329
rect 300994 233470 301022 237323
rect 301090 233484 301118 239691
rect 301846 239231 301898 239237
rect 301846 239173 301898 239179
rect 301462 237307 301514 237313
rect 301462 237249 301514 237255
rect 301474 233484 301502 237249
rect 301858 233484 301886 239173
rect 301954 234131 301982 246480
rect 302434 246415 302462 246573
rect 302422 246409 302474 246415
rect 302422 246351 302474 246357
rect 302326 244559 302378 244565
rect 302326 244501 302378 244507
rect 302338 242937 302366 244501
rect 302422 243301 302474 243307
rect 302422 243243 302474 243249
rect 302434 243011 302462 243243
rect 302422 243005 302474 243011
rect 302422 242947 302474 242953
rect 302326 242931 302378 242937
rect 302326 242873 302378 242879
rect 302530 239237 302558 246494
rect 303010 239681 303038 246494
rect 303394 243085 303422 246494
rect 303840 246480 304094 246508
rect 303382 243079 303434 243085
rect 303382 243021 303434 243027
rect 303478 243079 303530 243085
rect 303478 243021 303530 243027
rect 303094 242931 303146 242937
rect 303094 242873 303146 242879
rect 303106 240347 303134 242873
rect 303490 242419 303518 243021
rect 303478 242413 303530 242419
rect 303478 242355 303530 242361
rect 303094 240341 303146 240347
rect 303094 240283 303146 240289
rect 303574 239823 303626 239829
rect 303574 239765 303626 239771
rect 302806 239675 302858 239681
rect 302806 239617 302858 239623
rect 302998 239675 303050 239681
rect 302998 239617 303050 239623
rect 302518 239231 302570 239237
rect 302518 239173 302570 239179
rect 302230 237455 302282 237461
rect 302230 237397 302282 237403
rect 301942 234125 301994 234131
rect 301942 234067 301994 234073
rect 302242 233484 302270 237397
rect 301090 233456 301392 233484
rect 301474 233456 301728 233484
rect 301858 233456 302112 233484
rect 302242 233456 302496 233484
rect 302818 233470 302846 239617
rect 303190 239009 303242 239015
rect 303190 238951 303242 238957
rect 303202 233470 303230 238951
rect 303586 233470 303614 239765
rect 303670 237011 303722 237017
rect 303670 236953 303722 236959
rect 303682 233484 303710 236953
rect 304066 236721 304094 246480
rect 304306 246212 304334 246494
rect 304438 246483 304490 246489
rect 304438 246425 304490 246431
rect 304258 246184 304334 246212
rect 304150 239601 304202 239607
rect 304150 239543 304202 239549
rect 304054 236715 304106 236721
rect 304054 236657 304106 236663
rect 304162 233484 304190 239543
rect 304258 234427 304286 246184
rect 304450 246119 304478 246425
rect 304438 246113 304490 246119
rect 304438 246055 304490 246061
rect 304534 246113 304586 246119
rect 304534 246055 304586 246061
rect 304546 244565 304574 246055
rect 304534 244559 304586 244565
rect 304534 244501 304586 244507
rect 304438 240193 304490 240199
rect 304438 240135 304490 240141
rect 304246 234421 304298 234427
rect 304246 234363 304298 234369
rect 304450 233484 304478 240135
rect 304738 239015 304766 246494
rect 305122 243159 305150 246494
rect 305110 243153 305162 243159
rect 305110 243095 305162 243101
rect 305014 241895 305066 241901
rect 305014 241837 305066 241843
rect 304726 239009 304778 239015
rect 304726 238951 304778 238957
rect 303682 233456 303936 233484
rect 304162 233456 304320 233484
rect 304450 233456 304704 233484
rect 305026 233470 305054 241837
rect 305300 239418 305356 239427
rect 305300 239353 305356 239362
rect 305314 233484 305342 239353
rect 305602 233761 305630 246494
rect 305698 246480 306048 246508
rect 305698 234575 305726 246480
rect 306514 246212 306542 246494
rect 306658 246480 306912 246508
rect 306514 246184 306590 246212
rect 306454 243005 306506 243011
rect 306452 242970 306454 242979
rect 306506 242970 306508 242979
rect 306452 242905 306508 242914
rect 306562 240347 306590 246184
rect 306658 244639 306686 246480
rect 306646 244633 306698 244639
rect 306646 244575 306698 244581
rect 306742 244633 306794 244639
rect 306742 244575 306794 244581
rect 306754 244343 306782 244575
rect 306742 244337 306794 244343
rect 306742 244279 306794 244285
rect 307330 243899 307358 246494
rect 307318 243893 307370 243899
rect 307318 243835 307370 243841
rect 306550 240341 306602 240347
rect 306550 240283 306602 240289
rect 306646 239749 306698 239755
rect 306646 239691 306698 239697
rect 306262 238935 306314 238941
rect 306262 238877 306314 238883
rect 305782 238343 305834 238349
rect 305782 238285 305834 238291
rect 305878 238343 305930 238349
rect 305878 238285 305930 238291
rect 305686 234569 305738 234575
rect 305686 234511 305738 234517
rect 305590 233755 305642 233761
rect 305590 233697 305642 233703
rect 305314 233456 305424 233484
rect 305794 233470 305822 238285
rect 305890 237535 305918 238285
rect 305878 237529 305930 237535
rect 305878 237471 305930 237477
rect 305974 237529 306026 237535
rect 305974 237471 306026 237477
rect 305986 236795 306014 237471
rect 305974 236789 306026 236795
rect 305974 236731 306026 236737
rect 305878 236567 305930 236573
rect 305878 236509 305930 236515
rect 305890 233484 305918 236509
rect 306274 233484 306302 238877
rect 306658 233484 306686 239691
rect 307606 239675 307658 239681
rect 307606 239617 307658 239623
rect 307222 239231 307274 239237
rect 307222 239173 307274 239179
rect 305890 233456 306144 233484
rect 306274 233456 306528 233484
rect 306658 233456 306912 233484
rect 307234 233470 307262 239173
rect 307618 233470 307646 239617
rect 307810 239385 307838 246494
rect 307906 244491 307934 246776
rect 308470 246705 308522 246711
rect 350134 246705 350186 246711
rect 308470 246647 308522 246653
rect 308086 246631 308138 246637
rect 308086 246573 308138 246579
rect 308098 246341 308126 246573
rect 307990 246335 308042 246341
rect 307990 246277 308042 246283
rect 308086 246335 308138 246341
rect 308086 246277 308138 246283
rect 308002 246064 308030 246277
rect 308482 246193 308510 246647
rect 334870 246631 334922 246637
rect 334870 246573 334922 246579
rect 334966 246631 335018 246637
rect 335232 246628 335486 246656
rect 350134 246647 350186 246653
rect 352342 246705 352394 246711
rect 352342 246647 352394 246653
rect 362614 246705 362666 246711
rect 362614 246647 362666 246653
rect 334966 246573 335018 246579
rect 308640 246480 308894 246508
rect 308470 246187 308522 246193
rect 308470 246129 308522 246135
rect 308566 246187 308618 246193
rect 308566 246129 308618 246135
rect 308578 246064 308606 246129
rect 308002 246036 308606 246064
rect 307894 244485 307946 244491
rect 307894 244427 307946 244433
rect 308278 244485 308330 244491
rect 308278 244427 308330 244433
rect 307894 239675 307946 239681
rect 307894 239617 307946 239623
rect 307906 239459 307934 239617
rect 307894 239453 307946 239459
rect 307894 239395 307946 239401
rect 307798 239379 307850 239385
rect 307798 239321 307850 239327
rect 308182 239009 308234 239015
rect 308182 238951 308234 238957
rect 307990 236715 308042 236721
rect 307990 236657 308042 236663
rect 308002 233470 308030 236657
rect 308194 233484 308222 238951
rect 308290 236129 308318 244427
rect 308866 239607 308894 246480
rect 308962 246480 309120 246508
rect 308962 246119 308990 246480
rect 308950 246113 309002 246119
rect 308950 246055 309002 246061
rect 308950 242413 309002 242419
rect 308950 242355 309002 242361
rect 308962 241943 308990 242355
rect 308948 241934 309004 241943
rect 308948 241869 309004 241878
rect 308950 240341 309002 240347
rect 308950 240283 309002 240289
rect 308854 239601 308906 239607
rect 308854 239543 308906 239549
rect 308278 236123 308330 236129
rect 308278 236065 308330 236071
rect 308710 233755 308762 233761
rect 308710 233697 308762 233703
rect 308194 233456 308352 233484
rect 308722 233470 308750 233697
rect 308962 233484 308990 240283
rect 309538 239681 309566 246494
rect 309526 239675 309578 239681
rect 309526 239617 309578 239623
rect 309814 239379 309866 239385
rect 309814 239321 309866 239327
rect 309430 234347 309482 234353
rect 309430 234289 309482 234295
rect 308962 233456 309120 233484
rect 309442 233470 309470 234289
rect 309826 233470 309854 239321
rect 309922 236055 309950 246494
rect 310416 246480 310718 246508
rect 310486 244411 310538 244417
rect 310486 244353 310538 244359
rect 310498 243159 310526 244353
rect 310486 243153 310538 243159
rect 310486 243095 310538 243101
rect 310484 242526 310540 242535
rect 310210 242484 310484 242512
rect 310210 242387 310238 242484
rect 310484 242461 310540 242470
rect 310196 242378 310252 242387
rect 310196 242313 310252 242322
rect 310294 239675 310346 239681
rect 310294 239617 310346 239623
rect 310198 239601 310250 239607
rect 310198 239543 310250 239549
rect 309910 236049 309962 236055
rect 309910 235991 309962 235997
rect 310210 233470 310238 239543
rect 310306 233484 310334 239617
rect 310690 233484 310718 246480
rect 310834 246212 310862 246494
rect 310786 246184 310862 246212
rect 311266 246480 311328 246508
rect 311458 246480 311664 246508
rect 310786 244565 310814 246184
rect 310774 244559 310826 244565
rect 310774 244501 310826 244507
rect 311266 233484 311294 246480
rect 311458 236647 311486 246480
rect 312022 244559 312074 244565
rect 312022 244501 312074 244507
rect 311638 239009 311690 239015
rect 311638 238951 311690 238957
rect 311446 236641 311498 236647
rect 311446 236583 311498 236589
rect 310306 233456 310560 233484
rect 310690 233456 310944 233484
rect 311266 233456 311328 233484
rect 311650 233470 311678 238951
rect 312034 233470 312062 244501
rect 312130 240273 312158 246494
rect 312406 246483 312458 246489
rect 312406 246425 312458 246431
rect 312418 246119 312446 246425
rect 312406 246113 312458 246119
rect 312406 246055 312458 246061
rect 312214 244485 312266 244491
rect 312214 244427 312266 244433
rect 312226 243307 312254 244427
rect 312406 244337 312458 244343
rect 312406 244279 312458 244285
rect 312214 243301 312266 243307
rect 312214 243243 312266 243249
rect 312118 240267 312170 240273
rect 312118 240209 312170 240215
rect 312418 233470 312446 244279
rect 312610 242937 312638 246494
rect 312802 246480 313056 246508
rect 313186 246480 313440 246508
rect 312598 242931 312650 242937
rect 312598 242873 312650 242879
rect 312802 239755 312830 246480
rect 313186 240421 313214 246480
rect 313366 243893 313418 243899
rect 313366 243835 313418 243841
rect 313174 240415 313226 240421
rect 313174 240357 313226 240363
rect 312790 239749 312842 239755
rect 312790 239691 312842 239697
rect 312982 236049 313034 236055
rect 312982 235991 313034 235997
rect 312994 233484 313022 235991
rect 313378 233484 313406 243835
rect 313654 240341 313706 240347
rect 313654 240283 313706 240289
rect 313666 236647 313694 240283
rect 313750 240193 313802 240199
rect 313750 240135 313802 240141
rect 313654 236641 313706 236647
rect 313654 236583 313706 236589
rect 313762 233484 313790 240135
rect 313858 239903 313886 246494
rect 314338 242567 314366 246494
rect 314326 242561 314378 242567
rect 314326 242503 314378 242509
rect 314614 240267 314666 240273
rect 314614 240209 314666 240215
rect 314230 240119 314282 240125
rect 314230 240061 314282 240067
rect 313846 239897 313898 239903
rect 313846 239839 313898 239845
rect 313846 236641 313898 236647
rect 313846 236583 313898 236589
rect 312768 233456 313022 233484
rect 313152 233456 313406 233484
rect 313536 233456 313790 233484
rect 313858 233470 313886 236583
rect 314242 233470 314270 240061
rect 314626 233470 314654 240209
rect 314818 239977 314846 246494
rect 314914 246480 315168 246508
rect 315394 246480 315648 246508
rect 314914 242715 314942 246480
rect 314996 242822 315052 242831
rect 314996 242757 315052 242766
rect 315010 242715 315038 242757
rect 314902 242709 314954 242715
rect 314902 242651 314954 242657
rect 314998 242709 315050 242715
rect 314998 242651 315050 242657
rect 315190 240415 315242 240421
rect 315190 240357 315242 240363
rect 314806 239971 314858 239977
rect 314806 239913 314858 239919
rect 315202 233484 315230 240357
rect 315394 236277 315422 246480
rect 315574 239823 315626 239829
rect 315574 239765 315626 239771
rect 315382 236271 315434 236277
rect 315382 236213 315434 236219
rect 315586 233484 315614 239765
rect 316066 239311 316094 246494
rect 316162 246480 316464 246508
rect 316054 239305 316106 239311
rect 316054 239247 316106 239253
rect 315958 238639 316010 238645
rect 315958 238581 316010 238587
rect 316054 238639 316106 238645
rect 316054 238581 316106 238587
rect 315970 237091 315998 238581
rect 315958 237085 316010 237091
rect 315958 237027 316010 237033
rect 315958 236271 316010 236277
rect 315958 236213 316010 236219
rect 315970 233484 315998 236213
rect 314976 233456 315230 233484
rect 315360 233456 315614 233484
rect 315744 233456 315998 233484
rect 316066 233470 316094 238581
rect 316162 233983 316190 246480
rect 316532 243266 316588 243275
rect 316532 243201 316588 243210
rect 316546 242937 316574 243201
rect 316726 243005 316778 243011
rect 316724 242970 316726 242979
rect 316778 242970 316780 242979
rect 316534 242931 316586 242937
rect 316724 242905 316780 242914
rect 316534 242873 316586 242879
rect 316724 242822 316780 242831
rect 316724 242757 316780 242766
rect 316738 242715 316766 242757
rect 316726 242709 316778 242715
rect 316726 242651 316778 242657
rect 316438 238935 316490 238941
rect 316438 238877 316490 238883
rect 316150 233977 316202 233983
rect 316150 233919 316202 233925
rect 316450 233470 316478 238877
rect 316822 237455 316874 237461
rect 316822 237397 316874 237403
rect 316834 233470 316862 237397
rect 316930 233687 316958 246494
rect 317122 246480 317376 246508
rect 317602 246480 317856 246508
rect 317986 246480 318192 246508
rect 318466 246480 318672 246508
rect 317122 242863 317150 246480
rect 317110 242857 317162 242863
rect 317110 242799 317162 242805
rect 317494 242561 317546 242567
rect 317494 242503 317546 242509
rect 317398 237381 317450 237387
rect 317398 237323 317450 237329
rect 316918 233681 316970 233687
rect 316918 233623 316970 233629
rect 317410 233484 317438 237323
rect 317506 234279 317534 242503
rect 317602 237535 317630 246480
rect 317986 242567 318014 246480
rect 318262 244263 318314 244269
rect 318262 244205 318314 244211
rect 318070 244189 318122 244195
rect 318070 244131 318122 244137
rect 318082 243011 318110 244131
rect 318166 243967 318218 243973
rect 318166 243909 318218 243915
rect 318178 243233 318206 243909
rect 318274 243307 318302 244205
rect 318262 243301 318314 243307
rect 318262 243243 318314 243249
rect 318166 243227 318218 243233
rect 318166 243169 318218 243175
rect 318070 243005 318122 243011
rect 318070 242947 318122 242953
rect 317974 242561 318026 242567
rect 317974 242503 318026 242509
rect 317878 241895 317930 241901
rect 317878 241837 317930 241843
rect 317890 241013 317918 241837
rect 318260 241786 318316 241795
rect 318260 241721 318316 241730
rect 317974 241599 318026 241605
rect 317974 241541 318026 241547
rect 317878 241007 317930 241013
rect 317878 240949 317930 240955
rect 317878 239971 317930 239977
rect 317878 239913 317930 239919
rect 317590 237529 317642 237535
rect 317590 237471 317642 237477
rect 317686 237529 317738 237535
rect 317686 237471 317738 237477
rect 317698 237239 317726 237471
rect 317782 237307 317834 237313
rect 317782 237249 317834 237255
rect 317686 237233 317738 237239
rect 317686 237175 317738 237181
rect 317494 234273 317546 234279
rect 317494 234215 317546 234221
rect 317794 233484 317822 237249
rect 317184 233456 317438 233484
rect 317568 233456 317822 233484
rect 317890 233484 317918 239913
rect 317986 239311 318014 241541
rect 318166 241525 318218 241531
rect 318166 241467 318218 241473
rect 318070 241451 318122 241457
rect 318070 241393 318122 241399
rect 317974 239305 318026 239311
rect 317974 239247 318026 239253
rect 318082 239163 318110 241393
rect 318178 241013 318206 241467
rect 318166 241007 318218 241013
rect 318166 240949 318218 240955
rect 318274 239871 318302 241721
rect 318358 241377 318410 241383
rect 318358 241319 318410 241325
rect 318260 239862 318316 239871
rect 318260 239797 318316 239806
rect 318070 239157 318122 239163
rect 318070 239099 318122 239105
rect 318370 239089 318398 241319
rect 318358 239083 318410 239089
rect 318358 239025 318410 239031
rect 318358 238861 318410 238867
rect 318358 238803 318410 238809
rect 318166 238787 318218 238793
rect 318166 238729 318218 238735
rect 318070 238565 318122 238571
rect 318070 238507 318122 238513
rect 318082 236351 318110 238507
rect 318178 237239 318206 238729
rect 318262 238713 318314 238719
rect 318262 238655 318314 238661
rect 318166 237233 318218 237239
rect 318166 237175 318218 237181
rect 318274 237165 318302 238655
rect 318370 238571 318398 238803
rect 318358 238565 318410 238571
rect 318358 238507 318410 238513
rect 318466 237535 318494 246480
rect 318646 238861 318698 238867
rect 318646 238803 318698 238809
rect 318454 237529 318506 237535
rect 318454 237471 318506 237477
rect 318550 237529 318602 237535
rect 318550 237471 318602 237477
rect 318262 237159 318314 237165
rect 318262 237101 318314 237107
rect 318070 236345 318122 236351
rect 318070 236287 318122 236293
rect 318562 233484 318590 237471
rect 317890 233456 317952 233484
rect 318288 233456 318590 233484
rect 318658 233470 318686 238803
rect 319030 238713 319082 238719
rect 319030 238655 319082 238661
rect 319042 233470 319070 238655
rect 319138 234205 319166 246494
rect 319330 246480 319584 246508
rect 319968 246480 320126 246508
rect 319330 236795 319358 246480
rect 319810 244861 320030 244880
rect 319798 244855 320042 244861
rect 319850 244852 319990 244855
rect 319798 244797 319850 244803
rect 319990 244797 320042 244803
rect 319702 244633 319754 244639
rect 319702 244575 319754 244581
rect 319714 242715 319742 244575
rect 319798 244485 319850 244491
rect 319894 244485 319946 244491
rect 319850 244445 319894 244473
rect 319798 244427 319850 244433
rect 319894 244427 319946 244433
rect 320098 242789 320126 246480
rect 320386 243085 320414 246494
rect 320578 246480 320880 246508
rect 320374 243079 320426 243085
rect 320374 243021 320426 243027
rect 320086 242783 320138 242789
rect 320086 242725 320138 242731
rect 319702 242709 319754 242715
rect 319702 242651 319754 242657
rect 320470 241599 320522 241605
rect 320470 241541 320522 241547
rect 319510 241525 319562 241531
rect 319510 241467 319562 241473
rect 319522 237313 319550 241467
rect 319606 238639 319658 238645
rect 319606 238581 319658 238587
rect 319510 237307 319562 237313
rect 319510 237249 319562 237255
rect 319318 236789 319370 236795
rect 319318 236731 319370 236737
rect 319126 234199 319178 234205
rect 319126 234141 319178 234147
rect 319618 233484 319646 238581
rect 319702 237529 319754 237535
rect 319754 237489 319934 237517
rect 319702 237471 319754 237477
rect 319906 237480 319934 237489
rect 319906 237461 320030 237480
rect 319906 237455 320042 237461
rect 319906 237452 319990 237455
rect 319990 237397 320042 237403
rect 319894 237307 319946 237313
rect 319894 237249 319946 237255
rect 319906 237059 319934 237249
rect 319892 237050 319948 237059
rect 319892 236985 319948 236994
rect 320374 236493 320426 236499
rect 320374 236435 320426 236441
rect 319990 236419 320042 236425
rect 319990 236361 320042 236367
rect 320002 233484 320030 236361
rect 320386 233484 320414 236435
rect 319392 233456 319646 233484
rect 319776 233456 320030 233484
rect 320160 233456 320414 233484
rect 320482 233470 320510 241541
rect 320578 233909 320606 246480
rect 321346 244491 321374 246494
rect 321442 246480 321696 246508
rect 321922 246480 322176 246508
rect 321334 244485 321386 244491
rect 321334 244427 321386 244433
rect 320854 239675 320906 239681
rect 320854 239617 320906 239623
rect 320566 233903 320618 233909
rect 320566 233845 320618 233851
rect 320866 233470 320894 239617
rect 321238 239379 321290 239385
rect 321238 239321 321290 239327
rect 321250 233470 321278 239321
rect 321442 233835 321470 246480
rect 321814 237307 321866 237313
rect 321814 237249 321866 237255
rect 321430 233829 321482 233835
rect 321430 233771 321482 233777
rect 321826 233484 321854 237249
rect 321922 234501 321950 246480
rect 322006 246409 322058 246415
rect 322006 246351 322058 246357
rect 322018 246193 322046 246351
rect 322006 246187 322058 246193
rect 322006 246129 322058 246135
rect 322594 242641 322622 246494
rect 322786 246480 323088 246508
rect 322582 242635 322634 242641
rect 322582 242577 322634 242583
rect 322678 239749 322730 239755
rect 322678 239691 322730 239697
rect 322198 239527 322250 239533
rect 322198 239469 322250 239475
rect 321910 234495 321962 234501
rect 321910 234437 321962 234443
rect 322210 233484 322238 239469
rect 322486 236567 322538 236573
rect 322486 236509 322538 236515
rect 322498 233484 322526 236509
rect 321600 233456 321854 233484
rect 321984 233456 322238 233484
rect 322368 233456 322526 233484
rect 322690 233470 322718 239691
rect 322786 234649 322814 246480
rect 323458 242493 323486 246494
rect 323650 246480 323904 246508
rect 324130 246480 324384 246508
rect 323446 242487 323498 242493
rect 323446 242429 323498 242435
rect 323062 239601 323114 239607
rect 323062 239543 323114 239549
rect 322774 234643 322826 234649
rect 322774 234585 322826 234591
rect 323074 233470 323102 239543
rect 323446 239453 323498 239459
rect 323446 239395 323498 239401
rect 323458 233470 323486 239395
rect 323650 239015 323678 246480
rect 323638 239009 323690 239015
rect 323638 238951 323690 238957
rect 323734 239009 323786 239015
rect 323734 238951 323786 238957
rect 323746 238793 323774 238951
rect 323734 238787 323786 238793
rect 323734 238729 323786 238735
rect 324130 238571 324158 246480
rect 324406 239897 324458 239903
rect 324406 239839 324458 239845
rect 324118 238565 324170 238571
rect 324118 238507 324170 238513
rect 324022 236863 324074 236869
rect 324022 236805 324074 236811
rect 324034 233484 324062 236805
rect 324418 233484 324446 239839
rect 324706 239681 324734 246494
rect 325076 242970 325132 242979
rect 325076 242905 325078 242914
rect 325130 242905 325132 242914
rect 325078 242873 325130 242879
rect 325186 241679 325214 246494
rect 325474 246480 325680 246508
rect 325858 246480 326112 246508
rect 326496 246480 326750 246508
rect 325174 241673 325226 241679
rect 325174 241615 325226 241621
rect 325270 241673 325322 241679
rect 325270 241615 325322 241621
rect 325282 239829 325310 241615
rect 325270 239823 325322 239829
rect 325270 239765 325322 239771
rect 324694 239675 324746 239681
rect 324694 239617 324746 239623
rect 325474 239108 325502 246480
rect 325186 239080 325502 239108
rect 324790 236789 324842 236795
rect 324790 236731 324842 236737
rect 324802 233484 324830 236731
rect 325186 233484 325214 239080
rect 325858 237091 325886 246480
rect 326722 241383 326750 246480
rect 326710 241377 326762 241383
rect 326710 241319 326762 241325
rect 326914 241161 326942 246494
rect 327394 241457 327422 246494
rect 327874 241901 327902 246494
rect 327970 246480 328224 246508
rect 328450 246480 328704 246508
rect 327862 241895 327914 241901
rect 327862 241837 327914 241843
rect 327970 241827 327998 246480
rect 328150 242561 328202 242567
rect 328148 242526 328150 242535
rect 328202 242526 328204 242535
rect 328148 242461 328204 242470
rect 328054 241895 328106 241901
rect 328054 241837 328106 241843
rect 327958 241821 328010 241827
rect 327958 241763 328010 241769
rect 327862 241673 327914 241679
rect 328066 241624 328094 241837
rect 327914 241621 328094 241624
rect 327862 241615 328094 241621
rect 327874 241596 328094 241615
rect 327382 241451 327434 241457
rect 327382 241393 327434 241399
rect 326902 241155 326954 241161
rect 326902 241097 326954 241103
rect 326998 241155 327050 241161
rect 326998 241097 327050 241103
rect 327010 239977 327038 241097
rect 326998 239971 327050 239977
rect 326998 239913 327050 239919
rect 328246 239971 328298 239977
rect 328246 239913 328298 239919
rect 326230 239823 326282 239829
rect 326230 239765 326282 239771
rect 325846 237085 325898 237091
rect 325846 237027 325898 237033
rect 325654 236715 325706 236721
rect 325654 236657 325706 236663
rect 325270 236641 325322 236647
rect 325270 236583 325322 236589
rect 323808 233456 324062 233484
rect 324192 233456 324446 233484
rect 324576 233456 324830 233484
rect 324912 233456 325214 233484
rect 325282 233470 325310 236583
rect 325666 233470 325694 236657
rect 326242 233484 326270 239765
rect 326998 239749 327050 239755
rect 326998 239691 327050 239697
rect 326614 239231 326666 239237
rect 326614 239173 326666 239179
rect 326626 233484 326654 239173
rect 327010 233484 327038 239691
rect 327478 237085 327530 237091
rect 327478 237027 327530 237033
rect 327094 237011 327146 237017
rect 327094 236953 327146 236959
rect 326016 233456 326270 233484
rect 326400 233456 326654 233484
rect 326784 233456 327038 233484
rect 327106 233470 327134 236953
rect 327490 233470 327518 237027
rect 327862 236937 327914 236943
rect 327862 236879 327914 236885
rect 327874 233470 327902 236879
rect 328258 233484 328286 239913
rect 328450 236277 328478 246480
rect 328534 242561 328586 242567
rect 328534 242503 328586 242509
rect 328546 242387 328574 242503
rect 328532 242378 328588 242387
rect 328532 242313 328588 242322
rect 328726 241821 328778 241827
rect 328726 241763 328778 241769
rect 328738 237165 328766 241763
rect 328918 241377 328970 241383
rect 328918 241319 328970 241325
rect 329014 241377 329066 241383
rect 329014 241319 329066 241325
rect 328726 237159 328778 237165
rect 328726 237101 328778 237107
rect 328822 237159 328874 237165
rect 328822 237101 328874 237107
rect 328438 236271 328490 236277
rect 328438 236213 328490 236219
rect 328834 233484 328862 237101
rect 328224 233456 328286 233484
rect 328608 233456 328862 233484
rect 328930 233484 328958 241319
rect 329026 239829 329054 241319
rect 329122 240051 329150 246494
rect 329602 241531 329630 246494
rect 329686 246335 329738 246341
rect 329686 246277 329738 246283
rect 329698 246193 329726 246277
rect 329686 246187 329738 246193
rect 329686 246129 329738 246135
rect 329986 241753 330014 246494
rect 330178 246480 330432 246508
rect 330562 246480 330912 246508
rect 329974 241747 330026 241753
rect 329974 241689 330026 241695
rect 330070 241673 330122 241679
rect 330070 241615 330122 241621
rect 329590 241525 329642 241531
rect 329590 241467 329642 241473
rect 329110 240045 329162 240051
rect 329110 239987 329162 239993
rect 329686 240045 329738 240051
rect 329686 239987 329738 239993
rect 329302 239897 329354 239903
rect 329302 239839 329354 239845
rect 329014 239823 329066 239829
rect 329014 239765 329066 239771
rect 328930 233456 328992 233484
rect 329314 233470 329342 239839
rect 329698 233470 329726 239987
rect 329782 238565 329834 238571
rect 329782 238507 329834 238513
rect 329794 237979 329822 238507
rect 329782 237973 329834 237979
rect 329782 237915 329834 237921
rect 329782 237529 329834 237535
rect 329782 237471 329834 237477
rect 329794 236911 329822 237471
rect 329780 236902 329836 236911
rect 329780 236837 329836 236846
rect 330082 233470 330110 241615
rect 330178 241161 330206 246480
rect 330166 241155 330218 241161
rect 330166 241097 330218 241103
rect 330562 237239 330590 246480
rect 330742 246187 330794 246193
rect 330742 246129 330794 246135
rect 330754 245749 330782 246129
rect 330742 245743 330794 245749
rect 330742 245685 330794 245691
rect 330838 245743 330890 245749
rect 330838 245685 330890 245691
rect 330850 245305 330878 245685
rect 330838 245299 330890 245305
rect 330838 245241 330890 245247
rect 330934 245299 330986 245305
rect 330934 245241 330986 245247
rect 330946 244861 330974 245241
rect 330934 244855 330986 244861
rect 330934 244797 330986 244803
rect 331124 243266 331180 243275
rect 331124 243201 331180 243210
rect 331138 242863 331166 243201
rect 331126 242857 331178 242863
rect 331126 242799 331178 242805
rect 331030 241747 331082 241753
rect 331030 241689 331082 241695
rect 330550 237233 330602 237239
rect 330550 237175 330602 237181
rect 330646 237233 330698 237239
rect 330646 237175 330698 237181
rect 330658 233484 330686 237175
rect 331042 233484 331070 241689
rect 331222 238787 331274 238793
rect 331222 238729 331274 238735
rect 331234 233780 331262 238729
rect 331330 237461 331358 246494
rect 331510 241525 331562 241531
rect 331510 241467 331562 241473
rect 331318 237455 331370 237461
rect 331318 237397 331370 237403
rect 330432 233456 330686 233484
rect 330816 233456 331070 233484
rect 331186 233752 331262 233780
rect 331186 233470 331214 233752
rect 331522 233470 331550 241467
rect 331714 241013 331742 246494
rect 331702 241007 331754 241013
rect 331702 240949 331754 240955
rect 332194 238867 332222 246494
rect 332386 246480 332640 246508
rect 332770 246480 333024 246508
rect 332278 241155 332330 241161
rect 332278 241097 332330 241103
rect 332182 238861 332234 238867
rect 332182 238803 332234 238809
rect 332290 238627 332318 241097
rect 332386 238719 332414 246480
rect 332770 239311 332798 246480
rect 332950 241451 333002 241457
rect 332950 241393 333002 241399
rect 332758 239305 332810 239311
rect 332758 239247 332810 239253
rect 332470 238861 332522 238867
rect 332470 238803 332522 238809
rect 332374 238713 332426 238719
rect 332374 238655 332426 238661
rect 332002 238599 332318 238627
rect 331798 237529 331850 237535
rect 331798 237471 331850 237477
rect 331810 237313 331838 237471
rect 331798 237307 331850 237313
rect 331798 237249 331850 237255
rect 331894 237307 331946 237313
rect 331894 237249 331946 237255
rect 331906 233470 331934 237249
rect 332002 233484 332030 238599
rect 332482 238571 332510 238803
rect 332470 238565 332522 238571
rect 332470 238507 332522 238513
rect 332854 238491 332906 238497
rect 332854 238433 332906 238439
rect 332470 238343 332522 238349
rect 332758 238343 332810 238349
rect 332522 238303 332758 238331
rect 332470 238285 332522 238291
rect 332758 238285 332810 238291
rect 332098 238201 332606 238220
rect 332086 238195 332618 238201
rect 332138 238192 332566 238195
rect 332086 238137 332138 238143
rect 332566 238137 332618 238143
rect 332662 238047 332714 238053
rect 332662 237989 332714 237995
rect 332278 237973 332330 237979
rect 332278 237915 332330 237921
rect 332290 237776 332318 237915
rect 332674 237776 332702 237989
rect 332290 237748 332702 237776
rect 332866 233484 332894 238433
rect 332962 233780 332990 241393
rect 333442 238645 333470 246494
rect 333922 241827 333950 246494
rect 333910 241821 333962 241827
rect 333910 241763 333962 241769
rect 333718 241007 333770 241013
rect 333718 240949 333770 240955
rect 333430 238639 333482 238645
rect 333430 238581 333482 238587
rect 333622 238639 333674 238645
rect 333622 238581 333674 238587
rect 332962 233752 333038 233780
rect 332002 233456 332304 233484
rect 332640 233456 332894 233484
rect 333010 233470 333038 233752
rect 333634 233484 333662 238581
rect 333408 233456 333662 233484
rect 333730 233470 333758 240949
rect 334102 238713 334154 238719
rect 334102 238655 334154 238661
rect 334114 233470 334142 238655
rect 334402 236425 334430 246494
rect 334594 246480 334752 246508
rect 334486 241821 334538 241827
rect 334486 241763 334538 241769
rect 334390 236419 334442 236425
rect 334390 236361 334442 236367
rect 334498 233470 334526 241763
rect 334594 239163 334622 246480
rect 334774 246261 334826 246267
rect 334774 246203 334826 246209
rect 334882 246212 334910 246573
rect 334978 246489 335006 246573
rect 335350 246557 335402 246563
rect 335350 246499 335402 246505
rect 334966 246483 335018 246489
rect 334966 246425 335018 246431
rect 335158 246335 335210 246341
rect 335158 246277 335210 246283
rect 335170 246212 335198 246277
rect 334786 246064 334814 246203
rect 334882 246184 335198 246212
rect 335362 246064 335390 246499
rect 334786 246036 335390 246064
rect 335458 244288 335486 246628
rect 335266 244260 335486 244288
rect 334582 239157 334634 239163
rect 334582 239099 334634 239105
rect 334870 238565 334922 238571
rect 334870 238507 334922 238513
rect 334882 233484 334910 238507
rect 335266 236499 335294 244260
rect 335350 244115 335402 244121
rect 335350 244057 335402 244063
rect 335254 236493 335306 236499
rect 335254 236435 335306 236441
rect 334964 235126 335020 235135
rect 334964 235061 335020 235070
rect 334848 233456 334910 233484
rect 334978 233484 335006 235061
rect 335362 233484 335390 244057
rect 335650 236351 335678 246494
rect 336130 241605 336158 246494
rect 336310 244041 336362 244047
rect 336310 243983 336362 243989
rect 336118 241599 336170 241605
rect 336118 241541 336170 241547
rect 335638 236345 335690 236351
rect 335638 236287 335690 236293
rect 335926 235605 335978 235611
rect 335926 235547 335978 235553
rect 334978 233456 335232 233484
rect 335362 233456 335616 233484
rect 335938 233470 335966 235547
rect 336322 233470 336350 243983
rect 336514 239089 336542 246494
rect 336960 246480 337022 246508
rect 336502 239083 336554 239089
rect 336502 239025 336554 239031
rect 336994 238423 337022 246480
rect 337186 246480 337440 246508
rect 337078 243005 337130 243011
rect 337078 242947 337130 242953
rect 336982 238417 337034 238423
rect 336982 238359 337034 238365
rect 336694 235753 336746 235759
rect 336694 235695 336746 235701
rect 336706 233470 336734 235695
rect 337090 233484 337118 242947
rect 337186 239385 337214 246480
rect 337558 243227 337610 243233
rect 337558 243169 337610 243175
rect 337174 239379 337226 239385
rect 337174 239321 337226 239327
rect 337174 235531 337226 235537
rect 337174 235473 337226 235479
rect 337056 233456 337118 233484
rect 337186 233484 337214 235473
rect 337570 233484 337598 243169
rect 337858 241309 337886 246494
rect 337954 246480 338256 246508
rect 338626 246480 338736 246508
rect 338914 246480 339168 246508
rect 339394 246480 339648 246508
rect 339970 246480 340032 246508
rect 337846 241303 337898 241309
rect 337846 241245 337898 241251
rect 337954 237535 337982 246480
rect 338134 245891 338186 245897
rect 338134 245833 338186 245839
rect 338230 245891 338282 245897
rect 338230 245833 338282 245839
rect 338146 245324 338174 245833
rect 338242 245453 338270 245833
rect 338518 245521 338570 245527
rect 338518 245463 338570 245469
rect 338230 245447 338282 245453
rect 338230 245389 338282 245395
rect 338422 245373 338474 245379
rect 338146 245321 338422 245324
rect 338146 245315 338474 245321
rect 338146 245296 338462 245315
rect 338530 244935 338558 245463
rect 338518 244929 338570 244935
rect 338518 244871 338570 244877
rect 338626 244843 338654 246480
rect 338530 244815 338654 244843
rect 338530 244473 338558 244815
rect 338530 244445 338750 244473
rect 338518 242709 338570 242715
rect 338518 242651 338570 242657
rect 337942 237529 337994 237535
rect 337942 237471 337994 237477
rect 338134 237381 338186 237387
rect 338134 237323 338186 237329
rect 338146 237059 338174 237323
rect 338132 237050 338188 237059
rect 338132 236985 338188 236994
rect 338134 235679 338186 235685
rect 338134 235621 338186 235627
rect 337186 233456 337440 233484
rect 337570 233456 337824 233484
rect 338146 233470 338174 235621
rect 338530 233470 338558 242651
rect 338722 238275 338750 244445
rect 338914 239533 338942 246480
rect 338996 242378 339052 242387
rect 338996 242313 339052 242322
rect 338902 239527 338954 239533
rect 338902 239469 338954 239475
rect 338710 238269 338762 238275
rect 338710 238211 338762 238217
rect 338902 235827 338954 235833
rect 338902 235769 338954 235775
rect 338914 233470 338942 235769
rect 339010 233484 339038 242313
rect 339394 241235 339422 246480
rect 339862 244411 339914 244417
rect 339862 244353 339914 244359
rect 339766 244337 339818 244343
rect 339874 244288 339902 244353
rect 339818 244285 339902 244288
rect 339766 244279 339902 244285
rect 339778 244260 339902 244279
rect 339862 243153 339914 243159
rect 339862 243095 339914 243101
rect 339574 242931 339626 242937
rect 339574 242873 339626 242879
rect 339586 242387 339614 242873
rect 339764 242526 339820 242535
rect 339764 242461 339820 242470
rect 339778 242419 339806 242461
rect 339766 242413 339818 242419
rect 339572 242378 339628 242387
rect 339766 242355 339818 242361
rect 339572 242313 339628 242322
rect 339382 241229 339434 241235
rect 339382 241171 339434 241177
rect 339478 241229 339530 241235
rect 339478 241171 339530 241177
rect 339490 237313 339518 241171
rect 339766 237455 339818 237461
rect 339766 237397 339818 237403
rect 339478 237307 339530 237313
rect 339478 237249 339530 237255
rect 339778 236911 339806 237397
rect 339764 236902 339820 236911
rect 339764 236837 339820 236846
rect 339382 235975 339434 235981
rect 339382 235917 339434 235923
rect 339394 233484 339422 235917
rect 339874 233484 339902 243095
rect 339970 236573 339998 246480
rect 340450 238201 340478 246494
rect 340726 243301 340778 243307
rect 340726 243243 340778 243249
rect 340438 238195 340490 238201
rect 340438 238137 340490 238143
rect 339958 236567 340010 236573
rect 339958 236509 340010 236515
rect 340342 235901 340394 235907
rect 340342 235843 340394 235849
rect 339010 233456 339264 233484
rect 339394 233456 339648 233484
rect 339874 233456 340032 233484
rect 340354 233470 340382 235843
rect 340738 233470 340766 243243
rect 340930 239681 340958 246494
rect 341204 242674 341260 242683
rect 341204 242609 341260 242618
rect 340918 239675 340970 239681
rect 340918 239617 340970 239623
rect 341108 235274 341164 235283
rect 341108 235209 341164 235218
rect 341122 233470 341150 235209
rect 341218 233484 341246 242609
rect 341314 239607 341342 246494
rect 341506 246480 341760 246508
rect 341986 246480 342240 246508
rect 341302 239601 341354 239607
rect 341302 239543 341354 239549
rect 341506 238127 341534 246480
rect 341986 239459 342014 246480
rect 342068 242970 342124 242979
rect 342068 242905 342124 242914
rect 341974 239453 342026 239459
rect 341974 239395 342026 239401
rect 341494 238121 341546 238127
rect 341494 238063 341546 238069
rect 341588 235718 341644 235727
rect 341588 235653 341644 235662
rect 341602 233484 341630 235653
rect 342082 233484 342110 242905
rect 342658 240939 342686 246494
rect 342742 246113 342794 246119
rect 342742 246055 342794 246061
rect 342754 244639 342782 246055
rect 342742 244633 342794 244639
rect 342742 244575 342794 244581
rect 342932 242822 342988 242831
rect 342932 242757 342988 242766
rect 342646 240933 342698 240939
rect 342646 240875 342698 240881
rect 342548 235866 342604 235875
rect 342548 235801 342604 235810
rect 341218 233456 341472 233484
rect 341602 233456 341856 233484
rect 342082 233456 342240 233484
rect 342562 233470 342590 235801
rect 342946 233470 342974 242757
rect 343042 236869 343070 246494
rect 343412 242230 343468 242239
rect 343412 242165 343468 242174
rect 343030 236863 343082 236869
rect 343030 236805 343082 236811
rect 343316 235570 343372 235579
rect 343316 235505 343372 235514
rect 343330 233470 343358 235505
rect 343426 233484 343454 242165
rect 343522 238053 343550 246494
rect 343714 246480 343968 246508
rect 344194 246480 344448 246508
rect 343714 239829 343742 246480
rect 344194 240865 344222 246480
rect 344276 242378 344332 242387
rect 344276 242313 344332 242322
rect 344182 240859 344234 240865
rect 344182 240801 344234 240807
rect 343702 239823 343754 239829
rect 343702 239765 343754 239771
rect 343510 238047 343562 238053
rect 343510 237989 343562 237995
rect 343796 235422 343852 235431
rect 343796 235357 343852 235366
rect 343810 233484 343838 235357
rect 344290 233484 344318 242313
rect 344770 236795 344798 246494
rect 345142 243449 345194 243455
rect 345142 243391 345194 243397
rect 344758 236789 344810 236795
rect 344758 236731 344810 236737
rect 344756 236162 344812 236171
rect 344756 236097 344812 236106
rect 343426 233456 343680 233484
rect 343810 233456 344064 233484
rect 344290 233456 344448 233484
rect 344770 233470 344798 236097
rect 345154 233470 345182 243391
rect 345250 237979 345278 246494
rect 345622 243375 345674 243381
rect 345622 243317 345674 243323
rect 345238 237973 345290 237979
rect 345238 237915 345290 237921
rect 345526 234717 345578 234723
rect 345526 234659 345578 234665
rect 345538 233470 345566 234659
rect 345634 233484 345662 243317
rect 345730 240717 345758 246494
rect 345922 246480 346176 246508
rect 346306 246480 346560 246508
rect 345718 240711 345770 240717
rect 345718 240653 345770 240659
rect 345922 236647 345950 246480
rect 346306 240569 346334 246480
rect 346390 243523 346442 243529
rect 346390 243465 346442 243471
rect 346294 240563 346346 240569
rect 346294 240505 346346 240511
rect 345910 236641 345962 236647
rect 345910 236583 345962 236589
rect 346004 236014 346060 236023
rect 346004 235949 346060 235958
rect 346018 233484 346046 235949
rect 346402 233484 346430 243465
rect 346978 236721 347006 246494
rect 347350 243671 347402 243677
rect 347350 243613 347402 243619
rect 346966 236715 347018 236721
rect 346966 236657 347018 236663
rect 346966 234791 347018 234797
rect 346966 234733 347018 234739
rect 345634 233456 345888 233484
rect 346018 233456 346272 233484
rect 346402 233456 346656 233484
rect 346978 233470 347006 234733
rect 347362 233470 347390 243613
rect 347458 238867 347486 246494
rect 347830 241969 347882 241975
rect 347830 241911 347882 241917
rect 347446 238861 347498 238867
rect 347446 238803 347498 238809
rect 347732 234386 347788 234395
rect 347732 234321 347788 234330
rect 347746 233470 347774 234321
rect 347842 233484 347870 241911
rect 347938 241383 347966 246494
rect 348034 246480 348288 246508
rect 348610 246480 348768 246508
rect 347926 241377 347978 241383
rect 347926 241319 347978 241325
rect 348034 240643 348062 246480
rect 348406 241673 348458 241679
rect 348406 241615 348458 241621
rect 348418 241587 348446 241615
rect 348502 241599 348554 241605
rect 348418 241559 348502 241587
rect 348502 241541 348554 241547
rect 348022 240637 348074 240643
rect 348022 240579 348074 240585
rect 348610 239237 348638 246480
rect 348694 242117 348746 242123
rect 348694 242059 348746 242065
rect 348598 239231 348650 239237
rect 348598 239173 348650 239179
rect 348406 237455 348458 237461
rect 348502 237455 348554 237461
rect 348458 237415 348502 237443
rect 348406 237397 348458 237403
rect 348502 237397 348554 237403
rect 348212 234978 348268 234987
rect 348212 234913 348268 234922
rect 348226 233484 348254 234913
rect 348706 233484 348734 242059
rect 349186 237905 349214 246494
rect 349270 243597 349322 243603
rect 349270 243539 349322 243545
rect 349174 237899 349226 237905
rect 349174 237841 349226 237847
rect 349172 234534 349228 234543
rect 349172 234469 349228 234478
rect 347842 233456 348096 233484
rect 348226 233456 348480 233484
rect 348706 233456 348864 233484
rect 349186 233470 349214 234469
rect 349282 233484 349310 243539
rect 349570 239755 349598 246494
rect 349762 246480 350064 246508
rect 349558 239749 349610 239755
rect 349558 239691 349610 239697
rect 349762 237017 349790 246480
rect 350146 246119 350174 246647
rect 350242 246480 350496 246508
rect 350722 246480 350976 246508
rect 350134 246113 350186 246119
rect 350134 246055 350186 246061
rect 350038 242191 350090 242197
rect 350038 242133 350090 242139
rect 349750 237011 349802 237017
rect 349750 236953 349802 236959
rect 349942 235235 349994 235241
rect 349942 235177 349994 235183
rect 349282 233456 349584 233484
rect 349954 233470 349982 235177
rect 350050 233484 350078 242133
rect 350242 240495 350270 246480
rect 350230 240489 350282 240495
rect 350230 240431 350282 240437
rect 350722 237091 350750 246480
rect 350806 243745 350858 243751
rect 350806 243687 350858 243693
rect 350710 237085 350762 237091
rect 350710 237027 350762 237033
rect 350422 235087 350474 235093
rect 350422 235029 350474 235035
rect 350434 233484 350462 235029
rect 350818 233484 350846 243687
rect 351298 240019 351326 246494
rect 351490 246480 351792 246508
rect 351970 246480 352272 246508
rect 351284 240010 351340 240019
rect 351284 239945 351340 239954
rect 351380 239122 351436 239131
rect 351380 239057 351436 239066
rect 351394 238867 351422 239057
rect 351382 238861 351434 238867
rect 351382 238803 351434 238809
rect 351490 236943 351518 246480
rect 351766 242043 351818 242049
rect 351766 241985 351818 241991
rect 351478 236937 351530 236943
rect 351478 236879 351530 236885
rect 351382 234865 351434 234871
rect 351382 234807 351434 234813
rect 350050 233456 350304 233484
rect 350434 233456 350688 233484
rect 350818 233456 351072 233484
rect 351394 233470 351422 234807
rect 351778 233470 351806 241985
rect 351970 237757 351998 246480
rect 352354 246341 352382 246647
rect 353206 246631 353258 246637
rect 353206 246573 353258 246579
rect 353302 246631 353354 246637
rect 353302 246573 353354 246579
rect 352450 246480 352704 246508
rect 352834 246480 353088 246508
rect 352342 246335 352394 246341
rect 352342 246277 352394 246283
rect 352244 243118 352300 243127
rect 352244 243053 352300 243062
rect 351958 237751 352010 237757
rect 351958 237693 352010 237699
rect 352150 235161 352202 235167
rect 352150 235103 352202 235109
rect 352162 233470 352190 235103
rect 352258 233484 352286 243053
rect 352450 239977 352478 246480
rect 352834 240167 352862 246480
rect 353218 246415 353246 246573
rect 353206 246409 353258 246415
rect 353206 246351 353258 246357
rect 353314 246119 353342 246573
rect 353302 246113 353354 246119
rect 353302 246055 353354 246061
rect 353014 242265 353066 242271
rect 353014 242207 353066 242213
rect 352820 240158 352876 240167
rect 352820 240093 352876 240102
rect 352438 239971 352490 239977
rect 352438 239913 352490 239919
rect 352630 234939 352682 234945
rect 352630 234881 352682 234887
rect 352642 233484 352670 234881
rect 353026 233484 353054 242207
rect 353506 237165 353534 246494
rect 353590 244855 353642 244861
rect 353590 244797 353642 244803
rect 353602 237387 353630 244797
rect 353686 243819 353738 243825
rect 353686 243761 353738 243767
rect 353590 237381 353642 237387
rect 353590 237323 353642 237329
rect 353494 237159 353546 237165
rect 353494 237101 353546 237107
rect 353590 235383 353642 235389
rect 353590 235325 353642 235331
rect 352258 233456 352512 233484
rect 352642 233456 352896 233484
rect 353026 233456 353280 233484
rect 353602 233470 353630 235325
rect 353698 233484 353726 243761
rect 353986 237831 354014 246494
rect 354466 241647 354494 246494
rect 354562 246480 354816 246508
rect 355042 246480 355296 246508
rect 354452 241638 354508 241647
rect 354452 241573 354508 241582
rect 354562 239903 354590 246480
rect 354644 242082 354700 242091
rect 354644 242017 354700 242026
rect 354550 239897 354602 239903
rect 354550 239839 354602 239845
rect 353974 237825 354026 237831
rect 353974 237767 354026 237773
rect 354358 235013 354410 235019
rect 354358 234955 354410 234961
rect 353698 233456 354000 233484
rect 354370 233470 354398 234955
rect 354658 233780 354686 242017
rect 355042 237609 355070 246480
rect 355222 242339 355274 242345
rect 355222 242281 355274 242287
rect 355030 237603 355082 237609
rect 355030 237545 355082 237551
rect 355126 237603 355178 237609
rect 355126 237545 355178 237551
rect 355138 237313 355166 237545
rect 355126 237307 355178 237313
rect 355126 237249 355178 237255
rect 354838 235309 354890 235315
rect 354838 235251 354890 235257
rect 354658 233752 354734 233780
rect 354706 233470 354734 233752
rect 354850 233484 354878 235251
rect 355234 233484 355262 242281
rect 355714 240051 355742 246494
rect 355798 245447 355850 245453
rect 355798 245389 355850 245395
rect 355702 240045 355754 240051
rect 355702 239987 355754 239993
rect 354850 233456 355104 233484
rect 355234 233456 355488 233484
rect 355810 233470 355838 245389
rect 355894 244929 355946 244935
rect 355894 244871 355946 244877
rect 355906 233484 355934 244871
rect 356194 237683 356222 246494
rect 356278 245817 356330 245823
rect 356278 245759 356330 245765
rect 356182 237677 356234 237683
rect 356182 237619 356234 237625
rect 356290 233484 356318 245759
rect 356578 241605 356606 246494
rect 356770 246480 357024 246508
rect 357250 246480 357504 246508
rect 356770 241795 356798 246480
rect 357142 245743 357194 245749
rect 357142 245685 357194 245691
rect 356756 241786 356812 241795
rect 356756 241721 356812 241730
rect 356566 241599 356618 241605
rect 356566 241541 356618 241547
rect 356662 235457 356714 235463
rect 356662 235399 356714 235405
rect 356674 233484 356702 235399
rect 357154 233484 357182 245685
rect 357250 237239 357278 246480
rect 357430 245891 357482 245897
rect 357430 245833 357482 245839
rect 357238 237233 357290 237239
rect 357238 237175 357290 237181
rect 357442 233484 357470 245833
rect 357826 237207 357854 246494
rect 358006 246187 358058 246193
rect 358006 246129 358058 246135
rect 357812 237198 357868 237207
rect 357812 237133 357868 237142
rect 355906 233456 356208 233484
rect 356290 233456 356592 233484
rect 356674 233456 356928 233484
rect 357154 233456 357312 233484
rect 357442 233456 357696 233484
rect 358018 233470 358046 246129
rect 358102 245373 358154 245379
rect 358102 245315 358154 245321
rect 358114 233484 358142 245315
rect 358306 241753 358334 246494
rect 358582 245447 358634 245453
rect 358582 245389 358634 245395
rect 358486 245373 358538 245379
rect 358486 245315 358538 245321
rect 358294 241747 358346 241753
rect 358294 241689 358346 241695
rect 358498 237355 358526 245315
rect 358594 245231 358622 245389
rect 358582 245225 358634 245231
rect 358582 245167 358634 245173
rect 358786 238793 358814 246494
rect 358978 246480 359232 246508
rect 359362 246480 359616 246508
rect 358978 241351 359006 246480
rect 359362 241531 359390 246480
rect 359350 241525 359402 241531
rect 359350 241467 359402 241473
rect 358964 241342 359020 241351
rect 358964 241277 359020 241286
rect 358870 238861 358922 238867
rect 358870 238803 358922 238809
rect 358774 238787 358826 238793
rect 358774 238729 358826 238735
rect 358774 237381 358826 237387
rect 358484 237346 358540 237355
rect 358774 237323 358826 237329
rect 358484 237281 358540 237290
rect 358114 233456 358416 233484
rect 358786 233470 358814 237323
rect 358882 233484 358910 238803
rect 359830 237751 359882 237757
rect 359830 237693 359882 237699
rect 359252 236606 359308 236615
rect 359252 236541 359308 236550
rect 359266 233484 359294 236541
rect 358882 233456 359136 233484
rect 359266 233456 359520 233484
rect 298196 233433 298252 233442
rect 359842 233336 359870 237693
rect 360034 237503 360062 246494
rect 360514 241235 360542 246494
rect 360706 246480 361008 246508
rect 361090 246480 361344 246508
rect 361666 246480 361824 246508
rect 360502 241229 360554 241235
rect 360502 241171 360554 241177
rect 360214 240045 360266 240051
rect 360214 239987 360266 239993
rect 360020 237494 360076 237503
rect 360020 237429 360076 237438
rect 360226 233470 360254 239987
rect 360598 239305 360650 239311
rect 360598 239247 360650 239253
rect 360610 233470 360638 239247
rect 360706 238687 360734 246480
rect 360982 241599 361034 241605
rect 360982 241541 361034 241547
rect 360692 238678 360748 238687
rect 360692 238613 360748 238622
rect 360994 233470 361022 241541
rect 361090 241161 361118 246480
rect 361558 241747 361610 241753
rect 361558 241689 361610 241695
rect 361078 241155 361130 241161
rect 361078 241097 361130 241103
rect 361570 233484 361598 241689
rect 361666 241055 361694 246480
rect 361942 241525 361994 241531
rect 361942 241467 361994 241473
rect 361652 241046 361708 241055
rect 361652 240981 361708 240990
rect 361954 233484 361982 241467
rect 362242 238497 362270 246494
rect 362626 246397 362654 246647
rect 362806 246631 362858 246637
rect 362806 246573 362858 246579
rect 362818 246397 362846 246573
rect 362626 246369 362846 246397
rect 362914 245379 362942 246776
rect 385078 246779 385130 246785
rect 385078 246721 385130 246727
rect 386998 246779 387050 246785
rect 388532 246818 388588 246827
rect 387380 246753 387436 246762
rect 388054 246779 388106 246785
rect 386998 246721 387050 246727
rect 369142 246705 369194 246711
rect 368962 246653 369142 246656
rect 368962 246647 369194 246653
rect 368962 246637 369182 246647
rect 368950 246631 369182 246637
rect 369002 246628 369182 246631
rect 368950 246573 369002 246579
rect 362902 245373 362954 245379
rect 362902 245315 362954 245321
rect 362326 241377 362378 241383
rect 362326 241319 362378 241325
rect 362230 238491 362282 238497
rect 362230 238433 362282 238439
rect 362338 233484 362366 241319
rect 362422 241155 362474 241161
rect 362422 241097 362474 241103
rect 361344 233456 361598 233484
rect 361728 233456 361982 233484
rect 362112 233456 362366 233484
rect 362434 233470 362462 241097
rect 363106 240759 363134 246494
rect 363298 246480 363552 246508
rect 363874 246480 364032 246508
rect 363190 241673 363242 241679
rect 363190 241615 363242 241621
rect 363092 240750 363148 240759
rect 363092 240685 363148 240694
rect 362806 237899 362858 237905
rect 362806 237841 362858 237847
rect 362818 233470 362846 237841
rect 363202 233470 363230 241615
rect 363298 238645 363326 246480
rect 363766 241303 363818 241309
rect 363766 241245 363818 241251
rect 363286 238639 363338 238645
rect 363286 238581 363338 238587
rect 363778 233484 363806 241245
rect 363874 238539 363902 246480
rect 364150 241229 364202 241235
rect 364150 241171 364202 241177
rect 363860 238530 363916 238539
rect 363860 238465 363916 238474
rect 364162 233484 364190 241171
rect 364354 241013 364382 246494
rect 364534 241451 364586 241457
rect 364534 241393 364586 241399
rect 364342 241007 364394 241013
rect 364342 240949 364394 240955
rect 364546 233484 364574 241393
rect 364834 240611 364862 246494
rect 365014 240637 365066 240643
rect 364820 240602 364876 240611
rect 364630 240563 364682 240569
rect 365014 240579 365066 240585
rect 364820 240537 364876 240546
rect 364630 240505 364682 240511
rect 363552 233456 363806 233484
rect 363936 233456 364190 233484
rect 364320 233456 364574 233484
rect 364642 233470 364670 240505
rect 365026 233470 365054 240579
rect 365314 238719 365342 246494
rect 365760 246480 365822 246508
rect 365398 240933 365450 240939
rect 365398 240875 365450 240881
rect 365302 238713 365354 238719
rect 365302 238655 365354 238661
rect 365410 233470 365438 240875
rect 365794 238243 365822 246480
rect 365890 246480 366144 246508
rect 365890 241827 365918 246480
rect 365878 241821 365930 241827
rect 365878 241763 365930 241769
rect 365974 240859 366026 240865
rect 365974 240801 366026 240807
rect 365780 238234 365836 238243
rect 365780 238169 365836 238178
rect 365986 233484 366014 240801
rect 366358 240489 366410 240495
rect 366562 240463 366590 246494
rect 366742 240711 366794 240717
rect 366742 240653 366794 240659
rect 366358 240431 366410 240437
rect 366548 240454 366604 240463
rect 366370 233484 366398 240431
rect 366548 240389 366604 240398
rect 366754 233484 366782 240653
rect 367042 238571 367070 246494
rect 367522 246045 367550 246494
rect 367618 246480 367872 246508
rect 368098 246480 368352 246508
rect 367510 246039 367562 246045
rect 367510 245981 367562 245987
rect 367618 244565 367646 246480
rect 367702 246039 367754 246045
rect 367702 245981 367754 245987
rect 367714 244639 367742 245981
rect 368098 245971 368126 246480
rect 368086 245965 368138 245971
rect 368086 245907 368138 245913
rect 367702 244633 367754 244639
rect 367702 244575 367754 244581
rect 367606 244559 367658 244565
rect 367606 244501 367658 244507
rect 368770 244491 368798 246494
rect 369250 245601 369278 246494
rect 369238 245595 369290 245601
rect 369238 245537 369290 245543
rect 368758 244485 368810 244491
rect 368758 244427 368810 244433
rect 367222 241007 367274 241013
rect 367222 240949 367274 240955
rect 367030 238565 367082 238571
rect 367030 238507 367082 238513
rect 366838 238491 366890 238497
rect 366838 238433 366890 238439
rect 365760 233456 366014 233484
rect 366144 233456 366398 233484
rect 366528 233456 366782 233484
rect 366850 233470 366878 238433
rect 367234 233470 367262 240949
rect 367604 240454 367660 240463
rect 367604 240389 367660 240398
rect 367618 233470 367646 240389
rect 368182 238861 368234 238867
rect 368182 238803 368234 238809
rect 368194 233484 368222 238803
rect 368662 238787 368714 238793
rect 368662 238729 368714 238735
rect 368674 233780 368702 238729
rect 369430 238491 369482 238497
rect 369430 238433 369482 238439
rect 369046 237381 369098 237387
rect 369046 237323 369098 237329
rect 368950 236789 369002 236795
rect 368950 236731 369002 236737
rect 368578 233752 368702 233780
rect 368578 233484 368606 233752
rect 368962 233484 368990 236731
rect 367968 233456 368222 233484
rect 368352 233456 368606 233484
rect 368736 233456 368990 233484
rect 369058 233470 369086 237323
rect 369442 233470 369470 238433
rect 369634 236055 369662 246494
rect 369826 246480 370080 246508
rect 370306 246480 370560 246508
rect 369826 240315 369854 246480
rect 370306 243899 370334 246480
rect 370978 245675 371006 246494
rect 370966 245669 371018 245675
rect 370966 245611 371018 245617
rect 370294 243893 370346 243899
rect 370294 243835 370346 243841
rect 369812 240306 369868 240315
rect 369812 240241 369868 240250
rect 371362 240199 371390 246494
rect 371842 240347 371870 246494
rect 372034 246480 372288 246508
rect 372418 246480 372672 246508
rect 372898 246480 373152 246508
rect 372034 245231 372062 246480
rect 372022 245225 372074 245231
rect 372022 245167 372074 245173
rect 371830 240341 371882 240347
rect 371830 240283 371882 240289
rect 371350 240193 371402 240199
rect 371350 240135 371402 240141
rect 372418 240125 372446 246480
rect 372898 241499 372926 246480
rect 372884 241490 372940 241499
rect 372884 241425 372940 241434
rect 373570 240273 373598 246494
rect 374050 245083 374078 246494
rect 374038 245077 374090 245083
rect 374038 245019 374090 245025
rect 374434 240421 374462 246494
rect 374626 246480 374880 246508
rect 375106 246480 375360 246508
rect 374626 245009 374654 246480
rect 374614 245003 374666 245009
rect 374614 244945 374666 244951
rect 375106 241901 375134 246480
rect 375094 241895 375146 241901
rect 375094 241837 375146 241843
rect 375778 240791 375806 246494
rect 376162 241087 376190 246494
rect 376150 241081 376202 241087
rect 376150 241023 376202 241029
rect 375766 240785 375818 240791
rect 375766 240727 375818 240733
rect 374422 240415 374474 240421
rect 374422 240357 374474 240363
rect 373558 240267 373610 240273
rect 373558 240209 373610 240215
rect 376438 240267 376490 240273
rect 376438 240209 376490 240215
rect 372406 240119 372458 240125
rect 372406 240061 372458 240067
rect 376054 240119 376106 240125
rect 376054 240061 376106 240067
rect 375670 239971 375722 239977
rect 375670 239913 375722 239919
rect 374806 239675 374858 239681
rect 374806 239617 374858 239623
rect 373366 239157 373418 239163
rect 373366 239099 373418 239105
rect 370486 238639 370538 238645
rect 370486 238581 370538 238587
rect 370006 238565 370058 238571
rect 370006 238507 370058 238513
rect 369814 238417 369866 238423
rect 369814 238359 369866 238365
rect 369622 236049 369674 236055
rect 369622 235991 369674 235997
rect 369826 233470 369854 238359
rect 370018 237757 370046 238507
rect 370390 238269 370442 238275
rect 370390 238211 370442 238217
rect 370006 237751 370058 237757
rect 370006 237693 370058 237699
rect 370402 233484 370430 238211
rect 370498 237905 370526 238581
rect 372022 238195 372074 238201
rect 372022 238137 372074 238143
rect 371638 238121 371690 238127
rect 371638 238063 371690 238069
rect 371254 238047 371306 238053
rect 371254 237989 371306 237995
rect 371158 237973 371210 237979
rect 371158 237915 371210 237921
rect 370486 237899 370538 237905
rect 370486 237841 370538 237847
rect 370582 237899 370634 237905
rect 370582 237841 370634 237847
rect 370594 237609 370622 237841
rect 370774 237751 370826 237757
rect 370774 237693 370826 237699
rect 370582 237603 370634 237609
rect 370582 237545 370634 237551
rect 370786 233484 370814 237693
rect 371170 233484 371198 237915
rect 370176 233456 370430 233484
rect 370560 233456 370814 233484
rect 370944 233456 371198 233484
rect 371266 233470 371294 237989
rect 371650 233470 371678 238063
rect 372034 233470 372062 238137
rect 372598 237529 372650 237535
rect 372598 237471 372650 237477
rect 372610 233484 372638 237471
rect 372982 237455 373034 237461
rect 372982 237397 373034 237403
rect 372994 233484 373022 237397
rect 373378 233484 373406 239099
rect 373846 239083 373898 239089
rect 373846 239025 373898 239031
rect 373462 237677 373514 237683
rect 373462 237619 373514 237625
rect 372384 233456 372638 233484
rect 372768 233456 373022 233484
rect 373152 233456 373406 233484
rect 373474 233470 373502 237619
rect 373858 233470 373886 239025
rect 374230 237603 374282 237609
rect 374230 237545 374282 237551
rect 374242 233470 374270 237545
rect 374818 233484 374846 239617
rect 375190 239453 375242 239459
rect 375190 239395 375242 239401
rect 375202 233484 375230 239395
rect 375574 237825 375626 237831
rect 375574 237767 375626 237773
rect 375586 233484 375614 237767
rect 374592 233456 374846 233484
rect 374976 233456 375230 233484
rect 375360 233456 375614 233484
rect 375682 233470 375710 239913
rect 376066 233470 376094 240061
rect 376450 233470 376478 240209
rect 376642 239015 376670 246494
rect 376834 246480 377088 246508
rect 377314 246480 377568 246508
rect 376834 241203 376862 246480
rect 377206 241821 377258 241827
rect 377206 241763 377258 241769
rect 376820 241194 376876 241203
rect 376820 241129 376876 241138
rect 377014 240415 377066 240421
rect 377014 240357 377066 240363
rect 376630 239009 376682 239015
rect 376630 238951 376682 238957
rect 377026 233484 377054 240357
rect 377218 233780 377246 241763
rect 377314 238941 377342 246480
rect 377890 240907 377918 246494
rect 378166 241895 378218 241901
rect 378166 241837 378218 241843
rect 377876 240898 377932 240907
rect 377876 240833 377932 240842
rect 377782 240045 377834 240051
rect 377782 239987 377834 239993
rect 377302 238935 377354 238941
rect 377302 238877 377354 238883
rect 376800 233456 377054 233484
rect 377170 233752 377246 233780
rect 377170 233470 377198 233752
rect 377794 233484 377822 239987
rect 378178 233484 378206 241837
rect 378262 240341 378314 240347
rect 378262 240283 378314 240289
rect 377568 233456 377822 233484
rect 377904 233456 378206 233484
rect 378274 233470 378302 240283
rect 378370 237313 378398 246494
rect 378646 246409 378698 246415
rect 378646 246351 378698 246357
rect 378658 246267 378686 246351
rect 378646 246261 378698 246267
rect 378646 246203 378698 246209
rect 378646 239897 378698 239903
rect 378646 239839 378698 239845
rect 378358 237307 378410 237313
rect 378358 237249 378410 237255
rect 378658 233470 378686 239839
rect 378850 238391 378878 246494
rect 379042 246480 379296 246508
rect 379426 246480 379680 246508
rect 378836 238382 378892 238391
rect 378836 238317 378892 238326
rect 379042 237905 379070 246480
rect 379222 240785 379274 240791
rect 379222 240727 379274 240733
rect 379030 237899 379082 237905
rect 379030 237841 379082 237847
rect 379234 233484 379262 240727
rect 379426 234839 379454 246480
rect 379606 241081 379658 241087
rect 379606 241023 379658 241029
rect 379412 234830 379468 234839
rect 379412 234765 379468 234774
rect 379618 233484 379646 241023
rect 380098 239607 380126 246494
rect 380578 239829 380606 246494
rect 380566 239823 380618 239829
rect 380566 239765 380618 239771
rect 380086 239601 380138 239607
rect 380086 239543 380138 239549
rect 380854 239527 380906 239533
rect 380854 239469 380906 239475
rect 380086 239231 380138 239237
rect 380086 239173 380138 239179
rect 379990 237307 380042 237313
rect 379990 237249 380042 237255
rect 380002 233484 380030 237249
rect 379008 233456 379262 233484
rect 379392 233456 379646 233484
rect 379776 233456 380030 233484
rect 380098 233470 380126 239173
rect 380470 239009 380522 239015
rect 380470 238951 380522 238957
rect 380482 233470 380510 238951
rect 380866 233470 380894 239469
rect 380962 238571 380990 246494
rect 381154 246480 381408 246508
rect 381888 246480 382142 246508
rect 381046 238787 381098 238793
rect 381046 238729 381098 238735
rect 381058 238571 381086 238729
rect 380950 238565 381002 238571
rect 380950 238507 381002 238513
rect 381046 238565 381098 238571
rect 381046 238507 381098 238513
rect 381154 237757 381182 246480
rect 381814 240193 381866 240199
rect 381814 240135 381866 240141
rect 381430 238935 381482 238941
rect 381430 238877 381482 238883
rect 381142 237751 381194 237757
rect 381142 237693 381194 237699
rect 381442 233484 381470 238877
rect 381826 233484 381854 240135
rect 381910 235975 381962 235981
rect 381910 235917 381962 235923
rect 381216 233456 381470 233484
rect 381600 233456 381854 233484
rect 381922 233336 381950 235917
rect 382114 233484 382142 246480
rect 382306 238645 382334 246494
rect 382690 239681 382718 246494
rect 383074 246480 383184 246508
rect 383362 246480 383616 246508
rect 383842 246480 384096 246508
rect 382678 239675 382730 239681
rect 382678 239617 382730 239623
rect 383074 239108 383102 246480
rect 383254 239749 383306 239755
rect 383254 239691 383306 239697
rect 382978 239080 383102 239108
rect 382294 238639 382346 238645
rect 382294 238581 382346 238587
rect 382978 233484 383006 239080
rect 383266 233484 383294 239691
rect 383362 238719 383390 246480
rect 383842 239903 383870 246480
rect 384022 239971 384074 239977
rect 384022 239913 384074 239919
rect 383830 239897 383882 239903
rect 383830 239839 383882 239845
rect 383638 239675 383690 239681
rect 383638 239617 383690 239623
rect 383350 238713 383402 238719
rect 383350 238655 383402 238661
rect 383650 233484 383678 239617
rect 383734 239601 383786 239607
rect 383734 239543 383786 239549
rect 383746 233780 383774 239543
rect 384034 239089 384062 239913
rect 384418 239755 384446 246494
rect 384610 246480 384912 246508
rect 384406 239749 384458 239755
rect 384406 239691 384458 239697
rect 384022 239083 384074 239089
rect 384022 239025 384074 239031
rect 384610 238867 384638 246480
rect 385090 245971 385118 246721
rect 385078 245965 385130 245971
rect 385078 245907 385130 245913
rect 384886 239823 384938 239829
rect 384886 239765 384938 239771
rect 384598 238861 384650 238867
rect 384598 238803 384650 238809
rect 384406 237899 384458 237905
rect 384406 237841 384458 237847
rect 383746 233752 383822 233780
rect 382114 233456 382320 233484
rect 382704 233456 383006 233484
rect 383088 233456 383294 233484
rect 383424 233456 383678 233484
rect 383794 233470 383822 233752
rect 384418 233484 384446 237841
rect 384502 237751 384554 237757
rect 384502 237693 384554 237699
rect 384192 233456 384446 233484
rect 384514 233470 384542 237693
rect 384898 233470 384926 239765
rect 385270 238343 385322 238349
rect 385270 238285 385322 238291
rect 385282 233470 385310 238285
rect 385378 237313 385406 246494
rect 385570 246480 385824 246508
rect 385954 246480 386208 246508
rect 385570 239681 385598 246480
rect 385558 239675 385610 239681
rect 385558 239617 385610 239623
rect 385954 238571 385982 246480
rect 386626 239237 386654 246494
rect 387010 245749 387038 246721
rect 386998 245743 387050 245749
rect 386998 245685 387050 245691
rect 386614 239231 386666 239237
rect 386614 239173 386666 239179
rect 385942 238565 385994 238571
rect 385942 238507 385994 238513
rect 385366 237307 385418 237313
rect 385366 237249 385418 237255
rect 387106 236795 387134 246494
rect 387286 246335 387338 246341
rect 387286 246277 387338 246283
rect 387298 245897 387326 246277
rect 387394 246119 387422 246753
rect 388532 246753 388588 246762
rect 389492 246818 389548 246827
rect 389492 246753 389548 246762
rect 389780 246818 389836 246827
rect 405908 246818 405964 246827
rect 389780 246753 389836 246762
rect 390262 246779 390314 246785
rect 388054 246721 388106 246727
rect 387382 246113 387434 246119
rect 387382 246055 387434 246061
rect 387286 245891 387338 245897
rect 387286 245833 387338 245839
rect 387286 239749 387338 239755
rect 387286 239691 387338 239697
rect 387298 239459 387326 239691
rect 387286 239453 387338 239459
rect 387286 239395 387338 239401
rect 387586 239015 387614 246494
rect 387682 246480 387936 246508
rect 387574 239009 387626 239015
rect 387574 238951 387626 238957
rect 387682 237387 387710 246480
rect 388066 245823 388094 246721
rect 388162 246480 388416 246508
rect 388054 245817 388106 245823
rect 388054 245759 388106 245765
rect 388162 239533 388190 246480
rect 388546 246415 388574 246753
rect 389506 246711 389534 246753
rect 389494 246705 389546 246711
rect 389494 246647 389546 246653
rect 388534 246409 388586 246415
rect 388534 246351 388586 246357
rect 388150 239527 388202 239533
rect 388150 239469 388202 239475
rect 388834 238497 388862 246494
rect 388918 246335 388970 246341
rect 388918 246277 388970 246283
rect 388930 246119 388958 246277
rect 388918 246113 388970 246119
rect 388918 246055 388970 246061
rect 389218 238941 389246 246494
rect 389302 246187 389354 246193
rect 389302 246129 389354 246135
rect 389314 246045 389342 246129
rect 389302 246039 389354 246045
rect 389302 245981 389354 245987
rect 389302 244929 389354 244935
rect 389302 244871 389354 244877
rect 389314 243571 389342 244871
rect 389300 243562 389356 243571
rect 389300 243497 389356 243506
rect 389206 238935 389258 238941
rect 389206 238877 389258 238883
rect 388822 238491 388874 238497
rect 388822 238433 388874 238439
rect 389698 238423 389726 246494
rect 389794 246415 389822 246753
rect 390262 246721 390314 246727
rect 402166 246779 402218 246785
rect 405908 246753 405964 246762
rect 406100 246818 406156 246827
rect 406100 246753 406102 246762
rect 402166 246721 402218 246727
rect 389890 246480 390144 246508
rect 389782 246409 389834 246415
rect 389782 246351 389834 246357
rect 389890 240199 389918 246480
rect 390274 245749 390302 246721
rect 397654 246705 397706 246711
rect 397654 246647 397706 246653
rect 397666 246563 397694 246647
rect 402178 246637 402206 246721
rect 402070 246631 402122 246637
rect 402070 246573 402122 246579
rect 402166 246631 402218 246637
rect 402166 246573 402218 246579
rect 396790 246557 396842 246563
rect 390370 246480 390624 246508
rect 390262 245743 390314 245749
rect 390262 245685 390314 245691
rect 389878 240193 389930 240199
rect 389878 240135 389930 240141
rect 389686 238417 389738 238423
rect 389686 238359 389738 238365
rect 390370 238275 390398 246480
rect 390358 238269 390410 238275
rect 390358 238211 390410 238217
rect 387670 237381 387722 237387
rect 387670 237323 387722 237329
rect 387094 236789 387146 236795
rect 387094 236731 387146 236737
rect 390946 235981 390974 246494
rect 391426 238095 391454 246494
rect 391412 238086 391468 238095
rect 391412 238021 391468 238030
rect 391906 237979 391934 246494
rect 392098 246480 392352 246508
rect 392482 246480 392736 246508
rect 392098 239385 392126 246480
rect 392086 239379 392138 239385
rect 392086 239321 392138 239327
rect 392482 238053 392510 246480
rect 392470 238047 392522 238053
rect 392470 237989 392522 237995
rect 391894 237973 391946 237979
rect 393154 237947 393182 246494
rect 393634 238127 393662 246494
rect 394114 239311 394142 246494
rect 394210 246480 394464 246508
rect 394690 246480 394944 246508
rect 394102 239305 394154 239311
rect 394102 239247 394154 239253
rect 394210 238201 394238 246480
rect 394198 238195 394250 238201
rect 394198 238137 394250 238143
rect 393622 238121 393674 238127
rect 393622 238063 393674 238069
rect 391894 237915 391946 237921
rect 393140 237938 393196 237947
rect 393140 237873 393196 237882
rect 394690 237799 394718 246480
rect 394676 237790 394732 237799
rect 394676 237725 394732 237734
rect 395362 237535 395390 246494
rect 395842 241605 395870 246494
rect 395926 241821 395978 241827
rect 395926 241763 395978 241769
rect 395938 241605 395966 241763
rect 395830 241599 395882 241605
rect 395830 241541 395882 241547
rect 395926 241599 395978 241605
rect 395926 241541 395978 241547
rect 395350 237529 395402 237535
rect 395350 237471 395402 237477
rect 396226 237461 396254 246494
rect 396418 246480 396672 246508
rect 397654 246557 397706 246563
rect 396790 246499 396842 246505
rect 396418 241753 396446 246480
rect 396802 246193 396830 246499
rect 396898 246480 397152 246508
rect 397654 246499 397706 246505
rect 397366 246483 397418 246489
rect 396790 246187 396842 246193
rect 396790 246129 396842 246135
rect 396406 241747 396458 241753
rect 396406 241689 396458 241695
rect 396898 239163 396926 246480
rect 397366 246425 397418 246431
rect 397378 245823 397406 246425
rect 397366 245817 397418 245823
rect 397366 245759 397418 245765
rect 397474 241531 397502 246494
rect 397462 241525 397514 241531
rect 397462 241467 397514 241473
rect 396886 239157 396938 239163
rect 396886 239099 396938 239105
rect 397954 237683 397982 246494
rect 398434 241383 398462 246494
rect 398626 246480 398880 246508
rect 399010 246480 399264 246508
rect 398422 241377 398474 241383
rect 398422 241319 398474 241325
rect 398626 239977 398654 246480
rect 399010 241161 399038 246480
rect 398998 241155 399050 241161
rect 398998 241097 399050 241103
rect 398614 239971 398666 239977
rect 398614 239913 398666 239919
rect 397942 237677 397994 237683
rect 397942 237619 397994 237625
rect 399682 237609 399710 246494
rect 400162 241679 400190 246494
rect 400150 241673 400202 241679
rect 400150 241615 400202 241621
rect 400642 239755 400670 246494
rect 400738 246480 400992 246508
rect 401218 246480 401472 246508
rect 400738 241309 400766 246480
rect 400726 241303 400778 241309
rect 400726 241245 400778 241251
rect 400630 239749 400682 239755
rect 400630 239691 400682 239697
rect 401218 237831 401246 246480
rect 401890 241235 401918 246494
rect 402082 245749 402110 246573
rect 402070 245743 402122 245749
rect 402070 245685 402122 245691
rect 401878 241229 401930 241235
rect 401878 241171 401930 241177
rect 402370 239903 402398 246494
rect 402754 241457 402782 246494
rect 403200 246480 403262 246508
rect 402742 241451 402794 241457
rect 402742 241393 402794 241399
rect 403234 240125 403262 246480
rect 403426 246480 403680 246508
rect 403426 240569 403454 246480
rect 403414 240563 403466 240569
rect 403414 240505 403466 240511
rect 404098 240273 404126 246494
rect 404482 240643 404510 246494
rect 404470 240637 404522 240643
rect 404470 240579 404522 240585
rect 404962 240421 404990 246494
rect 405154 246480 405408 246508
rect 405538 246480 405792 246508
rect 405154 240939 405182 246480
rect 405538 241605 405566 246480
rect 405922 245453 405950 246753
rect 406154 246753 406156 246762
rect 406496 246758 406520 246834
rect 406598 246758 406612 246834
rect 406496 246744 406612 246758
rect 406772 246818 406828 246827
rect 406772 246753 406828 246762
rect 407060 246818 407116 246827
rect 407060 246753 407116 246762
rect 407252 246818 407308 246827
rect 407252 246753 407308 246762
rect 407636 246818 407692 246827
rect 407636 246753 407692 246762
rect 408116 246818 408172 246827
rect 408116 246753 408172 246762
rect 408596 246818 408652 246827
rect 408596 246753 408652 246762
rect 408788 246818 408844 246827
rect 408788 246753 408844 246762
rect 408980 246818 409036 246827
rect 408980 246753 408982 246762
rect 406102 246721 406154 246727
rect 406786 246637 406814 246753
rect 406774 246631 406826 246637
rect 406774 246573 406826 246579
rect 406114 246480 406272 246508
rect 405910 245447 405962 245453
rect 405910 245389 405962 245395
rect 405718 245151 405770 245157
rect 405718 245093 405770 245099
rect 405730 243571 405758 245093
rect 405716 243562 405772 243571
rect 405716 243497 405772 243506
rect 405526 241599 405578 241605
rect 405526 241541 405578 241547
rect 405142 240933 405194 240939
rect 405142 240875 405194 240881
rect 406114 240865 406142 246480
rect 406198 246187 406250 246193
rect 406198 246129 406250 246135
rect 406210 243571 406238 246129
rect 406196 243562 406252 243571
rect 406196 243497 406252 243506
rect 406102 240859 406154 240865
rect 406102 240801 406154 240807
rect 404950 240415 405002 240421
rect 404950 240357 405002 240363
rect 404086 240267 404138 240273
rect 404086 240209 404138 240215
rect 403222 240119 403274 240125
rect 403222 240061 403274 240067
rect 406690 240051 406718 246494
rect 407074 245749 407102 246753
rect 407062 245743 407114 245749
rect 407062 245685 407114 245691
rect 407170 240495 407198 246494
rect 407266 246489 407294 246753
rect 407254 246483 407306 246489
rect 407254 246425 407306 246431
rect 407554 241827 407582 246494
rect 407650 246341 407678 246753
rect 407746 246480 408000 246508
rect 407638 246335 407690 246341
rect 407638 246277 407690 246283
rect 407542 241821 407594 241827
rect 407542 241763 407594 241769
rect 407746 240717 407774 246480
rect 408130 244861 408158 246753
rect 408322 246480 408480 246508
rect 408118 244855 408170 244861
rect 408118 244797 408170 244803
rect 407734 240711 407786 240717
rect 407734 240653 407786 240659
rect 407158 240489 407210 240495
rect 407158 240431 407210 240437
rect 408322 240347 408350 246480
rect 408610 246415 408638 246753
rect 408802 246711 408830 246753
rect 409034 246753 409036 246762
rect 409172 246818 409228 246827
rect 409172 246753 409228 246762
rect 409364 246818 409420 246827
rect 409844 246818 409900 246827
rect 409364 246753 409366 246762
rect 408982 246721 409034 246727
rect 408790 246705 408842 246711
rect 408790 246647 408842 246653
rect 408598 246409 408650 246415
rect 408598 246351 408650 246357
rect 408898 241013 408926 246494
rect 409186 245971 409214 246753
rect 409418 246753 409420 246762
rect 409462 246779 409514 246785
rect 409366 246721 409418 246727
rect 409844 246753 409900 246762
rect 409462 246721 409514 246727
rect 409174 245965 409226 245971
rect 409174 245907 409226 245913
rect 408886 241007 408938 241013
rect 408886 240949 408938 240955
rect 409282 240791 409310 246494
rect 409474 245897 409502 246721
rect 409462 245891 409514 245897
rect 409462 245833 409514 245839
rect 409270 240785 409322 240791
rect 409270 240727 409322 240733
rect 409762 240463 409790 246494
rect 409858 246045 409886 246753
rect 412066 246563 412094 247197
rect 412162 246785 412190 247493
rect 412436 247410 412492 247419
rect 412436 247345 412492 247354
rect 412244 247114 412300 247123
rect 412244 247049 412300 247058
rect 412150 246779 412202 246785
rect 412150 246721 412202 246727
rect 412054 246557 412106 246563
rect 409954 246480 410208 246508
rect 410434 246480 410688 246508
rect 412054 246499 412106 246505
rect 409846 246039 409898 246045
rect 409846 245981 409898 245987
rect 409954 241087 409982 246480
rect 409942 241081 409994 241087
rect 409942 241023 409994 241029
rect 409748 240454 409804 240463
rect 409748 240389 409804 240398
rect 408310 240341 408362 240347
rect 408310 240283 408362 240289
rect 406678 240045 406730 240051
rect 406678 239987 406730 239993
rect 402358 239897 402410 239903
rect 402358 239839 402410 239845
rect 410434 237905 410462 246480
rect 410422 237899 410474 237905
rect 410422 237841 410474 237847
rect 401206 237825 401258 237831
rect 401206 237767 401258 237773
rect 411010 237757 411038 246494
rect 411490 245231 411518 246494
rect 411478 245225 411530 245231
rect 411478 245167 411530 245173
rect 410998 237751 411050 237757
rect 410998 237693 411050 237699
rect 411970 237651 411998 246494
rect 412258 246267 412286 247049
rect 412246 246261 412298 246267
rect 412246 246203 412298 246209
rect 412450 245453 412478 247345
rect 412438 245447 412490 245453
rect 412438 245389 412490 245395
rect 412642 238835 412670 247516
rect 505366 246113 505418 246119
rect 505366 246055 505418 246061
rect 463702 242709 463754 242715
rect 453620 242674 453676 242683
rect 453620 242609 453676 242618
rect 463700 242674 463702 242683
rect 483766 242709 483818 242715
rect 463754 242674 463756 242683
rect 483766 242651 483818 242657
rect 463700 242609 463756 242618
rect 453634 242567 453662 242609
rect 443638 242561 443690 242567
rect 430484 242526 430540 242535
rect 430484 242461 430540 242470
rect 443444 242526 443500 242535
rect 443444 242461 443500 242470
rect 443636 242526 443638 242535
rect 453622 242561 453674 242567
rect 443690 242526 443692 242535
rect 483778 242535 483806 242651
rect 453622 242503 453674 242509
rect 483764 242526 483820 242535
rect 443636 242461 443692 242470
rect 483764 242461 483820 242470
rect 489524 242526 489580 242535
rect 489580 242484 489758 242512
rect 489524 242461 489580 242470
rect 430498 242419 430526 242461
rect 443458 242419 443486 242461
rect 430486 242413 430538 242419
rect 430486 242355 430538 242361
rect 443446 242413 443498 242419
rect 489730 242387 489758 242484
rect 504022 242413 504074 242419
rect 443446 242355 443498 242361
rect 489716 242378 489772 242387
rect 489716 242313 489772 242322
rect 504020 242378 504022 242387
rect 504074 242378 504076 242387
rect 504020 242313 504076 242322
rect 412628 238826 412684 238835
rect 412628 238761 412684 238770
rect 497494 237677 497546 237683
rect 411956 237642 412012 237651
rect 399670 237603 399722 237609
rect 505378 237651 505406 246055
rect 511126 242413 511178 242419
rect 511126 242355 511178 242361
rect 511138 237799 511166 242355
rect 547522 238983 547550 257728
rect 576226 241943 576254 277856
rect 578530 275201 578558 277870
rect 579682 276015 579710 277870
rect 579670 276009 579722 276015
rect 579670 275951 579722 275957
rect 580930 275687 580958 277870
rect 580916 275678 580972 275687
rect 580916 275613 580972 275622
rect 578518 275195 578570 275201
rect 578518 275137 578570 275143
rect 582082 270359 582110 277870
rect 582068 270350 582124 270359
rect 582068 270285 582124 270294
rect 583234 270095 583262 277870
rect 584386 271099 584414 277870
rect 585634 275053 585662 277870
rect 585622 275047 585674 275053
rect 585622 274989 585674 274995
rect 584372 271090 584428 271099
rect 584372 271025 584428 271034
rect 583222 270089 583274 270095
rect 580244 270054 580300 270063
rect 583222 270031 583274 270037
rect 586786 270021 586814 277870
rect 587938 272389 587966 277870
rect 587926 272383 587978 272389
rect 587926 272325 587978 272331
rect 589186 270211 589214 277870
rect 590338 271353 590366 277870
rect 591586 272463 591614 277870
rect 592738 276427 592766 277870
rect 592724 276418 592780 276427
rect 592724 276353 592780 276362
rect 591574 272457 591626 272463
rect 591574 272399 591626 272405
rect 593986 271427 594014 277870
rect 595138 272611 595166 277870
rect 595126 272605 595178 272611
rect 595126 272547 595178 272553
rect 593974 271421 594026 271427
rect 593974 271363 594026 271369
rect 590326 271347 590378 271353
rect 590326 271289 590378 271295
rect 589172 270202 589228 270211
rect 589172 270137 589228 270146
rect 580244 269989 580300 269998
rect 586774 270015 586826 270021
rect 580258 268879 580286 269989
rect 586774 269957 586826 269963
rect 596386 268879 596414 277870
rect 597538 269725 597566 277870
rect 599842 276279 599870 277870
rect 599828 276270 599884 276279
rect 599828 276205 599884 276214
rect 601090 275719 601118 277870
rect 601078 275713 601130 275719
rect 601078 275655 601130 275661
rect 602242 275539 602270 277870
rect 602228 275530 602284 275539
rect 602228 275465 602284 275474
rect 603394 269915 603422 277870
rect 603380 269906 603436 269915
rect 603380 269841 603436 269850
rect 597526 269719 597578 269725
rect 597526 269661 597578 269667
rect 604642 269577 604670 277870
rect 605794 269767 605822 277870
rect 607042 272315 607070 277870
rect 607030 272309 607082 272315
rect 607030 272251 607082 272257
rect 605780 269758 605836 269767
rect 605780 269693 605836 269702
rect 604630 269571 604682 269577
rect 604630 269513 604682 269519
rect 580244 268870 580300 268879
rect 580244 268805 580300 268814
rect 596372 268870 596428 268879
rect 596372 268805 596428 268814
rect 608194 267357 608222 277870
rect 608182 267351 608234 267357
rect 608182 267293 608234 267299
rect 609442 266215 609470 277870
rect 610594 276131 610622 277870
rect 611842 276681 611870 277870
rect 611830 276675 611882 276681
rect 611830 276617 611882 276623
rect 610580 276122 610636 276131
rect 610580 276057 610636 276066
rect 612994 273573 613022 277870
rect 612982 273567 613034 273573
rect 612982 273509 613034 273515
rect 614242 267843 614270 277870
rect 614228 267834 614284 267843
rect 614228 267769 614284 267778
rect 609428 266206 609484 266215
rect 609428 266141 609484 266150
rect 615394 265137 615422 277870
rect 616546 275391 616574 277870
rect 617698 277019 617726 277870
rect 617684 277010 617740 277019
rect 617684 276945 617740 276954
rect 616532 275382 616588 275391
rect 616532 275317 616588 275326
rect 618850 272019 618878 277870
rect 618838 272013 618890 272019
rect 618838 271955 618890 271961
rect 620098 269619 620126 277870
rect 620084 269610 620140 269619
rect 620084 269545 620140 269554
rect 621250 267801 621278 277870
rect 622498 275423 622526 277870
rect 622486 275417 622538 275423
rect 622486 275359 622538 275365
rect 623650 275243 623678 277870
rect 624898 275983 624926 277870
rect 624884 275974 624940 275983
rect 624884 275909 624940 275918
rect 623636 275234 623692 275243
rect 623636 275169 623692 275178
rect 626050 268435 626078 277870
rect 627298 275095 627326 277870
rect 627284 275086 627340 275095
rect 627284 275021 627340 275030
rect 626036 268426 626092 268435
rect 626036 268361 626092 268370
rect 621238 267795 621290 267801
rect 621238 267737 621290 267743
rect 628450 265475 628478 277870
rect 628436 265466 628492 265475
rect 628436 265401 628492 265410
rect 615382 265131 615434 265137
rect 615382 265073 615434 265079
rect 629698 265063 629726 277870
rect 630742 273641 630794 273647
rect 630742 273583 630794 273589
rect 629686 265057 629738 265063
rect 629686 264999 629738 265005
rect 630754 257811 630782 273583
rect 630850 269471 630878 277870
rect 631810 277856 632112 277884
rect 630836 269462 630892 269471
rect 630836 269397 630892 269406
rect 631810 265919 631838 277856
rect 633154 275349 633182 277870
rect 633142 275343 633194 275349
rect 633142 275285 633194 275291
rect 634306 269323 634334 277870
rect 636706 276607 636734 277870
rect 636694 276601 636746 276607
rect 636694 276543 636746 276549
rect 637954 275835 637982 277870
rect 637940 275826 637996 275835
rect 637940 275761 637996 275770
rect 634292 269314 634348 269323
rect 634292 269249 634348 269258
rect 639106 267695 639134 277870
rect 639382 276823 639434 276829
rect 639382 276765 639434 276771
rect 639394 273647 639422 276765
rect 639382 273641 639434 273647
rect 639382 273583 639434 273589
rect 640354 269175 640382 277870
rect 641506 270655 641534 277870
rect 642754 276871 642782 277870
rect 642740 276862 642796 276871
rect 642740 276797 642796 276806
rect 642262 273567 642314 273573
rect 642262 273509 642314 273515
rect 641492 270646 641548 270655
rect 641492 270581 641548 270590
rect 640340 269166 640396 269175
rect 640340 269101 640396 269110
rect 639092 267686 639148 267695
rect 639092 267621 639148 267630
rect 631796 265910 631852 265919
rect 631796 265845 631852 265854
rect 642274 265008 642302 273509
rect 643906 272907 643934 277870
rect 645154 274947 645182 277870
rect 646306 276723 646334 277870
rect 646292 276714 646348 276723
rect 646292 276649 646348 276658
rect 647554 275127 647582 277870
rect 648034 277856 648720 277884
rect 647542 275121 647594 275127
rect 647542 275063 647594 275069
rect 645140 274938 645196 274947
rect 645140 274873 645196 274882
rect 643894 272901 643946 272907
rect 643894 272843 643946 272849
rect 642178 264980 642302 265008
rect 642178 259291 642206 264980
rect 632470 259285 632522 259291
rect 632470 259227 632522 259233
rect 642166 259285 642218 259291
rect 642166 259227 642218 259233
rect 616342 257805 616394 257811
rect 616342 257747 616394 257753
rect 630742 257805 630794 257811
rect 630742 257747 630794 257753
rect 616354 250633 616382 257747
rect 616342 250627 616394 250633
rect 616342 250569 616394 250575
rect 607702 250553 607754 250559
rect 607702 250495 607754 250501
rect 607714 244861 607742 250495
rect 632482 248117 632510 259227
rect 639286 256399 639338 256405
rect 639286 256341 639338 256347
rect 627862 248111 627914 248117
rect 627862 248053 627914 248059
rect 632470 248111 632522 248117
rect 632470 248053 632522 248059
rect 607702 244855 607754 244861
rect 607702 244797 607754 244803
rect 603094 244781 603146 244787
rect 603094 244723 603146 244729
rect 576212 241934 576268 241943
rect 576212 241869 576268 241878
rect 603106 239237 603134 244723
rect 627874 240495 627902 248053
rect 607606 240489 607658 240495
rect 607606 240431 607658 240437
rect 627862 240489 627914 240495
rect 627862 240431 627914 240437
rect 596182 239231 596234 239237
rect 596182 239173 596234 239179
rect 603094 239231 603146 239237
rect 603094 239173 603146 239179
rect 547508 238974 547564 238983
rect 547508 238909 547564 238918
rect 511124 237790 511180 237799
rect 511124 237725 511180 237734
rect 549238 237751 549290 237757
rect 497494 237619 497546 237625
rect 505364 237642 505420 237651
rect 411956 237577 412012 237586
rect 420598 237603 420650 237609
rect 399670 237545 399722 237551
rect 420598 237545 420650 237551
rect 396214 237455 396266 237461
rect 396214 237397 396266 237403
rect 400340 236754 400396 236763
rect 400340 236689 400342 236698
rect 400394 236689 400396 236698
rect 420404 236754 420460 236763
rect 420404 236689 420406 236698
rect 400342 236657 400394 236663
rect 420458 236689 420460 236698
rect 420406 236657 420458 236663
rect 420610 236467 420638 237545
rect 440660 236754 440716 236763
rect 440660 236689 440662 236698
rect 440714 236689 440716 236698
rect 460724 236754 460780 236763
rect 460724 236689 460726 236698
rect 440662 236657 440714 236663
rect 460778 236689 460780 236698
rect 480980 236754 481036 236763
rect 480980 236689 481036 236698
rect 460726 236657 460778 236663
rect 420596 236458 420652 236467
rect 420596 236393 420652 236402
rect 390934 235975 390986 235981
rect 390934 235917 390986 235923
rect 420610 233470 420638 236393
rect 480994 235759 481022 236689
rect 497506 235759 497534 237619
rect 505364 237577 505420 237586
rect 480982 235753 481034 235759
rect 480982 235695 481034 235701
rect 497494 235753 497546 235759
rect 497494 235695 497546 235701
rect 497506 233470 497534 235695
rect 505378 233484 505406 237577
rect 511138 233484 511166 237725
rect 549238 237693 549290 237699
rect 549250 236203 549278 237693
rect 596194 237683 596222 239173
rect 596182 237677 596234 237683
rect 596182 237619 596234 237625
rect 607618 237609 607646 240431
rect 607606 237603 607658 237609
rect 607606 237545 607658 237551
rect 638038 236567 638090 236573
rect 638038 236509 638090 236515
rect 637366 236493 637418 236499
rect 637366 236435 637418 236441
rect 547126 236197 547178 236203
rect 547126 236139 547178 236145
rect 549238 236197 549290 236203
rect 549238 236139 549290 236145
rect 547138 234691 547166 236139
rect 547124 234682 547180 234691
rect 547124 234617 547180 234626
rect 549250 233484 549278 236139
rect 637172 233646 637228 233655
rect 637172 233581 637228 233590
rect 505378 233456 505632 233484
rect 510384 233456 511166 233484
rect 549024 233456 549278 233484
rect 637186 233484 637214 233581
rect 637378 233484 637406 236435
rect 637942 236419 637994 236425
rect 637942 236361 637994 236367
rect 637186 233456 637406 233484
rect 637460 233498 637516 233507
rect 637954 233484 637982 236361
rect 638050 233951 638078 236509
rect 639190 236345 639242 236351
rect 638420 236310 638476 236319
rect 639298 236319 639326 256341
rect 648034 243719 648062 277856
rect 648020 243710 648076 243719
rect 648020 243645 648076 243654
rect 649378 237757 649406 995083
rect 650036 994514 650092 994523
rect 650036 994449 650092 994458
rect 649748 994218 649804 994227
rect 649748 994153 649804 994162
rect 649652 994070 649708 994079
rect 649652 994005 649708 994014
rect 649558 983597 649610 983603
rect 649558 983539 649610 983545
rect 649462 983523 649514 983529
rect 649462 983465 649514 983471
rect 649474 273647 649502 983465
rect 649570 276829 649598 983539
rect 649666 941835 649694 994005
rect 649652 941826 649708 941835
rect 649652 941761 649708 941770
rect 649654 927431 649706 927437
rect 649654 927373 649706 927379
rect 649558 276823 649610 276829
rect 649558 276765 649610 276771
rect 649462 273641 649514 273647
rect 649462 273583 649514 273589
rect 649366 237751 649418 237757
rect 649366 237693 649418 237699
rect 639190 236287 639242 236293
rect 639284 236310 639340 236319
rect 638420 236245 638476 236254
rect 638806 236271 638858 236277
rect 638036 233942 638092 233951
rect 638036 233877 638092 233886
rect 637516 233456 637982 233484
rect 637460 233433 637516 233442
rect 638050 233336 638078 233877
rect 638228 233498 638284 233507
rect 638434 233484 638462 236245
rect 638806 236213 638858 236219
rect 638818 233803 638846 236213
rect 638804 233794 638860 233803
rect 638804 233729 638860 233738
rect 638284 233470 638462 233484
rect 638818 233470 638846 233729
rect 638900 233646 638956 233655
rect 638900 233581 638956 233590
rect 638914 233484 638942 233581
rect 639202 233484 639230 236287
rect 649666 236277 649694 927373
rect 649762 848299 649790 994153
rect 649846 989295 649898 989301
rect 649846 989237 649898 989243
rect 649748 848290 649804 848299
rect 649748 848225 649804 848234
rect 649750 748869 649802 748875
rect 649750 748811 649802 748817
rect 639284 236245 639340 236254
rect 649654 236271 649706 236277
rect 649654 236213 649706 236219
rect 639766 236197 639818 236203
rect 639766 236139 639818 236145
rect 639778 233484 639806 236139
rect 638914 233470 639230 233484
rect 638284 233456 638448 233470
rect 638914 233456 639216 233470
rect 639552 233456 639806 233484
rect 638228 233433 638284 233442
rect 227362 233308 227424 233336
rect 359842 233308 359904 233336
rect 381922 233308 381984 233336
rect 638050 233308 638112 233336
rect 210274 62673 210398 62692
rect 210262 62667 210398 62673
rect 210314 62664 210398 62667
rect 210262 62609 210314 62615
rect 210164 62558 210220 62567
rect 210164 62493 210220 62502
rect 210260 58044 210316 58053
rect 210316 58002 210398 58030
rect 210260 57979 210316 57988
rect 210260 56934 210316 56943
rect 210260 56869 210316 56878
rect 210164 55306 210220 55315
rect 210164 55241 210220 55250
rect 210178 53719 210206 55241
rect 210274 54385 210302 56869
rect 210262 54379 210314 54385
rect 210262 54321 210314 54327
rect 210260 54122 210316 54131
rect 210260 54057 210316 54066
rect 210166 53713 210218 53719
rect 210166 53655 210218 53661
rect 210274 53349 210302 54057
rect 210370 53867 210398 58002
rect 217462 54305 217514 54311
rect 210452 54270 210508 54279
rect 210452 54205 210508 54214
rect 210644 54270 210700 54279
rect 210644 54205 210700 54214
rect 214772 54270 214828 54279
rect 214828 54228 214896 54256
rect 219382 54305 219434 54311
rect 217462 54247 217514 54253
rect 217474 54242 217502 54247
rect 219202 54237 219312 54256
rect 219382 54247 219434 54253
rect 219190 54231 219312 54237
rect 214772 54205 214828 54214
rect 210358 53861 210410 53867
rect 210358 53803 210410 53809
rect 210262 53343 210314 53349
rect 210262 53285 210314 53291
rect 210466 53201 210494 54205
rect 210658 53423 210686 54205
rect 219242 54228 219312 54231
rect 219190 54173 219242 54179
rect 213766 54157 213818 54163
rect 213766 54099 213818 54105
rect 216980 54122 217036 54131
rect 213778 54094 213806 54099
rect 217036 54080 217104 54108
rect 216980 54057 217036 54066
rect 218182 54009 218234 54015
rect 216980 53974 217036 53983
rect 214966 53935 215018 53941
rect 218182 53951 218234 53957
rect 218194 53946 218222 53951
rect 216980 53909 217036 53918
rect 214966 53877 215018 53883
rect 210646 53417 210698 53423
rect 210646 53359 210698 53365
rect 210454 53195 210506 53201
rect 210454 53137 210506 53143
rect 210070 48903 210122 48909
rect 210070 48845 210122 48851
rect 209206 48237 209258 48243
rect 209206 48179 209258 48185
rect 209302 48237 209354 48243
rect 209302 48179 209354 48185
rect 209218 46689 209246 48179
rect 209206 46683 209258 46689
rect 209206 46625 209258 46631
rect 208822 46461 208874 46467
rect 208822 46403 208874 46409
rect 208726 46387 208778 46393
rect 208726 46329 208778 46335
rect 208534 46313 208586 46319
rect 208534 46255 208586 46261
rect 206382 42023 207408 42051
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 211042 40663 211070 53650
rect 211200 53636 211262 53664
rect 211392 53636 211454 53664
rect 211234 52461 211262 53636
rect 211222 52455 211274 52461
rect 211222 52397 211274 52403
rect 211426 44987 211454 53636
rect 211570 53368 211598 53650
rect 211714 53636 211776 53664
rect 211906 53636 211968 53664
rect 211570 53340 211646 53368
rect 211618 52831 211646 53340
rect 211606 52825 211658 52831
rect 211606 52767 211658 52773
rect 211510 50457 211562 50463
rect 211510 50399 211562 50405
rect 211522 49649 211550 50399
rect 211510 49643 211562 49649
rect 211510 49585 211562 49591
rect 211414 44981 211466 44987
rect 211414 44923 211466 44929
rect 211714 44839 211742 53636
rect 211906 52059 211934 53636
rect 211892 52050 211948 52059
rect 211892 51985 211948 51994
rect 212098 45061 212126 53650
rect 212290 52535 212318 53650
rect 212278 52529 212330 52535
rect 212278 52471 212330 52477
rect 212086 45055 212138 45061
rect 212086 44997 212138 45003
rect 211702 44833 211754 44839
rect 211702 44775 211754 44781
rect 212482 44691 212510 53650
rect 212674 51911 212702 53650
rect 212660 51902 212716 51911
rect 212660 51837 212716 51846
rect 212866 44807 212894 53650
rect 213058 53539 213086 53650
rect 213044 53530 213100 53539
rect 213044 53465 213100 53474
rect 213250 45251 213278 53650
rect 213408 53636 213470 53664
rect 213600 53636 213662 53664
rect 213442 53201 213470 53636
rect 213430 53195 213482 53201
rect 213430 53137 213482 53143
rect 213430 52529 213482 52535
rect 213430 52471 213482 52477
rect 213442 51869 213470 52471
rect 213430 51863 213482 51869
rect 213430 51805 213482 51811
rect 213236 45242 213292 45251
rect 213236 45177 213292 45186
rect 212852 44798 212908 44807
rect 212852 44733 212908 44742
rect 212470 44685 212522 44691
rect 212470 44627 212522 44633
rect 213634 42249 213662 53636
rect 213922 53636 213984 53664
rect 214114 53636 214176 53664
rect 213814 52455 213866 52461
rect 213814 52397 213866 52403
rect 213826 51795 213854 52397
rect 213814 51789 213866 51795
rect 213814 51731 213866 51737
rect 213922 44913 213950 53636
rect 214114 51721 214142 53636
rect 214102 51715 214154 51721
rect 214102 51657 214154 51663
rect 213910 44907 213962 44913
rect 213910 44849 213962 44855
rect 213622 42243 213674 42249
rect 213622 42185 213674 42191
rect 214306 42175 214334 53650
rect 214498 51647 214526 53650
rect 214486 51641 214538 51647
rect 214486 51583 214538 51589
rect 214690 45103 214718 53650
rect 214978 53539 215006 53877
rect 215616 53784 215678 53812
rect 214964 53530 215020 53539
rect 214964 53465 215020 53474
rect 214676 45094 214732 45103
rect 214676 45029 214732 45038
rect 215074 43285 215102 53650
rect 215266 53571 215294 53650
rect 215254 53565 215306 53571
rect 215254 53507 215306 53513
rect 215458 44955 215486 53650
rect 215650 53275 215678 53784
rect 215794 53539 215822 53650
rect 215986 53539 216014 53650
rect 216130 53636 216192 53664
rect 215780 53530 215836 53539
rect 215780 53465 215836 53474
rect 215972 53530 216028 53539
rect 215972 53465 216028 53474
rect 215638 53269 215690 53275
rect 215638 53211 215690 53217
rect 216130 50611 216158 53636
rect 216370 53571 216398 53650
rect 216358 53565 216410 53571
rect 216358 53507 216410 53513
rect 216514 52757 216542 53650
rect 216706 53391 216734 53650
rect 216692 53382 216748 53391
rect 216692 53317 216748 53326
rect 216502 52751 216554 52757
rect 216502 52693 216554 52699
rect 216118 50605 216170 50611
rect 216118 50547 216170 50553
rect 216898 50537 216926 53650
rect 216994 53053 217022 53909
rect 217824 53784 217886 53812
rect 216982 53047 217034 53053
rect 216982 52989 217034 52995
rect 217282 52905 217310 53650
rect 217270 52899 217322 52905
rect 217270 52841 217322 52847
rect 216886 50531 216938 50537
rect 216886 50473 216938 50479
rect 217666 47651 217694 53650
rect 217858 53243 217886 53784
rect 219190 53787 219242 53793
rect 219190 53729 219242 53735
rect 218016 53636 218078 53664
rect 217844 53234 217900 53243
rect 217844 53169 217900 53178
rect 218050 47725 218078 53636
rect 218338 53636 218400 53664
rect 218038 47719 218090 47725
rect 218038 47661 218090 47667
rect 217654 47645 217706 47651
rect 217654 47587 217706 47593
rect 218338 47577 218366 53636
rect 218578 53368 218606 53650
rect 218578 53340 218654 53368
rect 218626 48983 218654 53340
rect 218614 48977 218666 48983
rect 218614 48919 218666 48925
rect 218326 47571 218378 47577
rect 218326 47513 218378 47519
rect 218722 47503 218750 53650
rect 218914 53497 218942 53650
rect 218902 53491 218954 53497
rect 218902 53433 218954 53439
rect 219106 48095 219134 53650
rect 219202 53497 219230 53729
rect 219190 53491 219242 53497
rect 219190 53433 219242 53439
rect 219394 53423 219422 54247
rect 221398 53861 221450 53867
rect 221398 53803 221450 53809
rect 219382 53417 219434 53423
rect 219382 53359 219434 53365
rect 219094 48089 219146 48095
rect 219094 48031 219146 48037
rect 219490 47873 219518 53650
rect 219682 53349 219710 53650
rect 219670 53343 219722 53349
rect 219670 53285 219722 53291
rect 219874 52239 219902 53650
rect 220032 53636 220094 53664
rect 219958 52825 220010 52831
rect 219958 52767 220010 52773
rect 219862 52233 219914 52239
rect 219862 52175 219914 52181
rect 219970 51869 219998 52767
rect 219958 51863 220010 51869
rect 219958 51805 220010 51811
rect 220066 48835 220094 53636
rect 220210 53368 220238 53650
rect 220402 53405 220430 53650
rect 220162 53340 220238 53368
rect 220354 53377 220430 53405
rect 220546 53636 220608 53664
rect 220738 53636 220800 53664
rect 220054 48829 220106 48835
rect 220054 48771 220106 48777
rect 219478 47867 219530 47873
rect 219478 47809 219530 47815
rect 220162 47799 220190 53340
rect 220354 53127 220382 53377
rect 220342 53121 220394 53127
rect 220342 53063 220394 53069
rect 220246 49051 220298 49057
rect 220246 48993 220298 48999
rect 220258 48835 220286 48993
rect 220246 48829 220298 48835
rect 220246 48771 220298 48777
rect 220546 47947 220574 53636
rect 220738 48909 220766 53636
rect 220930 52091 220958 53650
rect 221122 53539 221150 53650
rect 221108 53530 221164 53539
rect 221108 53465 221164 53474
rect 220918 52085 220970 52091
rect 220918 52027 220970 52033
rect 220726 48903 220778 48909
rect 220726 48845 220778 48851
rect 221314 48021 221342 53650
rect 221410 53349 221438 53803
rect 221398 53343 221450 53349
rect 221398 53285 221450 53291
rect 221506 50389 221534 53650
rect 221494 50383 221546 50389
rect 221494 50325 221546 50331
rect 221698 48761 221726 53650
rect 221890 52207 221918 53650
rect 221876 52198 221932 52207
rect 221876 52133 221932 52142
rect 221686 48755 221738 48761
rect 221686 48697 221738 48703
rect 222082 48169 222110 53650
rect 222240 53636 222302 53664
rect 222432 53636 222494 53664
rect 222274 48761 222302 53636
rect 222262 48755 222314 48761
rect 222262 48697 222314 48703
rect 222466 48687 222494 53636
rect 222610 53368 222638 53650
rect 222754 53636 222816 53664
rect 222946 53636 223008 53664
rect 222610 53340 222686 53368
rect 222658 51615 222686 53340
rect 222644 51606 222700 51615
rect 222644 51541 222700 51550
rect 222454 48681 222506 48687
rect 222454 48623 222506 48629
rect 222754 48243 222782 53636
rect 222946 48687 222974 53636
rect 222934 48681 222986 48687
rect 222934 48623 222986 48629
rect 222742 48237 222794 48243
rect 222742 48179 222794 48185
rect 222070 48163 222122 48169
rect 222070 48105 222122 48111
rect 221302 48015 221354 48021
rect 221302 47957 221354 47963
rect 220534 47941 220586 47947
rect 220534 47883 220586 47889
rect 220150 47793 220202 47799
rect 220150 47735 220202 47741
rect 218710 47497 218762 47503
rect 218710 47439 218762 47445
rect 223138 46689 223166 53650
rect 223330 52355 223358 53650
rect 223316 52346 223372 52355
rect 223316 52281 223372 52290
rect 223522 48835 223550 53650
rect 223714 51763 223742 53650
rect 223700 51754 223756 51763
rect 223700 51689 223756 51698
rect 223906 50093 223934 53650
rect 223894 50087 223946 50093
rect 223894 50029 223946 50035
rect 223510 48829 223562 48835
rect 223510 48771 223562 48777
rect 224098 48243 224126 53650
rect 224086 48237 224138 48243
rect 224086 48179 224138 48185
rect 223126 46683 223178 46689
rect 223126 46625 223178 46631
rect 224290 46319 224318 53650
rect 224640 53636 224702 53664
rect 224674 46467 224702 53636
rect 224962 53636 225024 53664
rect 224662 46461 224714 46467
rect 224662 46403 224714 46409
rect 224962 46393 224990 53636
rect 225172 53602 225228 54402
rect 225346 50019 225374 53650
rect 225540 53602 225596 54402
rect 225730 52313 225758 53650
rect 225908 53602 225964 54402
rect 225718 52307 225770 52313
rect 225718 52249 225770 52255
rect 225334 50013 225386 50019
rect 225334 49955 225386 49961
rect 226114 49797 226142 53650
rect 226276 53602 226332 54402
rect 261922 53941 262046 53960
rect 261910 53935 262046 53941
rect 261962 53932 262046 53935
rect 261910 53877 261962 53883
rect 262018 53867 262046 53932
rect 282166 53935 282218 53941
rect 282166 53877 282218 53883
rect 231766 53861 231818 53867
rect 231766 53803 231818 53809
rect 262006 53861 262058 53867
rect 262006 53803 262058 53809
rect 226102 49791 226154 49797
rect 226102 49733 226154 49739
rect 226498 49649 226526 53650
rect 226594 53636 226848 53664
rect 226978 53636 227232 53664
rect 226594 52387 226622 53636
rect 226582 52381 226634 52387
rect 226582 52323 226634 52329
rect 226978 52165 227006 53636
rect 226966 52159 227018 52165
rect 226966 52101 227018 52107
rect 227554 51943 227582 53650
rect 227542 51937 227594 51943
rect 227542 51879 227594 51885
rect 226486 49643 226538 49649
rect 226486 49585 226538 49591
rect 227938 46615 227966 53650
rect 228322 46763 228350 53650
rect 228706 50759 228734 53650
rect 228802 53636 229056 53664
rect 229186 53636 229440 53664
rect 228802 50833 228830 53636
rect 228790 50827 228842 50833
rect 228790 50769 228842 50775
rect 228694 50753 228746 50759
rect 228694 50695 228746 50701
rect 229186 50685 229214 53636
rect 229174 50679 229226 50685
rect 229174 50621 229226 50627
rect 229762 46911 229790 53650
rect 230146 50907 230174 53650
rect 230134 50901 230186 50907
rect 230134 50843 230186 50849
rect 229750 46905 229802 46911
rect 229750 46847 229802 46853
rect 230530 46837 230558 53650
rect 230914 50981 230942 53650
rect 231010 53636 231264 53664
rect 231394 53636 231648 53664
rect 231778 53645 231806 53803
rect 282178 53701 282206 53877
rect 282178 53673 282398 53701
rect 231766 53639 231818 53645
rect 230902 50975 230954 50981
rect 230902 50917 230954 50923
rect 231010 47207 231038 53636
rect 231394 51129 231422 53636
rect 231766 53581 231818 53587
rect 231382 51123 231434 51129
rect 231382 51065 231434 51071
rect 231970 51055 231998 53650
rect 232354 51203 232382 53650
rect 232342 51197 232394 51203
rect 232342 51139 232394 51145
rect 231958 51049 232010 51055
rect 231958 50991 232010 50997
rect 232738 50167 232766 53650
rect 232726 50161 232778 50167
rect 232726 50103 232778 50109
rect 230998 47201 231050 47207
rect 230998 47143 231050 47149
rect 230518 46831 230570 46837
rect 230518 46773 230570 46779
rect 228310 46757 228362 46763
rect 228310 46699 228362 46705
rect 227926 46609 227978 46615
rect 227926 46551 227978 46557
rect 233122 46541 233150 53650
rect 233314 53636 233472 53664
rect 233602 53636 233856 53664
rect 233314 47059 233342 53636
rect 233602 51499 233630 53636
rect 233590 51493 233642 51499
rect 233590 51435 233642 51441
rect 233302 47053 233354 47059
rect 233302 46995 233354 47001
rect 234178 46985 234206 53650
rect 234562 51425 234590 53650
rect 234550 51419 234602 51425
rect 234550 51361 234602 51367
rect 234946 50241 234974 53650
rect 235330 51277 235358 53650
rect 235426 53636 235680 53664
rect 235810 53636 236064 53664
rect 235318 51271 235370 51277
rect 235318 51213 235370 51219
rect 235426 50315 235454 53636
rect 235810 51351 235838 53636
rect 235798 51345 235850 51351
rect 235798 51287 235850 51293
rect 235414 50309 235466 50315
rect 235414 50251 235466 50257
rect 234934 50235 234986 50241
rect 234934 50177 234986 50183
rect 236386 47133 236414 53650
rect 236770 51023 236798 53650
rect 236756 51014 236812 51023
rect 236756 50949 236812 50958
rect 237154 49723 237182 53650
rect 237538 51319 237566 53650
rect 237634 53636 237888 53664
rect 238018 53636 238272 53664
rect 237524 51310 237580 51319
rect 237524 51245 237580 51254
rect 237634 51171 237662 53636
rect 237620 51162 237676 51171
rect 237620 51097 237676 51106
rect 237142 49717 237194 49723
rect 237142 49659 237194 49665
rect 238018 47429 238046 53636
rect 238006 47423 238058 47429
rect 238006 47365 238058 47371
rect 238594 47355 238622 53650
rect 238582 47349 238634 47355
rect 238582 47291 238634 47297
rect 238978 47281 239006 53650
rect 239362 48613 239390 53650
rect 239350 48607 239402 48613
rect 239350 48549 239402 48555
rect 239746 48465 239774 53650
rect 239842 53636 240096 53664
rect 240226 53636 240480 53664
rect 239734 48459 239786 48465
rect 239734 48401 239786 48407
rect 239842 48391 239870 53636
rect 240226 48539 240254 53636
rect 240214 48533 240266 48539
rect 240214 48475 240266 48481
rect 239830 48385 239882 48391
rect 239830 48327 239882 48333
rect 238966 47275 239018 47281
rect 238966 47217 239018 47223
rect 236374 47127 236426 47133
rect 236374 47069 236426 47075
rect 234166 46979 234218 46985
rect 234166 46921 234218 46927
rect 233110 46535 233162 46541
rect 233110 46477 233162 46483
rect 224950 46387 225002 46393
rect 224950 46329 225002 46335
rect 224278 46313 224330 46319
rect 224278 46255 224330 46261
rect 240802 46245 240830 53650
rect 241186 49945 241214 53650
rect 241174 49939 241226 49945
rect 241174 49881 241226 49887
rect 241570 48317 241598 53650
rect 241954 48359 241982 53650
rect 242050 53636 242304 53664
rect 242434 53636 242688 53664
rect 241940 48350 241996 48359
rect 241558 48311 241610 48317
rect 241940 48285 241996 48294
rect 241558 48253 241610 48259
rect 242050 48211 242078 53636
rect 242434 48655 242462 53636
rect 243010 48803 243038 53650
rect 242996 48794 243052 48803
rect 242996 48729 243052 48738
rect 242420 48646 242476 48655
rect 242420 48581 242476 48590
rect 243394 48507 243422 53650
rect 243778 51467 243806 53650
rect 243764 51458 243820 51467
rect 243764 51393 243820 51402
rect 244162 49871 244190 53650
rect 251926 53195 251978 53201
rect 251926 53137 251978 53143
rect 251938 52979 251966 53137
rect 251926 52973 251978 52979
rect 251926 52915 251978 52921
rect 244150 49865 244202 49871
rect 244150 49807 244202 49813
rect 243380 48498 243436 48507
rect 243380 48433 243436 48442
rect 242036 48202 242092 48211
rect 242036 48137 242092 48146
rect 240790 46239 240842 46245
rect 240790 46181 240842 46187
rect 215444 44946 215500 44955
rect 215444 44881 215500 44890
rect 215062 43279 215114 43285
rect 215062 43221 215114 43227
rect 214294 42169 214346 42175
rect 282370 42143 282398 53673
rect 351286 53565 351338 53571
rect 351286 53507 351338 53513
rect 315670 53269 315722 53275
rect 315670 53211 315722 53217
rect 315682 53053 315710 53211
rect 315670 53047 315722 53053
rect 315670 52989 315722 52995
rect 351298 49076 351326 53507
rect 384406 53491 384458 53497
rect 384406 53433 384458 53439
rect 368566 53269 368618 53275
rect 368618 53217 368702 53220
rect 368566 53211 368702 53217
rect 368578 53201 368702 53211
rect 368578 53195 368714 53201
rect 368578 53192 368662 53195
rect 368662 53137 368714 53143
rect 351298 49048 351422 49076
rect 297238 45055 297290 45061
rect 297238 44997 297290 45003
rect 297250 43179 297278 44997
rect 310102 44685 310154 44691
rect 310102 44627 310154 44633
rect 297236 43170 297292 43179
rect 297236 43105 297292 43114
rect 302420 43170 302476 43179
rect 302420 43105 302476 43114
rect 214294 42111 214346 42117
rect 282356 42134 282412 42143
rect 302434 42120 302462 43105
rect 306740 42134 306796 42143
rect 302434 42092 302688 42120
rect 282356 42069 282412 42078
rect 306796 42092 307008 42120
rect 310114 42106 310142 44627
rect 351394 43179 351422 49048
rect 384418 45431 384446 53433
rect 467446 53417 467498 53423
rect 408994 53340 409118 53368
rect 467446 53359 467498 53365
rect 469366 53417 469418 53423
rect 469366 53359 469418 53365
rect 501046 53417 501098 53423
rect 501046 53359 501098 53365
rect 408994 53275 409022 53340
rect 388822 53269 388874 53275
rect 388738 53217 388822 53220
rect 388738 53211 388874 53217
rect 408982 53269 409034 53275
rect 408982 53211 409034 53217
rect 388738 53201 388862 53211
rect 388726 53195 388862 53201
rect 388778 53192 388862 53195
rect 388726 53137 388778 53143
rect 409090 53053 409118 53340
rect 409078 53047 409130 53053
rect 409078 52989 409130 52995
rect 467458 49099 467486 53359
rect 469378 53201 469406 53359
rect 501058 53201 501086 53359
rect 501142 53343 501194 53349
rect 501142 53285 501194 53291
rect 469366 53195 469418 53201
rect 469366 53137 469418 53143
rect 501046 53195 501098 53201
rect 501046 53137 501098 53143
rect 467444 49090 467500 49099
rect 467444 49025 467500 49034
rect 501154 48909 501182 53285
rect 509686 53195 509738 53201
rect 509686 53137 509738 53143
rect 509698 49057 509726 53137
rect 639682 51721 639710 233456
rect 649762 233243 649790 748811
rect 649858 707551 649886 989237
rect 650050 754467 650078 994449
rect 650326 993513 650378 993519
rect 650326 993455 650378 993461
rect 650230 986705 650282 986711
rect 650230 986647 650282 986653
rect 650134 986631 650186 986637
rect 650134 986573 650186 986579
rect 650146 895215 650174 986573
rect 650132 895206 650188 895215
rect 650132 895141 650188 895150
rect 650242 801383 650270 986647
rect 650228 801374 650284 801383
rect 650228 801309 650284 801318
rect 650036 754458 650092 754467
rect 650036 754393 650092 754402
rect 649844 707542 649900 707551
rect 649844 707477 649900 707486
rect 649846 702767 649898 702773
rect 649846 702709 649898 702715
rect 649858 236351 649886 702709
rect 650338 660635 650366 993455
rect 658006 986557 658058 986563
rect 658006 986499 658058 986505
rect 655124 976754 655180 976763
rect 655124 976689 655180 976698
rect 655138 939129 655166 976689
rect 655220 965062 655276 965071
rect 655220 964997 655276 965006
rect 655234 939277 655262 964997
rect 655316 953370 655372 953379
rect 655316 953305 655372 953314
rect 655330 939425 655358 953305
rect 655318 939419 655370 939425
rect 655318 939361 655370 939367
rect 655222 939271 655274 939277
rect 655222 939213 655274 939219
rect 655126 939123 655178 939129
rect 655126 939065 655178 939071
rect 658018 936169 658046 986499
rect 658102 986483 658154 986489
rect 658102 986425 658154 986431
rect 658114 939573 658142 986425
rect 660886 986409 660938 986415
rect 660886 986351 660938 986357
rect 658102 939567 658154 939573
rect 658102 939509 658154 939515
rect 660898 938019 660926 986351
rect 674518 983745 674570 983751
rect 674518 983687 674570 983693
rect 674326 983671 674378 983677
rect 674326 983613 674378 983619
rect 674338 967587 674366 983613
rect 674324 967578 674380 967587
rect 674324 967513 674380 967522
rect 674530 967439 674558 983687
rect 674996 967578 675052 967587
rect 674996 967513 675052 967522
rect 674516 967430 674572 967439
rect 674516 967365 674572 967374
rect 675010 960573 675038 967513
rect 675202 966722 675408 966750
rect 675202 964923 675230 966722
rect 675778 965663 675806 966070
rect 675764 965654 675820 965663
rect 675764 965589 675820 965598
rect 675298 965421 675408 965449
rect 675298 965071 675326 965421
rect 675284 965062 675340 965071
rect 675284 964997 675340 965006
rect 675188 964914 675244 964923
rect 675188 964849 675244 964858
rect 675106 963581 675408 963609
rect 675106 962851 675134 963581
rect 675202 963022 675408 963050
rect 675092 962842 675148 962851
rect 675092 962777 675148 962786
rect 675202 962555 675230 963022
rect 675188 962546 675244 962555
rect 675188 962481 675244 962490
rect 675778 962259 675806 962399
rect 675764 962250 675820 962259
rect 675764 962185 675820 962194
rect 675394 961519 675422 961778
rect 675380 961510 675436 961519
rect 675380 961445 675436 961454
rect 675682 961075 675710 961186
rect 675668 961066 675724 961075
rect 675668 961001 675724 961010
rect 675010 960559 675792 960573
rect 675010 960545 675806 960559
rect 675778 960187 675806 960545
rect 675764 960178 675820 960187
rect 675764 960113 675820 960122
rect 675490 959151 675518 959262
rect 675476 959142 675532 959151
rect 675476 959077 675532 959086
rect 675394 958443 675422 958744
rect 675094 958437 675146 958443
rect 675094 958379 675146 958385
rect 675382 958437 675434 958443
rect 675382 958379 675434 958385
rect 669526 954737 669578 954743
rect 669526 954679 669578 954685
rect 660886 938013 660938 938019
rect 660886 937955 660938 937961
rect 658006 936163 658058 936169
rect 658006 936105 658058 936111
rect 654452 929838 654508 929847
rect 654452 929773 654508 929782
rect 654466 927511 654494 929773
rect 654454 927505 654506 927511
rect 654454 927447 654506 927453
rect 666742 927505 666794 927511
rect 666742 927447 666794 927453
rect 653972 918146 654028 918155
rect 653972 918081 654028 918090
rect 653986 915893 654014 918081
rect 653974 915887 654026 915893
rect 653974 915829 654026 915835
rect 660982 915887 661034 915893
rect 660982 915829 661034 915835
rect 654452 906454 654508 906463
rect 654452 906389 654508 906398
rect 654466 904423 654494 906389
rect 654454 904417 654506 904423
rect 654454 904359 654506 904365
rect 653972 882922 654028 882931
rect 653972 882857 654028 882866
rect 653986 881335 654014 882857
rect 653974 881329 654026 881335
rect 653974 881271 654026 881277
rect 660886 881329 660938 881335
rect 660886 881271 660938 881277
rect 654452 871230 654508 871239
rect 654452 871165 654508 871174
rect 654466 869865 654494 871165
rect 654454 869859 654506 869865
rect 654454 869801 654506 869807
rect 654164 859538 654220 859547
rect 654164 859473 654220 859482
rect 654178 858321 654206 859473
rect 654166 858315 654218 858321
rect 654166 858257 654218 858263
rect 653972 836006 654028 836015
rect 653972 835941 654028 835950
rect 653986 835233 654014 835941
rect 653974 835227 654026 835233
rect 653974 835169 654026 835175
rect 653972 824314 654028 824323
rect 653972 824249 654028 824258
rect 653986 823763 654014 824249
rect 653974 823757 654026 823763
rect 653974 823699 654026 823705
rect 654452 812622 654508 812631
rect 654452 812557 654508 812566
rect 654466 812219 654494 812557
rect 654454 812213 654506 812219
rect 654454 812155 654506 812161
rect 654068 789090 654124 789099
rect 654068 789025 654124 789034
rect 654082 786319 654110 789025
rect 654070 786313 654122 786319
rect 654070 786255 654122 786261
rect 654068 777398 654124 777407
rect 654068 777333 654124 777342
rect 654082 774775 654110 777333
rect 654070 774769 654122 774775
rect 654070 774711 654122 774717
rect 653972 765558 654028 765567
rect 653972 765493 654028 765502
rect 653986 763305 654014 765493
rect 653974 763299 654026 763305
rect 653974 763241 654026 763247
rect 653972 742174 654028 742183
rect 653972 742109 654028 742118
rect 653986 740217 654014 742109
rect 653974 740211 654026 740217
rect 653974 740153 654026 740159
rect 655220 730482 655276 730491
rect 655220 730417 655276 730426
rect 654260 718642 654316 718651
rect 654260 718577 654316 718586
rect 654274 717203 654302 718577
rect 654262 717197 654314 717203
rect 654262 717139 654314 717145
rect 654452 695258 654508 695267
rect 654452 695193 654508 695202
rect 654466 694115 654494 695193
rect 654454 694109 654506 694115
rect 654454 694051 654506 694057
rect 655124 683566 655180 683575
rect 655124 683501 655180 683510
rect 654452 671726 654508 671735
rect 654452 671661 654508 671670
rect 654466 671101 654494 671661
rect 654454 671095 654506 671101
rect 654454 671037 654506 671043
rect 650324 660626 650380 660635
rect 650324 660561 650380 660570
rect 649942 659551 649994 659557
rect 649942 659493 649994 659499
rect 649846 236345 649898 236351
rect 649846 236287 649898 236293
rect 645718 233237 645770 233243
rect 645718 233179 645770 233185
rect 649750 233237 649802 233243
rect 649750 233179 649802 233185
rect 645142 233089 645194 233095
rect 645142 233031 645194 233037
rect 645154 231139 645182 233031
rect 645334 233015 645386 233021
rect 645334 232957 645386 232963
rect 645238 232941 645290 232947
rect 645238 232883 645290 232889
rect 645250 231583 645278 232883
rect 645236 231574 645292 231583
rect 645236 231509 645292 231518
rect 645140 231130 645196 231139
rect 645140 231065 645196 231074
rect 645154 141113 645182 231065
rect 645250 141113 645278 231509
rect 645346 230695 645374 232957
rect 645730 232027 645758 233179
rect 649954 233169 649982 659493
rect 654260 648342 654316 648351
rect 654260 648277 654316 648286
rect 654274 648087 654302 648277
rect 654262 648081 654314 648087
rect 654262 648023 654314 648029
rect 654068 624810 654124 624819
rect 654068 624745 654124 624754
rect 654082 622187 654110 624745
rect 654070 622181 654122 622187
rect 654070 622123 654122 622129
rect 650038 613523 650090 613529
rect 650038 613465 650090 613471
rect 650050 236203 650078 613465
rect 654358 613449 654410 613455
rect 654358 613391 654410 613397
rect 654370 613127 654398 613391
rect 654356 613118 654412 613127
rect 654356 613053 654412 613062
rect 654452 601426 654508 601435
rect 654452 601361 654508 601370
rect 654466 599099 654494 601361
rect 654454 599093 654506 599099
rect 654454 599035 654506 599041
rect 654452 589586 654508 589595
rect 654452 589521 654508 589530
rect 654466 587555 654494 589521
rect 654454 587549 654506 587555
rect 654454 587491 654506 587497
rect 654452 577894 654508 577903
rect 654452 577829 654508 577838
rect 654466 576085 654494 577829
rect 654454 576079 654506 576085
rect 654454 576021 654506 576027
rect 650134 567421 650186 567427
rect 650134 567363 650186 567369
rect 650038 236197 650090 236203
rect 650038 236139 650090 236145
rect 645814 233163 645866 233169
rect 645814 233105 645866 233111
rect 649942 233163 649994 233169
rect 649942 233105 649994 233111
rect 645826 232767 645854 233105
rect 650146 233021 650174 567363
rect 654454 567347 654506 567353
rect 654454 567289 654506 567295
rect 654466 566211 654494 567289
rect 654452 566202 654508 566211
rect 654452 566137 654508 566146
rect 654452 554510 654508 554519
rect 654452 554445 654508 554454
rect 654466 552997 654494 554445
rect 654454 552991 654506 552997
rect 654454 552933 654506 552939
rect 654452 542670 654508 542679
rect 654452 542605 654508 542614
rect 654466 541527 654494 542605
rect 654454 541521 654506 541527
rect 654454 541463 654506 541469
rect 655138 535829 655166 683501
rect 655234 582005 655262 730417
rect 660898 717351 660926 881271
rect 660994 762935 661022 915829
rect 663958 904417 664010 904423
rect 663958 904359 664010 904365
rect 663766 869859 663818 869865
rect 663766 869801 663818 869807
rect 661078 858315 661130 858321
rect 661078 858257 661130 858263
rect 660982 762929 661034 762935
rect 660982 762871 661034 762877
rect 660982 737325 661034 737331
rect 660982 737267 661034 737273
rect 660886 717345 660938 717351
rect 660886 717287 660938 717293
rect 655316 636650 655372 636659
rect 655316 636585 655372 636594
rect 655222 581999 655274 582005
rect 655222 581941 655274 581947
rect 655126 535823 655178 535829
rect 655126 535765 655178 535771
rect 654068 530978 654124 530987
rect 654068 530913 654124 530922
rect 654082 529983 654110 530913
rect 654070 529977 654122 529983
rect 654070 529919 654122 529925
rect 650230 524353 650282 524359
rect 650230 524295 650282 524301
rect 650242 236499 650270 524295
rect 654454 519321 654506 519327
rect 654452 519286 654454 519295
rect 654506 519286 654508 519295
rect 654452 519221 654508 519230
rect 654452 507446 654508 507455
rect 654452 507381 654508 507390
rect 654466 506969 654494 507381
rect 654454 506963 654506 506969
rect 654454 506905 654506 506911
rect 654356 495754 654412 495763
rect 654356 495689 654412 495698
rect 654370 495425 654398 495689
rect 654358 495419 654410 495425
rect 654358 495361 654410 495367
rect 655330 492539 655358 636585
rect 660886 555877 660938 555883
rect 660886 555819 660938 555825
rect 655318 492533 655370 492539
rect 655318 492475 655370 492481
rect 654260 484062 654316 484071
rect 654260 483997 654316 484006
rect 654274 483881 654302 483997
rect 654262 483875 654314 483881
rect 654262 483817 654314 483823
rect 650326 479509 650378 479515
rect 650326 479451 650378 479457
rect 650230 236493 650282 236499
rect 650230 236435 650282 236441
rect 650338 236425 650366 479451
rect 654454 472257 654506 472263
rect 654452 472222 654454 472231
rect 654506 472222 654508 472231
rect 654452 472157 654508 472166
rect 654452 460530 654508 460539
rect 654452 460465 654508 460474
rect 654466 457981 654494 460465
rect 654454 457975 654506 457981
rect 654454 457917 654506 457923
rect 654356 448838 654412 448847
rect 654356 448773 654412 448782
rect 654370 446437 654398 448773
rect 654358 446431 654410 446437
rect 654358 446373 654410 446379
rect 654452 436998 654508 437007
rect 654452 436933 654508 436942
rect 654466 434967 654494 436933
rect 654454 434961 654506 434967
rect 654454 434903 654506 434909
rect 654454 426229 654506 426235
rect 654454 426171 654506 426177
rect 654466 425463 654494 426171
rect 654452 425454 654508 425463
rect 654452 425389 654508 425398
rect 653876 413614 653932 413623
rect 653876 413549 653932 413558
rect 653890 411879 653918 413549
rect 653878 411873 653930 411879
rect 653878 411815 653930 411821
rect 654452 401774 654508 401783
rect 654452 401709 654508 401718
rect 654466 400409 654494 401709
rect 654454 400403 654506 400409
rect 654454 400345 654506 400351
rect 650422 391819 650474 391825
rect 650422 391761 650474 391767
rect 650326 236419 650378 236425
rect 650326 236361 650378 236367
rect 650434 233095 650462 391761
rect 654452 390082 654508 390091
rect 654452 390017 654508 390026
rect 654466 388865 654494 390017
rect 654454 388859 654506 388865
rect 654454 388801 654506 388807
rect 654454 380127 654506 380133
rect 654454 380069 654506 380075
rect 654466 378547 654494 380069
rect 654452 378538 654508 378547
rect 654452 378473 654508 378482
rect 654452 366550 654508 366559
rect 654452 366485 654508 366494
rect 654466 365851 654494 366485
rect 654454 365845 654506 365851
rect 654454 365787 654506 365793
rect 655220 354858 655276 354867
rect 655220 354793 655276 354802
rect 650518 345643 650570 345649
rect 650518 345585 650570 345591
rect 650530 236573 650558 345585
rect 654452 343166 654508 343175
rect 654452 343101 654508 343110
rect 654466 342763 654494 343101
rect 654454 342757 654506 342763
rect 654454 342699 654506 342705
rect 654454 332323 654506 332329
rect 654454 332265 654506 332271
rect 654466 331631 654494 332265
rect 654452 331622 654508 331631
rect 654452 331557 654508 331566
rect 655124 319782 655180 319791
rect 655124 319717 655180 319726
rect 650614 302649 650666 302655
rect 650614 302591 650666 302597
rect 650518 236567 650570 236573
rect 650518 236509 650570 236515
rect 650422 233089 650474 233095
rect 650422 233031 650474 233037
rect 650134 233015 650186 233021
rect 650134 232957 650186 232963
rect 650626 232947 650654 302591
rect 654548 296250 654604 296259
rect 654548 296185 654604 296194
rect 654562 293849 654590 296185
rect 654550 293843 654602 293849
rect 654550 293785 654602 293791
rect 654070 284815 654122 284821
rect 654070 284757 654122 284763
rect 654082 284715 654110 284757
rect 654068 284706 654124 284715
rect 654068 284641 654124 284650
rect 650614 232941 650666 232947
rect 650614 232883 650666 232889
rect 645812 232758 645868 232767
rect 645812 232693 645868 232702
rect 645716 232018 645772 232027
rect 645716 231953 645772 231962
rect 645332 230686 645388 230695
rect 645332 230621 645388 230630
rect 645346 141155 645374 230621
rect 645430 216069 645482 216075
rect 645430 216011 645482 216017
rect 645442 207343 645470 216011
rect 645620 210410 645676 210419
rect 645620 210345 645676 210354
rect 645430 207337 645482 207343
rect 645430 207279 645482 207285
rect 645430 141255 645482 141261
rect 645430 141197 645482 141203
rect 645332 141146 645388 141155
rect 645142 141107 645194 141113
rect 645142 141049 645194 141055
rect 645238 141107 645290 141113
rect 645442 141113 645470 141197
rect 645332 141081 645388 141090
rect 645430 141107 645482 141113
rect 645238 141049 645290 141055
rect 645430 141049 645482 141055
rect 645332 140850 645388 140859
rect 645238 140811 645290 140817
rect 645332 140785 645388 140794
rect 645238 140753 645290 140759
rect 645142 140589 645194 140595
rect 645142 140531 645194 140537
rect 640726 76283 640778 76289
rect 640726 76225 640778 76231
rect 639670 51715 639722 51721
rect 639670 51657 639722 51663
rect 509686 49051 509738 49057
rect 509686 48993 509738 48999
rect 525910 49051 525962 49057
rect 525910 48993 525962 48999
rect 501142 48903 501194 48909
rect 501142 48845 501194 48851
rect 507094 48903 507146 48909
rect 507094 48845 507146 48851
rect 465814 46091 465866 46097
rect 465814 46033 465866 46039
rect 384406 45425 384458 45431
rect 384406 45367 384458 45373
rect 388822 45425 388874 45431
rect 388822 45367 388874 45373
rect 361750 44981 361802 44987
rect 361750 44923 361802 44929
rect 351380 43170 351436 43179
rect 351380 43105 351436 43114
rect 357140 43170 357196 43179
rect 357140 43105 357196 43114
rect 357154 42120 357182 43105
rect 357154 42092 357456 42120
rect 361762 42106 361790 44923
rect 362806 44833 362858 44839
rect 362806 44775 362858 44781
rect 362818 42143 362846 44775
rect 362804 42134 362860 42143
rect 306740 42069 306796 42078
rect 362804 42069 362860 42078
rect 364628 42134 364684 42143
rect 364684 42092 364944 42120
rect 364628 42069 364684 42078
rect 374324 41246 374380 41255
rect 374324 41181 374380 41190
rect 334100 40950 334156 40959
rect 334100 40885 334102 40894
rect 334154 40885 334156 40894
rect 344180 40950 344236 40959
rect 344180 40885 344182 40894
rect 334102 40853 334154 40859
rect 344234 40885 344236 40894
rect 344182 40853 344234 40859
rect 374338 40811 374366 41181
rect 374324 40802 374380 40811
rect 374324 40737 374380 40746
rect 211028 40654 211084 40663
rect 211028 40589 211084 40598
rect 388834 40325 388862 45367
rect 411092 45242 411148 45251
rect 411092 45177 411148 45186
rect 411106 44488 411134 45177
rect 455734 44907 455786 44913
rect 455734 44849 455786 44855
rect 416564 44798 416620 44807
rect 416564 44733 416620 44742
rect 411088 44460 411134 44488
rect 411088 44178 411116 44460
rect 405526 42317 405578 42323
rect 405526 42259 405578 42265
rect 405538 42106 405566 42259
rect 416578 42106 416606 44733
rect 455746 43179 455774 44849
rect 465826 44164 465854 46033
rect 507106 43359 507134 48845
rect 507094 43353 507146 43359
rect 521588 43318 521644 43327
rect 507094 43295 507146 43301
rect 518722 43285 518834 43304
rect 518710 43279 518834 43285
rect 518762 43276 518834 43279
rect 521588 43253 521644 43262
rect 518710 43221 518762 43227
rect 520342 43205 520394 43211
rect 455732 43170 455788 43179
rect 455732 43105 455788 43114
rect 463988 43170 464044 43179
rect 520342 43147 520394 43153
rect 463988 43105 464044 43114
rect 460054 42243 460106 42249
rect 460054 42185 460106 42191
rect 460066 42120 460094 42185
rect 460066 42092 460368 42120
rect 464002 42106 464030 43105
rect 514870 42169 514922 42175
rect 471092 42134 471148 42143
rect 471148 42092 471408 42120
rect 520354 42120 520382 43147
rect 521602 42120 521630 43253
rect 525922 42120 525950 48993
rect 640738 47577 640766 76225
rect 645154 48687 645182 140531
rect 645250 48761 645278 140753
rect 645238 48755 645290 48761
rect 645238 48697 645290 48703
rect 645142 48681 645194 48687
rect 645142 48623 645194 48629
rect 645346 48243 645374 140785
rect 645526 126677 645578 126683
rect 645526 126619 645578 126625
rect 645538 106555 645566 126619
rect 645526 106549 645578 106555
rect 645526 106491 645578 106497
rect 645430 104551 645482 104557
rect 645430 104493 645482 104499
rect 645442 104303 645470 104493
rect 645428 104294 645484 104303
rect 645428 104229 645484 104238
rect 645428 87718 645484 87727
rect 645428 87653 645484 87662
rect 645442 87093 645470 87653
rect 645430 87087 645482 87093
rect 645430 87029 645482 87035
rect 645430 86939 645482 86945
rect 645430 86881 645482 86887
rect 645442 86427 645470 86881
rect 645430 86421 645482 86427
rect 645430 86363 645482 86369
rect 645430 85237 645482 85243
rect 645430 85179 645482 85185
rect 645442 85063 645470 85179
rect 645428 85054 645484 85063
rect 645428 84989 645484 84998
rect 645430 83461 645482 83467
rect 645430 83403 645482 83409
rect 645442 83287 645470 83403
rect 645428 83278 645484 83287
rect 645428 83213 645484 83222
rect 645428 82538 645484 82547
rect 645428 82473 645484 82482
rect 645442 81913 645470 82473
rect 645430 81907 645482 81913
rect 645430 81849 645482 81855
rect 645428 81354 645484 81363
rect 645428 81289 645430 81298
rect 645482 81289 645484 81298
rect 645430 81257 645482 81263
rect 645430 80205 645482 80211
rect 645430 80147 645482 80153
rect 645442 80031 645470 80147
rect 645428 80022 645484 80031
rect 645428 79957 645484 79966
rect 645430 78947 645482 78953
rect 645430 78889 645482 78895
rect 645442 78699 645470 78889
rect 645428 78690 645484 78699
rect 645428 78625 645484 78634
rect 645430 77689 645482 77695
rect 645428 77654 645430 77663
rect 645482 77654 645484 77663
rect 645428 77589 645484 77598
rect 645430 77319 645482 77325
rect 645430 77261 645482 77267
rect 645442 77071 645470 77261
rect 645428 77062 645484 77071
rect 645428 76997 645484 77006
rect 645430 76949 645482 76955
rect 645430 76891 645482 76897
rect 645442 76775 645470 76891
rect 645428 76766 645484 76775
rect 645428 76701 645484 76710
rect 645430 75543 645482 75549
rect 645430 75485 645482 75491
rect 645442 75443 645470 75485
rect 645428 75434 645484 75443
rect 645428 75369 645484 75378
rect 645428 74398 645484 74407
rect 645428 74333 645484 74342
rect 645442 73033 645470 74333
rect 645430 73027 645482 73033
rect 645430 72969 645482 72975
rect 645428 72918 645484 72927
rect 645428 72853 645484 72862
rect 645442 72145 645470 72853
rect 645430 72139 645482 72145
rect 645430 72081 645482 72087
rect 645526 66293 645578 66299
rect 645526 66235 645578 66241
rect 645538 51869 645566 66235
rect 645526 51863 645578 51869
rect 645526 51805 645578 51811
rect 645634 48983 645662 210345
rect 645730 51795 645758 231953
rect 645826 216075 645854 232693
rect 645814 216069 645866 216075
rect 645814 216011 645866 216017
rect 647924 210410 647980 210419
rect 647924 210345 647980 210354
rect 647938 210303 647966 210345
rect 647926 210297 647978 210303
rect 647926 210239 647978 210245
rect 645814 207337 645866 207343
rect 645814 207279 645866 207285
rect 645826 141261 645854 207279
rect 646870 167451 646922 167457
rect 646870 167393 646922 167399
rect 646294 167229 646346 167235
rect 646294 167171 646346 167177
rect 646306 166315 646334 167171
rect 646292 166306 646348 166315
rect 646292 166241 646348 166250
rect 646882 166019 646910 167393
rect 647926 167155 647978 167161
rect 647926 167097 647978 167103
rect 647938 167055 647966 167097
rect 647924 167046 647980 167055
rect 647924 166981 647980 166990
rect 646868 166010 646924 166019
rect 646868 165945 646924 165954
rect 645814 141255 645866 141261
rect 645814 141197 645866 141203
rect 645814 141107 645866 141113
rect 645814 141049 645866 141055
rect 645826 126683 645854 141049
rect 655138 132677 655166 319717
rect 655234 178705 655262 354793
rect 655316 307942 655372 307951
rect 655316 307877 655372 307886
rect 655222 178699 655274 178705
rect 655222 178641 655274 178647
rect 655330 132825 655358 307877
rect 660898 284821 660926 555819
rect 660994 472263 661022 737267
rect 661090 716907 661118 858257
rect 661174 763299 661226 763305
rect 661174 763241 661226 763247
rect 661078 716901 661130 716907
rect 661078 716843 661130 716849
rect 661078 671095 661130 671101
rect 661078 671037 661130 671043
rect 661090 536643 661118 671037
rect 661186 626923 661214 763241
rect 663778 717943 663806 869801
rect 663862 780541 663914 780547
rect 663862 780483 663914 780489
rect 663766 717937 663818 717943
rect 663766 717879 663818 717885
rect 661174 626917 661226 626923
rect 661174 626859 661226 626865
rect 663766 601979 663818 601985
rect 663766 601921 663818 601927
rect 661078 536637 661130 536643
rect 661078 536579 661130 536585
rect 661174 495419 661226 495425
rect 661174 495361 661226 495367
rect 660982 472257 661034 472263
rect 660982 472199 661034 472205
rect 660982 457975 661034 457981
rect 660982 457917 661034 457923
rect 660886 284815 660938 284821
rect 660886 284757 660938 284763
rect 660994 269799 661022 457917
rect 661078 365845 661130 365851
rect 661078 365787 661130 365793
rect 660982 269793 661034 269799
rect 660982 269735 661034 269741
rect 661090 179371 661118 365787
rect 661186 315087 661214 495361
rect 663778 332329 663806 601921
rect 663874 519327 663902 780483
rect 663970 762047 663998 904359
rect 666646 864087 666698 864093
rect 666646 864029 666698 864035
rect 664054 812213 664106 812219
rect 664054 812155 664106 812161
rect 663958 762041 664010 762047
rect 663958 761983 664010 761989
rect 663958 740211 664010 740217
rect 663958 740153 664010 740159
rect 663970 582079 663998 740153
rect 664066 671619 664094 812155
rect 664054 671613 664106 671619
rect 664054 671555 664106 671561
rect 664054 648081 664106 648087
rect 664054 648023 664106 648029
rect 663958 582073 664010 582079
rect 663958 582015 664010 582021
rect 663862 519321 663914 519327
rect 663862 519263 663914 519269
rect 663862 506963 663914 506969
rect 663862 506905 663914 506911
rect 663766 332323 663818 332329
rect 663766 332265 663818 332271
rect 661174 315081 661226 315087
rect 661174 315023 661226 315029
rect 663874 314791 663902 506905
rect 664066 492983 664094 648023
rect 666658 567353 666686 864029
rect 666754 762343 666782 927447
rect 666838 835227 666890 835233
rect 666838 835169 666890 835175
rect 666742 762337 666794 762343
rect 666742 762279 666794 762285
rect 666850 672211 666878 835169
rect 666934 717197 666986 717203
rect 666934 717139 666986 717145
rect 666838 672205 666890 672211
rect 666838 672147 666890 672153
rect 666742 645195 666794 645201
rect 666742 645137 666794 645143
rect 666646 567347 666698 567353
rect 666646 567289 666698 567295
rect 666646 552991 666698 552997
rect 666646 552933 666698 552939
rect 664054 492977 664106 492983
rect 664054 492919 664106 492925
rect 663958 434961 664010 434967
rect 663958 434903 664010 434909
rect 663862 314785 663914 314791
rect 663862 314727 663914 314733
rect 663766 293843 663818 293849
rect 663766 293785 663818 293791
rect 661078 179365 661130 179371
rect 661078 179307 661130 179313
rect 663778 133639 663806 293785
rect 663970 269207 663998 434903
rect 666658 359783 666686 552933
rect 666754 380133 666782 645137
rect 666838 587549 666890 587555
rect 666838 587491 666890 587497
rect 666850 405515 666878 587491
rect 666946 581635 666974 717139
rect 669538 613455 669566 954679
rect 674134 953923 674186 953929
rect 674134 953865 674186 953871
rect 674038 952073 674090 952079
rect 674038 952015 674090 952021
rect 673844 939162 673900 939171
rect 673844 939097 673900 939106
rect 673366 866973 673418 866979
rect 673366 866915 673418 866921
rect 669814 823757 669866 823763
rect 669814 823699 669866 823705
rect 669718 786313 669770 786319
rect 669718 786255 669770 786261
rect 669622 686265 669674 686271
rect 669622 686207 669674 686213
rect 669526 613449 669578 613455
rect 669526 613391 669578 613397
rect 669526 599093 669578 599099
rect 669526 599035 669578 599041
rect 666934 581629 666986 581635
rect 666934 581571 666986 581577
rect 666934 483875 666986 483881
rect 666934 483817 666986 483823
rect 666838 405509 666890 405515
rect 666838 405451 666890 405457
rect 666838 400403 666890 400409
rect 666838 400345 666890 400351
rect 666742 380127 666794 380133
rect 666742 380069 666794 380075
rect 666646 359777 666698 359783
rect 666646 359719 666698 359725
rect 666646 342757 666698 342763
rect 666646 342699 666698 342705
rect 663958 269201 664010 269207
rect 663958 269143 664010 269149
rect 666658 178853 666686 342699
rect 666850 225103 666878 400345
rect 666946 314051 666974 483817
rect 669538 404775 669566 599035
rect 669634 426235 669662 686207
rect 669730 627367 669758 786255
rect 669826 672729 669854 823699
rect 672502 783501 672554 783507
rect 672502 783443 672554 783449
rect 672406 774769 672458 774775
rect 672406 774711 672458 774717
rect 672310 760487 672362 760493
rect 672310 760429 672362 760435
rect 672322 716315 672350 760429
rect 672310 716309 672362 716315
rect 672310 716251 672362 716257
rect 669814 672723 669866 672729
rect 669814 672665 669866 672671
rect 671734 648303 671786 648309
rect 671734 648245 671786 648251
rect 669718 627361 669770 627367
rect 669718 627303 669770 627309
rect 670966 625215 671018 625221
rect 670966 625157 671018 625163
rect 670978 580895 671006 625157
rect 670966 580889 671018 580895
rect 670966 580831 671018 580837
rect 669718 576079 669770 576085
rect 669718 576021 669770 576027
rect 669622 426229 669674 426235
rect 669622 426171 669674 426177
rect 669622 411873 669674 411879
rect 669622 411815 669674 411821
rect 669526 404769 669578 404775
rect 669526 404711 669578 404717
rect 669526 388859 669578 388865
rect 669526 388801 669578 388807
rect 666934 314045 666986 314051
rect 666934 313987 666986 313993
rect 666838 225097 666890 225103
rect 666838 225039 666890 225045
rect 669538 224067 669566 388801
rect 669634 224363 669662 411815
rect 669730 404479 669758 576021
rect 671746 574531 671774 648245
rect 672310 648081 672362 648087
rect 672310 648023 672362 648029
rect 672214 644603 672266 644609
rect 672214 644545 672266 644551
rect 671926 622255 671978 622261
rect 671926 622197 671978 622203
rect 671830 599093 671882 599099
rect 671830 599035 671882 599041
rect 671734 574525 671786 574531
rect 671734 574467 671786 574473
rect 671842 528651 671870 599035
rect 671938 588813 671966 622197
rect 672118 604125 672170 604131
rect 672118 604067 672170 604073
rect 672022 603311 672074 603317
rect 672022 603253 672074 603259
rect 671926 588807 671978 588813
rect 671926 588749 671978 588755
rect 671926 580075 671978 580081
rect 671926 580017 671978 580023
rect 671938 536791 671966 580017
rect 671926 536785 671978 536791
rect 671926 536727 671978 536733
rect 672034 529539 672062 603253
rect 672130 529909 672158 604067
rect 672226 573125 672254 644545
rect 672214 573119 672266 573125
rect 672214 573061 672266 573067
rect 672322 572903 672350 648023
rect 672418 627811 672446 774711
rect 672514 709803 672542 783443
rect 672982 783131 673034 783137
rect 672982 783073 673034 783079
rect 672886 779357 672938 779363
rect 672886 779299 672938 779305
rect 672598 777655 672650 777661
rect 672598 777597 672650 777603
rect 672502 709797 672554 709803
rect 672502 709739 672554 709745
rect 672610 709211 672638 777597
rect 672790 738139 672842 738145
rect 672790 738081 672842 738087
rect 672694 737917 672746 737923
rect 672694 737859 672746 737865
rect 672598 709205 672650 709211
rect 672598 709147 672650 709153
rect 672502 694109 672554 694115
rect 672502 694051 672554 694057
rect 672406 627805 672458 627811
rect 672406 627747 672458 627753
rect 672406 602201 672458 602207
rect 672406 602143 672458 602149
rect 672310 572897 672362 572903
rect 672310 572839 672362 572845
rect 672418 564319 672446 602143
rect 672406 564313 672458 564319
rect 672406 564255 672458 564261
rect 672406 541521 672458 541527
rect 672406 541463 672458 541469
rect 672118 529903 672170 529909
rect 672118 529845 672170 529851
rect 672022 529533 672074 529539
rect 672022 529475 672074 529481
rect 671830 528645 671882 528651
rect 671830 528587 671882 528593
rect 669718 404473 669770 404479
rect 669718 404415 669770 404421
rect 672418 360079 672446 541463
rect 672514 538567 672542 694051
rect 672706 665255 672734 737859
rect 672802 699887 672830 738081
rect 672898 708693 672926 779299
rect 672994 745989 673022 783073
rect 673270 782983 673322 782989
rect 673270 782925 673322 782931
rect 673078 779801 673130 779807
rect 673078 779743 673130 779749
rect 672982 745983 673034 745989
rect 672982 745925 673034 745931
rect 672982 733625 673034 733631
rect 672982 733567 673034 733573
rect 672886 708687 672938 708693
rect 672886 708629 672938 708635
rect 672790 699881 672842 699887
rect 672790 699823 672842 699829
rect 672790 692925 672842 692931
rect 672790 692867 672842 692873
rect 672694 665249 672746 665255
rect 672694 665191 672746 665197
rect 672598 644085 672650 644091
rect 672598 644027 672650 644033
rect 672610 573495 672638 644027
rect 672694 622181 672746 622187
rect 672694 622123 672746 622129
rect 672598 573489 672650 573495
rect 672598 573431 672650 573437
rect 672502 538561 672554 538567
rect 672502 538503 672554 538509
rect 672598 529977 672650 529983
rect 672598 529919 672650 529925
rect 672502 446431 672554 446437
rect 672502 446373 672554 446379
rect 672406 360073 672458 360079
rect 672406 360015 672458 360021
rect 672514 270687 672542 446373
rect 672610 359043 672638 529919
rect 672706 492465 672734 622123
rect 672802 619227 672830 692867
rect 672994 662369 673022 733567
rect 673090 707551 673118 779743
rect 673174 778617 673226 778623
rect 673174 778559 673226 778565
rect 673076 707542 673132 707551
rect 673076 707477 673132 707486
rect 673186 707107 673214 778559
rect 673282 708143 673310 782925
rect 673378 752099 673406 866915
rect 673858 761275 673886 939097
rect 674050 934731 674078 952015
rect 674146 936951 674174 953865
rect 675106 953527 675134 958379
rect 675490 957671 675518 958078
rect 675476 957662 675532 957671
rect 675476 957597 675532 957606
rect 675490 957037 675518 957412
rect 675190 957031 675242 957037
rect 675190 956973 675242 956979
rect 675478 957031 675530 957037
rect 675478 956973 675530 956979
rect 675092 953518 675148 953527
rect 675092 953453 675148 953462
rect 675202 953379 675230 956973
rect 675490 956043 675518 956228
rect 675476 956034 675532 956043
rect 675476 955969 675532 955978
rect 675394 954743 675422 955044
rect 675382 954737 675434 954743
rect 675382 954679 675434 954685
rect 675490 953929 675518 954378
rect 675478 953923 675530 953929
rect 675478 953865 675530 953871
rect 675188 953370 675244 953379
rect 675188 953305 675244 953314
rect 675490 952079 675518 952528
rect 675478 952073 675530 952079
rect 675478 952015 675530 952021
rect 676820 940938 676876 940947
rect 676820 940873 676876 940882
rect 674612 939902 674668 939911
rect 674612 939837 674668 939846
rect 674420 939606 674476 939615
rect 674420 939541 674422 939550
rect 674474 939541 674476 939550
rect 674422 939509 674474 939515
rect 674626 939425 674654 939837
rect 674614 939419 674666 939425
rect 674614 939361 674666 939367
rect 676834 939277 676862 940873
rect 676916 940494 676972 940503
rect 676916 940429 676972 940438
rect 676822 939271 676874 939277
rect 676822 939213 676874 939219
rect 676930 939129 676958 940429
rect 676918 939123 676970 939129
rect 676918 939065 676970 939071
rect 676820 938274 676876 938283
rect 676820 938209 676876 938218
rect 674422 938013 674474 938019
rect 674420 937978 674422 937987
rect 674474 937978 674476 937987
rect 674420 937913 674476 937922
rect 674132 936942 674188 936951
rect 674132 936877 674188 936886
rect 676834 936169 676862 938209
rect 676822 936163 676874 936169
rect 676822 936105 676874 936111
rect 674036 934722 674092 934731
rect 674036 934657 674092 934666
rect 677012 929542 677068 929551
rect 677012 929477 677068 929486
rect 676820 928950 676876 928959
rect 676820 928885 676876 928894
rect 676834 928515 676862 928885
rect 677026 928515 677054 929477
rect 676820 928506 676876 928515
rect 676820 928441 676876 928450
rect 677012 928506 677068 928515
rect 677012 928441 677068 928450
rect 677026 927437 677054 928441
rect 677014 927431 677066 927437
rect 677014 927373 677066 927379
rect 675394 877011 675422 877523
rect 675380 877002 675436 877011
rect 675380 876937 675436 876946
rect 675394 876567 675422 876900
rect 675380 876558 675436 876567
rect 675380 876493 675436 876502
rect 675284 875966 675340 875975
rect 675284 875901 675340 875910
rect 675092 875670 675148 875679
rect 675092 875605 675148 875614
rect 674614 872153 674666 872159
rect 674614 872095 674666 872101
rect 674422 869045 674474 869051
rect 674422 868987 674474 868993
rect 674326 865049 674378 865055
rect 674326 864991 674378 864997
rect 674134 773659 674186 773665
rect 674134 773601 674186 773607
rect 673844 761266 673900 761275
rect 673844 761201 673900 761210
rect 673844 760674 673900 760683
rect 673844 760609 673900 760618
rect 673858 760493 673886 760609
rect 673846 760487 673898 760493
rect 673846 760429 673898 760435
rect 673364 752090 673420 752099
rect 673364 752025 673420 752034
rect 674146 745471 674174 773601
rect 674338 773115 674366 864991
rect 674434 862095 674462 868987
rect 674518 866529 674570 866535
rect 674518 866471 674570 866477
rect 674422 862089 674474 862095
rect 674422 862031 674474 862037
rect 674530 777555 674558 866471
rect 674516 777546 674572 777555
rect 674516 777481 674572 777490
rect 674626 776963 674654 872095
rect 675106 871512 675134 875605
rect 674818 871493 675134 871512
rect 675298 872030 675326 875901
rect 675394 875827 675422 876234
rect 675380 875818 675436 875827
rect 675380 875753 675436 875762
rect 675490 874199 675518 874384
rect 675476 874190 675532 874199
rect 675476 874125 675532 874134
rect 675394 873459 675422 873866
rect 675380 873450 675436 873459
rect 675380 873385 675436 873394
rect 675394 872867 675422 873200
rect 675380 872858 675436 872867
rect 675380 872793 675436 872802
rect 675490 872159 675518 872534
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 675298 872002 675408 872030
rect 674818 871487 675146 871493
rect 674818 871484 675094 871487
rect 674818 864556 674846 871484
rect 675094 871429 675146 871435
rect 675298 871216 675326 872002
rect 675382 871487 675434 871493
rect 675382 871429 675434 871435
rect 675394 871350 675422 871429
rect 675106 871188 675326 871216
rect 675106 869440 675134 871188
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675298 869560 675422 869588
rect 675298 869514 675326 869560
rect 675010 869412 675134 869440
rect 675202 869486 675326 869514
rect 675394 869500 675422 869560
rect 675010 864852 675038 869412
rect 675202 869051 675230 869486
rect 675190 869045 675242 869051
rect 675190 868987 675242 868993
rect 675106 868861 675408 868889
rect 675106 865055 675134 868861
rect 675202 868228 675408 868256
rect 675202 866979 675230 868228
rect 675190 866973 675242 866979
rect 675190 866915 675242 866921
rect 675394 866535 675422 867058
rect 675382 866529 675434 866535
rect 675382 866471 675434 866477
rect 675202 865825 675408 865853
rect 675094 865049 675146 865055
rect 675094 864991 675146 864997
rect 675010 864824 675134 864852
rect 674818 864528 675038 864556
rect 674900 862202 674956 862211
rect 674818 862160 674900 862188
rect 674612 776954 674668 776963
rect 674612 776889 674668 776898
rect 674422 775509 674474 775515
rect 674422 775451 674474 775457
rect 674324 773106 674380 773115
rect 674324 773041 674380 773050
rect 674326 762929 674378 762935
rect 674324 762894 674326 762903
rect 674378 762894 674380 762903
rect 674324 762829 674380 762838
rect 674326 762337 674378 762343
rect 674324 762302 674326 762311
rect 674378 762302 674380 762311
rect 674324 762237 674380 762246
rect 674134 745465 674186 745471
rect 674134 745407 674186 745413
rect 674230 735475 674282 735481
rect 674230 735417 674282 735423
rect 673366 734957 673418 734963
rect 673366 734899 673418 734905
rect 673268 708134 673324 708143
rect 673268 708069 673324 708078
rect 673172 707098 673228 707107
rect 673172 707033 673228 707042
rect 673174 699881 673226 699887
rect 673174 699823 673226 699829
rect 673186 693005 673214 699823
rect 673174 692999 673226 693005
rect 673174 692941 673226 692947
rect 673078 688633 673130 688639
rect 673078 688575 673130 688581
rect 672982 662363 673034 662369
rect 672982 662305 673034 662311
rect 672886 643419 672938 643425
rect 672886 643361 672938 643367
rect 672790 619221 672842 619227
rect 672790 619163 672842 619169
rect 672790 597169 672842 597175
rect 672790 597111 672842 597117
rect 672802 529613 672830 597111
rect 672898 571867 672926 643361
rect 673090 616827 673118 688575
rect 673186 653785 673214 692941
rect 673270 689817 673322 689823
rect 673270 689759 673322 689765
rect 673174 653779 673226 653785
rect 673174 653721 673226 653727
rect 673282 617419 673310 689759
rect 673378 662411 673406 734899
rect 674242 728969 674270 735417
rect 674230 728963 674282 728969
rect 674230 728905 674282 728911
rect 674434 728840 674462 775451
rect 674818 774868 674846 862160
rect 674900 862137 674956 862146
rect 674902 862089 674954 862095
rect 674902 862031 674954 862037
rect 674914 776223 674942 862031
rect 675010 861133 675038 864528
rect 674998 861127 675050 861133
rect 674998 861069 675050 861075
rect 674998 800669 675050 800675
rect 674998 800611 675050 800617
rect 675010 782545 675038 800611
rect 675106 783137 675134 864824
rect 675202 864093 675230 865825
rect 675394 864727 675422 865208
rect 675380 864718 675436 864727
rect 675380 864653 675436 864662
rect 675190 864087 675242 864093
rect 675190 864029 675242 864035
rect 675202 863344 675408 863372
rect 675202 862211 675230 863344
rect 675188 862202 675244 862211
rect 675188 862137 675244 862146
rect 675190 861127 675242 861133
rect 675190 861069 675242 861075
rect 675202 800675 675230 861069
rect 675190 800669 675242 800675
rect 675190 800611 675242 800617
rect 675778 788063 675806 788322
rect 675764 788054 675820 788063
rect 675764 787989 675820 787998
rect 675490 787175 675518 787656
rect 675476 787166 675532 787175
rect 675476 787101 675532 787110
rect 675778 786731 675806 787035
rect 675764 786722 675820 786731
rect 675764 786657 675820 786666
rect 675778 784955 675806 785214
rect 675764 784946 675820 784955
rect 675764 784881 675820 784890
rect 675682 784215 675710 784622
rect 675668 784206 675724 784215
rect 675668 784141 675724 784150
rect 675394 783507 675422 783999
rect 675382 783501 675434 783507
rect 675382 783443 675434 783449
rect 675094 783131 675146 783137
rect 675094 783073 675146 783079
rect 675394 782989 675422 783364
rect 675478 783131 675530 783137
rect 675478 783073 675530 783079
rect 675382 782983 675434 782989
rect 675382 782925 675434 782931
rect 675490 782803 675518 783073
rect 674998 782539 675050 782545
rect 674998 782481 675050 782487
rect 675478 782539 675530 782545
rect 675478 782481 675530 782487
rect 675490 782194 675518 782481
rect 675490 782180 675792 782194
rect 675504 782166 675806 782180
rect 675778 781995 675806 782166
rect 675764 781986 675820 781995
rect 675764 781921 675820 781930
rect 675778 780663 675806 780848
rect 675764 780654 675820 780663
rect 675764 780589 675820 780598
rect 675094 780541 675146 780547
rect 675094 780483 675146 780489
rect 675106 777069 675134 780483
rect 675394 779807 675422 780330
rect 675382 779801 675434 779807
rect 675382 779743 675434 779749
rect 675490 779363 675518 779664
rect 675478 779357 675530 779363
rect 675478 779299 675530 779305
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675490 777661 675518 777814
rect 675478 777655 675530 777661
rect 675478 777597 675530 777603
rect 675094 777063 675146 777069
rect 675094 777005 675146 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 674900 776214 674956 776223
rect 674900 776149 674956 776158
rect 675394 775515 675422 775995
rect 675382 775509 675434 775515
rect 675382 775451 675434 775457
rect 674900 774882 674956 774891
rect 674818 774840 674900 774868
rect 674900 774817 674956 774826
rect 675490 773665 675518 774155
rect 675478 773659 675530 773665
rect 675478 773601 675530 773607
rect 674614 762041 674666 762047
rect 674612 762006 674614 762015
rect 674666 762006 674668 762015
rect 674612 761941 674668 761950
rect 677876 760378 677932 760387
rect 677876 760313 677932 760322
rect 677890 759943 677918 760313
rect 677876 759934 677932 759943
rect 677876 759869 677932 759878
rect 676916 759786 676972 759795
rect 676916 759721 676972 759730
rect 676930 756095 676958 759721
rect 677588 759342 677644 759351
rect 677588 759277 677644 759286
rect 676916 756086 676972 756095
rect 676916 756021 676972 756030
rect 677602 753431 677630 759277
rect 677588 753422 677644 753431
rect 677588 753357 677644 753366
rect 677012 751202 677068 751211
rect 677012 751137 677068 751146
rect 677026 750619 677054 751137
rect 676820 750610 676876 750619
rect 676820 750545 676876 750554
rect 677012 750610 677068 750619
rect 677012 750545 677068 750554
rect 676834 750175 676862 750545
rect 676820 750166 676876 750175
rect 676820 750101 676876 750110
rect 677026 748875 677054 750545
rect 677014 748869 677066 748875
rect 677014 748811 677066 748817
rect 675094 745983 675146 745989
rect 675094 745925 675146 745931
rect 674518 745465 674570 745471
rect 674518 745407 674570 745413
rect 674146 728812 674462 728840
rect 673748 715682 673804 715691
rect 673748 715617 673804 715626
rect 673762 671143 673790 715617
rect 674146 713619 674174 728812
rect 674230 728741 674282 728747
rect 674230 728683 674282 728689
rect 674132 713610 674188 713619
rect 674132 713545 674188 713554
rect 673748 671134 673804 671143
rect 673748 671069 673804 671078
rect 674242 666703 674270 728683
rect 674326 728667 674378 728673
rect 674326 728609 674378 728615
rect 674338 713596 674366 728609
rect 674530 728123 674558 745407
rect 675106 738145 675134 745925
rect 675394 743219 675422 743330
rect 675380 743210 675436 743219
rect 675380 743145 675436 743154
rect 675490 742479 675518 742664
rect 675476 742470 675532 742479
rect 675476 742405 675532 742414
rect 675490 741739 675518 742035
rect 675476 741730 675532 741739
rect 675476 741665 675532 741674
rect 675188 740398 675244 740407
rect 675188 740333 675244 740342
rect 675094 738139 675146 738145
rect 675094 738081 675146 738087
rect 675202 737701 675230 740333
rect 675394 740111 675422 740222
rect 675380 740102 675436 740111
rect 675380 740037 675436 740046
rect 675490 739223 675518 739630
rect 675476 739214 675532 739223
rect 675476 739149 675532 739158
rect 675394 738631 675422 738999
rect 675380 738622 675436 738631
rect 675380 738557 675436 738566
rect 675394 737923 675422 738372
rect 675478 738139 675530 738145
rect 675478 738081 675530 738087
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 675490 737780 675518 738081
rect 675190 737695 675242 737701
rect 675190 737637 675242 737643
rect 675382 737695 675434 737701
rect 675382 737637 675434 737643
rect 675202 737572 675230 737637
rect 675010 737544 675230 737572
rect 674902 732367 674954 732373
rect 674902 732309 674954 732315
rect 674614 730517 674666 730523
rect 674614 730459 674666 730465
rect 674516 728114 674572 728123
rect 674516 728049 674572 728058
rect 674422 717937 674474 717943
rect 674420 717902 674422 717911
rect 674474 717902 674476 717911
rect 674420 717837 674476 717846
rect 674422 717345 674474 717351
rect 674420 717310 674422 717319
rect 674474 717310 674476 717319
rect 674420 717245 674476 717254
rect 674422 716901 674474 716907
rect 674420 716866 674422 716875
rect 674474 716866 674476 716875
rect 674420 716801 674476 716810
rect 674422 716309 674474 716315
rect 674420 716274 674422 716283
rect 674474 716274 674476 716283
rect 674420 716209 674476 716218
rect 674338 713568 674558 713596
rect 674422 709797 674474 709803
rect 674420 709762 674422 709771
rect 674474 709762 674476 709771
rect 674420 709697 674476 709706
rect 674422 709205 674474 709211
rect 674420 709170 674422 709179
rect 674474 709170 674476 709179
rect 674420 709105 674476 709114
rect 674422 708687 674474 708693
rect 674420 708652 674422 708661
rect 674474 708652 674476 708661
rect 674420 708587 674476 708596
rect 674326 685525 674378 685531
rect 674326 685467 674378 685473
rect 674228 666694 674284 666703
rect 674228 666629 674284 666638
rect 673846 665249 673898 665255
rect 673846 665191 673898 665197
rect 673858 662855 673886 665191
rect 673844 662846 673900 662855
rect 673844 662781 673900 662790
rect 673364 662402 673420 662411
rect 673364 662337 673420 662346
rect 673846 662363 673898 662369
rect 673846 662305 673898 662311
rect 673858 661819 673886 662305
rect 673844 661810 673900 661819
rect 673844 661745 673900 661754
rect 674230 646453 674282 646459
rect 674230 646395 674282 646401
rect 673366 642309 673418 642315
rect 673366 642251 673418 642257
rect 673268 617410 673324 617419
rect 673268 617345 673324 617354
rect 673076 616818 673132 616827
rect 673076 616753 673132 616762
rect 673270 602719 673322 602725
rect 673270 602661 673322 602667
rect 673174 601757 673226 601763
rect 673174 601699 673226 601705
rect 673078 599611 673130 599617
rect 673078 599553 673130 599559
rect 672982 598427 673034 598433
rect 672982 598369 673034 598375
rect 672886 571861 672938 571867
rect 672886 571803 672938 571809
rect 672790 529607 672842 529613
rect 672790 529549 672842 529555
rect 672994 526695 673022 598369
rect 673090 527139 673118 599553
rect 673186 590441 673214 601699
rect 673174 590435 673226 590441
rect 673174 590377 673226 590383
rect 673174 553953 673226 553959
rect 673174 553895 673226 553901
rect 673076 527130 673132 527139
rect 673076 527065 673132 527074
rect 672980 526686 673036 526695
rect 672980 526621 673036 526630
rect 672694 492459 672746 492465
rect 672694 492401 672746 492407
rect 673186 484219 673214 553895
rect 673282 527731 673310 602661
rect 673378 573759 673406 642251
rect 674132 630730 674188 630739
rect 674132 630665 674188 630674
rect 673846 627805 673898 627811
rect 673844 627770 673846 627779
rect 673898 627770 673900 627779
rect 673844 627705 673900 627714
rect 673750 622107 673802 622113
rect 673750 622049 673802 622055
rect 673462 602127 673514 602133
rect 673462 602069 673514 602075
rect 673364 573750 673420 573759
rect 673364 573685 673420 573694
rect 673474 563949 673502 602069
rect 673762 601763 673790 622049
rect 674146 619935 674174 630665
rect 674132 619926 674188 619935
rect 674132 619861 674188 619870
rect 673846 619221 673898 619227
rect 673846 619163 673898 619169
rect 673858 617863 673886 619163
rect 673844 617854 673900 617863
rect 673844 617789 673900 617798
rect 674242 613455 674270 646395
rect 674338 623339 674366 685467
rect 674422 672723 674474 672729
rect 674420 672688 674422 672697
rect 674474 672688 674476 672697
rect 674420 672623 674476 672632
rect 674422 672205 674474 672211
rect 674420 672170 674422 672179
rect 674474 672170 674476 672179
rect 674420 672105 674476 672114
rect 674422 671613 674474 671619
rect 674420 671578 674422 671587
rect 674474 671578 674476 671587
rect 674420 671513 674476 671522
rect 674530 666407 674558 713568
rect 674626 668627 674654 730459
rect 674914 684125 674942 732309
rect 675010 725787 675038 737544
rect 675094 737325 675146 737331
rect 675094 737267 675146 737273
rect 675106 732077 675134 737267
rect 675394 737159 675422 737637
rect 675490 735481 675518 735856
rect 675478 735475 675530 735481
rect 675478 735417 675530 735423
rect 675394 734963 675422 735338
rect 675382 734957 675434 734963
rect 675382 734899 675434 734905
rect 675394 734487 675422 734672
rect 675380 734478 675436 734487
rect 675380 734413 675436 734422
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675094 732071 675146 732077
rect 675094 732013 675146 732019
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 674998 725781 675050 725787
rect 674998 725723 675050 725729
rect 675382 725781 675434 725787
rect 675382 725723 675434 725729
rect 675394 705659 675422 725723
rect 677012 706210 677068 706219
rect 677012 706145 677068 706154
rect 675190 705653 675242 705659
rect 675190 705595 675242 705601
rect 675382 705653 675434 705659
rect 677026 705627 677054 706145
rect 675382 705595 675434 705601
rect 676820 705618 676876 705627
rect 675094 693517 675146 693523
rect 675094 693459 675146 693465
rect 674998 690705 675050 690711
rect 674998 690647 675050 690653
rect 675010 684125 675038 690647
rect 675106 688311 675134 693459
rect 675202 692709 675230 705595
rect 676820 705553 676876 705562
rect 677012 705618 677068 705627
rect 677012 705553 677068 705562
rect 676834 705183 676862 705553
rect 676820 705174 676876 705183
rect 676820 705109 676876 705118
rect 677026 702773 677054 705553
rect 677014 702767 677066 702773
rect 677014 702709 677066 702715
rect 675490 697931 675518 698338
rect 675476 697922 675532 697931
rect 675476 697857 675532 697866
rect 675778 697339 675806 697672
rect 675764 697330 675820 697339
rect 675764 697265 675820 697274
rect 675394 696895 675422 697035
rect 675380 696886 675436 696895
rect 675380 696821 675436 696830
rect 675682 694823 675710 695195
rect 675668 694814 675724 694823
rect 675668 694749 675724 694758
rect 675490 694379 675518 694638
rect 675476 694370 675532 694379
rect 675476 694305 675532 694314
rect 675490 693523 675518 693972
rect 675478 693517 675530 693523
rect 675478 693459 675530 693465
rect 675394 692931 675422 693380
rect 675478 692999 675530 693005
rect 675478 692941 675530 692947
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 692788 675518 692941
rect 675190 692703 675242 692709
rect 675190 692645 675242 692651
rect 675382 692703 675434 692709
rect 675382 692645 675434 692651
rect 675394 692173 675422 692645
rect 675394 692159 675792 692173
rect 675408 692145 675806 692159
rect 675778 692011 675806 692145
rect 675764 692002 675820 692011
rect 675764 691937 675820 691946
rect 675490 690711 675518 690864
rect 675478 690705 675530 690711
rect 675478 690647 675530 690653
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675778 689199 675806 689680
rect 675764 689190 675820 689199
rect 675764 689125 675820 689134
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 675092 688302 675148 688311
rect 675092 688237 675148 688246
rect 675490 687381 675518 687830
rect 675094 687375 675146 687381
rect 675094 687317 675146 687323
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 674902 684119 674954 684125
rect 674902 684061 674954 684067
rect 674998 684119 675050 684125
rect 674998 684061 675050 684067
rect 675106 683996 675134 687317
rect 675394 686271 675422 686646
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 674818 683968 675134 683996
rect 674612 668618 674668 668627
rect 674612 668553 674668 668562
rect 674516 666398 674572 666407
rect 674516 666333 674572 666342
rect 674422 661031 674474 661037
rect 674422 660973 674474 660979
rect 674324 623330 674380 623339
rect 674324 623265 674380 623274
rect 674434 621119 674462 660973
rect 674614 655259 674666 655265
rect 674614 655201 674666 655207
rect 674518 647119 674570 647125
rect 674518 647061 674570 647067
rect 674420 621110 674476 621119
rect 674420 621045 674476 621054
rect 674230 613449 674282 613455
rect 674230 613391 674282 613397
rect 674530 602133 674558 647061
rect 674626 645275 674654 655201
rect 674614 645269 674666 645275
rect 674614 645211 674666 645217
rect 674614 627361 674666 627367
rect 674612 627326 674614 627335
rect 674666 627326 674668 627335
rect 674612 627261 674668 627270
rect 674614 626917 674666 626923
rect 674612 626882 674614 626891
rect 674666 626882 674668 626891
rect 674612 626817 674668 626826
rect 674612 625254 674668 625263
rect 674612 625189 674614 625198
rect 674666 625189 674668 625198
rect 674614 625157 674666 625163
rect 674818 619172 674846 683968
rect 674998 683897 675050 683903
rect 674998 683839 675050 683845
rect 674902 683823 674954 683829
rect 674902 683765 674954 683771
rect 674914 664187 674942 683765
rect 675010 681017 675038 683839
rect 675490 683681 675518 684130
rect 675094 683675 675146 683681
rect 675094 683617 675146 683623
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 674998 681011 675050 681017
rect 674998 680953 675050 680959
rect 674900 664178 674956 664187
rect 674900 664113 674956 664122
rect 675106 661037 675134 683617
rect 675190 681011 675242 681017
rect 675190 680953 675242 680959
rect 675094 661031 675146 661037
rect 675094 660973 675146 660979
rect 674900 660922 674956 660931
rect 674900 660857 674956 660866
rect 674914 660487 674942 660857
rect 674900 660478 674956 660487
rect 674900 660413 674956 660422
rect 675092 660478 675148 660487
rect 675092 660413 675148 660422
rect 674914 659557 674942 660413
rect 675106 659895 675134 660413
rect 675092 659886 675148 659895
rect 675092 659821 675148 659830
rect 674902 659551 674954 659557
rect 674902 659493 674954 659499
rect 675202 655265 675230 680953
rect 675190 655259 675242 655265
rect 675190 655201 675242 655207
rect 675190 653779 675242 653785
rect 675190 653721 675242 653727
rect 675092 653670 675148 653679
rect 675092 653605 675148 653614
rect 675106 646459 675134 653605
rect 675202 647125 675230 653721
rect 675394 652643 675422 653124
rect 675380 652634 675436 652643
rect 675380 652569 675436 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675490 651459 675518 651835
rect 675476 651450 675532 651459
rect 675476 651385 675532 651394
rect 675394 649683 675422 650016
rect 675380 649674 675436 649683
rect 675380 649609 675436 649618
rect 675490 648943 675518 649424
rect 675476 648934 675532 648943
rect 675476 648869 675532 648878
rect 675394 648309 675422 648799
rect 675382 648303 675434 648309
rect 675382 648245 675434 648251
rect 675394 648087 675422 648166
rect 675382 648081 675434 648087
rect 675382 648023 675434 648029
rect 675394 647125 675422 647603
rect 675190 647119 675242 647125
rect 675190 647061 675242 647067
rect 675382 647119 675434 647125
rect 675382 647061 675434 647067
rect 675394 646459 675422 646982
rect 675094 646453 675146 646459
rect 675094 646395 675146 646401
rect 675382 646453 675434 646459
rect 675382 646395 675434 646401
rect 675778 645391 675806 645650
rect 675764 645382 675820 645391
rect 675764 645317 675820 645326
rect 674902 645269 674954 645275
rect 674902 645211 674954 645217
rect 674914 622007 674942 645211
rect 675094 645195 675146 645201
rect 675094 645137 675146 645143
rect 675106 641871 675134 645137
rect 675490 644609 675518 645132
rect 675478 644603 675530 644609
rect 675478 644545 675530 644551
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675094 641865 675146 641871
rect 675094 641807 675146 641813
rect 675382 641865 675434 641871
rect 675382 641807 675434 641813
rect 675394 641432 675422 641807
rect 675394 640359 675422 640795
rect 675380 640350 675436 640359
rect 675380 640285 675436 640294
rect 675778 638583 675806 638955
rect 675764 638574 675820 638583
rect 675764 638509 675820 638518
rect 674996 630730 675052 630739
rect 674996 630665 675052 630674
rect 674900 621998 674956 622007
rect 674900 621933 674956 621942
rect 675010 620823 675038 630665
rect 677204 624662 677260 624671
rect 677204 624597 677260 624606
rect 676820 624070 676876 624079
rect 676820 624005 676876 624014
rect 676834 622113 676862 624005
rect 677218 622261 677246 624597
rect 677206 622255 677258 622261
rect 677206 622197 677258 622203
rect 676822 622107 676874 622113
rect 676822 622049 676874 622055
rect 674996 620814 675052 620823
rect 674996 620749 675052 620758
rect 674900 619186 674956 619195
rect 674818 619144 674900 619172
rect 674900 619121 674956 619130
rect 677108 615930 677164 615939
rect 677108 615865 677164 615874
rect 677122 615347 677150 615865
rect 676916 615338 676972 615347
rect 676916 615273 676972 615282
rect 677108 615338 677164 615347
rect 677108 615273 677164 615282
rect 676930 614903 676958 615273
rect 676916 614894 676972 614903
rect 676916 614829 676972 614838
rect 677122 613529 677150 615273
rect 677110 613523 677162 613529
rect 677110 613465 677162 613471
rect 675190 613449 675242 613455
rect 675190 613391 675242 613397
rect 675202 602207 675230 613391
rect 675394 607799 675422 608132
rect 675380 607790 675436 607799
rect 675380 607725 675436 607734
rect 675490 607207 675518 607466
rect 675476 607198 675532 607207
rect 675476 607133 675532 607142
rect 675490 606467 675518 606835
rect 675476 606458 675532 606467
rect 675476 606393 675532 606402
rect 675394 604839 675422 604995
rect 675380 604830 675436 604839
rect 675380 604765 675436 604774
rect 675490 604131 675518 604432
rect 675478 604125 675530 604131
rect 675478 604067 675530 604073
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675394 602725 675422 603174
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 675190 602201 675242 602207
rect 675190 602143 675242 602149
rect 675382 602201 675434 602207
rect 675382 602143 675434 602149
rect 674518 602127 674570 602133
rect 674518 602069 674570 602075
rect 675094 601979 675146 601985
rect 675394 601959 675422 602143
rect 675490 602133 675518 602582
rect 675478 602127 675530 602133
rect 675478 602069 675530 602075
rect 675094 601921 675146 601927
rect 673750 601757 673802 601763
rect 673750 601699 673802 601705
rect 674614 600425 674666 600431
rect 674614 600367 674666 600373
rect 674626 590483 674654 600367
rect 675106 596879 675134 601921
rect 675490 600431 675518 600658
rect 675478 600425 675530 600431
rect 675478 600367 675530 600373
rect 675394 599617 675422 600140
rect 675382 599611 675434 599617
rect 675382 599553 675434 599559
rect 675394 599099 675422 599474
rect 675382 599093 675434 599099
rect 675382 599035 675434 599041
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 675094 596873 675146 596879
rect 675094 596815 675146 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675092 595506 675148 595515
rect 675092 595441 675148 595450
rect 674900 590622 674956 590631
rect 674900 590557 674956 590566
rect 674612 590474 674668 590483
rect 673846 590435 673898 590441
rect 674612 590409 674668 590418
rect 673846 590377 673898 590383
rect 673858 587555 673886 590377
rect 674914 590187 674942 590557
rect 675106 590515 675134 595441
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 675094 590509 675146 590515
rect 675094 590451 675146 590457
rect 675478 590509 675530 590515
rect 675478 590451 675530 590457
rect 675490 590335 675518 590451
rect 675476 590326 675532 590335
rect 675476 590261 675532 590270
rect 674900 590178 674956 590187
rect 674900 590113 674956 590122
rect 676918 588807 676970 588813
rect 676918 588749 676970 588755
rect 673846 587549 673898 587555
rect 673846 587491 673898 587497
rect 676822 587549 676874 587555
rect 676822 587491 676874 587497
rect 674612 582186 674668 582195
rect 674612 582121 674668 582130
rect 674422 582073 674474 582079
rect 674422 582015 674474 582021
rect 674434 581973 674462 582015
rect 674626 582005 674654 582121
rect 674614 581999 674666 582005
rect 674420 581964 674476 581973
rect 674614 581941 674666 581947
rect 674420 581899 674476 581908
rect 674614 581629 674666 581635
rect 674612 581594 674614 581603
rect 674666 581594 674668 581603
rect 674612 581529 674668 581538
rect 674422 580889 674474 580895
rect 674420 580854 674422 580863
rect 674474 580854 674476 580863
rect 674420 580789 674476 580798
rect 674612 580114 674668 580123
rect 674612 580049 674614 580058
rect 674666 580049 674668 580058
rect 674614 580017 674666 580023
rect 676834 579531 676862 587491
rect 676930 580123 676958 588749
rect 676916 580114 676972 580123
rect 676916 580049 676972 580058
rect 676820 579522 676876 579531
rect 676820 579457 676876 579466
rect 674614 574525 674666 574531
rect 674612 574490 674614 574499
rect 674666 574490 674668 574499
rect 674612 574425 674668 574434
rect 674614 573489 674666 573495
rect 674612 573454 674614 573463
rect 674666 573454 674668 573463
rect 674612 573389 674668 573398
rect 673750 573119 673802 573125
rect 673750 573061 673802 573067
rect 673762 572131 673790 573061
rect 674614 572897 674666 572903
rect 674612 572862 674614 572871
rect 674666 572862 674668 572871
rect 674612 572797 674668 572806
rect 673748 572122 673804 572131
rect 673748 572057 673804 572066
rect 674614 571861 674666 571867
rect 674612 571826 674614 571835
rect 674666 571826 674668 571835
rect 674612 571761 674668 571770
rect 677012 570790 677068 570799
rect 677012 570725 677068 570734
rect 677026 570207 677054 570725
rect 676820 570198 676876 570207
rect 676820 570133 676876 570142
rect 677012 570198 677068 570207
rect 677012 570133 677068 570142
rect 676834 569763 676862 570133
rect 676820 569754 676876 569763
rect 676820 569689 676876 569698
rect 677026 567427 677054 570133
rect 677014 567421 677066 567427
rect 677014 567363 677066 567369
rect 675094 564313 675146 564319
rect 675094 564255 675146 564261
rect 673462 563943 673514 563949
rect 673462 563885 673514 563891
rect 674614 559429 674666 559435
rect 674614 559371 674666 559377
rect 673462 557653 673514 557659
rect 673462 557595 673514 557601
rect 673366 553213 673418 553219
rect 673366 553155 673418 553161
rect 673268 527722 673324 527731
rect 673268 527657 673324 527666
rect 673172 484210 673228 484219
rect 673172 484145 673228 484154
rect 673378 482591 673406 553155
rect 673474 483775 673502 557595
rect 674422 555285 674474 555291
rect 674422 555227 674474 555233
rect 674326 551955 674378 551961
rect 674326 551897 674378 551903
rect 673750 538561 673802 538567
rect 673750 538503 673802 538509
rect 673762 536907 673790 538503
rect 673748 536898 673804 536907
rect 673748 536833 673804 536842
rect 673750 536785 673802 536791
rect 673750 536727 673802 536733
rect 673762 535871 673790 536727
rect 673748 535862 673804 535871
rect 673748 535797 673804 535806
rect 673748 529942 673804 529951
rect 673748 529877 673750 529886
rect 673802 529877 673804 529886
rect 673750 529845 673802 529851
rect 673750 529607 673802 529613
rect 673750 529549 673802 529555
rect 673762 528767 673790 529549
rect 673748 528758 673804 528767
rect 673748 528693 673804 528702
rect 673750 528645 673802 528651
rect 673750 528587 673802 528593
rect 673762 528323 673790 528587
rect 673748 528314 673804 528323
rect 673748 528249 673804 528258
rect 674338 499736 674366 551897
rect 674242 499708 674366 499736
rect 673846 492459 673898 492465
rect 673846 492401 673898 492407
rect 673858 492359 673886 492401
rect 673844 492350 673900 492359
rect 673844 492285 673900 492294
rect 674242 484811 674270 499708
rect 674326 492977 674378 492983
rect 674324 492942 674326 492951
rect 674378 492942 674380 492951
rect 674324 492877 674380 492886
rect 674434 487475 674462 555227
rect 674518 548255 674570 548261
rect 674518 548197 674570 548203
rect 674530 536440 674558 548197
rect 674626 536791 674654 559371
rect 674902 558097 674954 558103
rect 674902 558039 674954 558045
rect 674914 550111 674942 558039
rect 675106 557141 675134 564255
rect 675190 563943 675242 563949
rect 675190 563885 675242 563891
rect 675202 557881 675230 563885
rect 675490 562511 675518 562918
rect 675476 562502 675532 562511
rect 675476 562437 675532 562446
rect 675490 562067 675518 562252
rect 675476 562058 675532 562067
rect 675476 561993 675532 562002
rect 675394 561475 675422 561660
rect 675380 561466 675436 561475
rect 675380 561401 675436 561410
rect 675394 559435 675422 559810
rect 675382 559429 675434 559435
rect 675382 559371 675434 559377
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675190 557875 675242 557881
rect 675190 557817 675242 557823
rect 675382 557875 675434 557881
rect 675382 557817 675434 557823
rect 675394 557403 675422 557817
rect 675490 557659 675518 557960
rect 675478 557653 675530 557659
rect 675478 557595 675530 557601
rect 675094 557135 675146 557141
rect 675094 557077 675146 557083
rect 675478 557135 675530 557141
rect 675478 557077 675530 557083
rect 675490 556776 675518 557077
rect 675094 555877 675146 555883
rect 675094 555819 675146 555825
rect 675106 551665 675134 555819
rect 675490 555291 675518 555444
rect 675478 555285 675530 555291
rect 675478 555227 675530 555233
rect 675778 554519 675806 554926
rect 675764 554510 675820 554519
rect 675764 554445 675820 554454
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675094 551659 675146 551665
rect 675094 551601 675146 551607
rect 675382 551659 675434 551665
rect 675382 551601 675434 551607
rect 675394 551226 675422 551601
rect 675490 550111 675518 550595
rect 674902 550105 674954 550111
rect 674902 550047 674954 550053
rect 675094 550105 675146 550111
rect 675094 550047 675146 550053
rect 675478 550105 675530 550111
rect 675478 550047 675530 550053
rect 674902 549883 674954 549889
rect 674902 549825 674954 549831
rect 674914 549760 674942 549825
rect 674818 549732 674942 549760
rect 674614 536785 674666 536791
rect 674614 536727 674666 536733
rect 674614 536637 674666 536643
rect 674612 536602 674614 536611
rect 674666 536602 674668 536611
rect 674612 536537 674668 536546
rect 674530 536412 674654 536440
rect 674518 536341 674570 536347
rect 674518 536283 674570 536289
rect 674530 489399 674558 536283
rect 674626 499717 674654 536412
rect 674614 499711 674666 499717
rect 674614 499653 674666 499659
rect 674612 493238 674668 493247
rect 674612 493173 674668 493182
rect 674626 492539 674654 493173
rect 674614 492533 674666 492539
rect 674614 492475 674666 492481
rect 674516 489390 674572 489399
rect 674516 489325 674572 489334
rect 674420 487466 674476 487475
rect 674420 487401 674476 487410
rect 674818 485528 674846 549732
rect 674902 536785 674954 536791
rect 674902 536727 674954 536733
rect 674914 529909 674942 536727
rect 675106 536347 675134 550047
rect 675490 548261 675518 548755
rect 675478 548255 675530 548261
rect 675478 548197 675530 548203
rect 676820 537194 676876 537203
rect 676820 537129 676876 537138
rect 675094 536341 675146 536347
rect 675094 536283 675146 536289
rect 676834 535829 676862 537129
rect 676822 535823 676874 535829
rect 676822 535765 676874 535771
rect 677396 534974 677452 534983
rect 677396 534909 677452 534918
rect 677204 534530 677260 534539
rect 677204 534465 677260 534474
rect 677012 533938 677068 533947
rect 677012 533873 677068 533882
rect 674902 529903 674954 529909
rect 674902 529845 674954 529851
rect 675190 529903 675242 529909
rect 675190 529845 675242 529851
rect 674902 529533 674954 529539
rect 674900 529498 674902 529507
rect 674954 529498 674956 529507
rect 674900 529433 674956 529442
rect 675202 524156 675230 529845
rect 676820 525206 676876 525215
rect 676820 525141 676876 525150
rect 676834 524771 676862 525141
rect 676820 524762 676876 524771
rect 676820 524697 676876 524706
rect 675106 524128 675230 524156
rect 675106 514147 675134 524128
rect 674902 514141 674954 514147
rect 674902 514083 674954 514089
rect 675094 514141 675146 514147
rect 675094 514083 675146 514089
rect 674914 504051 674942 514083
rect 677026 509800 677054 533873
rect 677108 525798 677164 525807
rect 677108 525733 677164 525742
rect 677122 525215 677150 525733
rect 677108 525206 677164 525215
rect 677108 525141 677164 525150
rect 677122 524359 677150 525141
rect 677110 524353 677162 524359
rect 677110 524295 677162 524301
rect 676834 509772 677054 509800
rect 674900 504042 674956 504051
rect 674900 503977 674956 503986
rect 675092 504042 675148 504051
rect 675092 503977 675148 503986
rect 674998 499711 675050 499717
rect 674998 499653 675050 499659
rect 675010 487179 675038 499653
rect 675106 496017 675134 503977
rect 675094 496011 675146 496017
rect 675094 495953 675146 495959
rect 675382 496011 675434 496017
rect 675382 495953 675434 495959
rect 675394 488363 675422 495953
rect 676834 490583 676862 509772
rect 677218 491175 677246 534465
rect 677410 492211 677438 534909
rect 677396 492202 677452 492211
rect 677396 492137 677452 492146
rect 677204 491166 677260 491175
rect 677204 491101 677260 491110
rect 676820 490574 676876 490583
rect 676820 490509 676876 490518
rect 675380 488354 675436 488363
rect 675380 488289 675436 488298
rect 674996 487170 675052 487179
rect 674996 487105 675052 487114
rect 674900 485542 674956 485551
rect 674818 485500 674900 485528
rect 674900 485477 674956 485486
rect 674228 484802 674284 484811
rect 674228 484737 674284 484746
rect 673460 483766 673516 483775
rect 673460 483701 673516 483710
rect 673364 482582 673420 482591
rect 673364 482517 673420 482526
rect 677012 481694 677068 481703
rect 677012 481629 677068 481638
rect 677026 481259 677054 481629
rect 676820 481250 676876 481259
rect 676820 481185 676876 481194
rect 677012 481250 677068 481259
rect 677012 481185 677068 481194
rect 676834 480815 676862 481185
rect 676820 480806 676876 480815
rect 676820 480741 676876 480750
rect 677026 479515 677054 481185
rect 677014 479509 677066 479515
rect 677014 479451 677066 479457
rect 674710 405509 674762 405515
rect 674708 405474 674710 405483
rect 674762 405474 674764 405483
rect 674708 405409 674764 405418
rect 674422 404769 674474 404775
rect 674420 404734 674422 404743
rect 674474 404734 674476 404743
rect 674420 404669 674476 404678
rect 674710 404473 674762 404479
rect 674708 404438 674710 404447
rect 674762 404438 674764 404447
rect 674708 404373 674764 404382
rect 673652 403106 673708 403115
rect 673652 403041 673708 403050
rect 673462 400551 673514 400557
rect 673462 400493 673514 400499
rect 673366 400477 673418 400483
rect 673366 400419 673418 400425
rect 673378 374403 673406 400419
rect 673364 374394 673420 374403
rect 673364 374329 673420 374338
rect 673474 373071 673502 400493
rect 673666 400409 673694 403041
rect 677300 402366 677356 402375
rect 677300 402301 677356 402310
rect 677108 401774 677164 401783
rect 677108 401709 677164 401718
rect 674900 401330 674956 401339
rect 674900 401265 674956 401274
rect 673654 400403 673706 400409
rect 673654 400345 673706 400351
rect 673846 400403 673898 400409
rect 673846 400345 673898 400351
rect 673460 373062 673516 373071
rect 673460 372997 673516 373006
rect 672598 359037 672650 359043
rect 672598 358979 672650 358985
rect 673858 358419 673886 400345
rect 674516 399702 674572 399711
rect 674516 399637 674572 399646
rect 674420 397630 674476 397639
rect 674420 397565 674476 397574
rect 673940 396594 673996 396603
rect 673940 396529 673996 396538
rect 673954 375767 673982 396529
rect 674228 394374 674284 394383
rect 674228 394309 674284 394318
rect 674242 376877 674270 394309
rect 674434 382353 674462 397565
rect 674530 383167 674558 399637
rect 674612 395854 674668 395863
rect 674612 395789 674668 395798
rect 674518 383161 674570 383167
rect 674518 383103 674570 383109
rect 674422 382347 674474 382353
rect 674422 382289 674474 382295
rect 674626 377617 674654 395789
rect 674708 395114 674764 395123
rect 674708 395049 674764 395058
rect 674722 385239 674750 395049
rect 674804 394670 674860 394679
rect 674804 394605 674860 394614
rect 674710 385233 674762 385239
rect 674710 385175 674762 385181
rect 674818 378209 674846 394605
rect 674914 384869 674942 401265
rect 677122 400483 677150 401709
rect 677314 400557 677342 402301
rect 677302 400551 677354 400557
rect 677302 400493 677354 400499
rect 677110 400477 677162 400483
rect 677110 400419 677162 400425
rect 674996 400146 675052 400155
rect 674996 400081 675052 400090
rect 675010 386201 675038 400081
rect 675188 397926 675244 397935
rect 675188 397861 675244 397870
rect 675092 396890 675148 396899
rect 675092 396825 675148 396834
rect 674998 386195 675050 386201
rect 674998 386137 675050 386143
rect 675106 385443 675134 396825
rect 675202 385535 675230 397861
rect 677108 393486 677164 393495
rect 677108 393421 677164 393430
rect 677122 393051 677150 393421
rect 676916 393042 676972 393051
rect 676916 392977 676972 392986
rect 677108 393042 677164 393051
rect 677108 392977 677164 392986
rect 676930 392607 676958 392977
rect 676916 392598 676972 392607
rect 676916 392533 676972 392542
rect 677122 391825 677150 392977
rect 677110 391819 677162 391825
rect 677110 391761 677162 391767
rect 675382 386195 675434 386201
rect 675382 386137 675434 386143
rect 675394 385723 675422 386137
rect 675190 385529 675242 385535
rect 675190 385471 675242 385477
rect 675478 385455 675530 385461
rect 675106 385415 675230 385443
rect 674998 385233 675050 385239
rect 674998 385175 675050 385181
rect 674902 384863 674954 384869
rect 674902 384805 674954 384811
rect 675010 381040 675038 385175
rect 675202 381410 675230 385415
rect 675478 385397 675530 385403
rect 675490 385096 675518 385397
rect 675382 384863 675434 384869
rect 675382 384805 675434 384811
rect 675394 384430 675422 384805
rect 675382 383161 675434 383167
rect 675382 383103 675434 383109
rect 675394 382580 675422 383103
rect 675478 382347 675530 382353
rect 675478 382289 675530 382295
rect 675490 382062 675518 382289
rect 675202 381382 675408 381410
rect 675010 381012 675422 381040
rect 675394 380730 675422 381012
rect 675106 380198 675408 380226
rect 674806 378203 674858 378209
rect 674806 378145 674858 378151
rect 674614 377611 674666 377617
rect 674614 377553 674666 377559
rect 674230 376871 674282 376877
rect 674230 376813 674282 376819
rect 673942 375761 673994 375767
rect 673942 375703 673994 375709
rect 675106 374551 675134 380198
rect 675202 379532 675408 379560
rect 675092 374542 675148 374551
rect 675092 374477 675148 374486
rect 675202 374107 675230 379532
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675382 378203 675434 378209
rect 675382 378145 675434 378151
rect 675394 377696 675422 378145
rect 675382 377611 675434 377617
rect 675382 377553 675434 377559
rect 675394 377075 675422 377553
rect 675478 376871 675530 376877
rect 675478 376813 675530 376819
rect 675490 376438 675518 376813
rect 675478 375761 675530 375767
rect 675478 375703 675530 375709
rect 675490 375254 675518 375703
rect 675188 374098 675244 374107
rect 675188 374033 675244 374042
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675380 372026 675436 372035
rect 675380 371961 675436 371970
rect 675394 371554 675422 371961
rect 674422 360073 674474 360079
rect 674420 360038 674422 360047
rect 674474 360038 674476 360047
rect 674420 359973 674476 359982
rect 674710 359777 674762 359783
rect 674708 359742 674710 359751
rect 674762 359742 674764 359751
rect 674708 359677 674764 359686
rect 674422 359037 674474 359043
rect 674420 359002 674422 359011
rect 674474 359002 674476 359011
rect 674420 358937 674476 358946
rect 673844 358410 673900 358419
rect 673844 358345 673900 358354
rect 674420 356338 674476 356347
rect 674420 356273 674476 356282
rect 673940 354118 673996 354127
rect 673940 354053 673996 354062
rect 673954 333587 673982 354053
rect 674324 350862 674380 350871
rect 674324 350797 674380 350806
rect 674228 349752 674284 349761
rect 674228 349687 674284 349696
rect 674036 349234 674092 349243
rect 674036 349169 674092 349178
rect 673942 333581 673994 333587
rect 673942 333523 673994 333529
rect 674050 331589 674078 349169
rect 674242 332995 674270 349687
rect 674230 332989 674282 332995
rect 674230 332931 674282 332937
rect 674338 332255 674366 350797
rect 674434 339581 674462 356273
rect 674804 355006 674860 355015
rect 674804 354941 674860 354950
rect 674612 354414 674668 354423
rect 674612 354349 674668 354358
rect 674516 352194 674572 352203
rect 674516 352129 674572 352138
rect 674422 339575 674474 339581
rect 674422 339517 674474 339523
rect 674530 337287 674558 352129
rect 674626 339803 674654 354349
rect 674708 350122 674764 350131
rect 674708 350057 674764 350066
rect 674614 339797 674666 339803
rect 674614 339739 674666 339745
rect 674518 337281 674570 337287
rect 674518 337223 674570 337229
rect 674722 335569 674750 350057
rect 674818 341653 674846 354941
rect 677012 353230 677068 353239
rect 677012 353165 677068 353174
rect 674900 352786 674956 352795
rect 674900 352721 674956 352730
rect 674806 341647 674858 341653
rect 674806 341589 674858 341595
rect 674914 341357 674942 352721
rect 674996 351750 675052 351759
rect 674996 351685 675052 351694
rect 674902 341351 674954 341357
rect 674902 341293 674954 341299
rect 675010 336492 675038 351685
rect 676820 351158 676876 351167
rect 676820 351093 676876 351102
rect 676834 345543 676862 351093
rect 676916 347754 676972 347763
rect 676916 347689 676972 347698
rect 676930 347319 676958 347689
rect 676916 347310 676972 347319
rect 676916 347245 676972 347254
rect 676820 345534 676876 345543
rect 676820 345469 676876 345478
rect 677026 345395 677054 353165
rect 677108 348346 677164 348355
rect 677108 348281 677164 348290
rect 677122 347763 677150 348281
rect 677108 347754 677164 347763
rect 677108 347689 677164 347698
rect 677122 345649 677150 347689
rect 677110 345643 677162 345649
rect 677110 345585 677162 345591
rect 677012 345386 677068 345395
rect 677012 345321 677068 345330
rect 675190 341647 675242 341653
rect 675190 341589 675242 341595
rect 675094 341351 675146 341357
rect 675094 341293 675146 341299
rect 675106 339896 675134 341293
rect 675202 340562 675230 341589
rect 675202 340534 675326 340562
rect 675298 340488 675326 340534
rect 675394 340488 675422 340548
rect 675298 340460 675422 340488
rect 675106 339868 675408 339896
rect 675094 339797 675146 339803
rect 675094 339739 675146 339745
rect 675106 337409 675134 339739
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675106 337381 675408 337409
rect 675094 337281 675146 337287
rect 675094 337223 675146 337229
rect 675106 336862 675134 337223
rect 675106 336834 675408 336862
rect 675010 336464 675422 336492
rect 675394 336182 675422 336464
rect 674722 335541 675408 335569
rect 675284 335026 675340 335035
rect 675202 334984 675284 335012
rect 674326 332249 674378 332255
rect 674326 332191 674378 332197
rect 674038 331583 674090 331589
rect 674038 331525 674090 331531
rect 675202 329559 675230 334984
rect 675340 334984 675408 335012
rect 675284 334961 675340 334970
rect 675298 334901 675326 334961
rect 675490 333851 675518 334332
rect 675476 333842 675532 333851
rect 675476 333777 675532 333786
rect 675382 333581 675434 333587
rect 675382 333523 675434 333529
rect 675394 333074 675422 333523
rect 675382 332989 675434 332995
rect 675382 332931 675434 332937
rect 675394 332519 675422 332931
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 675382 331583 675434 331589
rect 675382 331525 675434 331531
rect 675394 331224 675422 331525
rect 675764 330586 675820 330595
rect 675764 330521 675820 330530
rect 675778 330040 675806 330521
rect 675188 329550 675244 329559
rect 675188 329485 675244 329494
rect 675380 328366 675436 328375
rect 675380 328301 675436 328310
rect 675394 328190 675422 328301
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 674422 315081 674474 315087
rect 674420 315046 674422 315055
rect 674474 315046 674476 315055
rect 674420 314981 674476 314990
rect 674710 314785 674762 314791
rect 674708 314750 674710 314759
rect 674762 314750 674764 314759
rect 674708 314685 674764 314694
rect 674422 314045 674474 314051
rect 674420 314010 674422 314019
rect 674474 314010 674476 314019
rect 674420 313945 674476 313954
rect 673940 311346 673996 311355
rect 673940 311281 673996 311290
rect 673954 294589 673982 311281
rect 674708 310014 674764 310023
rect 674708 309949 674764 309958
rect 674324 309644 674380 309653
rect 674324 309579 674380 309588
rect 674036 305870 674092 305879
rect 674036 305805 674092 305814
rect 673942 294583 673994 294589
rect 673942 294525 673994 294531
rect 674050 287263 674078 305805
rect 674228 304242 674284 304251
rect 674228 304177 674284 304186
rect 674038 287257 674090 287263
rect 674038 287199 674090 287205
rect 674242 286819 674270 304177
rect 674338 292961 674366 309579
rect 674612 305130 674668 305139
rect 674612 305065 674668 305074
rect 674516 304538 674572 304547
rect 674516 304473 674572 304482
rect 674420 303650 674476 303659
rect 674420 303585 674476 303594
rect 674434 302655 674462 303585
rect 674422 302649 674474 302655
rect 674420 302614 674422 302623
rect 674474 302614 674476 302623
rect 674420 302549 674476 302558
rect 674530 300676 674558 304473
rect 674434 300648 674558 300676
rect 674326 292955 674378 292961
rect 674326 292897 674378 292903
rect 674434 287781 674462 300648
rect 674518 300577 674570 300583
rect 674518 300519 674570 300525
rect 674530 295995 674558 300519
rect 674518 295989 674570 295995
rect 674518 295931 674570 295937
rect 674626 291111 674654 305065
rect 674722 300583 674750 309949
rect 674996 308830 675052 308839
rect 674996 308765 675052 308774
rect 674900 307794 674956 307803
rect 674900 307729 674956 307738
rect 674804 306758 674860 306767
rect 674804 306693 674860 306702
rect 674710 300577 674762 300583
rect 674710 300519 674762 300525
rect 674818 291777 674846 306693
rect 674914 295403 674942 307729
rect 674902 295397 674954 295403
rect 674902 295339 674954 295345
rect 674806 291771 674858 291777
rect 674806 291713 674858 291719
rect 674614 291105 674666 291111
rect 674614 291047 674666 291053
rect 675010 288595 675038 308765
rect 677012 308238 677068 308247
rect 677012 308173 677068 308182
rect 675092 307202 675148 307211
rect 675092 307137 675148 307146
rect 675106 291870 675134 307137
rect 676916 306018 676972 306027
rect 676916 305953 676972 305962
rect 676820 302762 676876 302771
rect 676820 302697 676876 302706
rect 676834 302327 676862 302697
rect 676820 302318 676876 302327
rect 676820 302253 676876 302262
rect 676930 299515 676958 305953
rect 676916 299506 676972 299515
rect 676916 299441 676972 299450
rect 677026 299367 677054 308173
rect 677012 299358 677068 299367
rect 677012 299293 677068 299302
rect 675382 295989 675434 295995
rect 675382 295931 675434 295937
rect 675394 295523 675422 295931
rect 675478 295397 675530 295403
rect 675478 295339 675530 295345
rect 675490 294890 675518 295339
rect 675382 294583 675434 294589
rect 675382 294525 675434 294531
rect 675394 294224 675422 294525
rect 675382 292955 675434 292961
rect 675382 292897 675434 292903
rect 675394 292374 675422 292897
rect 675106 291842 675408 291870
rect 675094 291771 675146 291777
rect 675094 291713 675146 291719
rect 675106 291204 675134 291713
rect 675106 291176 675408 291204
rect 675094 291105 675146 291111
rect 675094 291047 675146 291053
rect 675106 290569 675134 291047
rect 675106 290541 675408 290569
rect 675284 290034 675340 290043
rect 675106 289992 675284 290020
rect 674998 288589 675050 288595
rect 674998 288531 675050 288537
rect 674422 287775 674474 287781
rect 674422 287717 674474 287723
rect 674230 286813 674282 286819
rect 674230 286755 674282 286761
rect 675106 284863 675134 289992
rect 675340 289992 675408 290020
rect 675284 289969 675340 289978
rect 675298 289909 675326 289969
rect 675476 289590 675532 289599
rect 675476 289525 675532 289534
rect 675298 289400 675422 289428
rect 675298 289354 675326 289400
rect 675202 289326 675326 289354
rect 675394 289354 675422 289400
rect 675490 289354 675518 289525
rect 675394 289340 675518 289354
rect 675408 289326 675504 289340
rect 675202 285011 675230 289326
rect 675478 288589 675530 288595
rect 675478 288531 675530 288537
rect 675490 288082 675518 288531
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675478 287257 675530 287263
rect 675478 287199 675530 287205
rect 675490 286898 675518 287199
rect 675382 286813 675434 286819
rect 675382 286755 675434 286761
rect 675394 286232 675422 286755
rect 675188 285002 675244 285011
rect 675188 284937 675244 284946
rect 675778 284863 675806 285048
rect 675092 284854 675148 284863
rect 675092 284789 675148 284798
rect 675764 284854 675820 284863
rect 675764 284789 675820 284798
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675764 281894 675820 281903
rect 675764 281829 675820 281838
rect 675778 281348 675806 281829
rect 673556 276418 673612 276427
rect 673612 276376 673670 276404
rect 673556 276353 673612 276362
rect 672502 270681 672554 270687
rect 672502 270623 672554 270629
rect 673846 270681 673898 270687
rect 673846 270623 673898 270629
rect 673858 270063 673886 270623
rect 673844 270054 673900 270063
rect 673844 269989 673900 269998
rect 674710 269793 674762 269799
rect 674708 269758 674710 269767
rect 674762 269758 674764 269767
rect 674708 269693 674764 269702
rect 674710 269201 674762 269207
rect 674708 269166 674710 269175
rect 674762 269166 674764 269175
rect 674708 269101 674764 269110
rect 674612 266058 674668 266067
rect 674612 265993 674668 266002
rect 674420 264652 674476 264661
rect 674420 264587 674476 264596
rect 674324 262506 674380 262515
rect 674324 262441 674380 262450
rect 674132 261322 674188 261331
rect 674132 261257 674188 261266
rect 674036 259250 674092 259259
rect 674036 259185 674092 259194
rect 674050 241605 674078 259185
rect 674038 241599 674090 241605
rect 674038 241541 674090 241547
rect 674146 240569 674174 261257
rect 674338 247081 674366 262441
rect 674434 247969 674462 264587
rect 674626 256572 674654 265993
rect 677204 265466 677260 265475
rect 677204 265401 677260 265410
rect 674900 265022 674956 265031
rect 674900 264957 674956 264966
rect 674708 261766 674764 261775
rect 674708 261701 674764 261710
rect 674530 256544 674654 256572
rect 674530 252779 674558 256544
rect 674614 256473 674666 256479
rect 674614 256415 674666 256421
rect 674626 253445 674654 256415
rect 674614 253439 674666 253445
rect 674614 253381 674666 253387
rect 674518 252773 674570 252779
rect 674518 252715 674570 252721
rect 674422 247963 674474 247969
rect 674422 247905 674474 247911
rect 674326 247075 674378 247081
rect 674326 247017 674378 247023
rect 674722 246785 674750 261701
rect 674804 260138 674860 260147
rect 674804 260073 674860 260082
rect 674710 246779 674762 246785
rect 674710 246721 674762 246727
rect 674818 246119 674846 260073
rect 674914 256479 674942 264957
rect 675188 262802 675244 262811
rect 675188 262737 675244 262746
rect 674996 259546 675052 259555
rect 674996 259481 675052 259490
rect 674902 256473 674954 256479
rect 674902 256415 674954 256421
rect 674806 246113 674858 246119
rect 674806 246055 674858 246061
rect 675010 243011 675038 259481
rect 675094 252773 675146 252779
rect 675094 252715 675146 252721
rect 675106 249246 675134 252715
rect 675202 249912 675230 262737
rect 677108 258362 677164 258371
rect 677108 258297 677164 258306
rect 676916 257770 676972 257779
rect 676916 257705 676972 257714
rect 676930 257335 676958 257705
rect 677122 257335 677150 258297
rect 676916 257326 676972 257335
rect 676916 257261 676972 257270
rect 677108 257326 677164 257335
rect 677108 257261 677164 257270
rect 677122 256405 677150 257261
rect 677110 256399 677162 256405
rect 677110 256341 677162 256347
rect 675286 253439 675338 253445
rect 675286 253381 675338 253387
rect 675298 250537 675326 253381
rect 677218 251563 677246 265401
rect 677588 263246 677644 263255
rect 677588 263181 677644 263190
rect 677602 251711 677630 263181
rect 677588 251702 677644 251711
rect 677588 251637 677644 251646
rect 677204 251554 677260 251563
rect 677204 251489 677260 251498
rect 675298 250509 675408 250537
rect 675202 249884 675326 249912
rect 675298 249764 675326 249884
rect 675394 249764 675422 249898
rect 675298 249736 675422 249764
rect 675106 249218 675408 249246
rect 675478 247963 675530 247969
rect 675478 247905 675530 247911
rect 675490 247382 675518 247905
rect 675478 247075 675530 247081
rect 675478 247017 675530 247023
rect 675490 246864 675518 247017
rect 675382 246779 675434 246785
rect 675382 246721 675434 246727
rect 675394 246198 675422 246721
rect 675382 246113 675434 246119
rect 675382 246055 675434 246061
rect 675188 245930 675244 245939
rect 675188 245865 675244 245874
rect 675202 244362 675230 245865
rect 675394 245532 675422 246055
rect 675394 244755 675422 245014
rect 675380 244746 675436 244755
rect 675380 244681 675436 244690
rect 675202 244334 675408 244362
rect 674998 243005 675050 243011
rect 674998 242947 675050 242953
rect 674134 240563 674186 240569
rect 674134 240505 674186 240511
rect 675202 238983 675230 244334
rect 675476 243562 675532 243571
rect 675476 243497 675532 243506
rect 675490 243090 675518 243497
rect 675382 243005 675434 243011
rect 675382 242947 675434 242953
rect 675394 242498 675422 242947
rect 675380 242082 675436 242091
rect 675380 242017 675436 242026
rect 675394 241875 675422 242017
rect 675478 241599 675530 241605
rect 675478 241541 675530 241547
rect 675490 241240 675518 241541
rect 675478 240563 675530 240569
rect 675478 240505 675530 240511
rect 675490 240056 675518 240505
rect 675188 238974 675244 238983
rect 675188 238909 675244 238918
rect 675764 238678 675820 238687
rect 675764 238613 675820 238622
rect 675778 238206 675806 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 674710 225097 674762 225103
rect 674708 225062 674710 225071
rect 674762 225062 674764 225071
rect 674708 224997 674764 225006
rect 669622 224357 669674 224363
rect 674422 224357 674474 224363
rect 669622 224299 669674 224305
rect 674420 224322 674422 224331
rect 674474 224322 674476 224331
rect 674420 224257 674476 224266
rect 669526 224061 669578 224067
rect 674710 224061 674762 224067
rect 669526 224003 669578 224009
rect 674708 224026 674710 224035
rect 674762 224026 674764 224035
rect 674708 223961 674764 223970
rect 674996 220918 675052 220927
rect 674996 220853 675052 220862
rect 674900 217070 674956 217079
rect 674900 217005 674956 217014
rect 674516 216478 674572 216487
rect 674516 216413 674572 216422
rect 674530 216001 674558 216413
rect 674134 215995 674186 216001
rect 674134 215937 674186 215943
rect 674518 215995 674570 216001
rect 674518 215937 674570 215943
rect 674146 201349 674174 215937
rect 674516 215442 674572 215451
rect 674516 215377 674572 215386
rect 674134 201343 674186 201349
rect 674134 201285 674186 201291
rect 674530 197057 674558 215377
rect 674804 214850 674860 214859
rect 674804 214785 674860 214794
rect 674708 214406 674764 214415
rect 674708 214341 674764 214350
rect 674612 213814 674668 213823
rect 674612 213749 674668 213758
rect 674518 197051 674570 197057
rect 674518 196993 674570 196999
rect 674626 196613 674654 213749
rect 674722 197649 674750 214341
rect 674818 200369 674846 214785
rect 674914 201664 674942 217005
rect 675010 204457 675038 220853
rect 675476 219734 675532 219743
rect 675476 219669 675532 219678
rect 675092 219290 675148 219299
rect 675092 219225 675148 219234
rect 675106 204624 675134 219225
rect 675284 217662 675340 217671
rect 675284 217597 675340 217606
rect 675298 210840 675326 217597
rect 675202 210812 675326 210840
rect 675202 204698 675230 210812
rect 675490 210692 675518 219669
rect 677108 218698 677164 218707
rect 677108 218633 677164 218642
rect 676916 216034 676972 216043
rect 676916 215969 676972 215978
rect 676820 212630 676876 212639
rect 676820 212565 676876 212574
rect 676834 212195 676862 212565
rect 676820 212186 676876 212195
rect 676820 212121 676876 212130
rect 675298 210664 675518 210692
rect 675298 205808 675326 210664
rect 676930 207459 676958 215969
rect 677012 213222 677068 213231
rect 677012 213157 677068 213166
rect 677026 212047 677054 213157
rect 677012 212038 677068 212047
rect 677012 211973 677068 211982
rect 677026 210303 677054 211973
rect 677014 210297 677066 210303
rect 677014 210239 677066 210245
rect 677122 207755 677150 218633
rect 677204 218106 677260 218115
rect 677204 218041 677260 218050
rect 677108 207746 677164 207755
rect 677108 207681 677164 207690
rect 677218 207607 677246 218041
rect 677204 207598 677260 207607
rect 677204 207533 677260 207542
rect 676916 207450 676972 207459
rect 676916 207385 676972 207394
rect 675298 205780 675518 205808
rect 675490 205350 675518 205780
rect 675202 204670 675408 204698
rect 675106 204596 675230 204624
rect 674998 204451 675050 204457
rect 674998 204393 675050 204399
rect 675202 202182 675230 204596
rect 675382 204451 675434 204457
rect 675382 204393 675434 204399
rect 675394 204018 675422 204393
rect 675298 202228 675422 202256
rect 675298 202182 675326 202228
rect 675202 202154 675326 202182
rect 675394 202168 675422 202228
rect 674914 201636 675408 201664
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674818 200341 675408 200369
rect 675380 200050 675436 200059
rect 675380 199985 675436 199994
rect 675394 199814 675422 199985
rect 675106 199800 675422 199814
rect 675106 199786 675408 199800
rect 674710 197643 674762 197649
rect 674710 197585 674762 197591
rect 674614 196607 674666 196613
rect 674614 196549 674666 196555
rect 675106 193103 675134 199786
rect 675476 199606 675532 199615
rect 675476 199541 675532 199550
rect 675490 199134 675518 199541
rect 675764 198422 675820 198431
rect 675764 198357 675820 198366
rect 675778 197876 675806 198357
rect 675382 197643 675434 197649
rect 675382 197585 675434 197591
rect 675394 197319 675422 197585
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675764 195314 675820 195323
rect 675764 195249 675820 195258
rect 675778 194842 675806 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675092 193094 675148 193103
rect 675092 193029 675148 193038
rect 675394 192992 675422 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 674612 179626 674668 179635
rect 674612 179561 674668 179570
rect 674422 179365 674474 179371
rect 674420 179330 674422 179339
rect 674474 179330 674476 179339
rect 674420 179265 674476 179274
rect 666646 178847 666698 178853
rect 674422 178847 674474 178853
rect 666646 178789 666698 178795
rect 674420 178812 674422 178821
rect 674474 178812 674476 178821
rect 674420 178747 674476 178756
rect 674626 178705 674654 179561
rect 674614 178699 674666 178705
rect 674614 178641 674666 178647
rect 675092 175926 675148 175935
rect 675092 175861 675148 175870
rect 674036 173854 674092 173863
rect 674036 173789 674092 173798
rect 673940 170598 673996 170607
rect 673940 170533 673996 170542
rect 673954 152065 673982 170533
rect 674050 153397 674078 173789
rect 674996 172078 675052 172087
rect 674996 172013 675052 172022
rect 674900 171486 674956 171495
rect 674900 171421 674956 171430
rect 674420 170154 674476 170163
rect 674420 170089 674476 170098
rect 674228 169562 674284 169571
rect 674228 169497 674284 169506
rect 674132 168970 674188 168979
rect 674132 168905 674188 168914
rect 674038 153391 674090 153397
rect 674038 153333 674090 153339
rect 673942 152059 673994 152065
rect 673942 152001 673994 152007
rect 674146 151547 674174 168905
rect 674242 152805 674270 169497
rect 674434 155369 674462 170089
rect 674708 168230 674764 168239
rect 674708 168165 674764 168174
rect 674612 167638 674668 167647
rect 674612 167573 674668 167582
rect 674626 167161 674654 167573
rect 674722 167457 674750 168165
rect 674710 167451 674762 167457
rect 674710 167393 674762 167399
rect 674710 167229 674762 167235
rect 674708 167194 674710 167203
rect 674762 167194 674764 167203
rect 674614 167155 674666 167161
rect 674708 167129 674764 167138
rect 674614 167097 674666 167103
rect 674914 156006 674942 171421
rect 675010 156672 675038 172013
rect 675106 159613 675134 175861
rect 676916 175186 676972 175195
rect 676916 175121 676972 175130
rect 675476 174742 675532 174751
rect 675476 174677 675532 174686
rect 675188 174298 675244 174307
rect 675188 174233 675244 174242
rect 675094 159607 675146 159613
rect 675094 159549 675146 159555
rect 675202 159484 675230 174233
rect 675284 172670 675340 172679
rect 675284 172605 675340 172614
rect 675298 159706 675326 172605
rect 675490 161019 675518 174677
rect 676820 173114 676876 173123
rect 676820 173049 676876 173058
rect 676834 161431 676862 173049
rect 676930 161579 676958 175121
rect 676916 161570 676972 161579
rect 676916 161505 676972 161514
rect 676820 161422 676876 161431
rect 676820 161357 676876 161366
rect 675478 161013 675530 161019
rect 675478 160955 675530 160961
rect 675478 160791 675530 160797
rect 675478 160733 675530 160739
rect 675490 160323 675518 160733
rect 675298 159678 675408 159706
rect 675286 159607 675338 159613
rect 675286 159549 675338 159555
rect 675106 159456 675230 159484
rect 675106 157190 675134 159456
rect 675298 159040 675326 159549
rect 675298 159012 675408 159040
rect 675106 157162 675326 157190
rect 675298 157116 675326 157162
rect 675490 157116 675518 157176
rect 675298 157088 675518 157116
rect 675010 156644 675326 156672
rect 675298 156524 675326 156644
rect 675394 156524 675422 156658
rect 675298 156496 675422 156524
rect 674914 155978 675408 156006
rect 674434 155341 675408 155369
rect 675284 155206 675340 155215
rect 675284 155141 675340 155150
rect 675298 154822 675326 155141
rect 675298 154794 675408 154822
rect 675476 154466 675532 154475
rect 675476 154401 675532 154410
rect 675490 154142 675518 154401
rect 675478 153391 675530 153397
rect 675478 153333 675530 153339
rect 675490 152884 675518 153333
rect 674230 152799 674282 152805
rect 674230 152741 674282 152747
rect 675382 152799 675434 152805
rect 675382 152741 675434 152747
rect 675394 152292 675422 152741
rect 675478 152059 675530 152065
rect 675478 152001 675530 152007
rect 675490 151700 675518 152001
rect 674134 151541 674186 151547
rect 674134 151483 674186 151489
rect 675382 151541 675434 151547
rect 675382 151483 675434 151489
rect 675394 151034 675422 151483
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675764 148546 675820 148555
rect 675764 148481 675820 148490
rect 675778 148000 675806 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 676916 134338 676972 134347
rect 676916 134273 676972 134282
rect 676820 133894 676876 133903
rect 676820 133829 676876 133838
rect 663766 133633 663818 133639
rect 674422 133633 674474 133639
rect 663766 133575 663818 133581
rect 674420 133598 674422 133607
rect 674474 133598 674476 133607
rect 674420 133533 674476 133542
rect 655318 132819 655370 132825
rect 655318 132761 655370 132767
rect 676834 132677 676862 133829
rect 676930 132825 676958 134273
rect 676918 132819 676970 132825
rect 676918 132761 676970 132767
rect 655126 132671 655178 132677
rect 655126 132613 655178 132619
rect 676822 132671 676874 132677
rect 676822 132613 676874 132619
rect 674420 132562 674476 132571
rect 647638 132523 647690 132529
rect 674420 132497 674422 132506
rect 647638 132465 647690 132471
rect 674474 132497 674476 132506
rect 674422 132465 674474 132471
rect 645814 126677 645866 126683
rect 645814 126619 645866 126625
rect 645908 121462 645964 121471
rect 645908 121397 645964 121406
rect 645814 121275 645866 121281
rect 645814 121217 645866 121223
rect 645826 121175 645854 121217
rect 645922 121207 645950 121397
rect 645910 121201 645962 121207
rect 645812 121166 645868 121175
rect 645910 121143 645962 121149
rect 645812 121101 645868 121110
rect 646006 121127 646058 121133
rect 646006 121069 646058 121075
rect 646018 120879 646046 121069
rect 646004 120870 646060 120879
rect 646004 120805 646060 120814
rect 647650 120435 647678 132465
rect 674516 130638 674572 130647
rect 674516 130573 674572 130582
rect 674324 129306 674380 129315
rect 674324 129241 674380 129250
rect 674228 127086 674284 127095
rect 674228 127021 674284 127030
rect 673940 125458 673996 125467
rect 673940 125393 673996 125402
rect 647636 120426 647692 120435
rect 647636 120361 647692 120370
rect 673954 106925 673982 125393
rect 674242 111883 674270 127021
rect 674338 113659 674366 129241
rect 674420 123830 674476 123839
rect 674420 123765 674476 123774
rect 674326 113653 674378 113659
rect 674326 113595 674378 113601
rect 674230 111877 674282 111883
rect 674230 111819 674282 111825
rect 673942 106919 673994 106925
rect 673942 106861 673994 106867
rect 645910 106549 645962 106555
rect 668182 106549 668234 106555
rect 645910 106491 645962 106497
rect 668180 106514 668182 106523
rect 668234 106514 668236 106523
rect 645812 88162 645868 88171
rect 645812 88097 645868 88106
rect 645826 87019 645854 88097
rect 645814 87013 645866 87019
rect 645814 86955 645866 86961
rect 645922 86945 645950 106491
rect 668180 106449 668236 106458
rect 674434 106407 674462 123765
rect 674530 114177 674558 130573
rect 677108 130046 677164 130055
rect 677108 129981 677164 129990
rect 675188 129602 675244 129611
rect 675188 129537 675244 129546
rect 675092 127382 675148 127391
rect 675092 127317 675148 127326
rect 674612 126346 674668 126355
rect 674612 126281 674668 126290
rect 674626 115232 674654 126281
rect 674804 124718 674860 124727
rect 674804 124653 674860 124662
rect 674708 121906 674764 121915
rect 674708 121841 674764 121850
rect 674722 121207 674750 121841
rect 674710 121201 674762 121207
rect 674710 121143 674762 121149
rect 674626 115204 674750 115232
rect 674518 114171 674570 114177
rect 674518 114113 674570 114119
rect 674722 111365 674750 115204
rect 674710 111359 674762 111365
rect 674710 111301 674762 111307
rect 674818 111291 674846 124653
rect 674900 124126 674956 124135
rect 674900 124061 674956 124070
rect 674806 111285 674858 111291
rect 674806 111227 674858 111233
rect 674914 107591 674942 124061
rect 675106 114492 675134 127317
rect 675202 115158 675230 129537
rect 677012 127826 677068 127835
rect 677012 127761 677068 127770
rect 676820 122942 676876 122951
rect 676820 122877 676876 122886
rect 676834 121281 676862 122877
rect 676916 122350 676972 122359
rect 676916 122285 676972 122294
rect 676822 121275 676874 121281
rect 676822 121217 676874 121223
rect 676930 121133 676958 122285
rect 676918 121127 676970 121133
rect 676918 121069 676970 121075
rect 677026 118067 677054 127761
rect 677012 118058 677068 118067
rect 677012 117993 677068 118002
rect 677122 117919 677150 129981
rect 677108 117910 677164 117919
rect 677108 117845 677164 117854
rect 675202 115130 675326 115158
rect 675298 115084 675326 115130
rect 675394 115084 675422 115144
rect 675298 115056 675422 115084
rect 675106 114464 675408 114492
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675094 113653 675146 113659
rect 675094 113595 675146 113601
rect 675106 112009 675134 113595
rect 675106 111981 675408 112009
rect 675094 111877 675146 111883
rect 675094 111819 675146 111825
rect 675106 111458 675134 111819
rect 675106 111430 675408 111458
rect 675382 111359 675434 111365
rect 675382 111301 675434 111307
rect 675094 111285 675146 111291
rect 675094 111227 675146 111233
rect 675106 110169 675134 111227
rect 675394 110778 675422 111301
rect 675106 110141 675408 110169
rect 675380 110066 675436 110075
rect 675380 110001 675436 110010
rect 675394 109594 675422 110001
rect 675476 109326 675532 109335
rect 675476 109261 675532 109270
rect 675490 108973 675518 109261
rect 675106 108959 675518 108973
rect 675106 108945 675504 108959
rect 674902 107585 674954 107591
rect 674902 107527 674954 107533
rect 675106 106555 675134 108945
rect 675380 108142 675436 108151
rect 675380 108077 675436 108086
rect 675394 107670 675422 108077
rect 675382 107585 675434 107591
rect 675382 107527 675434 107533
rect 675394 107119 675422 107527
rect 675478 106919 675530 106925
rect 675478 106861 675530 106867
rect 675094 106549 675146 106555
rect 675094 106491 675146 106497
rect 675490 106486 675518 106861
rect 674422 106401 674474 106407
rect 674422 106343 674474 106349
rect 675382 106401 675434 106407
rect 675382 106343 675434 106349
rect 675394 105820 675422 106343
rect 665300 105182 665356 105191
rect 665300 105117 665356 105126
rect 675380 105182 675436 105191
rect 675380 105117 675436 105126
rect 665204 104590 665260 104599
rect 665204 104525 665206 104534
rect 665258 104525 665260 104534
rect 665206 104493 665258 104499
rect 665314 104483 665342 105117
rect 675394 104636 675422 105117
rect 659542 104477 659594 104483
rect 659542 104419 659594 104425
rect 665302 104477 665354 104483
rect 665302 104419 665354 104425
rect 659554 93753 659582 104419
rect 675764 103258 675820 103267
rect 675764 103193 675820 103202
rect 675778 102786 675806 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 651286 93747 651338 93753
rect 651286 93689 651338 93695
rect 659542 93747 659594 93753
rect 659542 93689 659594 93695
rect 646390 92711 646442 92717
rect 646390 92653 646442 92659
rect 646198 92563 646250 92569
rect 646198 92505 646250 92511
rect 645910 86939 645962 86945
rect 645910 86881 645962 86887
rect 645812 86682 645868 86691
rect 645812 86617 645868 86626
rect 645826 86501 645854 86617
rect 645814 86495 645866 86501
rect 645814 86437 645866 86443
rect 646102 86421 646154 86427
rect 646102 86363 646154 86369
rect 645812 84166 645868 84175
rect 645812 84101 645868 84110
rect 645826 81839 645854 84101
rect 645814 81833 645866 81839
rect 645814 81775 645866 81781
rect 646004 80170 646060 80179
rect 646004 80105 646060 80114
rect 645812 79282 645868 79291
rect 645812 79217 645868 79226
rect 645826 78435 645854 79217
rect 645910 79095 645962 79101
rect 645910 79037 645962 79043
rect 645922 78551 645950 79037
rect 645908 78542 645964 78551
rect 645908 78477 645964 78486
rect 645814 78429 645866 78435
rect 645814 78371 645866 78377
rect 646018 78065 646046 80105
rect 646006 78059 646058 78065
rect 646006 78001 646058 78007
rect 645910 77023 645962 77029
rect 645910 76965 645962 76971
rect 645814 76727 645866 76733
rect 645814 76669 645866 76675
rect 645826 76035 645854 76669
rect 645812 76026 645868 76035
rect 645812 75961 645868 75970
rect 645922 75295 645950 76965
rect 645908 75286 645964 75295
rect 645908 75221 645964 75230
rect 645812 73806 645868 73815
rect 645812 73741 645868 73750
rect 645826 72367 645854 73741
rect 645814 72361 645866 72367
rect 645814 72303 645866 72309
rect 646114 66299 646142 86363
rect 646210 80919 646238 92505
rect 646196 80910 646252 80919
rect 646196 80845 646252 80854
rect 646402 72779 646430 92653
rect 647446 92637 647498 92643
rect 647446 92579 647498 92585
rect 647254 92341 647306 92347
rect 647254 92283 647306 92289
rect 646678 92193 646730 92199
rect 646678 92135 646730 92141
rect 646388 72770 646444 72779
rect 646388 72705 646444 72714
rect 646690 72187 646718 92135
rect 647266 85803 647294 92283
rect 647252 85794 647308 85803
rect 647252 85729 647308 85738
rect 647458 82251 647486 92579
rect 647830 92415 647882 92421
rect 647830 92357 647882 92363
rect 647734 92267 647786 92273
rect 647734 92209 647786 92215
rect 647540 89050 647596 89059
rect 647540 88985 647596 88994
rect 647444 82242 647500 82251
rect 647444 82177 647500 82186
rect 647554 81691 647582 88985
rect 647636 87422 647692 87431
rect 647636 87357 647692 87366
rect 647542 81685 647594 81691
rect 647542 81627 647594 81633
rect 647650 77769 647678 87357
rect 647746 85507 647774 92209
rect 647842 86247 647870 92357
rect 650614 87383 650666 87389
rect 650614 87325 650666 87331
rect 647828 86238 647884 86247
rect 647828 86173 647884 86182
rect 647732 85498 647788 85507
rect 647732 85433 647788 85442
rect 650626 83879 650654 87325
rect 650998 87013 651050 87019
rect 650900 86978 650956 86987
rect 650998 86955 651050 86961
rect 650900 86913 650956 86922
rect 650914 85243 650942 86913
rect 651010 85359 651038 86955
rect 651094 86495 651146 86501
rect 651094 86437 651146 86443
rect 650996 85350 651052 85359
rect 650996 85285 651052 85294
rect 650902 85237 650954 85243
rect 650902 85179 650954 85185
rect 650996 84314 651052 84323
rect 650996 84249 651052 84258
rect 650612 83870 650668 83879
rect 650612 83805 650668 83814
rect 650900 82686 650956 82695
rect 650900 82621 650956 82630
rect 647638 77763 647690 77769
rect 647638 77705 647690 77711
rect 650914 76733 650942 82621
rect 651010 77695 651038 84249
rect 651106 83435 651134 86437
rect 651188 86238 651244 86247
rect 651188 86173 651244 86182
rect 651092 83426 651148 83435
rect 651092 83361 651148 83370
rect 651202 79101 651230 86173
rect 651190 79095 651242 79101
rect 651190 79037 651242 79043
rect 650998 77689 651050 77695
rect 650998 77631 651050 77637
rect 650902 76727 650954 76733
rect 650902 76669 650954 76675
rect 651298 76289 651326 93689
rect 659830 92711 659882 92717
rect 659830 92653 659882 92659
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 658882 87986 658910 92135
rect 659842 88000 659870 92653
rect 661750 92637 661802 92643
rect 661750 92579 661802 92585
rect 660694 92563 660746 92569
rect 660694 92505 660746 92511
rect 659842 87972 660144 88000
rect 660706 87986 660734 92505
rect 661174 92341 661226 92347
rect 661174 92283 661226 92289
rect 661186 88000 661214 92283
rect 661762 88000 661790 92579
rect 663094 92415 663146 92421
rect 663094 92357 663146 92363
rect 662518 92267 662570 92273
rect 662518 92209 662570 92215
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 92209
rect 663106 87986 663134 92357
rect 659362 87389 659616 87408
rect 659350 87383 659616 87389
rect 659402 87380 659616 87383
rect 659350 87325 659402 87331
rect 658006 87309 658058 87315
rect 656866 87232 657792 87260
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 651286 76283 651338 76289
rect 651286 76225 651338 76231
rect 656866 75549 656894 87232
rect 657046 87161 657098 87167
rect 657046 87103 657098 87109
rect 657058 83467 657086 87103
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 663298 85211 663326 87029
rect 663476 85646 663532 85655
rect 663476 85581 663532 85590
rect 663284 85202 663340 85211
rect 663284 85137 663340 85146
rect 663380 84758 663436 84767
rect 663202 84716 663380 84744
rect 657046 83461 657098 83467
rect 657046 83403 657098 83409
rect 661078 81685 661130 81691
rect 661130 81633 661440 81636
rect 661078 81627 661440 81633
rect 661090 81608 661440 81627
rect 657538 81321 657792 81340
rect 657526 81315 657792 81321
rect 657578 81312 657792 81315
rect 657526 81257 657578 81263
rect 662900 81206 662956 81215
rect 662900 81141 662956 81150
rect 656962 81016 657216 81044
rect 656962 80211 656990 81016
rect 656950 80205 657002 80211
rect 656950 80147 657002 80153
rect 658306 76955 658334 81030
rect 658882 78953 658910 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658870 78947 658922 78953
rect 658870 78889 658922 78895
rect 659458 77769 659486 80665
rect 659446 77763 659498 77769
rect 659446 77705 659498 77711
rect 658294 76949 658346 76955
rect 658294 76891 658346 76897
rect 656854 75543 656906 75549
rect 656854 75485 656906 75491
rect 660130 72367 660158 81030
rect 660706 78065 660734 81030
rect 661762 81016 662016 81044
rect 660694 78059 660746 78065
rect 660694 78001 660746 78007
rect 661762 77029 661790 81016
rect 662530 78435 662558 81030
rect 662518 78429 662570 78435
rect 662518 78371 662570 78377
rect 662914 77325 662942 81141
rect 662902 77319 662954 77325
rect 662902 77261 662954 77267
rect 661750 77023 661802 77029
rect 661750 76965 661802 76971
rect 660118 72361 660170 72367
rect 660118 72303 660170 72309
rect 646676 72178 646732 72187
rect 663202 72145 663230 84716
rect 663380 84693 663436 84702
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663490 80600 663518 85581
rect 663394 80572 663518 80600
rect 663394 73033 663422 80572
rect 663382 73027 663434 73033
rect 663382 72969 663434 72975
rect 646676 72113 646732 72122
rect 663190 72139 663242 72145
rect 663190 72081 663242 72087
rect 646102 66293 646154 66299
rect 646102 66235 646154 66241
rect 645718 51789 645770 51795
rect 645718 51731 645770 51737
rect 645622 48977 645674 48983
rect 645622 48919 645674 48925
rect 645334 48237 645386 48243
rect 645334 48179 645386 48185
rect 623446 47571 623498 47577
rect 623446 47513 623498 47519
rect 640726 47571 640778 47577
rect 640726 47513 640778 47519
rect 529268 43318 529324 43327
rect 529268 43253 529324 43262
rect 514922 42117 515136 42120
rect 514870 42111 515136 42117
rect 514882 42092 515136 42111
rect 520354 42092 520656 42120
rect 521602 42092 521856 42120
rect 525922 42092 526176 42120
rect 529282 42106 529310 43253
rect 471092 42069 471148 42078
rect 404374 41577 404426 41583
rect 404374 41519 404426 41525
rect 388822 40319 388874 40325
rect 388822 40261 388874 40267
rect 394582 40319 394634 40325
rect 394582 40261 394634 40267
rect 142100 40210 142156 40219
rect 142100 40145 142156 40154
rect 394594 37439 394622 40261
rect 404386 37439 404414 41519
rect 443444 40654 443500 40663
rect 443444 40589 443500 40598
rect 453524 40654 453580 40663
rect 453524 40589 453580 40598
rect 443458 40367 443486 40589
rect 453538 40367 453566 40589
rect 623458 40515 623486 47513
rect 623444 40506 623500 40515
rect 623444 40441 623500 40450
rect 443444 40358 443500 40367
rect 443444 40293 443500 40302
rect 453524 40358 453580 40367
rect 453524 40293 453580 40302
rect 394582 37433 394634 37439
rect 394582 37375 394634 37381
rect 404374 37433 404426 37439
rect 404374 37375 404426 37381
<< via2 >>
rect 92276 1016658 92332 1016714
rect 81044 995790 81100 995846
rect 148532 1015918 148588 1015974
rect 353396 1015918 353452 1015974
rect 145364 1007926 145420 1007982
rect 148532 1007926 148588 1007982
rect 85940 995642 85996 995698
rect 42068 968706 42124 968762
rect 41780 967078 41836 967134
rect 42068 965006 42124 965062
rect 41780 963970 41836 964026
rect 41780 963230 41836 963286
rect 42836 963230 42892 963286
rect 41780 962638 41836 962694
rect 41876 962046 41932 962102
rect 42164 960418 42220 960474
rect 41780 959678 41836 959734
rect 41780 959086 41836 959142
rect 41780 958494 41836 958550
rect 41876 957754 41932 957810
rect 42164 955830 42220 955886
rect 40340 942954 40396 943010
rect 35156 932594 35212 932650
rect 35156 932150 35212 932206
rect 40148 927266 40204 927322
rect 39860 927118 39916 927174
rect 42434 950088 42494 950148
rect 42356 940290 42412 940346
rect 42164 938070 42220 938126
rect 41684 818782 41740 818838
rect 40340 817154 40396 817210
rect 40244 816710 40300 816766
rect 35156 806794 35212 806850
rect 35156 806350 35212 806406
rect 41780 814934 41836 814990
rect 41684 813306 41740 813362
rect 37364 802058 37420 802114
rect 41972 812714 42028 812770
rect 41876 812270 41932 812326
rect 42068 811086 42124 811142
rect 42164 810494 42220 810550
rect 42068 800430 42124 800486
rect 41972 800282 42028 800338
rect 42356 809458 42412 809514
rect 42356 799690 42412 799746
rect 42644 944878 42700 944934
rect 42644 944303 42700 944342
rect 42644 944286 42646 944303
rect 42646 944286 42698 944303
rect 42698 944286 42700 944303
rect 42834 950090 42894 950150
rect 42740 943768 42796 943824
rect 42644 942697 42646 942714
rect 42646 942697 42698 942714
rect 42698 942697 42700 942714
rect 42644 942658 42700 942697
rect 42644 942179 42646 942196
rect 42646 942179 42698 942196
rect 42698 942179 42700 942196
rect 42644 942140 42700 942179
rect 42644 932167 42700 932206
rect 42644 932150 42646 932167
rect 42646 932150 42698 932167
rect 42698 932150 42700 932167
rect 42644 819117 42646 819134
rect 42646 819117 42698 819134
rect 42698 819117 42700 819134
rect 42644 819078 42700 819117
rect 42644 818081 42646 818098
rect 42646 818081 42698 818098
rect 42698 818081 42700 818098
rect 42644 818042 42700 818081
rect 43220 817450 43276 817506
rect 42644 814342 42700 814398
rect 43028 810346 43084 810402
rect 42740 809236 42796 809292
rect 42836 808126 42892 808182
rect 42452 797618 42508 797674
rect 42452 797470 42508 797526
rect 42548 797026 42604 797082
rect 43124 808718 43180 808774
rect 42548 792586 42604 792642
rect 42356 791846 42412 791902
rect 42068 791254 42124 791310
rect 42164 791106 42220 791162
rect 42452 791698 42508 791754
rect 42452 776049 42454 776066
rect 42454 776049 42506 776066
rect 42506 776049 42508 776066
rect 42452 776010 42508 776049
rect 42836 775309 42838 775326
rect 42838 775309 42890 775326
rect 42890 775309 42892 775326
rect 42836 775270 42892 775309
rect 42836 774791 42838 774808
rect 42838 774791 42890 774808
rect 42890 774791 42892 774808
rect 42836 774752 42892 774791
rect 44564 806498 44620 806554
rect 43412 774234 43468 774290
rect 43220 773642 43276 773698
rect 43028 772014 43084 772070
rect 42068 771126 42124 771182
rect 40244 770682 40300 770738
rect 35156 763578 35212 763634
rect 35156 763134 35212 763190
rect 41684 769498 41740 769554
rect 41588 764762 41644 764818
rect 40244 760174 40300 760230
rect 41588 757362 41644 757418
rect 41876 766242 41932 766298
rect 41780 765798 41836 765854
rect 42836 770386 42892 770442
rect 42356 769054 42412 769110
rect 42164 767870 42220 767926
rect 42068 760174 42124 760230
rect 41876 757066 41932 757122
rect 42164 757066 42220 757122
rect 42932 767722 42988 767778
rect 42836 759138 42892 759194
rect 42068 754846 42124 754902
rect 43124 767130 43180 767186
rect 43028 751886 43084 751942
rect 42068 751738 42124 751794
rect 42740 751590 42796 751646
rect 41876 750998 41932 751054
rect 42164 750554 42220 750610
rect 41972 748630 42028 748686
rect 41780 747150 41836 747206
rect 43028 750258 43084 750314
rect 42836 749666 42892 749722
rect 42740 746114 42796 746170
rect 43124 746854 43180 746910
rect 42740 732685 42742 732702
rect 42742 732685 42794 732702
rect 42794 732685 42796 732702
rect 42740 732646 42796 732685
rect 42740 732093 42742 732110
rect 42742 732093 42794 732110
rect 42794 732093 42796 732110
rect 42740 732054 42796 732093
rect 42356 731797 42358 731814
rect 42358 731797 42410 731814
rect 42410 731797 42412 731814
rect 42356 731758 42412 731797
rect 43700 731018 43756 731074
rect 43412 730426 43468 730482
rect 41588 728650 41644 728706
rect 40724 724210 40780 724266
rect 35156 720362 35212 720418
rect 35156 719918 35212 719974
rect 41492 723026 41548 723082
rect 41876 727910 41932 727966
rect 41684 726874 41740 726930
rect 41588 714294 41644 714350
rect 41780 726282 41836 726338
rect 40724 714146 40780 714202
rect 41492 714146 41548 714202
rect 42356 725838 42412 725894
rect 42164 723618 42220 723674
rect 41876 713850 41932 713906
rect 42164 713850 42220 713906
rect 43028 722878 43084 722934
rect 42740 721768 42796 721824
rect 42068 711630 42124 711686
rect 43028 711630 43084 711686
rect 42740 711482 42796 711538
rect 42452 711186 42508 711242
rect 42164 709854 42220 709910
rect 43220 711334 43276 711390
rect 43028 710890 43084 710946
rect 41780 707338 41836 707394
rect 42452 707190 42508 707246
rect 42356 705118 42412 705174
rect 42164 704526 42220 704582
rect 41780 704082 41836 704138
rect 42068 700530 42124 700586
rect 43124 706450 43180 706506
rect 42452 703342 42508 703398
rect 43220 689469 43222 689486
rect 43222 689469 43274 689486
rect 43274 689469 43276 689486
rect 43220 689430 43276 689469
rect 43124 688986 43180 689042
rect 42836 688433 42838 688450
rect 42838 688433 42890 688450
rect 42890 688433 42892 688450
rect 42836 688394 42892 688433
rect 43412 687802 43468 687858
rect 42068 685434 42124 685490
rect 41876 684842 41932 684898
rect 41012 681438 41068 681494
rect 35156 677146 35212 677202
rect 35156 676702 35212 676758
rect 41780 678774 41836 678830
rect 41684 675518 41740 675574
rect 41012 670930 41068 670986
rect 41684 670930 41740 670986
rect 41972 679810 42028 679866
rect 42356 682622 42412 682678
rect 42164 680402 42220 680458
rect 42068 670634 42124 670690
rect 43220 681290 43276 681346
rect 43124 679810 43180 679866
rect 42932 670930 42988 670986
rect 43508 687654 43564 687710
rect 43700 683658 43756 683714
rect 42164 665306 42220 665362
rect 42164 664714 42220 664770
rect 43028 670634 43084 670690
rect 42644 663974 42700 664030
rect 42356 662790 42412 662846
rect 42068 662198 42124 662254
rect 41876 661014 41932 661070
rect 43028 662346 43084 662402
rect 43124 660866 43180 660922
rect 42932 646214 42988 646270
rect 42356 645474 42412 645530
rect 43220 645178 43276 645234
rect 43796 647102 43852 647158
rect 43604 646954 43660 647010
rect 43316 644438 43372 644494
rect 43988 644586 44044 644642
rect 43796 643550 43852 643606
rect 43604 642958 43660 643014
rect 43508 642070 43564 642126
rect 41780 641626 41836 641682
rect 41012 640442 41068 640498
rect 35156 633930 35212 633986
rect 35156 633486 35212 633542
rect 41588 639998 41644 640054
rect 41492 638370 41548 638426
rect 41492 627714 41548 627770
rect 41876 639406 41932 639462
rect 41972 637778 42028 637834
rect 43220 637186 43276 637242
rect 42164 636742 42220 636798
rect 42068 636150 42124 636206
rect 42356 635114 42412 635170
rect 42164 628158 42220 628214
rect 42068 627566 42124 627622
rect 41972 627418 42028 627474
rect 42644 628158 42700 628214
rect 42356 626974 42412 627030
rect 42452 624458 42508 624514
rect 42452 622090 42508 622146
rect 42356 619574 42412 619630
rect 42164 618242 42220 618298
rect 41972 617650 42028 617706
rect 42644 621498 42700 621554
rect 43316 635558 43372 635614
rect 42452 617206 42508 617262
rect 42356 616466 42412 616522
rect 42452 602850 42508 602906
rect 42356 602110 42412 602166
rect 43220 602406 43276 602462
rect 43220 601370 43276 601426
rect 43124 598706 43180 598762
rect 41588 597226 41644 597282
rect 41780 596782 41836 596838
rect 41684 594562 41740 594618
rect 41876 596190 41932 596246
rect 41972 595154 42028 595210
rect 42932 594340 42988 594396
rect 42068 593526 42124 593582
rect 41972 584202 42028 584258
rect 43028 592712 43084 592768
rect 42452 581242 42508 581298
rect 42164 578874 42220 578930
rect 41972 575914 42028 575970
rect 42068 574582 42124 574638
rect 41780 574434 41836 574490
rect 42932 576950 42988 577006
rect 42452 573102 42508 573158
rect 43124 573842 43180 573898
rect 42548 559486 42604 559542
rect 42452 559059 42508 559098
rect 42452 559042 42454 559059
rect 42454 559042 42506 559059
rect 42506 559042 42508 559059
rect 42932 558746 42988 558802
rect 43988 601222 44044 601278
rect 43796 600334 43852 600390
rect 43412 600038 43468 600094
rect 43604 600038 43660 600094
rect 43796 570290 43852 570346
rect 43796 570142 43852 570198
rect 43508 560522 43564 560578
rect 43412 558450 43468 558506
rect 43220 558006 43276 558062
rect 41684 555786 41740 555842
rect 35156 547498 35212 547554
rect 35156 547054 35212 547110
rect 41972 555194 42028 555250
rect 41780 554010 41836 554066
rect 41876 551346 41932 551402
rect 41780 549718 41836 549774
rect 41684 541282 41740 541338
rect 41780 541134 41836 541190
rect 41876 540986 41932 541042
rect 42932 553862 42988 553918
rect 42452 552974 42508 553030
rect 42068 551938 42124 551994
rect 42164 550310 42220 550366
rect 42836 549496 42892 549552
rect 43028 551124 43084 551180
rect 43028 548978 43084 549034
rect 42932 541578 42988 541634
rect 42164 540690 42220 540746
rect 42452 540690 42508 540746
rect 42452 536842 42508 536898
rect 42356 533290 42412 533346
rect 42164 532698 42220 532754
rect 42164 531810 42220 531866
rect 41780 531662 41836 531718
rect 42356 531218 42412 531274
rect 43028 535658 43084 535714
rect 42932 534326 42988 534382
rect 42932 530626 42988 530682
rect 42836 432245 42838 432262
rect 42838 432245 42890 432262
rect 42890 432245 42892 432262
rect 42836 432206 42892 432245
rect 42836 431727 42838 431744
rect 42838 431727 42890 431744
rect 42890 431727 42892 431744
rect 42836 431688 42892 431727
rect 42356 431318 42412 431374
rect 43220 430578 43276 430634
rect 42836 429581 42838 429598
rect 42838 429581 42890 429598
rect 42890 429581 42892 429598
rect 42836 429542 42892 429581
rect 42836 427914 42892 427970
rect 41876 425398 41932 425454
rect 40244 423326 40300 423382
rect 39956 422734 40012 422790
rect 35156 419922 35212 419978
rect 35156 419478 35212 419534
rect 40052 422142 40108 422198
rect 40148 421550 40204 421606
rect 42356 420514 42412 420570
rect 42356 419478 42412 419534
rect 42932 421402 42988 421458
rect 41780 406010 41836 406066
rect 41876 405122 41932 405178
rect 41780 404382 41836 404438
rect 42164 403050 42220 403106
rect 42164 402606 42220 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 42356 389325 42358 389342
rect 42358 389325 42410 389342
rect 42410 389325 42412 389342
rect 42356 389286 42412 389325
rect 42356 388733 42358 388750
rect 42358 388733 42410 388750
rect 42410 388733 42412 388750
rect 42356 388694 42412 388733
rect 42740 387993 42742 388010
rect 42742 387993 42794 388010
rect 42794 387993 42796 388010
rect 42740 387954 42796 387993
rect 43412 430134 43468 430190
rect 43604 556822 43660 556878
rect 43508 428950 43564 429006
rect 43316 387214 43372 387270
rect 43220 387066 43276 387122
rect 42164 384402 42220 384458
rect 40052 381146 40108 381202
rect 39956 380110 40012 380166
rect 39860 378926 39916 378982
rect 35156 376706 35212 376762
rect 35156 376262 35212 376318
rect 40148 380554 40204 380610
rect 40052 375078 40108 375134
rect 40244 378334 40300 378390
rect 40148 372858 40204 372914
rect 42356 382182 42412 382238
rect 42548 379518 42604 379574
rect 43124 378186 43180 378242
rect 42644 377594 42700 377650
rect 42644 376575 42700 376614
rect 42644 376558 42646 376575
rect 42646 376558 42698 376575
rect 42698 376558 42700 376575
rect 41780 362794 41836 362850
rect 42068 360870 42124 360926
rect 41972 360574 42028 360630
rect 42164 359834 42220 359890
rect 42068 359390 42124 359446
rect 41780 358650 41836 358706
rect 41780 356874 41836 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 42452 346109 42454 346126
rect 42454 346109 42506 346126
rect 42506 346109 42508 346126
rect 42452 346070 42508 346109
rect 42452 345517 42454 345534
rect 42454 345517 42506 345534
rect 42506 345517 42508 345534
rect 42452 345478 42508 345517
rect 42932 344777 42934 344794
rect 42934 344777 42986 344794
rect 42986 344777 42988 344794
rect 42932 344738 42988 344777
rect 43124 343998 43180 344054
rect 43220 343702 43276 343758
rect 42932 341482 42988 341538
rect 41876 338966 41932 339022
rect 40148 337338 40204 337394
rect 39956 336894 40012 336950
rect 39860 335118 39916 335174
rect 35156 333490 35212 333546
rect 35156 333046 35212 333102
rect 40052 336302 40108 336358
rect 40244 335710 40300 335766
rect 40148 329790 40204 329846
rect 42836 333359 42892 333398
rect 42836 333342 42838 333359
rect 42838 333342 42890 333359
rect 42890 333342 42892 333359
rect 42356 326534 42412 326590
rect 43028 334970 43084 335026
rect 42452 320910 42508 320966
rect 41780 319726 41836 319782
rect 41972 318690 42028 318746
rect 41972 317802 42028 317858
rect 42068 316618 42124 316674
rect 42068 316026 42124 316082
rect 41780 315434 41836 315490
rect 41876 313658 41932 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 42548 302893 42550 302910
rect 42550 302893 42602 302910
rect 42602 302893 42604 302910
rect 42548 302854 42604 302893
rect 42548 302301 42550 302318
rect 42550 302301 42602 302318
rect 42602 302301 42604 302318
rect 42548 302262 42604 302301
rect 42548 301857 42550 301874
rect 42550 301857 42602 301874
rect 42602 301857 42604 301874
rect 42548 301818 42604 301857
rect 43316 300930 43372 300986
rect 43220 300486 43276 300542
rect 41204 297970 41260 298026
rect 40244 294122 40300 294178
rect 40148 293678 40204 293734
rect 39860 292494 39916 292550
rect 35156 290422 35212 290478
rect 35156 289830 35212 289886
rect 40052 292050 40108 292106
rect 40244 285094 40300 285150
rect 41972 295750 42028 295806
rect 42932 291754 42988 291810
rect 42548 289847 42604 289886
rect 42548 289830 42550 289847
rect 42550 289830 42602 289847
rect 42602 289830 42604 289847
rect 42164 277990 42220 278046
rect 41780 276510 41836 276566
rect 41972 275474 42028 275530
rect 42164 274734 42220 274790
rect 43124 274734 43180 274790
rect 41780 273550 41836 273606
rect 42068 272958 42124 273014
rect 41780 272218 41836 272274
rect 41780 270590 41836 270646
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 42452 259677 42454 259694
rect 42454 259677 42506 259694
rect 42506 259677 42508 259694
rect 42452 259638 42508 259677
rect 42836 258937 42838 258954
rect 42838 258937 42890 258954
rect 42890 258937 42892 258954
rect 42836 258898 42892 258937
rect 42452 258641 42454 258658
rect 42454 258641 42506 258658
rect 42506 258641 42508 258658
rect 42452 258602 42508 258641
rect 42452 257418 42508 257474
rect 42164 255938 42220 255994
rect 41876 252534 41932 252590
rect 40148 250906 40204 250962
rect 39956 249870 40012 249926
rect 39860 249278 39916 249334
rect 35156 247206 35212 247262
rect 35156 246762 35212 246818
rect 40052 248834 40108 248890
rect 40244 250462 40300 250518
rect 40148 244838 40204 244894
rect 42068 248242 42124 248298
rect 43028 255050 43084 255106
rect 42452 246762 42508 246818
rect 42164 242470 42220 242526
rect 42068 242026 42124 242082
rect 42452 242026 42508 242082
rect 42548 238326 42604 238382
rect 43220 257566 43276 257622
rect 43124 243802 43180 243858
rect 42068 234034 42124 234090
rect 41780 233294 41836 233350
rect 41780 231666 41836 231722
rect 41972 231074 42028 231130
rect 41780 230334 41836 230390
rect 41780 229742 41836 229798
rect 41780 229002 41836 229058
rect 41780 227226 41836 227282
rect 41780 226634 41836 226690
rect 41780 225894 41836 225950
rect 42452 216461 42454 216478
rect 42454 216461 42506 216478
rect 42506 216461 42508 216478
rect 42452 216422 42508 216461
rect 42836 215721 42838 215738
rect 42838 215721 42890 215738
rect 42890 215721 42892 215738
rect 42836 215682 42892 215721
rect 42836 215203 42838 215220
rect 42838 215203 42890 215220
rect 42890 215203 42892 215220
rect 42836 215164 42892 215203
rect 47444 941622 47500 941678
rect 44564 246170 44620 246226
rect 43220 214054 43276 214110
rect 43508 242470 43564 242526
rect 43412 213610 43468 213666
rect 43316 213018 43372 213074
rect 42452 211686 42508 211742
rect 42068 209466 42124 209522
rect 40052 207246 40108 207302
rect 39956 206062 40012 206118
rect 35156 203990 35212 204046
rect 35156 203546 35212 203602
rect 40148 206654 40204 206710
rect 40244 205618 40300 205674
rect 41121 197767 41181 197827
rect 42452 204451 42508 204490
rect 42452 204434 42454 204451
rect 42454 204434 42506 204451
rect 42506 204434 42508 204451
rect 42452 203990 42508 204046
rect 43028 205322 43084 205378
rect 42164 190966 42220 191022
rect 41780 190078 41836 190134
rect 41780 189042 41836 189098
rect 41972 188302 42028 188358
rect 44852 547350 44908 547406
rect 46196 256678 46252 256734
rect 59444 975366 59500 975422
rect 53300 763282 53356 763338
rect 53396 720066 53452 720122
rect 53300 247650 53356 247706
rect 53588 676850 53644 676906
rect 85364 995346 85420 995402
rect 86420 995198 86476 995254
rect 87764 995050 87820 995106
rect 88724 993866 88780 993922
rect 84500 993718 84556 993774
rect 106292 999381 106294 999398
rect 106294 999381 106346 999398
rect 106346 999381 106348 999398
rect 106292 999342 106348 999381
rect 99572 995938 99628 995994
rect 102932 995955 102988 995994
rect 102932 995938 102934 995955
rect 102934 995938 102986 995955
rect 102986 995938 102988 995955
rect 94964 995790 95020 995846
rect 62036 963230 62092 963286
rect 61844 961898 61900 961954
rect 59540 960862 59596 960918
rect 59540 946654 59596 946710
rect 59540 932150 59596 932206
rect 59540 917794 59596 917850
rect 59540 903438 59596 903494
rect 59540 889082 59596 889138
rect 59540 874726 59596 874782
rect 58580 860370 58636 860426
rect 59540 846014 59596 846070
rect 59540 831658 59596 831714
rect 59540 817302 59596 817358
rect 59540 802798 59596 802854
rect 59540 788590 59596 788646
rect 59540 774086 59596 774142
rect 59540 759730 59596 759786
rect 59540 745522 59596 745578
rect 59540 731018 59596 731074
rect 59540 716662 59596 716718
rect 59540 702306 59596 702362
rect 59540 687950 59596 688006
rect 59540 673594 59596 673650
rect 59540 659238 59596 659294
rect 59540 644882 59596 644938
rect 56084 633930 56140 633986
rect 53780 590566 53836 590622
rect 59540 630526 59596 630582
rect 59540 616170 59596 616226
rect 59540 601853 59542 601870
rect 59542 601853 59594 601870
rect 59594 601853 59596 601870
rect 59540 601814 59596 601853
rect 58772 587458 58828 587514
rect 59540 572954 59596 573010
rect 59540 558911 59596 558950
rect 59540 558894 59542 558911
rect 59542 558894 59594 558911
rect 59594 558894 59596 558911
rect 59540 544390 59596 544446
rect 59540 530034 59596 530090
rect 59540 515678 59596 515734
rect 59540 501191 59596 501230
rect 59540 501174 59542 501191
rect 59542 501174 59594 501191
rect 59594 501174 59596 501191
rect 58580 486818 58636 486874
rect 59540 472462 59596 472518
rect 59540 458106 59596 458162
rect 59540 443750 59596 443806
rect 59540 429394 59596 429450
rect 58388 415038 58444 415094
rect 58388 400682 58444 400738
rect 59252 386326 59308 386382
rect 59540 371822 59596 371878
rect 59540 357614 59596 357670
rect 58388 343110 58444 343166
rect 57812 328754 57868 328810
rect 58004 314546 58060 314602
rect 59444 300042 59500 300098
rect 58100 285834 58156 285890
rect 53588 246466 53644 246522
rect 97940 995807 97996 995846
rect 97940 995790 97942 995807
rect 97942 995790 97994 995807
rect 97994 995790 97996 995807
rect 98996 995659 99052 995698
rect 98996 995642 98998 995659
rect 98998 995642 99050 995659
rect 99050 995642 99052 995659
rect 97844 995494 97900 995550
rect 93812 995346 93868 995402
rect 102452 995790 102508 995846
rect 104468 995790 104524 995846
rect 99572 995198 99628 995254
rect 97844 994902 97900 994958
rect 108980 995977 108982 995994
rect 108982 995977 109034 995994
rect 109034 995977 109036 995994
rect 108980 995938 109036 995977
rect 109556 995938 109612 995994
rect 107924 995790 107980 995846
rect 107540 995494 107596 995550
rect 105908 995346 105964 995402
rect 105332 995198 105388 995254
rect 104468 993718 104524 993774
rect 106964 995198 107020 995254
rect 109172 995494 109228 995550
rect 109364 995050 109420 995106
rect 126644 995790 126700 995846
rect 134324 995790 134380 995846
rect 110228 995198 110284 995254
rect 131828 994162 131884 994218
rect 133652 994458 133708 994514
rect 132788 994310 132844 994366
rect 136148 995790 136204 995846
rect 139220 995494 139276 995550
rect 135188 994014 135244 994070
rect 140372 993718 140428 993774
rect 144116 995790 144172 995846
rect 144692 995346 144748 995402
rect 144692 994310 144748 994366
rect 349652 1007778 349708 1007834
rect 353300 1007778 353356 1007834
rect 299156 1005854 299212 1005910
rect 302996 1005854 303052 1005910
rect 160436 1003207 160492 1003246
rect 160436 1003190 160438 1003207
rect 160438 1003190 160490 1003207
rect 160490 1003190 160492 1003207
rect 161492 1003153 161548 1003209
rect 151124 1002467 151180 1002506
rect 151124 1002450 151126 1002467
rect 151126 1002450 151178 1002467
rect 151178 1002450 151180 1002467
rect 152756 1002341 152758 1002358
rect 152758 1002341 152810 1002358
rect 152810 1002341 152812 1002358
rect 152756 1002302 152812 1002341
rect 157652 1000839 157708 1000878
rect 157652 1000822 157654 1000839
rect 157654 1000822 157706 1000839
rect 157706 1000822 157708 1000839
rect 155540 999507 155596 999546
rect 155540 999490 155542 999507
rect 155542 999490 155594 999507
rect 155594 999490 155596 999507
rect 156020 996547 156076 996586
rect 156020 996530 156022 996547
rect 156022 996530 156074 996547
rect 156074 996530 156076 996547
rect 159188 996103 159244 996142
rect 159188 996086 159190 996103
rect 159190 996086 159242 996103
rect 159242 996086 159244 996103
rect 159764 996125 159766 996142
rect 159766 996125 159818 996142
rect 159818 996125 159820 996142
rect 159764 996086 159820 996125
rect 152084 995955 152140 995994
rect 152084 995938 152086 995955
rect 152086 995938 152138 995955
rect 152138 995938 152140 995955
rect 160436 995977 160438 995994
rect 160438 995977 160490 995994
rect 160490 995977 160492 995994
rect 160436 995938 160492 995977
rect 151700 995790 151756 995846
rect 154868 995807 154924 995846
rect 154868 995790 154870 995807
rect 154870 995790 154922 995807
rect 154922 995790 154924 995807
rect 146804 994458 146860 994514
rect 146900 994310 146956 994366
rect 146900 994014 146956 994070
rect 158228 995790 158284 995846
rect 161492 995790 161548 995846
rect 154772 995346 154828 995402
rect 149684 995198 149740 995254
rect 157268 995198 157324 995254
rect 154772 994162 154828 994218
rect 161684 995198 161740 995254
rect 213812 1005114 213868 1005170
rect 218804 1005153 218806 1005170
rect 218806 1005153 218858 1005170
rect 218858 1005153 218860 1005170
rect 218804 1005114 218860 1005153
rect 211796 1003207 211852 1003246
rect 211796 1003190 211798 1003207
rect 211798 1003190 211850 1003207
rect 211850 1003190 211852 1003207
rect 209108 1000839 209164 1000878
rect 209108 1000822 209110 1000839
rect 209110 1000822 209162 1000839
rect 209162 1000822 209164 1000839
rect 188756 995790 188812 995846
rect 189428 995790 189484 995846
rect 206900 999381 206902 999398
rect 206902 999381 206954 999398
rect 206954 999381 206956 999398
rect 206900 999342 206956 999381
rect 205268 996547 205324 996586
rect 205268 996530 205270 996547
rect 205270 996530 205322 996547
rect 205322 996530 205324 996547
rect 188084 995494 188140 995550
rect 190580 995346 190636 995402
rect 185780 994310 185836 994366
rect 187316 994310 187372 994366
rect 204020 996125 204022 996142
rect 204022 996125 204074 996142
rect 204074 996125 204076 996142
rect 204020 996086 204076 996125
rect 210164 996103 210220 996142
rect 210164 996086 210166 996103
rect 210166 996086 210218 996103
rect 210218 996086 210220 996103
rect 253844 1002319 253900 1002358
rect 253844 1002302 253846 1002319
rect 253846 1002302 253898 1002319
rect 253898 1002302 253900 1002319
rect 255476 1002341 255478 1002358
rect 255478 1002341 255530 1002358
rect 255530 1002341 255532 1002358
rect 255476 1002302 255532 1002341
rect 198644 995938 198700 995994
rect 207380 995938 207436 995994
rect 210644 995977 210646 995994
rect 210646 995977 210698 995994
rect 210698 995977 210700 995994
rect 210644 995938 210700 995977
rect 211796 995955 211852 995994
rect 211796 995938 211798 995955
rect 211798 995938 211850 995955
rect 211850 995938 211852 995955
rect 198644 995829 198646 995846
rect 198646 995829 198698 995846
rect 198698 995829 198700 995846
rect 198644 995790 198700 995829
rect 202484 995829 202486 995846
rect 202486 995829 202538 995846
rect 202538 995829 202540 995846
rect 202484 995790 202540 995829
rect 202964 995790 203020 995846
rect 205652 995807 205708 995846
rect 205652 995790 205654 995807
rect 205654 995790 205706 995807
rect 205706 995790 205708 995807
rect 197204 995642 197260 995698
rect 191540 994014 191596 994070
rect 198452 995494 198508 995550
rect 198644 995533 198646 995550
rect 198646 995533 198698 995550
rect 198698 995533 198700 995550
rect 198644 995494 198700 995533
rect 198644 995198 198700 995254
rect 219092 995938 219148 995994
rect 213332 995790 213388 995846
rect 208148 995198 208204 995254
rect 208724 995198 208780 995254
rect 209780 995198 209836 995254
rect 207380 994310 207436 994366
rect 216020 995642 216076 995698
rect 243188 995790 243244 995846
rect 243956 995790 244012 995846
rect 258836 999655 258892 999694
rect 258836 999638 258838 999655
rect 258838 999638 258890 999655
rect 258890 999638 258892 999655
rect 241844 995642 241900 995698
rect 232532 994310 232588 994366
rect 236468 995494 236524 995550
rect 246932 995938 246988 995994
rect 246836 995790 246892 995846
rect 238964 995346 239020 995402
rect 237524 994162 237580 994218
rect 258356 999529 258358 999546
rect 258358 999529 258410 999546
rect 258410 999529 258412 999546
rect 258356 999490 258412 999529
rect 260468 999507 260524 999546
rect 260468 999490 260470 999507
rect 260470 999490 260522 999507
rect 260522 999490 260524 999507
rect 259988 996547 260044 996586
rect 259988 996530 259990 996547
rect 259990 996530 260042 996547
rect 260042 996530 260044 996547
rect 247028 995346 247084 995402
rect 262100 996234 262156 996290
rect 262004 996103 262060 996142
rect 263060 996125 263062 996142
rect 263062 996125 263114 996142
rect 263114 996125 263116 996142
rect 262004 996086 262006 996103
rect 262006 996086 262058 996103
rect 262058 996086 262060 996103
rect 263060 996086 263116 996125
rect 254516 995938 254572 995994
rect 257684 995938 257740 995994
rect 263252 995977 263254 995994
rect 263254 995977 263306 995994
rect 263306 995977 263308 995994
rect 263252 995938 263308 995977
rect 256148 995790 256204 995846
rect 259412 995790 259468 995846
rect 270740 995790 270796 995846
rect 247604 995681 247606 995698
rect 247606 995681 247658 995698
rect 247658 995681 247660 995698
rect 247604 995642 247660 995681
rect 247796 995642 247852 995698
rect 247604 995346 247660 995402
rect 250484 995198 250540 995254
rect 267956 995642 268012 995698
rect 267860 995494 267916 995550
rect 298162 997468 298222 997528
rect 280244 997122 280300 997178
rect 298100 997139 298156 997178
rect 298100 997122 298102 997139
rect 298102 997122 298154 997139
rect 298154 997122 298156 997139
rect 298164 996680 298224 996740
rect 290516 995790 290572 995846
rect 288020 994606 288076 994662
rect 286004 994458 286060 994514
rect 288020 994162 288076 994218
rect 292532 995642 292588 995698
rect 298388 995790 298444 995846
rect 293588 995494 293644 995550
rect 288980 994606 289036 994662
rect 316436 1003190 316492 1003246
rect 308852 1002911 308908 1002950
rect 308852 1002894 308854 1002911
rect 308854 1002894 308906 1002911
rect 308906 1002894 308908 1002911
rect 308276 1002763 308332 1002802
rect 308276 1002746 308278 1002763
rect 308278 1002746 308330 1002763
rect 308330 1002746 308332 1002763
rect 309332 1002785 309334 1002802
rect 309334 1002785 309386 1002802
rect 309386 1002785 309388 1002802
rect 309332 1002746 309388 1002785
rect 310484 999507 310540 999546
rect 310484 999490 310486 999507
rect 310486 999490 310538 999507
rect 310538 999490 310540 999507
rect 312116 999529 312118 999546
rect 312118 999529 312170 999546
rect 312170 999529 312172 999546
rect 312116 999490 312172 999529
rect 309908 999381 309910 999398
rect 309910 999381 309962 999398
rect 309962 999381 309964 999398
rect 309908 999342 309964 999381
rect 304340 999233 304342 999250
rect 304342 999233 304394 999250
rect 304394 999233 304396 999250
rect 304340 999194 304396 999233
rect 304916 999233 304918 999250
rect 304918 999233 304970 999250
rect 304970 999233 304972 999250
rect 304916 999194 304972 999233
rect 314804 997731 314860 997770
rect 314804 997714 314806 997731
rect 314806 997714 314858 997731
rect 314858 997714 314860 997731
rect 313748 997139 313804 997178
rect 313748 997122 313750 997139
rect 313750 997122 313802 997139
rect 313802 997122 313804 997139
rect 313172 996103 313228 996142
rect 313172 996086 313174 996103
rect 313174 996086 313226 996103
rect 313226 996086 313228 996103
rect 314804 996125 314806 996142
rect 314806 996125 314858 996142
rect 314858 996125 314860 996142
rect 314804 996086 314860 996125
rect 303956 995938 304012 995994
rect 304340 995938 304396 995994
rect 311540 995938 311596 995994
rect 319604 995938 319660 995994
rect 306068 995807 306124 995846
rect 306068 995790 306070 995807
rect 306070 995790 306122 995807
rect 306122 995790 306124 995807
rect 306548 995790 306604 995846
rect 306452 995681 306454 995698
rect 306454 995681 306506 995698
rect 306506 995681 306508 995698
rect 306452 995642 306508 995681
rect 308084 994606 308140 994662
rect 308084 994310 308140 994366
rect 294548 994162 294604 994218
rect 312788 995346 312844 995402
rect 319700 995642 319756 995698
rect 359060 1003207 359116 1003246
rect 359060 1003190 359062 1003207
rect 359062 1003190 359114 1003207
rect 359114 1003190 359116 1003207
rect 362516 1003207 362572 1003246
rect 362516 1003190 362518 1003207
rect 362518 1003190 362570 1003207
rect 362570 1003190 362572 1003207
rect 361268 1002615 361324 1002654
rect 361268 1002598 361270 1002615
rect 361270 1002598 361322 1002615
rect 361322 1002598 361324 1002615
rect 361844 1002489 361846 1002506
rect 361846 1002489 361898 1002506
rect 361898 1002489 361900 1002506
rect 361844 1002450 361900 1002489
rect 362900 1002319 362956 1002358
rect 362900 1002302 362902 1002319
rect 362902 1002302 362954 1002319
rect 362954 1002302 362956 1002319
rect 363476 1002341 363478 1002358
rect 363478 1002341 363530 1002358
rect 363530 1002341 363532 1002358
rect 363476 1002302 363532 1002341
rect 356372 1000861 356374 1000878
rect 356374 1000861 356426 1000878
rect 356426 1000861 356428 1000878
rect 356372 1000822 356428 1000861
rect 360212 1000839 360268 1000878
rect 360212 1000822 360214 1000839
rect 360214 1000822 360266 1000839
rect 360266 1000822 360268 1000839
rect 357044 999342 357100 999398
rect 364532 999211 364588 999250
rect 364532 999194 364534 999211
rect 364534 999194 364586 999211
rect 364586 999194 364588 999211
rect 365204 997731 365260 997770
rect 365204 997714 365206 997731
rect 365206 997714 365258 997731
rect 365258 997714 365260 997731
rect 363956 995977 363958 995994
rect 363958 995977 364010 995994
rect 364010 995977 364012 995994
rect 363956 995938 364012 995977
rect 358100 995790 358156 995846
rect 366164 995790 366220 995846
rect 366740 995807 366796 995846
rect 366740 995790 366742 995807
rect 366742 995790 366794 995807
rect 366794 995790 366796 995807
rect 358196 995642 358252 995698
rect 371540 995790 371596 995846
rect 368660 995642 368716 995698
rect 365780 995494 365836 995550
rect 358484 994754 358540 994810
rect 358100 994458 358156 994514
rect 362900 993313 362902 993330
rect 362902 993313 362954 993330
rect 362954 993313 362956 993330
rect 362900 993274 362956 993313
rect 383060 995790 383116 995846
rect 377204 995642 377260 995698
rect 426068 1003207 426124 1003246
rect 426068 1003190 426070 1003207
rect 426070 1003190 426122 1003207
rect 426122 1003190 426124 1003207
rect 429236 1003207 429292 1003246
rect 429236 1003190 429238 1003207
rect 429238 1003190 429290 1003207
rect 429290 1003190 429292 1003207
rect 425396 1003059 425452 1003098
rect 425396 1003042 425398 1003059
rect 425398 1003042 425450 1003059
rect 425450 1003042 425452 1003059
rect 430292 1003059 430348 1003098
rect 430292 1003042 430294 1003059
rect 430294 1003042 430346 1003059
rect 430346 1003042 430348 1003059
rect 424340 1002933 424342 1002950
rect 424342 1002933 424394 1002950
rect 424394 1002933 424396 1002950
rect 424340 1002894 424396 1002933
rect 428756 1002911 428812 1002950
rect 428756 1002894 428758 1002911
rect 428758 1002894 428810 1002911
rect 428810 1002894 428812 1002911
rect 423764 1002763 423820 1002802
rect 423764 1002746 423766 1002763
rect 423766 1002746 423818 1002763
rect 423818 1002746 423820 1002763
rect 428276 1002785 428278 1002802
rect 428278 1002785 428330 1002802
rect 428330 1002785 428332 1002802
rect 428276 1002746 428332 1002785
rect 424820 1002637 424822 1002654
rect 424822 1002637 424874 1002654
rect 424874 1002637 424876 1002654
rect 424820 1002598 424876 1002637
rect 427700 1002615 427756 1002654
rect 427700 1002598 427702 1002615
rect 427702 1002598 427754 1002615
rect 427754 1002598 427756 1002615
rect 426644 1002489 426646 1002506
rect 426646 1002489 426698 1002506
rect 426698 1002489 426700 1002506
rect 426644 1002450 426700 1002489
rect 427124 1002467 427180 1002506
rect 427124 1002450 427126 1002467
rect 427126 1002450 427178 1002467
rect 427178 1002450 427180 1002467
rect 435188 1005854 435244 1005910
rect 465716 1005854 465772 1005910
rect 435092 1005114 435148 1005170
rect 431924 1002341 431926 1002358
rect 431926 1002341 431978 1002358
rect 431978 1002341 431980 1002358
rect 431924 1002302 431980 1002341
rect 429908 1000861 429910 1000878
rect 429910 1000861 429962 1000878
rect 429962 1000861 429964 1000878
rect 429908 1000822 429964 1000861
rect 430964 1000839 431020 1000878
rect 430964 1000822 430966 1000839
rect 430966 1000822 431018 1000839
rect 431018 1000822 431020 1000839
rect 432596 996251 432652 996290
rect 432596 996234 432598 996251
rect 432598 996234 432650 996251
rect 432650 996234 432652 996251
rect 432500 996125 432502 996142
rect 432502 996125 432554 996142
rect 432554 996125 432556 996142
rect 432500 996086 432556 996125
rect 443540 1005114 443596 1005170
rect 430964 995977 430966 995994
rect 430966 995977 431018 995994
rect 431018 995977 431020 995994
rect 430964 995938 431020 995977
rect 437876 995938 437932 995994
rect 393716 995790 393772 995846
rect 422132 995790 422188 995846
rect 387476 995642 387532 995698
rect 377108 995050 377164 995106
rect 382964 993313 382966 993330
rect 382966 993313 383018 993330
rect 383018 993313 383020 993330
rect 388340 994902 388396 994958
rect 389396 994754 389452 994810
rect 391124 995346 391180 995402
rect 390836 994310 390892 994366
rect 395156 994606 395212 994662
rect 393044 994458 393100 994514
rect 396980 995050 397036 995106
rect 396308 994310 396364 994366
rect 382964 993274 383020 993313
rect 437780 995642 437836 995698
rect 423380 993587 423436 993626
rect 423380 993570 423382 993587
rect 423382 993570 423434 993587
rect 423434 993570 423436 993587
rect 437972 995494 438028 995550
rect 463700 996086 463756 996142
rect 463796 995642 463852 995698
rect 465332 995494 465388 995550
rect 467828 995938 467884 995994
rect 501332 1003059 501388 1003098
rect 501332 1003042 501334 1003059
rect 501334 1003042 501386 1003059
rect 501386 1003042 501388 1003059
rect 502388 1003081 502390 1003098
rect 502390 1003081 502442 1003098
rect 502442 1003081 502444 1003098
rect 502388 1003042 502444 1003081
rect 502964 1003081 502966 1003098
rect 502966 1003081 503018 1003098
rect 503018 1003081 503020 1003098
rect 502964 1003042 503020 1003081
rect 504020 1003059 504076 1003098
rect 504020 1003042 504022 1003059
rect 504022 1003042 504074 1003059
rect 504074 1003042 504076 1003059
rect 503444 1002341 503446 1002358
rect 503446 1002341 503498 1002358
rect 503498 1002341 503500 1002358
rect 503444 1002302 503500 1002341
rect 472244 995790 472300 995846
rect 476468 995790 476524 995846
rect 481460 995790 481516 995846
rect 482036 995790 482092 995846
rect 477716 995642 477772 995698
rect 482708 995642 482764 995698
rect 478100 995198 478156 995254
rect 472148 995050 472204 995106
rect 467060 994902 467116 994958
rect 464756 994754 464812 994810
rect 478100 994606 478156 994662
rect 481076 995050 481132 995106
rect 484148 994902 484204 994958
rect 479828 994606 479884 994662
rect 485972 994754 486028 994810
rect 485588 994458 485644 994514
rect 443444 993570 443500 993626
rect 506228 1001453 506230 1001470
rect 506230 1001453 506282 1001470
rect 506282 1001453 506284 1001470
rect 506228 1001414 506284 1001453
rect 507860 1000987 507916 1001026
rect 507860 1000970 507862 1000987
rect 507862 1000970 507914 1000987
rect 507914 1000970 507916 1000987
rect 512660 1000987 512716 1001026
rect 512660 1000970 512662 1000987
rect 512662 1000970 512714 1000987
rect 512714 1000970 512716 1000987
rect 500756 1000839 500812 1000878
rect 500756 1000822 500758 1000839
rect 500758 1000822 500810 1000839
rect 500810 1000822 500812 1000839
rect 514004 1000822 514060 1000878
rect 506900 1000691 506956 1000730
rect 506900 1000674 506902 1000691
rect 506902 1000674 506954 1000691
rect 506954 1000674 506956 1000691
rect 512084 1000691 512140 1000730
rect 512084 1000674 512086 1000691
rect 512086 1000674 512138 1000691
rect 512138 1000674 512140 1000691
rect 518420 999786 518476 999842
rect 502004 999677 502006 999694
rect 502006 999677 502058 999694
rect 502058 999677 502060 999694
rect 502004 999638 502060 999677
rect 512084 999677 512086 999694
rect 512086 999677 512138 999694
rect 512138 999677 512140 999694
rect 512084 999638 512140 999677
rect 504692 999529 504694 999546
rect 504694 999529 504746 999546
rect 504746 999529 504748 999546
rect 504692 999490 504748 999529
rect 512084 999529 512086 999546
rect 512086 999529 512138 999546
rect 512138 999529 512140 999546
rect 512084 999490 512140 999529
rect 500180 999381 500182 999398
rect 500182 999381 500234 999398
rect 500234 999381 500236 999398
rect 500180 999342 500236 999381
rect 505652 996547 505708 996586
rect 505652 996530 505654 996547
rect 505654 996530 505706 996547
rect 505706 996530 505708 996547
rect 507284 996569 507286 996586
rect 507286 996569 507338 996586
rect 507338 996569 507340 996586
rect 507284 996530 507340 996569
rect 508340 996251 508396 996290
rect 508340 996234 508342 996251
rect 508342 996234 508394 996251
rect 508394 996234 508396 996251
rect 508532 996103 508588 996142
rect 508532 996086 508534 996103
rect 508534 996086 508586 996103
rect 508586 996086 508588 996103
rect 509588 996125 509590 996142
rect 509590 996125 509642 996142
rect 509642 996125 509644 996142
rect 509588 996086 509644 996125
rect 510548 995955 510604 995994
rect 510548 995938 510550 995955
rect 510550 995938 510602 995955
rect 510602 995938 510604 995955
rect 515540 995938 515596 995994
rect 511124 995807 511180 995846
rect 511124 995790 511126 995807
rect 511126 995790 511178 995807
rect 511178 995790 511180 995807
rect 518516 999342 518572 999398
rect 518420 995642 518476 995698
rect 554900 1002933 554902 1002950
rect 554902 1002933 554954 1002950
rect 554954 1002933 554956 1002950
rect 554900 1002894 554956 1002933
rect 554324 1002785 554326 1002802
rect 554326 1002785 554378 1002802
rect 554378 1002785 554380 1002802
rect 554324 1002746 554380 1002785
rect 553748 1002615 553804 1002654
rect 553748 1002598 553750 1002615
rect 553750 1002598 553802 1002615
rect 553802 1002598 553804 1002615
rect 553268 1002341 553270 1002358
rect 553270 1002341 553322 1002358
rect 553322 1002341 553324 1002358
rect 553268 1002302 553324 1002341
rect 555380 1002319 555436 1002358
rect 555380 1002302 555382 1002319
rect 555382 1002302 555434 1002319
rect 555434 1002302 555436 1002319
rect 557780 1001305 557782 1001322
rect 557782 1001305 557834 1001322
rect 557834 1001305 557836 1001322
rect 557780 1001266 557836 1001305
rect 523796 1000970 523852 1001026
rect 523508 1000822 523564 1000878
rect 521204 995790 521260 995846
rect 521300 995494 521356 995550
rect 523700 999638 523756 999694
rect 523604 999342 523660 999398
rect 523508 995642 523564 995698
rect 552308 1000861 552310 1000878
rect 552310 1000861 552362 1000878
rect 552362 1000861 552364 1000878
rect 552308 1000822 552364 1000861
rect 552884 1000822 552940 1000878
rect 523988 1000674 524044 1000730
rect 523892 999786 523948 999842
rect 524084 999490 524140 999546
rect 557204 999085 557206 999102
rect 557206 999085 557258 999102
rect 557258 999085 557260 999102
rect 557204 999046 557260 999085
rect 558836 998937 558838 998954
rect 558838 998937 558890 998954
rect 558890 998937 558892 998954
rect 558836 998898 558892 998937
rect 555956 997731 556012 997770
rect 555956 997714 555958 997731
rect 555958 997714 556010 997731
rect 556010 997714 556012 997731
rect 558164 997435 558220 997474
rect 558164 997418 558166 997435
rect 558166 997418 558218 997435
rect 558218 997418 558220 997435
rect 559412 997309 559414 997326
rect 559414 997309 559466 997326
rect 559466 997309 559468 997326
rect 559412 997270 559468 997309
rect 561044 996125 561046 996142
rect 561046 996125 561098 996142
rect 561098 996125 561100 996142
rect 561044 996086 561100 996125
rect 529076 995642 529132 995698
rect 532244 995790 532300 995846
rect 550484 995790 550540 995846
rect 559796 995807 559852 995846
rect 559796 995790 559798 995807
rect 559798 995790 559850 995807
rect 559850 995790 559852 995807
rect 561908 995955 561964 995994
rect 561908 995938 561910 995955
rect 561910 995938 561962 995955
rect 561962 995938 561964 995955
rect 555380 995642 555436 995698
rect 560180 995659 560236 995698
rect 560180 995642 560182 995659
rect 560182 995642 560234 995659
rect 560234 995642 560236 995659
rect 524084 994645 524086 994662
rect 524086 994645 524138 994662
rect 524138 994645 524140 994662
rect 524084 994606 524140 994645
rect 536756 994606 536812 994662
rect 550484 995494 550540 995550
rect 561620 995346 561676 995402
rect 569684 995642 569740 995698
rect 565844 995494 565900 995550
rect 569876 995790 569932 995846
rect 573044 995494 573100 995550
rect 573236 995198 573292 995254
rect 573812 995642 573868 995698
rect 634004 995642 634060 995698
rect 630932 995494 630988 995550
rect 575156 995346 575212 995402
rect 573524 995050 573580 995106
rect 572948 994902 573004 994958
rect 572852 994754 572908 994810
rect 604628 994310 604684 994366
rect 576308 993866 576364 993922
rect 634580 995346 634636 995402
rect 636116 995198 636172 995254
rect 635252 994902 635308 994958
rect 637364 994754 637420 994810
rect 634292 994606 634348 994662
rect 639188 995050 639244 995106
rect 638516 993866 638572 993922
rect 642260 993866 642316 993922
rect 641108 993718 641164 993774
rect 204500 278434 204556 278490
rect 70580 272662 70636 272718
rect 69428 272366 69484 272422
rect 71732 272070 71788 272126
rect 65108 246318 65164 246374
rect 60500 246061 60502 246078
rect 60502 246061 60554 246078
rect 60554 246061 60556 246078
rect 60500 246022 60556 246061
rect 66260 246061 66262 246078
rect 66262 246061 66314 246078
rect 66314 246061 66316 246078
rect 66260 246022 66316 246061
rect 74900 273106 74956 273162
rect 74900 272366 74956 272422
rect 74132 272218 74188 272274
rect 76340 272662 76396 272718
rect 76532 272662 76588 272718
rect 76340 271626 76396 271682
rect 72980 271330 73036 271386
rect 78932 272810 78988 272866
rect 77780 270886 77836 270942
rect 81332 272958 81388 273014
rect 83636 273550 83692 273606
rect 86036 273254 86092 273310
rect 82580 271182 82636 271238
rect 88436 273402 88492 273458
rect 90836 271922 90892 271978
rect 94868 273106 94924 273162
rect 94772 272514 94828 272570
rect 93236 271774 93292 271830
rect 94868 272366 94924 272422
rect 94772 271626 94828 271682
rect 87188 271034 87244 271090
rect 96788 271626 96844 271682
rect 100820 271643 100876 271682
rect 100820 271626 100822 271643
rect 100822 271626 100874 271643
rect 100874 271626 100876 271643
rect 100724 271478 100780 271534
rect 114644 276658 114700 276714
rect 115220 273106 115276 273162
rect 115316 272514 115372 272570
rect 115220 272366 115276 272422
rect 115316 270738 115372 270794
rect 120788 271643 120844 271682
rect 120788 271626 120790 271643
rect 120790 271626 120842 271643
rect 120842 271626 120844 271643
rect 120980 271665 120982 271682
rect 120982 271665 121034 271682
rect 121034 271665 121036 271682
rect 120980 271626 121036 271665
rect 135284 273106 135340 273162
rect 135284 272366 135340 272422
rect 141044 271665 141046 271682
rect 141046 271665 141098 271682
rect 141098 271665 141100 271682
rect 141044 271626 141100 271665
rect 141332 271665 141334 271682
rect 141334 271665 141386 271682
rect 141386 271665 141388 271682
rect 141332 271626 141388 271665
rect 141140 271517 141142 271534
rect 141142 271517 141194 271534
rect 141194 271517 141196 271534
rect 141140 271478 141196 271517
rect 141620 271517 141622 271534
rect 141622 271517 141674 271534
rect 141674 271517 141676 271534
rect 141620 271478 141676 271517
rect 141140 271330 141196 271386
rect 141620 271330 141676 271386
rect 146132 240546 146188 240602
rect 144116 238622 144172 238678
rect 142484 237586 142540 237642
rect 144020 236254 144076 236310
rect 144020 233590 144076 233646
rect 144116 232110 144172 232166
rect 144020 231370 144076 231426
rect 144212 230186 144268 230242
rect 144116 228410 144172 228466
rect 144020 227818 144076 227874
rect 144404 223674 144460 223730
rect 144404 220122 144460 220178
rect 144212 215238 144268 215294
rect 145364 210502 145420 210558
rect 144980 203250 145036 203306
rect 145076 198958 145132 199014
rect 144596 196590 144652 196646
rect 144404 194814 144460 194870
rect 42932 188302 42988 188358
rect 41780 187118 41836 187174
rect 41780 186378 41836 186434
rect 41780 185786 41836 185842
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 144020 181790 144076 181846
rect 144116 176758 144172 176814
rect 144212 163586 144268 163642
rect 144020 159886 144076 159942
rect 144116 158110 144172 158166
rect 144308 155594 144364 155650
rect 144308 144346 144364 144402
rect 144308 142422 144364 142478
rect 144308 141255 144364 141294
rect 144308 141238 144310 141255
rect 144310 141238 144362 141255
rect 144362 141238 144364 141255
rect 144308 139462 144364 139518
rect 144308 137538 144364 137594
rect 144308 134726 144364 134782
rect 144308 132802 144364 132858
rect 144308 129990 144364 130046
rect 144308 129250 144364 129306
rect 39860 125293 39862 125310
rect 39862 125293 39914 125310
rect 39914 125293 39916 125310
rect 39860 125254 39916 125293
rect 141044 104090 141100 104146
rect 141044 103794 141100 103850
rect 144308 126734 144364 126790
rect 144500 183270 144556 183326
rect 144500 151598 144556 151654
rect 144500 145974 144556 146030
rect 144500 143162 144556 143218
rect 144500 133986 144556 134042
rect 144500 131026 144556 131082
rect 144404 125106 144460 125162
rect 144308 124514 144364 124570
rect 144308 124366 144364 124422
rect 144404 122590 144460 122646
rect 144308 121554 144364 121610
rect 144404 119038 144460 119094
rect 144308 118189 144310 118206
rect 144310 118189 144362 118206
rect 144362 118189 144364 118206
rect 144308 118150 144364 118189
rect 144308 116670 144364 116726
rect 144308 115930 144364 115986
rect 144404 114154 144460 114210
rect 144308 113266 144364 113322
rect 144308 113118 144364 113174
rect 144308 112417 144310 112434
rect 144310 112417 144362 112434
rect 144362 112417 144364 112434
rect 144308 112378 144364 112417
rect 144404 111194 144460 111250
rect 144308 109714 144364 109770
rect 144308 107494 144364 107550
rect 144404 106754 144460 106810
rect 144212 87810 144268 87866
rect 144116 87070 144172 87126
rect 144020 75121 144022 75138
rect 144022 75121 144074 75138
rect 144074 75121 144076 75138
rect 144020 75082 144076 75121
rect 144020 69754 144076 69810
rect 144020 56473 144022 56490
rect 144022 56473 144074 56490
rect 144074 56473 144076 56490
rect 144020 56434 144076 56473
rect 144404 77450 144460 77506
rect 144404 72714 144460 72770
rect 144980 174390 145036 174446
rect 144788 173354 144844 173410
rect 144788 168322 144844 168378
rect 144788 166546 144844 166602
rect 144884 162846 144940 162902
rect 144980 161366 145036 161422
rect 144884 159294 144940 159350
rect 144884 156334 144940 156390
rect 144788 154410 144844 154466
rect 144884 152930 144940 152986
rect 144884 150858 144940 150914
rect 144788 149674 144844 149730
rect 144692 146862 144748 146918
rect 144884 147898 144940 147954
rect 144596 120814 144652 120870
rect 144596 108234 144652 108290
rect 144596 80706 144652 80762
rect 144788 54675 144844 54714
rect 144788 54658 144790 54675
rect 144790 54658 144842 54675
rect 144842 54658 144844 54675
rect 144500 54105 144502 54122
rect 144502 54105 144554 54122
rect 144554 54105 144556 54122
rect 144500 54066 144556 54105
rect 145268 179718 145324 179774
rect 145268 172022 145324 172078
rect 145172 164770 145228 164826
rect 145076 106606 145132 106662
rect 145076 84110 145132 84166
rect 145460 207986 145516 208042
rect 145556 205618 145612 205674
rect 145748 205026 145804 205082
rect 145652 201326 145708 201382
rect 145844 193630 145900 193686
rect 145940 190078 145996 190134
rect 145844 69014 145900 69070
rect 146036 189338 146092 189394
rect 146612 239806 146668 239862
rect 149588 245726 149644 245782
rect 146324 236846 146380 236902
rect 146228 185194 146284 185250
rect 146132 99798 146188 99854
rect 146132 89586 146188 89642
rect 146132 83518 146188 83574
rect 146516 235070 146572 235126
rect 146420 186378 146476 186434
rect 146324 144790 146380 144846
rect 146324 138278 146380 138334
rect 146324 104682 146380 104738
rect 146324 102758 146380 102814
rect 146324 99058 146380 99114
rect 146324 96246 146380 96302
rect 146324 94322 146380 94378
rect 146324 91362 146380 91418
rect 146324 79374 146380 79430
rect 146324 75674 146380 75730
rect 146804 226634 146860 226690
rect 146804 225006 146860 225062
rect 146804 222934 146860 222990
rect 146708 221750 146764 221806
rect 146804 218198 146860 218254
rect 146804 213314 146860 213370
rect 146804 211686 146860 211742
rect 146708 209762 146764 209818
rect 146804 207411 146860 207450
rect 146804 207394 146806 207411
rect 146806 207394 146858 207411
rect 146858 207394 146860 207411
rect 146804 202066 146860 202122
rect 146804 199550 146860 199606
rect 146804 197774 146860 197830
rect 146708 192890 146764 192946
rect 146804 191706 146860 191762
rect 146804 188154 146860 188210
rect 146804 184454 146860 184510
rect 146612 180458 146668 180514
rect 146516 127622 146572 127678
rect 146516 106475 146572 106514
rect 146516 106458 146518 106475
rect 146518 106458 146570 106475
rect 146570 106458 146572 106475
rect 146516 104090 146572 104146
rect 146516 101591 146572 101630
rect 146516 101574 146518 101591
rect 146518 101574 146570 101591
rect 146570 101574 146572 101591
rect 146516 98061 146518 98078
rect 146518 98061 146570 98078
rect 146570 98061 146572 98078
rect 146516 98022 146572 98061
rect 146516 95506 146572 95562
rect 146516 92694 146572 92750
rect 146516 90770 146572 90826
rect 146516 85886 146572 85942
rect 146516 82334 146572 82390
rect 146516 78634 146572 78690
rect 146804 178573 146806 178590
rect 146806 178573 146858 178590
rect 146858 178573 146860 178590
rect 146804 178534 146860 178573
rect 146804 176018 146860 176074
rect 146804 171282 146860 171338
rect 146708 170098 146764 170154
rect 146804 167582 146860 167638
rect 146708 73898 146764 73954
rect 146708 70955 146764 70994
rect 146708 70938 146710 70955
rect 146710 70938 146762 70955
rect 146762 70938 146764 70955
rect 146708 67403 146764 67442
rect 146708 67386 146710 67403
rect 146710 67386 146762 67403
rect 146762 67386 146764 67403
rect 146900 136058 146956 136114
rect 146996 126899 147052 126938
rect 146996 126882 146998 126899
rect 146998 126882 147050 126899
rect 147050 126882 147052 126899
rect 146804 66350 146860 66406
rect 146708 65462 146764 65518
rect 146804 64761 146806 64778
rect 146806 64761 146858 64778
rect 146858 64761 146860 64778
rect 146804 64722 146860 64761
rect 146804 62519 146860 62558
rect 146804 62502 146806 62519
rect 146806 62502 146858 62519
rect 146858 62502 146860 62519
rect 146900 62354 146956 62410
rect 146900 60726 146956 60782
rect 146804 59581 146806 59598
rect 146806 59581 146858 59598
rect 146858 59581 146860 59598
rect 146804 59542 146860 59581
rect 146804 58654 146860 58710
rect 146804 57065 146806 57082
rect 146806 57065 146858 57082
rect 146858 57065 146860 57082
rect 146804 57026 146860 57065
rect 155348 245430 155404 245486
rect 156884 273106 156940 273162
rect 156980 272514 157036 272570
rect 156884 272366 156940 272422
rect 156980 270738 157036 270794
rect 160820 271774 160876 271830
rect 161204 271774 161260 271830
rect 161108 271665 161110 271682
rect 161110 271665 161162 271682
rect 161162 271665 161164 271682
rect 161108 271626 161164 271665
rect 158324 245134 158380 245190
rect 161108 244986 161164 245042
rect 157748 237734 157804 237790
rect 163988 247206 164044 247262
rect 166868 244838 166924 244894
rect 177044 273106 177100 273162
rect 177140 272514 177196 272570
rect 177044 272366 177100 272422
rect 177140 270738 177196 270794
rect 175508 247502 175564 247558
rect 172724 246614 172780 246670
rect 168404 48738 168460 48794
rect 171284 48590 171340 48646
rect 178388 243506 178444 243562
rect 174164 48442 174220 48498
rect 165524 48146 165580 48202
rect 181268 247354 181324 247410
rect 181460 247206 181516 247262
rect 187028 246022 187084 246078
rect 190004 247058 190060 247114
rect 187700 246466 187756 246522
rect 187700 245578 187756 245634
rect 198740 273698 198796 273754
rect 197204 273106 197260 273162
rect 197396 272514 197452 272570
rect 197204 272366 197260 272422
rect 196340 270590 196396 270646
rect 197396 270738 197452 270794
rect 263732 278434 263788 278490
rect 196820 247650 196876 247706
rect 197204 247206 197260 247262
rect 197588 246170 197644 246226
rect 197204 246022 197260 246078
rect 196820 242174 196876 242230
rect 193652 66202 193708 66258
rect 196052 219382 196108 219438
rect 194420 90030 194476 90086
rect 194708 98614 194764 98670
rect 195476 93730 195532 93786
rect 194804 92250 194860 92306
rect 196052 83518 196108 83574
rect 194516 78634 194572 78690
rect 196916 75230 196972 75286
rect 195476 68866 195532 68922
rect 196244 68274 196300 68330
rect 195476 63407 195532 63446
rect 195476 63390 195478 63407
rect 195478 63390 195530 63407
rect 195530 63390 195532 63407
rect 195476 60726 195532 60782
rect 199700 223970 199756 224026
rect 198836 221158 198892 221214
rect 197300 90622 197356 90678
rect 198356 100390 198412 100446
rect 197876 86774 197932 86830
rect 197780 85738 197836 85794
rect 198740 84702 198796 84758
rect 197396 79226 197452 79282
rect 198548 65610 198604 65666
rect 198356 59098 198412 59154
rect 201716 223378 201772 223434
rect 201620 222786 201676 222842
rect 201812 221750 201868 221806
rect 201716 220122 201772 220178
rect 201620 219530 201676 219586
rect 200660 218494 200716 218550
rect 201716 217902 201772 217958
rect 201620 216866 201676 216922
rect 201716 215238 201772 215294
rect 200180 91214 200236 91270
rect 201716 99354 201772 99410
rect 200564 97765 200566 97782
rect 200566 97765 200618 97782
rect 200618 97765 200620 97782
rect 200564 97726 200620 97765
rect 201044 97134 201100 97190
rect 200756 96098 200812 96154
rect 201716 95506 201772 95562
rect 201716 94470 201772 94526
rect 201620 92842 201676 92898
rect 201716 89586 201772 89642
rect 201332 88402 201388 88458
rect 201716 88994 201772 89050
rect 201620 87958 201676 88014
rect 201812 87366 201868 87422
rect 201620 86330 201676 86386
rect 201716 85146 201772 85202
rect 201812 84110 201868 84166
rect 201716 83074 201772 83130
rect 201620 82482 201676 82538
rect 201716 81890 201772 81946
rect 201812 81446 201868 81502
rect 201524 80854 201580 80910
rect 200276 80114 200332 80170
rect 200276 75970 200332 76026
rect 201716 77598 201772 77654
rect 201716 77006 201772 77062
rect 201620 75378 201676 75434
rect 201716 74342 201772 74398
rect 201620 73750 201676 73806
rect 201812 72714 201868 72770
rect 201524 72122 201580 72178
rect 201716 71086 201772 71142
rect 201620 70494 201676 70550
rect 200372 69902 200428 69958
rect 201812 69458 201868 69514
rect 201716 67830 201772 67886
rect 201620 67238 201676 67294
rect 201812 66646 201868 66702
rect 201716 65018 201772 65074
rect 201716 64574 201772 64630
rect 201812 63982 201868 64038
rect 201716 62946 201772 63002
rect 201620 62354 201676 62410
rect 201524 61762 201580 61818
rect 201812 61318 201868 61374
rect 201716 60134 201772 60190
rect 204692 232110 204748 232166
rect 204788 231518 204844 231574
rect 204884 230926 204940 230982
rect 204596 228262 204652 228318
rect 204500 227670 204556 227726
rect 205076 232702 205132 232758
rect 204980 225006 205036 225062
rect 205172 226634 205228 226690
rect 205460 230482 205516 230538
rect 205364 226042 205420 226098
rect 205652 227226 205708 227282
rect 205556 225598 205612 225654
rect 203060 93878 203116 93934
rect 204596 102018 204652 102074
rect 204692 101574 204748 101630
rect 204500 100982 204556 101038
rect 204596 98762 204652 98818
rect 203156 80262 203212 80318
rect 206036 229298 206092 229354
rect 205940 214498 205996 214554
rect 211700 271182 211756 271238
rect 211508 268666 211564 268722
rect 211124 268074 211180 268130
rect 211028 267778 211084 267834
rect 207188 261266 207244 261322
rect 206996 249278 207052 249334
rect 206612 243358 206668 243414
rect 206420 214646 206476 214702
rect 206324 213610 206380 213666
rect 206324 213018 206380 213074
rect 206132 212722 206188 212778
rect 206804 224414 206860 224470
rect 206708 216274 206764 216330
rect 206612 211982 206668 212038
rect 207092 229742 207148 229798
rect 206996 222342 207052 222398
rect 206900 211390 206956 211446
rect 205748 202658 205804 202714
rect 207188 97874 207244 97930
rect 206996 57470 207052 57526
rect 206900 55842 206956 55898
rect 202964 48294 203020 48350
rect 209876 247058 209932 247114
rect 209780 246318 209836 246374
rect 209972 246762 210028 246818
rect 210260 246762 210316 246818
rect 209972 245578 210028 245634
rect 210548 245430 210604 245486
rect 210260 245134 210316 245190
rect 210068 245003 210124 245042
rect 210068 244986 210070 245003
rect 210070 244986 210122 245003
rect 210122 244986 210124 245003
rect 210068 244855 210124 244894
rect 210068 244838 210070 244855
rect 210070 244838 210122 244855
rect 210122 244838 210124 244855
rect 209972 243654 210028 243710
rect 210644 243210 210700 243266
rect 209780 243062 209836 243118
rect 209396 239066 209452 239122
rect 209588 237586 209644 237642
rect 207956 232110 208012 232166
rect 208052 97874 208108 97930
rect 209300 231518 209356 231574
rect 209204 202658 209260 202714
rect 209492 230482 209548 230538
rect 209492 62798 209548 62854
rect 209684 236698 209740 236754
rect 210836 245765 210838 245782
rect 210838 245765 210890 245782
rect 210890 245765 210892 245782
rect 210836 245726 210892 245765
rect 210164 234774 210220 234830
rect 210066 233751 210126 233811
rect 209972 71643 209974 71660
rect 209974 71643 210026 71660
rect 210026 71643 210028 71660
rect 209972 71604 210028 71643
rect 209972 59616 210028 59672
rect 209972 56360 210028 56416
rect 210164 228854 210220 228910
rect 210164 220640 210220 220696
rect 210164 217384 210220 217440
rect 210164 215756 210220 215812
rect 210164 205026 210220 205082
rect 210164 164178 210220 164234
rect 210164 125106 210220 125162
rect 210164 121258 210220 121314
rect 210164 99872 210220 99928
rect 210164 96616 210220 96672
rect 210164 94988 210220 95044
rect 210164 91732 210220 91788
rect 210164 78116 210220 78172
rect 210164 76488 210220 76544
rect 210164 73232 210220 73288
rect 211028 246466 211084 246522
rect 211028 243654 211084 243710
rect 211508 267778 211564 267834
rect 211124 241878 211180 241934
rect 211604 247058 211660 247114
rect 211604 246614 211660 246670
rect 212084 271034 212140 271090
rect 217364 273106 217420 273162
rect 217460 272514 217516 272570
rect 217364 272366 217420 272422
rect 217460 270738 217516 270794
rect 221780 271626 221836 271682
rect 221780 271182 221836 271238
rect 241556 271478 241612 271534
rect 242036 271478 242092 271534
rect 241652 271330 241708 271386
rect 241940 271330 241996 271386
rect 246164 271626 246220 271682
rect 246164 271182 246220 271238
rect 250676 274142 250732 274198
rect 250292 268518 250348 268574
rect 251828 274290 251884 274346
rect 252404 274438 252460 274494
rect 252020 268814 252076 268870
rect 254132 274734 254188 274790
rect 253940 274586 253996 274642
rect 253364 270442 253420 270498
rect 252884 268962 252940 269018
rect 256820 273846 256876 273902
rect 254612 267926 254668 267982
rect 259604 273106 259660 273162
rect 257396 268666 257452 268722
rect 257300 268074 257356 268130
rect 259316 271034 259372 271090
rect 258932 268370 258988 268426
rect 261620 275622 261676 275678
rect 260660 270738 260716 270794
rect 260564 269110 260620 269166
rect 261332 268518 261388 268574
rect 261140 268222 261196 268278
rect 261332 268222 261388 268278
rect 262004 267778 262060 267834
rect 262868 274882 262924 274938
rect 262196 271626 262252 271682
rect 263348 273994 263404 274050
rect 264404 275474 264460 275530
rect 265940 275326 265996 275382
rect 265460 271182 265516 271238
rect 264884 269702 264940 269758
rect 265076 268666 265132 268722
rect 266612 269554 266668 269610
rect 267092 275178 267148 275234
rect 267188 275030 267244 275086
rect 267668 269406 267724 269462
rect 267380 267778 267436 267834
rect 268148 269258 268204 269314
rect 267764 267778 267820 267834
rect 268052 267778 268108 267834
rect 268244 267778 268300 267834
rect 269204 269850 269260 269906
rect 273524 271034 273580 271090
rect 277844 268666 277900 268722
rect 277652 268074 277708 268130
rect 277844 268074 277900 268130
rect 280820 269110 280876 269166
rect 280820 268666 280876 268722
rect 282164 271626 282220 271682
rect 282260 268962 282316 269018
rect 288020 269998 288076 270054
rect 288308 268666 288364 268722
rect 288020 268370 288076 268426
rect 288308 268370 288364 268426
rect 287540 267778 287596 267834
rect 288500 267778 288556 267834
rect 291860 268666 291916 268722
rect 291860 268074 291916 268130
rect 303380 278286 303436 278342
rect 296756 271034 296812 271090
rect 296660 269110 296716 269166
rect 304532 278138 304588 278194
rect 305204 277842 305260 277898
rect 304916 270146 304972 270202
rect 307124 277694 307180 277750
rect 308372 277546 308428 277602
rect 308084 269998 308140 270054
rect 308084 268370 308140 268426
rect 309524 277398 309580 277454
rect 309428 276954 309484 277010
rect 309620 276806 309676 276862
rect 310964 277250 311020 277306
rect 312404 277102 312460 277158
rect 312116 267795 312172 267834
rect 312116 267778 312118 267795
rect 312118 267778 312170 267795
rect 312170 267778 312172 267795
rect 315092 276510 315148 276566
rect 312692 268074 312748 268130
rect 315092 270886 315148 270942
rect 315572 270294 315628 270350
rect 315572 268666 315628 268722
rect 315764 268666 315820 268722
rect 316532 271330 316588 271386
rect 316724 271330 316780 271386
rect 316628 271034 316684 271090
rect 317108 277990 317164 278046
rect 316532 269998 316588 270054
rect 316724 269850 316780 269906
rect 373172 278582 373228 278638
rect 373364 278582 373420 278638
rect 318356 276954 318412 277010
rect 318452 276806 318508 276862
rect 318644 276362 318700 276418
rect 317108 270590 317164 270646
rect 317108 270146 317164 270202
rect 317492 270886 317548 270942
rect 317972 270590 318028 270646
rect 317972 270294 318028 270350
rect 317588 268962 317644 269018
rect 317588 268074 317644 268130
rect 317780 268962 317836 269018
rect 318164 270294 318220 270350
rect 319604 276214 319660 276270
rect 319508 271034 319564 271090
rect 319412 270146 319468 270202
rect 319508 269998 319564 270054
rect 321428 276954 321484 277010
rect 320852 276066 320908 276122
rect 319700 269998 319756 270054
rect 320180 269850 320236 269906
rect 322100 276658 322156 276714
rect 322388 271034 322444 271090
rect 322580 271034 322636 271090
rect 323924 275918 323980 275974
rect 325076 276806 325132 276862
rect 325556 276658 325612 276714
rect 327860 267795 327916 267834
rect 327860 267778 327862 267795
rect 327862 267778 327914 267795
rect 327914 267778 327916 267795
rect 328532 275770 328588 275826
rect 328532 271330 328588 271386
rect 328628 270886 328684 270942
rect 328436 269998 328492 270054
rect 328628 269998 328684 270054
rect 332276 271034 332332 271090
rect 334100 271330 334156 271386
rect 334100 269110 334156 269166
rect 336212 268074 336268 268130
rect 336404 268091 336460 268130
rect 336404 268074 336406 268091
rect 336406 268074 336458 268091
rect 336458 268074 336460 268091
rect 336980 268113 336982 268130
rect 336982 268113 337034 268130
rect 337034 268113 337036 268130
rect 336980 268074 337036 268113
rect 338516 270294 338572 270350
rect 338036 269998 338092 270054
rect 347252 269110 347308 269166
rect 347540 269110 347596 269166
rect 348020 269110 348076 269166
rect 348596 268370 348652 268426
rect 267570 264862 267630 264922
rect 349172 272514 349228 272570
rect 349460 272366 349516 272422
rect 357044 271330 357100 271386
rect 358292 272366 358348 272422
rect 358484 272366 358540 272422
rect 358484 272070 358540 272126
rect 358676 272070 358732 272126
rect 367124 271221 367126 271238
rect 367126 271221 367178 271238
rect 367178 271221 367180 271238
rect 367124 271182 367180 271221
rect 367124 271034 367180 271090
rect 367124 269110 367180 269166
rect 368660 271330 368716 271386
rect 368564 270886 368620 270942
rect 369236 274882 369292 274938
rect 368468 270607 368524 270646
rect 368468 270590 368470 270607
rect 368470 270590 368522 270607
rect 368522 270590 368524 270607
rect 369428 270590 369484 270646
rect 368756 269110 368812 269166
rect 369812 270590 369868 270646
rect 370004 270590 370060 270646
rect 373364 276510 373420 276566
rect 373940 276510 373996 276566
rect 374324 273550 374380 273606
rect 374132 273402 374188 273458
rect 374708 273254 374764 273310
rect 374708 272662 374764 272718
rect 375188 272070 375244 272126
rect 374324 270886 374380 270942
rect 374900 271922 374956 271978
rect 376532 272958 376588 273014
rect 375668 272514 375724 272570
rect 376532 272218 376588 272274
rect 377492 274882 377548 274938
rect 377300 273402 377356 273458
rect 377300 272958 377356 273014
rect 377492 273402 377548 273458
rect 377300 271182 377356 271238
rect 376916 269110 376972 269166
rect 377108 269110 377164 269166
rect 376820 267778 376876 267834
rect 377204 267926 377260 267982
rect 384020 278582 384076 278638
rect 377684 273402 377740 273458
rect 377012 267778 377068 267834
rect 379028 274882 379084 274938
rect 379412 274882 379468 274938
rect 378260 273846 378316 273902
rect 378452 273846 378508 273902
rect 378260 273402 378316 273458
rect 378164 272070 378220 272126
rect 378164 271182 378220 271238
rect 379028 272070 379084 272126
rect 377972 267817 377974 267834
rect 377974 267817 378026 267834
rect 378026 267817 378028 267834
rect 377972 267778 378028 267817
rect 378164 268370 378220 268426
rect 379220 269110 379276 269166
rect 378740 267778 378796 267834
rect 379316 267778 379372 267834
rect 379604 272514 379660 272570
rect 379988 274882 380044 274938
rect 380180 274882 380236 274938
rect 380084 272958 380140 273014
rect 380276 272958 380332 273014
rect 380180 272514 380236 272570
rect 380276 272070 380332 272126
rect 380084 269110 380140 269166
rect 381140 272810 381196 272866
rect 381332 272810 381388 272866
rect 382964 273994 383020 274050
rect 383156 273994 383212 274050
rect 382772 273550 382828 273606
rect 382964 273550 383020 273606
rect 383060 272810 383116 272866
rect 382292 272662 382348 272718
rect 381812 272218 381868 272274
rect 381620 271922 381676 271978
rect 381812 271922 381868 271978
rect 383060 272218 383116 272274
rect 383828 273254 383884 273310
rect 383444 267778 383500 267834
rect 384884 272810 384940 272866
rect 384116 272366 384172 272422
rect 384404 271922 384460 271978
rect 385364 272662 385420 272718
rect 387860 276510 387916 276566
rect 385940 272810 385996 272866
rect 386612 272810 386668 272866
rect 386324 271922 386380 271978
rect 387764 271182 387820 271238
rect 598484 278434 598540 278490
rect 467540 278286 467596 278342
rect 474740 278138 474796 278194
rect 488948 277990 489004 278046
rect 388340 273254 388396 273310
rect 388148 271774 388204 271830
rect 388628 273994 388684 274050
rect 389108 271774 389164 271830
rect 388628 268370 388684 268426
rect 388820 268370 388876 268426
rect 389300 271626 389356 271682
rect 389204 268370 389260 268426
rect 389684 271626 389740 271682
rect 389396 268370 389452 268426
rect 389876 271478 389932 271534
rect 391412 273698 391468 273754
rect 390836 273254 390892 273310
rect 390932 272366 390988 272422
rect 397364 273550 397420 273606
rect 392852 273402 392908 273458
rect 393140 273402 393196 273458
rect 391604 270886 391660 270942
rect 392948 270886 393004 270942
rect 388979 264909 389039 264913
rect 394484 272958 394540 273014
rect 395636 272958 395692 273014
rect 394292 272514 394348 272570
rect 395636 272662 395692 272718
rect 395828 272662 395884 272718
rect 394004 272366 394060 272422
rect 394484 272070 394540 272126
rect 395156 271478 395212 271534
rect 394484 271034 394540 271090
rect 394388 270738 394444 270794
rect 395444 267926 395500 267982
rect 396308 271922 396364 271978
rect 396884 271182 396940 271238
rect 397748 271034 397804 271090
rect 397556 267943 397612 267982
rect 397556 267926 397558 267943
rect 397558 267926 397610 267943
rect 397610 267926 397612 267943
rect 397844 267778 397900 267834
rect 398420 272366 398476 272422
rect 399476 270886 399532 270942
rect 400148 272218 400204 272274
rect 401204 270738 401260 270794
rect 402740 272070 402796 272126
rect 401876 271922 401932 271978
rect 401684 267926 401740 267982
rect 403700 268370 403756 268426
rect 403892 268370 403948 268426
rect 404756 267926 404812 267982
rect 406676 271922 406732 271978
rect 405620 267926 405676 267982
rect 406100 268370 406156 268426
rect 406676 271182 406732 271238
rect 408980 270738 409036 270794
rect 408980 269998 409036 270054
rect 408596 267926 408652 267982
rect 408788 267943 408844 267982
rect 408788 267926 408790 267943
rect 408790 267926 408842 267943
rect 408842 267926 408844 267943
rect 408788 267778 408844 267834
rect 388979 264857 388983 264909
rect 388983 264857 389035 264909
rect 389035 264857 389039 264909
rect 388979 264853 389039 264857
rect 393014 264839 393074 264899
rect 407103 264880 407163 264940
rect 407706 264874 407766 264934
rect 408114 264873 408174 264933
rect 409996 264861 410056 264921
rect 410533 264881 410593 264941
rect 412052 264522 412108 264578
rect 211988 255346 212044 255402
rect 412148 247502 412204 247558
rect 412916 267778 412972 267834
rect 418964 270294 419020 270350
rect 418964 267926 419020 267982
rect 414932 267630 414988 267686
rect 415124 267630 415180 267686
rect 413684 266150 413740 266206
rect 419156 270738 419212 270794
rect 419156 270294 419212 270350
rect 428180 270886 428236 270942
rect 428948 270146 429004 270202
rect 429236 270146 429292 270202
rect 438932 270294 438988 270350
rect 439124 267965 439126 267982
rect 439126 267965 439178 267982
rect 439178 267965 439180 267982
rect 439124 267926 439180 267965
rect 439316 267926 439372 267982
rect 446324 270886 446380 270942
rect 449300 271182 449356 271238
rect 449588 271182 449644 271238
rect 449204 270294 449260 270350
rect 449204 269998 449260 270054
rect 449204 267926 449260 267982
rect 452180 271051 452236 271090
rect 452180 271034 452182 271051
rect 452182 271034 452234 271051
rect 452234 271034 452236 271051
rect 452180 270903 452236 270942
rect 452180 270886 452182 270903
rect 452182 270886 452234 270903
rect 452234 270886 452236 270903
rect 452180 270755 452236 270794
rect 452180 270738 452182 270755
rect 452182 270738 452234 270755
rect 452234 270738 452236 270755
rect 452468 270903 452524 270942
rect 452468 270886 452470 270903
rect 452470 270886 452522 270903
rect 452522 270886 452524 270903
rect 452660 270755 452716 270794
rect 452660 270738 452662 270755
rect 452662 270738 452714 270755
rect 452714 270738 452716 270755
rect 469460 271051 469516 271090
rect 469460 271034 469462 271051
rect 469462 271034 469514 271051
rect 469514 271034 469516 271051
rect 469460 270294 469516 270350
rect 469460 267926 469516 267982
rect 414932 265854 414988 265910
rect 480980 271221 480982 271238
rect 480982 271221 481034 271238
rect 481034 271221 481036 271238
rect 480980 271182 481036 271221
rect 481844 277842 481900 277898
rect 491636 274142 491692 274198
rect 489524 270294 489580 270350
rect 488084 268222 488140 268278
rect 489524 267926 489580 267982
rect 496148 277694 496204 277750
rect 498836 274290 498892 274346
rect 501044 271221 501046 271238
rect 501046 271221 501098 271238
rect 501098 271221 501100 271238
rect 501044 271182 501100 271221
rect 507092 277546 507148 277602
rect 505940 274438 505996 274494
rect 513044 270442 513100 270498
rect 509492 268814 509548 268870
rect 502292 268518 502348 268574
rect 517748 277398 517804 277454
rect 520148 274734 520204 274790
rect 516596 274586 516652 274642
rect 412916 265410 412972 265466
rect 528500 277250 528556 277306
rect 412820 265262 412876 265318
rect 527348 265262 527404 265318
rect 412724 265114 412780 265170
rect 530900 265114 530956 265170
rect 412628 264983 412684 265022
rect 412628 264966 412630 264983
rect 412630 264966 412682 264983
rect 412682 264966 412684 264983
rect 539252 277102 539308 277158
rect 539924 270146 539980 270202
rect 540020 269998 540076 270054
rect 539924 268814 539980 268870
rect 540020 268518 540076 268574
rect 538004 264966 538060 265022
rect 489524 264818 489580 264874
rect 449396 264709 449398 264726
rect 449398 264709 449450 264726
rect 449450 264709 449452 264726
rect 449396 264670 449452 264709
rect 469364 264709 469366 264726
rect 469366 264709 469418 264726
rect 469418 264709 469420 264726
rect 469364 264670 469420 264709
rect 475796 264709 475798 264726
rect 475798 264709 475850 264726
rect 475850 264709 475852 264726
rect 475796 264670 475852 264709
rect 552308 273994 552364 274050
rect 548564 270481 548566 270498
rect 548566 270481 548618 270498
rect 548618 270481 548620 270498
rect 548564 270442 548620 270481
rect 559412 271330 559468 271386
rect 560180 270146 560236 270202
rect 560084 269998 560140 270054
rect 560180 268814 560236 268870
rect 560084 268518 560140 268574
rect 563060 273106 563116 273162
rect 564500 271051 564556 271090
rect 564500 271034 564502 271051
rect 564502 271034 564554 271051
rect 564554 271034 564556 271051
rect 575924 270442 575980 270498
rect 574868 268962 574924 269018
rect 567764 268666 567820 268722
rect 560660 268074 560716 268130
rect 555860 264522 555916 264578
rect 412052 247206 412108 247262
rect 226388 246762 226444 246818
rect 211508 243654 211564 243710
rect 211316 238918 211372 238974
rect 211220 238770 211276 238826
rect 212180 236698 212236 236754
rect 211303 233751 211363 233811
rect 212372 235070 212428 235126
rect 212564 233886 212620 233942
rect 212276 233738 212332 233794
rect 212084 233590 212140 233646
rect 211700 233442 211756 233498
rect 212564 233590 212620 233646
rect 213236 242914 213292 242970
rect 214196 234922 214252 234978
rect 214964 243062 215020 243118
rect 215828 238178 215884 238234
rect 215252 238030 215308 238086
rect 214868 237882 214924 237938
rect 214772 237586 214828 237642
rect 214772 236550 214828 236606
rect 214292 233442 214348 233498
rect 216212 237586 216268 237642
rect 217172 242026 217228 242082
rect 216692 237734 216748 237790
rect 218900 242766 218956 242822
rect 218228 235218 218284 235274
rect 221204 243210 221260 243266
rect 220820 242618 220876 242674
rect 219764 235662 219820 235718
rect 221396 243210 221452 243266
rect 221300 235810 221356 235866
rect 223700 242174 223756 242230
rect 223028 235514 223084 235570
rect 224468 235366 224524 235422
rect 226004 243654 226060 243710
rect 227348 246762 227404 246818
rect 237044 246762 237100 246818
rect 227444 243654 227500 243710
rect 227732 242322 227788 242378
rect 227348 242026 227404 242082
rect 225812 236106 225868 236162
rect 227444 236698 227500 236754
rect 227636 236698 227692 236754
rect 228212 243210 228268 243266
rect 228212 242026 228268 242082
rect 229556 235958 229612 236014
rect 237716 246762 237772 246818
rect 240020 246762 240076 246818
rect 240500 246762 240556 246818
rect 241748 246762 241804 246818
rect 242516 246762 242572 246818
rect 252500 246762 252556 246818
rect 252692 246762 252748 246818
rect 266708 246762 266764 246818
rect 268628 246762 268684 246818
rect 237716 242766 237772 242822
rect 237428 242618 237484 242674
rect 238676 234330 238732 234386
rect 238964 234478 239020 234534
rect 240980 240398 241036 240454
rect 241364 238474 241420 238530
rect 241748 240546 241804 240602
rect 242324 238474 242380 238530
rect 243188 240990 243244 241046
rect 242708 240694 242764 240750
rect 243092 237290 243148 237346
rect 243572 238622 243628 238678
rect 244532 241286 244588 241342
rect 243956 237438 244012 237494
rect 245396 241730 245452 241786
rect 245300 237142 245356 237198
rect 246740 241582 246796 241638
rect 247508 242487 247564 242526
rect 247508 242470 247510 242487
rect 247510 242470 247562 242487
rect 247562 242470 247564 242487
rect 247700 242470 247756 242526
rect 247700 240102 247756 240158
rect 247988 239954 248044 240010
rect 256052 243358 256108 243414
rect 256244 243358 256300 243414
rect 256244 243227 256300 243266
rect 256244 243210 256246 243227
rect 256246 243210 256298 243227
rect 256298 243210 256300 243227
rect 256532 243210 256588 243266
rect 256340 243062 256396 243118
rect 256724 243062 256780 243118
rect 258644 238326 258700 238382
rect 259028 240842 259084 240898
rect 259604 241138 259660 241194
rect 259124 236698 259180 236754
rect 259124 236254 259180 236310
rect 261236 241434 261292 241490
rect 262964 240250 263020 240306
rect 269300 239806 269356 239862
rect 271508 241286 271564 241342
rect 271316 240990 271372 241046
rect 271508 240990 271564 241046
rect 271124 240398 271180 240454
rect 271316 240398 271372 240454
rect 271124 239658 271180 239714
rect 276404 243210 276460 243266
rect 286100 246762 286156 246818
rect 286292 246762 286348 246818
rect 288884 246762 288940 246818
rect 291956 246762 292012 246818
rect 292244 246762 292300 246818
rect 292628 246762 292684 246818
rect 277748 241730 277804 241786
rect 277748 241286 277804 241342
rect 278036 240694 278092 240750
rect 277556 240398 277612 240454
rect 278228 239806 278284 239862
rect 277940 239510 277996 239566
rect 279764 239510 279820 239566
rect 287732 241878 287788 241934
rect 287636 239510 287692 239566
rect 289652 241286 289708 241342
rect 289844 241286 289900 241342
rect 288980 236271 289036 236310
rect 288980 236254 288982 236271
rect 288982 236254 289034 236271
rect 289034 236254 289036 236271
rect 289844 240694 289900 240750
rect 289652 239806 289708 239862
rect 290900 233442 290956 233498
rect 293396 239362 293452 239418
rect 293780 239510 293836 239566
rect 293972 239214 294028 239270
rect 294068 236271 294124 236310
rect 294068 236254 294070 236271
rect 294070 236254 294122 236271
rect 294122 236254 294124 236271
rect 296276 239214 296332 239270
rect 297812 241286 297868 241342
rect 298004 241286 298060 241342
rect 298004 240990 298060 241046
rect 298196 240990 298252 241046
rect 298004 240398 298060 240454
rect 298004 239658 298060 239714
rect 298196 233442 298252 233498
rect 305300 239362 305356 239418
rect 306452 242953 306454 242970
rect 306454 242953 306506 242970
rect 306506 242953 306508 242970
rect 306452 242914 306508 242953
rect 308948 241878 309004 241934
rect 310484 242470 310540 242526
rect 310196 242322 310252 242378
rect 314996 242766 315052 242822
rect 316532 243210 316588 243266
rect 316724 242953 316726 242970
rect 316726 242953 316778 242970
rect 316778 242953 316780 242970
rect 316724 242914 316780 242953
rect 316724 242766 316780 242822
rect 318260 241730 318316 241786
rect 318260 239806 318316 239862
rect 319892 236994 319948 237050
rect 325076 242931 325132 242970
rect 325076 242914 325078 242931
rect 325078 242914 325130 242931
rect 325130 242914 325132 242931
rect 328148 242509 328150 242526
rect 328150 242509 328202 242526
rect 328202 242509 328204 242526
rect 328148 242470 328204 242509
rect 328532 242322 328588 242378
rect 329780 236846 329836 236902
rect 331124 243210 331180 243266
rect 334964 235070 335020 235126
rect 338132 236994 338188 237050
rect 338996 242322 339052 242378
rect 339764 242470 339820 242526
rect 339572 242322 339628 242378
rect 339764 236846 339820 236902
rect 341204 242618 341260 242674
rect 341108 235218 341164 235274
rect 342068 242914 342124 242970
rect 341588 235662 341644 235718
rect 342932 242766 342988 242822
rect 342548 235810 342604 235866
rect 343412 242174 343468 242230
rect 343316 235514 343372 235570
rect 344276 242322 344332 242378
rect 343796 235366 343852 235422
rect 344756 236106 344812 236162
rect 346004 235958 346060 236014
rect 347732 234330 347788 234386
rect 348212 234922 348268 234978
rect 349172 234478 349228 234534
rect 351284 239954 351340 240010
rect 351380 239066 351436 239122
rect 352244 243062 352300 243118
rect 352820 240102 352876 240158
rect 354452 241582 354508 241638
rect 354644 242026 354700 242082
rect 356756 241730 356812 241786
rect 357812 237142 357868 237198
rect 358964 241286 359020 241342
rect 358484 237290 358540 237346
rect 359252 236550 359308 236606
rect 360020 237438 360076 237494
rect 360692 238622 360748 238678
rect 361652 240990 361708 241046
rect 387380 246762 387436 246818
rect 363092 240694 363148 240750
rect 363860 238474 363916 238530
rect 364820 240546 364876 240602
rect 365780 238178 365836 238234
rect 366548 240398 366604 240454
rect 367604 240398 367660 240454
rect 369812 240250 369868 240306
rect 372884 241434 372940 241490
rect 376820 241138 376876 241194
rect 377876 240842 377932 240898
rect 378836 238326 378892 238382
rect 379412 234774 379468 234830
rect 388532 246762 388588 246818
rect 389492 246762 389548 246818
rect 389780 246762 389836 246818
rect 389300 243506 389356 243562
rect 405908 246762 405964 246818
rect 406100 246779 406156 246818
rect 406100 246762 406102 246779
rect 406102 246762 406154 246779
rect 406154 246762 406156 246779
rect 391412 238030 391468 238086
rect 393140 237882 393196 237938
rect 394676 237734 394732 237790
rect 406520 246830 406598 246834
rect 406520 246778 406524 246830
rect 406524 246778 406576 246830
rect 406576 246778 406598 246830
rect 406520 246758 406598 246778
rect 406772 246762 406828 246818
rect 407060 246762 407116 246818
rect 407252 246762 407308 246818
rect 407636 246762 407692 246818
rect 408116 246762 408172 246818
rect 408596 246762 408652 246818
rect 408788 246762 408844 246818
rect 408980 246779 409036 246818
rect 408980 246762 408982 246779
rect 408982 246762 409034 246779
rect 409034 246762 409036 246779
rect 405716 243506 405772 243562
rect 406196 243506 406252 243562
rect 409172 246762 409228 246818
rect 409364 246779 409420 246818
rect 409364 246762 409366 246779
rect 409366 246762 409418 246779
rect 409418 246762 409420 246779
rect 409844 246762 409900 246818
rect 412436 247354 412492 247410
rect 412244 247058 412300 247114
rect 409748 240398 409804 240454
rect 453620 242618 453676 242674
rect 463700 242657 463702 242674
rect 463702 242657 463754 242674
rect 463754 242657 463756 242674
rect 463700 242618 463756 242657
rect 430484 242470 430540 242526
rect 443444 242470 443500 242526
rect 443636 242509 443638 242526
rect 443638 242509 443690 242526
rect 443690 242509 443692 242526
rect 443636 242470 443692 242509
rect 483764 242470 483820 242526
rect 489524 242470 489580 242526
rect 489716 242322 489772 242378
rect 504020 242361 504022 242378
rect 504022 242361 504074 242378
rect 504074 242361 504076 242378
rect 504020 242322 504076 242361
rect 412628 238770 412684 238826
rect 411956 237586 412012 237642
rect 580916 275622 580972 275678
rect 582068 270294 582124 270350
rect 584372 271034 584428 271090
rect 580244 269998 580300 270054
rect 592724 276362 592780 276418
rect 589172 270146 589228 270202
rect 599828 276214 599884 276270
rect 602228 275474 602284 275530
rect 603380 269850 603436 269906
rect 605780 269702 605836 269758
rect 580244 268814 580300 268870
rect 596372 268814 596428 268870
rect 610580 276066 610636 276122
rect 614228 267778 614284 267834
rect 609428 266150 609484 266206
rect 617684 276954 617740 277010
rect 616532 275326 616588 275382
rect 620084 269554 620140 269610
rect 624884 275918 624940 275974
rect 623636 275178 623692 275234
rect 627284 275030 627340 275086
rect 626036 268370 626092 268426
rect 628436 265410 628492 265466
rect 630836 269406 630892 269462
rect 637940 275770 637996 275826
rect 634292 269258 634348 269314
rect 642740 276806 642796 276862
rect 641492 270590 641548 270646
rect 640340 269110 640396 269166
rect 639092 267630 639148 267686
rect 631796 265854 631852 265910
rect 646292 276658 646348 276714
rect 645140 274882 645196 274938
rect 576212 241878 576268 241934
rect 547508 238918 547564 238974
rect 511124 237734 511180 237790
rect 400340 236715 400396 236754
rect 400340 236698 400342 236715
rect 400342 236698 400394 236715
rect 400394 236698 400396 236715
rect 420404 236715 420460 236754
rect 420404 236698 420406 236715
rect 420406 236698 420458 236715
rect 420458 236698 420460 236715
rect 440660 236715 440716 236754
rect 440660 236698 440662 236715
rect 440662 236698 440714 236715
rect 440714 236698 440716 236715
rect 460724 236715 460780 236754
rect 460724 236698 460726 236715
rect 460726 236698 460778 236715
rect 460778 236698 460780 236715
rect 480980 236698 481036 236754
rect 420596 236402 420652 236458
rect 505364 237586 505420 237642
rect 547124 234626 547180 234682
rect 637172 233590 637228 233646
rect 637460 233442 637516 233498
rect 638420 236254 638476 236310
rect 648020 243654 648076 243710
rect 650036 994458 650092 994514
rect 649748 994162 649804 994218
rect 649652 994014 649708 994070
rect 649652 941770 649708 941826
rect 638036 233886 638092 233942
rect 638228 233442 638284 233498
rect 638804 233738 638860 233794
rect 638900 233590 638956 233646
rect 639284 236254 639340 236310
rect 649748 848234 649804 848290
rect 210164 62502 210220 62558
rect 210260 57988 210316 58044
rect 210260 56878 210316 56934
rect 210164 55250 210220 55306
rect 210260 54066 210316 54122
rect 210452 54214 210508 54270
rect 210644 54214 210700 54270
rect 214772 54214 214828 54270
rect 216980 54066 217036 54122
rect 216980 53918 217036 53974
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 211892 51994 211948 52050
rect 212660 51846 212716 51902
rect 213044 53474 213100 53530
rect 213236 45186 213292 45242
rect 212852 44742 212908 44798
rect 214964 53474 215020 53530
rect 214676 45038 214732 45094
rect 215780 53474 215836 53530
rect 215972 53474 216028 53530
rect 216692 53326 216748 53382
rect 217844 53178 217900 53234
rect 221108 53474 221164 53530
rect 221876 52142 221932 52198
rect 222644 51550 222700 51606
rect 223316 52290 223372 52346
rect 223700 51698 223756 51754
rect 236756 50958 236812 51014
rect 237524 51254 237580 51310
rect 237620 51106 237676 51162
rect 241940 48294 241996 48350
rect 242996 48738 243052 48794
rect 242420 48590 242476 48646
rect 243764 51402 243820 51458
rect 243380 48442 243436 48498
rect 242036 48146 242092 48202
rect 215444 44890 215500 44946
rect 297236 43114 297292 43170
rect 302420 43114 302476 43170
rect 282356 42078 282412 42134
rect 306740 42078 306796 42134
rect 467444 49034 467500 49090
rect 650132 895150 650188 895206
rect 650228 801318 650284 801374
rect 650036 754402 650092 754458
rect 649844 707486 649900 707542
rect 655124 976698 655180 976754
rect 655220 965006 655276 965062
rect 655316 953314 655372 953370
rect 674324 967522 674380 967578
rect 674996 967522 675052 967578
rect 674516 967374 674572 967430
rect 675764 965598 675820 965654
rect 675284 965006 675340 965062
rect 675188 964858 675244 964914
rect 675092 962786 675148 962842
rect 675188 962490 675244 962546
rect 675764 962194 675820 962250
rect 675380 961454 675436 961510
rect 675668 961010 675724 961066
rect 675764 960122 675820 960178
rect 675476 959086 675532 959142
rect 654452 929782 654508 929838
rect 653972 918090 654028 918146
rect 654452 906398 654508 906454
rect 653972 882866 654028 882922
rect 654452 871174 654508 871230
rect 654164 859482 654220 859538
rect 653972 835950 654028 836006
rect 653972 824258 654028 824314
rect 654452 812566 654508 812622
rect 654068 789034 654124 789090
rect 654068 777342 654124 777398
rect 653972 765502 654028 765558
rect 653972 742118 654028 742174
rect 655220 730426 655276 730482
rect 654260 718586 654316 718642
rect 654452 695202 654508 695258
rect 655124 683510 655180 683566
rect 654452 671670 654508 671726
rect 650324 660570 650380 660626
rect 645236 231518 645292 231574
rect 645140 231074 645196 231130
rect 654260 648286 654316 648342
rect 654068 624754 654124 624810
rect 654356 613062 654412 613118
rect 654452 601370 654508 601426
rect 654452 589530 654508 589586
rect 654452 577838 654508 577894
rect 654452 566146 654508 566202
rect 654452 554454 654508 554510
rect 654452 542614 654508 542670
rect 655316 636594 655372 636650
rect 654068 530922 654124 530978
rect 654452 519269 654454 519286
rect 654454 519269 654506 519286
rect 654506 519269 654508 519286
rect 654452 519230 654508 519269
rect 654452 507390 654508 507446
rect 654356 495698 654412 495754
rect 654260 484006 654316 484062
rect 654452 472205 654454 472222
rect 654454 472205 654506 472222
rect 654506 472205 654508 472222
rect 654452 472166 654508 472205
rect 654452 460474 654508 460530
rect 654356 448782 654412 448838
rect 654452 436942 654508 436998
rect 654452 425398 654508 425454
rect 653876 413558 653932 413614
rect 654452 401718 654508 401774
rect 654452 390026 654508 390082
rect 654452 378482 654508 378538
rect 654452 366494 654508 366550
rect 655220 354802 655276 354858
rect 654452 343110 654508 343166
rect 654452 331566 654508 331622
rect 655124 319726 655180 319782
rect 654548 296194 654604 296250
rect 654068 284650 654124 284706
rect 645812 232702 645868 232758
rect 645716 231962 645772 232018
rect 645332 230630 645388 230686
rect 645620 210354 645676 210410
rect 645332 141090 645388 141146
rect 645332 140794 645388 140850
rect 351380 43114 351436 43170
rect 357140 43114 357196 43170
rect 362804 42078 362860 42134
rect 364628 42078 364684 42134
rect 374324 41190 374380 41246
rect 334100 40911 334156 40950
rect 334100 40894 334102 40911
rect 334102 40894 334154 40911
rect 334154 40894 334156 40911
rect 344180 40911 344236 40950
rect 344180 40894 344182 40911
rect 344182 40894 344234 40911
rect 344234 40894 344236 40911
rect 374324 40746 374380 40802
rect 211028 40598 211084 40654
rect 411092 45186 411148 45242
rect 416564 44742 416620 44798
rect 521588 43262 521644 43318
rect 455732 43114 455788 43170
rect 463988 43114 464044 43170
rect 471092 42078 471148 42134
rect 645428 104238 645484 104294
rect 645428 87662 645484 87718
rect 645428 84998 645484 85054
rect 645428 83222 645484 83278
rect 645428 82482 645484 82538
rect 645428 81315 645484 81354
rect 645428 81298 645430 81315
rect 645430 81298 645482 81315
rect 645482 81298 645484 81315
rect 645428 79966 645484 80022
rect 645428 78634 645484 78690
rect 645428 77637 645430 77654
rect 645430 77637 645482 77654
rect 645482 77637 645484 77654
rect 645428 77598 645484 77637
rect 645428 77006 645484 77062
rect 645428 76710 645484 76766
rect 645428 75378 645484 75434
rect 645428 74342 645484 74398
rect 645428 72862 645484 72918
rect 647924 210354 647980 210410
rect 646292 166250 646348 166306
rect 647924 166990 647980 167046
rect 646868 165954 646924 166010
rect 655316 307886 655372 307942
rect 673844 939106 673900 939162
rect 673076 707486 673132 707542
rect 675476 957606 675532 957662
rect 675092 953462 675148 953518
rect 675476 955978 675532 956034
rect 675188 953314 675244 953370
rect 676820 940882 676876 940938
rect 674612 939846 674668 939902
rect 674420 939567 674476 939606
rect 674420 939550 674422 939567
rect 674422 939550 674474 939567
rect 674474 939550 674476 939567
rect 676916 940438 676972 940494
rect 676820 938218 676876 938274
rect 674420 937961 674422 937978
rect 674422 937961 674474 937978
rect 674474 937961 674476 937978
rect 674420 937922 674476 937961
rect 674132 936886 674188 936942
rect 674036 934666 674092 934722
rect 677012 929486 677068 929542
rect 676820 928894 676876 928950
rect 676820 928450 676876 928506
rect 677012 928450 677068 928506
rect 675380 876946 675436 877002
rect 675380 876502 675436 876558
rect 675284 875910 675340 875966
rect 675092 875614 675148 875670
rect 673844 761210 673900 761266
rect 673844 760618 673900 760674
rect 673364 752034 673420 752090
rect 674516 777490 674572 777546
rect 675380 875762 675436 875818
rect 675476 874134 675532 874190
rect 675380 873394 675436 873450
rect 675380 872802 675436 872858
rect 675380 869842 675436 869898
rect 674612 776898 674668 776954
rect 674324 773050 674380 773106
rect 674324 762877 674326 762894
rect 674326 762877 674378 762894
rect 674378 762877 674380 762894
rect 674324 762838 674380 762877
rect 674324 762285 674326 762302
rect 674326 762285 674378 762302
rect 674378 762285 674380 762302
rect 674324 762246 674380 762285
rect 673268 708078 673324 708134
rect 673172 707042 673228 707098
rect 674900 862146 674956 862202
rect 675380 864662 675436 864718
rect 675188 862146 675244 862202
rect 675764 787998 675820 788054
rect 675476 787110 675532 787166
rect 675764 786666 675820 786722
rect 675764 784890 675820 784946
rect 675668 784150 675724 784206
rect 675764 781930 675820 781986
rect 675764 780598 675820 780654
rect 674900 776158 674956 776214
rect 674900 774826 674956 774882
rect 674612 761989 674614 762006
rect 674614 761989 674666 762006
rect 674666 761989 674668 762006
rect 674612 761950 674668 761989
rect 677876 760322 677932 760378
rect 677876 759878 677932 759934
rect 676916 759730 676972 759786
rect 677588 759286 677644 759342
rect 676916 756030 676972 756086
rect 677588 753366 677644 753422
rect 677012 751146 677068 751202
rect 676820 750554 676876 750610
rect 677012 750554 677068 750610
rect 676820 750110 676876 750166
rect 673748 715626 673804 715682
rect 674132 713554 674188 713610
rect 673748 671078 673804 671134
rect 675380 743154 675436 743210
rect 675476 742414 675532 742470
rect 675476 741674 675532 741730
rect 675188 740342 675244 740398
rect 675380 740046 675436 740102
rect 675476 739158 675532 739214
rect 675380 738566 675436 738622
rect 674516 728058 674572 728114
rect 674420 717885 674422 717902
rect 674422 717885 674474 717902
rect 674474 717885 674476 717902
rect 674420 717846 674476 717885
rect 674420 717293 674422 717310
rect 674422 717293 674474 717310
rect 674474 717293 674476 717310
rect 674420 717254 674476 717293
rect 674420 716849 674422 716866
rect 674422 716849 674474 716866
rect 674474 716849 674476 716866
rect 674420 716810 674476 716849
rect 674420 716257 674422 716274
rect 674422 716257 674474 716274
rect 674474 716257 674476 716274
rect 674420 716218 674476 716257
rect 674420 709745 674422 709762
rect 674422 709745 674474 709762
rect 674474 709745 674476 709762
rect 674420 709706 674476 709745
rect 674420 709153 674422 709170
rect 674422 709153 674474 709170
rect 674474 709153 674476 709170
rect 674420 709114 674476 709153
rect 674420 708635 674422 708652
rect 674422 708635 674474 708652
rect 674474 708635 674476 708652
rect 674420 708596 674476 708635
rect 674228 666638 674284 666694
rect 673844 662790 673900 662846
rect 673364 662346 673420 662402
rect 673844 661754 673900 661810
rect 673268 617354 673324 617410
rect 673076 616762 673132 616818
rect 673076 527074 673132 527130
rect 672980 526630 673036 526686
rect 674132 630674 674188 630730
rect 673844 627753 673846 627770
rect 673846 627753 673898 627770
rect 673898 627753 673900 627770
rect 673844 627714 673900 627753
rect 673364 573694 673420 573750
rect 674132 619870 674188 619926
rect 673844 617798 673900 617854
rect 674420 672671 674422 672688
rect 674422 672671 674474 672688
rect 674474 672671 674476 672688
rect 674420 672632 674476 672671
rect 674420 672153 674422 672170
rect 674422 672153 674474 672170
rect 674474 672153 674476 672170
rect 674420 672114 674476 672153
rect 674420 671561 674422 671578
rect 674422 671561 674474 671578
rect 674474 671561 674476 671578
rect 674420 671522 674476 671561
rect 675380 734422 675436 734478
rect 677012 706154 677068 706210
rect 676820 705562 676876 705618
rect 677012 705562 677068 705618
rect 676820 705118 676876 705174
rect 675476 697866 675532 697922
rect 675764 697274 675820 697330
rect 675380 696830 675436 696886
rect 675668 694758 675724 694814
rect 675476 694314 675532 694370
rect 675764 691946 675820 692002
rect 675764 689134 675820 689190
rect 675092 688246 675148 688302
rect 674612 668562 674668 668618
rect 674516 666342 674572 666398
rect 674324 623274 674380 623330
rect 674420 621054 674476 621110
rect 674612 627309 674614 627326
rect 674614 627309 674666 627326
rect 674666 627309 674668 627326
rect 674612 627270 674668 627309
rect 674612 626865 674614 626882
rect 674614 626865 674666 626882
rect 674666 626865 674668 626882
rect 674612 626826 674668 626865
rect 674612 625215 674668 625254
rect 674612 625198 674614 625215
rect 674614 625198 674666 625215
rect 674666 625198 674668 625215
rect 674900 664122 674956 664178
rect 674900 660866 674956 660922
rect 674900 660422 674956 660478
rect 675092 660422 675148 660478
rect 675092 659830 675148 659886
rect 675092 653614 675148 653670
rect 675380 652578 675436 652634
rect 675476 652134 675532 652190
rect 675476 651394 675532 651450
rect 675380 649618 675436 649674
rect 675476 648878 675532 648934
rect 675764 645326 675820 645382
rect 675380 640294 675436 640350
rect 675764 638518 675820 638574
rect 674996 630674 675052 630730
rect 674900 621942 674956 621998
rect 677204 624606 677260 624662
rect 676820 624014 676876 624070
rect 674996 620758 675052 620814
rect 674900 619130 674956 619186
rect 677108 615874 677164 615930
rect 676916 615282 676972 615338
rect 677108 615282 677164 615338
rect 676916 614838 676972 614894
rect 675380 607734 675436 607790
rect 675476 607142 675532 607198
rect 675476 606402 675532 606458
rect 675380 604774 675436 604830
rect 675092 595450 675148 595506
rect 674900 590566 674956 590622
rect 674612 590418 674668 590474
rect 675764 595302 675820 595358
rect 675764 593378 675820 593434
rect 675476 590270 675532 590326
rect 674900 590122 674956 590178
rect 674612 582130 674668 582186
rect 674420 581908 674476 581964
rect 674612 581577 674614 581594
rect 674614 581577 674666 581594
rect 674666 581577 674668 581594
rect 674612 581538 674668 581577
rect 674420 580837 674422 580854
rect 674422 580837 674474 580854
rect 674474 580837 674476 580854
rect 674420 580798 674476 580837
rect 674612 580075 674668 580114
rect 674612 580058 674614 580075
rect 674614 580058 674666 580075
rect 674666 580058 674668 580075
rect 676916 580058 676972 580114
rect 676820 579466 676876 579522
rect 674612 574473 674614 574490
rect 674614 574473 674666 574490
rect 674666 574473 674668 574490
rect 674612 574434 674668 574473
rect 674612 573437 674614 573454
rect 674614 573437 674666 573454
rect 674666 573437 674668 573454
rect 674612 573398 674668 573437
rect 674612 572845 674614 572862
rect 674614 572845 674666 572862
rect 674666 572845 674668 572862
rect 674612 572806 674668 572845
rect 673748 572066 673804 572122
rect 674612 571809 674614 571826
rect 674614 571809 674666 571826
rect 674666 571809 674668 571826
rect 674612 571770 674668 571809
rect 677012 570734 677068 570790
rect 676820 570142 676876 570198
rect 677012 570142 677068 570198
rect 676820 569698 676876 569754
rect 673268 527666 673324 527722
rect 673172 484154 673228 484210
rect 673748 536842 673804 536898
rect 673748 535806 673804 535862
rect 673748 529903 673804 529942
rect 673748 529886 673750 529903
rect 673750 529886 673802 529903
rect 673802 529886 673804 529903
rect 673748 528702 673804 528758
rect 673748 528258 673804 528314
rect 673844 492294 673900 492350
rect 674324 492925 674326 492942
rect 674326 492925 674378 492942
rect 674378 492925 674380 492942
rect 674324 492886 674380 492925
rect 675476 562446 675532 562502
rect 675476 562002 675532 562058
rect 675380 561410 675436 561466
rect 675476 558894 675532 558950
rect 675764 554454 675820 554510
rect 674612 536585 674614 536602
rect 674614 536585 674666 536602
rect 674666 536585 674668 536602
rect 674612 536546 674668 536585
rect 674612 493182 674668 493238
rect 674516 489334 674572 489390
rect 674420 487410 674476 487466
rect 676820 537138 676876 537194
rect 677396 534918 677452 534974
rect 677204 534474 677260 534530
rect 677012 533882 677068 533938
rect 674900 529481 674902 529498
rect 674902 529481 674954 529498
rect 674954 529481 674956 529498
rect 674900 529442 674956 529481
rect 676820 525150 676876 525206
rect 676820 524706 676876 524762
rect 677108 525742 677164 525798
rect 677108 525150 677164 525206
rect 674900 503986 674956 504042
rect 675092 503986 675148 504042
rect 677396 492146 677452 492202
rect 677204 491110 677260 491166
rect 676820 490518 676876 490574
rect 675380 488298 675436 488354
rect 674996 487114 675052 487170
rect 674900 485486 674956 485542
rect 674228 484746 674284 484802
rect 673460 483710 673516 483766
rect 673364 482526 673420 482582
rect 677012 481638 677068 481694
rect 676820 481194 676876 481250
rect 677012 481194 677068 481250
rect 676820 480750 676876 480806
rect 674708 405457 674710 405474
rect 674710 405457 674762 405474
rect 674762 405457 674764 405474
rect 674708 405418 674764 405457
rect 674420 404717 674422 404734
rect 674422 404717 674474 404734
rect 674474 404717 674476 404734
rect 674420 404678 674476 404717
rect 674708 404421 674710 404438
rect 674710 404421 674762 404438
rect 674762 404421 674764 404438
rect 674708 404382 674764 404421
rect 673652 403050 673708 403106
rect 673364 374338 673420 374394
rect 677300 402310 677356 402366
rect 677108 401718 677164 401774
rect 674900 401274 674956 401330
rect 673460 373006 673516 373062
rect 674516 399646 674572 399702
rect 674420 397574 674476 397630
rect 673940 396538 673996 396594
rect 674228 394318 674284 394374
rect 674612 395798 674668 395854
rect 674708 395058 674764 395114
rect 674804 394614 674860 394670
rect 674996 400090 675052 400146
rect 675188 397870 675244 397926
rect 675092 396834 675148 396890
rect 677108 393430 677164 393486
rect 676916 392986 676972 393042
rect 677108 392986 677164 393042
rect 676916 392542 676972 392598
rect 675092 374486 675148 374542
rect 675476 378778 675532 378834
rect 675188 374042 675244 374098
rect 675476 373894 675532 373950
rect 675380 371970 675436 372026
rect 674420 360021 674422 360038
rect 674422 360021 674474 360038
rect 674474 360021 674476 360038
rect 674420 359982 674476 360021
rect 674708 359725 674710 359742
rect 674710 359725 674762 359742
rect 674762 359725 674764 359742
rect 674708 359686 674764 359725
rect 674420 358985 674422 359002
rect 674422 358985 674474 359002
rect 674474 358985 674476 359002
rect 674420 358946 674476 358985
rect 673844 358354 673900 358410
rect 674420 356282 674476 356338
rect 673940 354062 673996 354118
rect 674324 350806 674380 350862
rect 674228 349696 674284 349752
rect 674036 349178 674092 349234
rect 674804 354950 674860 355006
rect 674612 354358 674668 354414
rect 674516 352138 674572 352194
rect 674708 350066 674764 350122
rect 677012 353174 677068 353230
rect 674900 352730 674956 352786
rect 674996 351694 675052 351750
rect 676820 351102 676876 351158
rect 676916 347698 676972 347754
rect 676916 347254 676972 347310
rect 676820 345478 676876 345534
rect 677108 348290 677164 348346
rect 677108 347698 677164 347754
rect 677012 345330 677068 345386
rect 675284 334970 675340 335026
rect 675476 333786 675532 333842
rect 675764 330530 675820 330586
rect 675188 329494 675244 329550
rect 675380 328310 675436 328366
rect 675764 326830 675820 326886
rect 674420 315029 674422 315046
rect 674422 315029 674474 315046
rect 674474 315029 674476 315046
rect 674420 314990 674476 315029
rect 674708 314733 674710 314750
rect 674710 314733 674762 314750
rect 674762 314733 674764 314750
rect 674708 314694 674764 314733
rect 674420 313993 674422 314010
rect 674422 313993 674474 314010
rect 674474 313993 674476 314010
rect 674420 313954 674476 313993
rect 673940 311290 673996 311346
rect 674708 309958 674764 310014
rect 674324 309588 674380 309644
rect 674036 305814 674092 305870
rect 674228 304186 674284 304242
rect 674612 305074 674668 305130
rect 674516 304482 674572 304538
rect 674420 303594 674476 303650
rect 674420 302597 674422 302614
rect 674422 302597 674474 302614
rect 674474 302597 674476 302614
rect 674420 302558 674476 302597
rect 674996 308774 675052 308830
rect 674900 307738 674956 307794
rect 674804 306702 674860 306758
rect 677012 308182 677068 308238
rect 675092 307146 675148 307202
rect 676916 305962 676972 306018
rect 676820 302706 676876 302762
rect 676820 302262 676876 302318
rect 676916 299450 676972 299506
rect 677012 299302 677068 299358
rect 675284 289978 675340 290034
rect 675476 289534 675532 289590
rect 675188 284946 675244 285002
rect 675092 284798 675148 284854
rect 675764 284798 675820 284854
rect 675380 283614 675436 283670
rect 675764 281838 675820 281894
rect 673556 276362 673612 276418
rect 673844 269998 673900 270054
rect 674708 269741 674710 269758
rect 674710 269741 674762 269758
rect 674762 269741 674764 269758
rect 674708 269702 674764 269741
rect 674708 269149 674710 269166
rect 674710 269149 674762 269166
rect 674762 269149 674764 269166
rect 674708 269110 674764 269149
rect 674612 266002 674668 266058
rect 674420 264596 674476 264652
rect 674324 262450 674380 262506
rect 674132 261266 674188 261322
rect 674036 259194 674092 259250
rect 677204 265410 677260 265466
rect 674900 264966 674956 265022
rect 674708 261710 674764 261766
rect 674804 260082 674860 260138
rect 675188 262746 675244 262802
rect 674996 259490 675052 259546
rect 677108 258306 677164 258362
rect 676916 257714 676972 257770
rect 676916 257270 676972 257326
rect 677108 257270 677164 257326
rect 677588 263190 677644 263246
rect 677588 251646 677644 251702
rect 677204 251498 677260 251554
rect 675188 245874 675244 245930
rect 675380 244690 675436 244746
rect 675476 243506 675532 243562
rect 675380 242026 675436 242082
rect 675188 238918 675244 238974
rect 675764 238622 675820 238678
rect 675764 236846 675820 236902
rect 674708 225045 674710 225062
rect 674710 225045 674762 225062
rect 674762 225045 674764 225062
rect 674708 225006 674764 225045
rect 674420 224305 674422 224322
rect 674422 224305 674474 224322
rect 674474 224305 674476 224322
rect 674420 224266 674476 224305
rect 674708 224009 674710 224026
rect 674710 224009 674762 224026
rect 674762 224009 674764 224026
rect 674708 223970 674764 224009
rect 674996 220862 675052 220918
rect 674900 217014 674956 217070
rect 674516 216422 674572 216478
rect 674516 215386 674572 215442
rect 674804 214794 674860 214850
rect 674708 214350 674764 214406
rect 674612 213758 674668 213814
rect 675476 219678 675532 219734
rect 675092 219234 675148 219290
rect 675284 217606 675340 217662
rect 677108 218642 677164 218698
rect 676916 215978 676972 216034
rect 676820 212574 676876 212630
rect 676820 212130 676876 212186
rect 677012 213166 677068 213222
rect 677012 211982 677068 212038
rect 677204 218050 677260 218106
rect 677108 207690 677164 207746
rect 677204 207542 677260 207598
rect 676916 207394 676972 207450
rect 675380 199994 675436 200050
rect 675476 199550 675532 199606
rect 675764 198366 675820 198422
rect 675764 195258 675820 195314
rect 675380 193482 675436 193538
rect 675092 193038 675148 193094
rect 675764 191558 675820 191614
rect 674612 179570 674668 179626
rect 674420 179313 674422 179330
rect 674422 179313 674474 179330
rect 674474 179313 674476 179330
rect 674420 179274 674476 179313
rect 674420 178795 674422 178812
rect 674422 178795 674474 178812
rect 674474 178795 674476 178812
rect 674420 178756 674476 178795
rect 675092 175870 675148 175926
rect 674036 173798 674092 173854
rect 673940 170542 673996 170598
rect 674996 172022 675052 172078
rect 674900 171430 674956 171486
rect 674420 170098 674476 170154
rect 674228 169506 674284 169562
rect 674132 168914 674188 168970
rect 674708 168174 674764 168230
rect 674612 167582 674668 167638
rect 674708 167177 674710 167194
rect 674710 167177 674762 167194
rect 674762 167177 674764 167194
rect 674708 167138 674764 167177
rect 676916 175130 676972 175186
rect 675476 174686 675532 174742
rect 675188 174242 675244 174298
rect 675284 172614 675340 172670
rect 676820 173058 676876 173114
rect 676916 161514 676972 161570
rect 676820 161366 676876 161422
rect 675284 155150 675340 155206
rect 675476 154410 675532 154466
rect 675476 150266 675532 150322
rect 675764 148490 675820 148546
rect 675764 146566 675820 146622
rect 676916 134282 676972 134338
rect 676820 133838 676876 133894
rect 674420 133581 674422 133598
rect 674422 133581 674474 133598
rect 674474 133581 674476 133598
rect 674420 133542 674476 133581
rect 674420 132523 674476 132562
rect 674420 132506 674422 132523
rect 674422 132506 674474 132523
rect 674474 132506 674476 132523
rect 645908 121406 645964 121462
rect 645812 121110 645868 121166
rect 646004 120814 646060 120870
rect 674516 130582 674572 130638
rect 674324 129250 674380 129306
rect 674228 127030 674284 127086
rect 673940 125402 673996 125458
rect 647636 120370 647692 120426
rect 674420 123774 674476 123830
rect 668180 106497 668182 106514
rect 668182 106497 668234 106514
rect 668234 106497 668236 106514
rect 645812 88106 645868 88162
rect 668180 106458 668236 106497
rect 677108 129990 677164 130046
rect 675188 129546 675244 129602
rect 675092 127326 675148 127382
rect 674612 126290 674668 126346
rect 674804 124662 674860 124718
rect 674708 121850 674764 121906
rect 674900 124070 674956 124126
rect 677012 127770 677068 127826
rect 676820 122886 676876 122942
rect 676916 122294 676972 122350
rect 677012 118002 677068 118058
rect 677108 117854 677164 117910
rect 675380 110010 675436 110066
rect 675476 109270 675532 109326
rect 675380 108086 675436 108142
rect 665300 105126 665356 105182
rect 675380 105126 675436 105182
rect 665204 104551 665260 104590
rect 665204 104534 665206 104551
rect 665206 104534 665258 104551
rect 665258 104534 665260 104551
rect 675764 103202 675820 103258
rect 675764 101426 675820 101482
rect 645812 86626 645868 86682
rect 645812 84110 645868 84166
rect 646004 80114 646060 80170
rect 645812 79226 645868 79282
rect 645908 78486 645964 78542
rect 645812 75970 645868 76026
rect 645908 75230 645964 75286
rect 645812 73750 645868 73806
rect 646196 80854 646252 80910
rect 646388 72714 646444 72770
rect 647252 85738 647308 85794
rect 647540 88994 647596 89050
rect 647444 82186 647500 82242
rect 647636 87366 647692 87422
rect 647828 86182 647884 86238
rect 647732 85442 647788 85498
rect 650900 86922 650956 86978
rect 650996 85294 651052 85350
rect 650996 84258 651052 84314
rect 650612 83814 650668 83870
rect 650900 82630 650956 82686
rect 651188 86182 651244 86238
rect 651092 83370 651148 83426
rect 663476 85590 663532 85646
rect 663284 85146 663340 85202
rect 662900 81150 662956 81206
rect 646676 72122 646732 72178
rect 663380 84702 663436 84758
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 529268 43262 529324 43318
rect 142100 40154 142156 40210
rect 443444 40598 443500 40654
rect 453524 40598 453580 40654
rect 623444 40450 623500 40506
rect 443444 40302 443500 40358
rect 453524 40302 453580 40358
<< metal3 >>
rect 125334 1031610 125934 1031616
rect 121358 1022708 121958 1031418
rect 92271 1016716 92337 1016719
rect 92271 1016714 104382 1016716
rect 92271 1016658 92276 1016714
rect 92332 1016658 104382 1016714
rect 92271 1016656 104382 1016658
rect 92271 1016653 92337 1016656
rect 98562 1015916 99486 1015976
rect 98562 1015680 98622 1015916
rect 99426 1015798 99486 1015916
rect 104322 1015798 104382 1016656
rect 98400 1015650 98622 1015680
rect 98370 1015620 98622 1015650
rect 60236 1000288 62784 1000294
rect 60236 1000238 62792 1000288
rect 60236 999438 60258 1000238
rect 62730 999438 62792 1000238
rect 60236 999380 62792 999438
rect 60236 997622 62784 999380
rect 60236 996948 60276 997622
rect 62750 996948 62784 997622
rect 60236 996908 62784 996948
rect 81039 995848 81105 995851
rect 94959 995848 95025 995851
rect 81039 995846 95025 995848
rect 81039 995790 81044 995846
rect 81100 995790 94964 995846
rect 95020 995790 95025 995846
rect 97935 995848 98001 995851
rect 98370 995848 98430 1015620
rect 106287 999400 106353 999403
rect 106287 999398 106464 999400
rect 106287 999342 106292 999398
rect 106348 999342 106464 999398
rect 106287 999340 106464 999342
rect 106287 999337 106353 999340
rect 121358 997559 121958 1022108
rect 122816 1022042 123416 1031150
rect 122816 997633 123416 1021442
rect 124006 1030858 124606 1031398
rect 121353 996961 121359 997559
rect 121957 996961 121963 997559
rect 122811 997035 122817 997633
rect 123415 997035 123421 997633
rect 124006 997605 124606 1030258
rect 125334 997663 125934 1031010
rect 173268 1022788 173868 1031494
rect 148527 1015976 148593 1015979
rect 148527 1015974 150846 1015976
rect 148527 1015918 148532 1015974
rect 148588 1015918 150846 1015974
rect 148527 1015916 150846 1015918
rect 148527 1015913 148593 1015916
rect 149730 1015798 149790 1015916
rect 150786 1015798 150846 1015916
rect 145359 1007984 145425 1007987
rect 148527 1007984 148593 1007987
rect 145359 1007982 148593 1007984
rect 145359 1007926 145364 1007982
rect 145420 1007926 148532 1007982
rect 148588 1007926 148593 1007982
rect 145359 1007924 148593 1007926
rect 145359 1007921 145425 1007924
rect 148527 1007921 148593 1007924
rect 161184 1005408 161598 1005468
rect 160431 1003248 160497 1003251
rect 160032 1003246 160497 1003248
rect 160032 1003190 160436 1003246
rect 160492 1003190 160497 1003246
rect 161538 1003214 161598 1005408
rect 160032 1003188 160497 1003190
rect 160431 1003185 160497 1003188
rect 161487 1003209 161598 1003214
rect 161487 1003153 161492 1003209
rect 161548 1003153 161598 1003209
rect 161487 1003151 161598 1003153
rect 161487 1003148 161553 1003151
rect 151119 1002508 151185 1002511
rect 151119 1002506 151392 1002508
rect 151119 1002450 151124 1002506
rect 151180 1002450 151392 1002506
rect 151119 1002448 151392 1002450
rect 151119 1002445 151185 1002448
rect 152751 1002360 152817 1002363
rect 152751 1002358 153024 1002360
rect 152751 1002302 152756 1002358
rect 152812 1002302 153024 1002358
rect 152751 1002300 153024 1002302
rect 152751 1002297 152817 1002300
rect 157647 1000880 157713 1000883
rect 157647 1000878 157920 1000880
rect 157647 1000822 157652 1000878
rect 157708 1000822 157920 1000878
rect 157647 1000820 157920 1000822
rect 157647 1000817 157713 1000820
rect 155535 999548 155601 999551
rect 155535 999546 155712 999548
rect 155535 999490 155540 999546
rect 155596 999490 155712 999546
rect 155535 999488 155712 999490
rect 155535 999485 155601 999488
rect 122816 997034 123416 997035
rect 124001 997007 124007 997605
rect 124605 997007 124611 997605
rect 125329 997065 125335 997663
rect 125933 997065 125939 997663
rect 173268 997623 173868 1022188
rect 174520 1022050 175120 1031360
rect 125334 997064 125934 997065
rect 173263 997025 173269 997623
rect 173867 997025 173873 997623
rect 174520 997529 175120 1021450
rect 173268 997024 173868 997025
rect 124006 997006 124606 997007
rect 121358 996960 121958 996961
rect 174520 996931 174521 997529
rect 175119 996931 175120 997529
rect 176204 1021268 176804 1031398
rect 176204 997437 176804 1020668
rect 177460 1020702 178060 1031868
rect 174520 996930 175120 996931
rect 174521 996925 175119 996930
rect 176199 996839 176205 997437
rect 176803 996839 176809 997437
rect 177460 997433 178060 1020102
rect 223906 1022792 224506 1030706
rect 200610 1015916 201726 1015976
rect 200610 1015798 200670 1015916
rect 201666 1015798 201726 1015916
rect 213807 1005172 213873 1005175
rect 218799 1005172 218865 1005175
rect 213807 1005170 218865 1005172
rect 213807 1005114 213812 1005170
rect 213868 1005114 218804 1005170
rect 218860 1005114 218865 1005170
rect 213807 1005112 218865 1005114
rect 213807 1005109 213873 1005112
rect 218799 1005109 218865 1005112
rect 211791 1003248 211857 1003251
rect 211488 1003246 211857 1003248
rect 211488 1003190 211796 1003246
rect 211852 1003190 211857 1003246
rect 211488 1003188 211857 1003190
rect 211791 1003185 211857 1003188
rect 209103 1000880 209169 1000883
rect 209103 1000878 209376 1000880
rect 209103 1000822 209108 1000878
rect 209164 1000822 209376 1000878
rect 209103 1000820 209376 1000822
rect 209103 1000817 209169 1000820
rect 206895 999400 206961 999403
rect 206895 999398 207168 999400
rect 206895 999342 206900 999398
rect 206956 999342 207168 999398
rect 206895 999340 207168 999342
rect 206895 999337 206961 999340
rect 176204 996838 176804 996839
rect 177455 996835 177461 997433
rect 178059 996835 178065 997433
rect 223906 997395 224506 1022192
rect 225484 1022096 226084 1030950
rect 177460 996834 178060 996835
rect 223901 996797 223907 997395
rect 224505 996797 224511 997395
rect 225484 997305 226084 1021496
rect 227324 1021398 227924 1030600
rect 227324 997481 227924 1020798
rect 228774 1020614 229374 1030600
rect 228774 997579 229374 1020014
rect 274880 1022726 275480 1031902
rect 251970 1015916 252798 1015976
rect 251970 1015798 252030 1015916
rect 252738 1015828 252798 1015916
rect 252738 1015768 253152 1015828
rect 253839 1002360 253905 1002363
rect 255471 1002360 255537 1002363
rect 253839 1002358 254208 1002360
rect 253839 1002302 253844 1002358
rect 253900 1002302 254208 1002358
rect 253839 1002300 254208 1002302
rect 255471 1002358 255840 1002360
rect 255471 1002302 255476 1002358
rect 255532 1002302 255840 1002358
rect 255471 1002300 255840 1002302
rect 253839 1002297 253905 1002300
rect 255471 1002297 255537 1002300
rect 258831 999696 258897 999699
rect 258831 999694 259104 999696
rect 258831 999638 258836 999694
rect 258892 999638 259104 999694
rect 258831 999636 259104 999638
rect 258831 999633 258897 999636
rect 258351 999548 258417 999551
rect 260463 999548 260529 999551
rect 258351 999546 258528 999548
rect 258351 999490 258356 999546
rect 258412 999490 258528 999546
rect 258351 999488 258528 999490
rect 260463 999546 260736 999548
rect 260463 999490 260468 999546
rect 260524 999490 260736 999546
rect 260463 999488 260736 999490
rect 258351 999485 258417 999488
rect 260463 999485 260529 999488
rect 223906 996796 224506 996797
rect 225479 996707 225485 997305
rect 226083 996707 226089 997305
rect 227319 996883 227325 997481
rect 227923 996883 227929 997481
rect 228769 996981 228775 997579
rect 229373 996981 229379 997579
rect 274880 997463 275480 1022126
rect 276374 1022110 276974 1031770
rect 276374 997551 276974 1021510
rect 277780 1021316 278380 1031858
rect 277780 997595 278380 1020716
rect 278922 1020656 279522 1031990
rect 278922 997595 279522 1020056
rect 327774 1022684 328374 1030212
rect 299151 1005912 299217 1005915
rect 302991 1005912 303057 1005915
rect 299151 1005910 303057 1005912
rect 299151 1005854 299156 1005910
rect 299212 1005854 302996 1005910
rect 303052 1005854 303057 1005910
rect 299151 1005852 303057 1005854
rect 299151 1005849 299217 1005852
rect 302991 1005849 303057 1005852
rect 316431 1003248 316497 1003251
rect 316128 1003246 316497 1003248
rect 316128 1003190 316436 1003246
rect 316492 1003190 316497 1003246
rect 316128 1003188 316497 1003190
rect 316431 1003185 316497 1003188
rect 308847 1002952 308913 1002955
rect 308847 1002950 309024 1002952
rect 308847 1002894 308852 1002950
rect 308908 1002894 309024 1002950
rect 308847 1002892 309024 1002894
rect 308847 1002889 308913 1002892
rect 308271 1002804 308337 1002807
rect 309327 1002804 309393 1002807
rect 308271 1002802 308448 1002804
rect 308271 1002746 308276 1002802
rect 308332 1002746 308448 1002802
rect 308271 1002744 308448 1002746
rect 309327 1002802 309600 1002804
rect 309327 1002746 309332 1002802
rect 309388 1002746 309600 1002802
rect 309327 1002744 309600 1002746
rect 308271 1002741 308337 1002744
rect 309327 1002741 309393 1002744
rect 310479 999548 310545 999551
rect 312111 999548 312177 999551
rect 310479 999546 310656 999548
rect 310479 999490 310484 999546
rect 310540 999490 310656 999546
rect 310479 999488 310656 999490
rect 312111 999546 312288 999548
rect 312111 999490 312116 999546
rect 312172 999490 312288 999546
rect 312111 999488 312288 999490
rect 310479 999485 310545 999488
rect 312111 999485 312177 999488
rect 309903 999400 309969 999403
rect 309903 999398 310176 999400
rect 309903 999342 309908 999398
rect 309964 999342 310176 999398
rect 309903 999340 310176 999342
rect 309903 999337 309969 999340
rect 304335 999252 304401 999255
rect 304128 999250 304401 999252
rect 304128 999194 304340 999250
rect 304396 999194 304401 999250
rect 304128 999192 304401 999194
rect 304335 999189 304401 999192
rect 304911 999252 304977 999255
rect 304911 999250 305184 999252
rect 304911 999194 304916 999250
rect 304972 999194 305184 999250
rect 304911 999192 305184 999194
rect 304911 999189 304977 999192
rect 314799 997772 314865 997775
rect 314496 997770 314865 997772
rect 314496 997714 314804 997770
rect 314860 997714 314865 997770
rect 314496 997712 314865 997714
rect 314799 997709 314865 997712
rect 228774 996980 229374 996981
rect 227324 996882 227924 996883
rect 274875 996865 274881 997463
rect 275479 996865 275485 997463
rect 276369 996953 276375 997551
rect 276973 996953 276979 997551
rect 277775 996997 277781 997595
rect 278379 996997 278385 997595
rect 278917 996997 278923 997595
rect 279521 996997 279527 997595
rect 327774 997589 328374 1022084
rect 329332 1021934 329932 1030860
rect 298142 997533 298244 997550
rect 298142 997463 298157 997533
rect 298227 997463 298244 997533
rect 298142 997450 298244 997463
rect 280239 997180 280305 997183
rect 298095 997180 298161 997183
rect 280239 997178 298161 997180
rect 280239 997122 280244 997178
rect 280300 997122 298100 997178
rect 298156 997122 298161 997178
rect 280239 997120 298161 997122
rect 280239 997117 280305 997120
rect 298095 997117 298161 997120
rect 313743 997180 313809 997183
rect 313743 997178 313920 997180
rect 313743 997122 313748 997178
rect 313804 997122 313920 997178
rect 313743 997120 313920 997122
rect 313743 997117 313809 997120
rect 277780 996996 278380 996997
rect 278922 996996 279522 996997
rect 327769 996991 327775 997589
rect 328373 996991 328379 997589
rect 329332 997441 329932 1021334
rect 330888 1021362 331488 1031066
rect 330888 997545 331488 1020762
rect 332436 1020700 333036 1031066
rect 332436 997603 333036 1020100
rect 377196 1022758 377796 1030722
rect 353391 1015976 353457 1015979
rect 353391 1015974 355326 1015976
rect 353391 1015918 353396 1015974
rect 353452 1015918 355326 1015974
rect 353391 1015916 355326 1015918
rect 353391 1015913 353457 1015916
rect 354498 1015798 354558 1015916
rect 355266 1015828 355326 1015916
rect 355266 1015768 355680 1015828
rect 349647 1007836 349713 1007839
rect 353295 1007836 353361 1007839
rect 349647 1007834 353361 1007836
rect 349647 1007778 349652 1007834
rect 349708 1007778 353300 1007834
rect 353356 1007778 353361 1007834
rect 349647 1007776 353361 1007778
rect 349647 1007773 349713 1007776
rect 353295 1007773 353361 1007776
rect 359055 1003248 359121 1003251
rect 362511 1003248 362577 1003251
rect 358944 1003246 359121 1003248
rect 358944 1003190 359060 1003246
rect 359116 1003190 359121 1003246
rect 358944 1003188 359121 1003190
rect 362208 1003246 362577 1003248
rect 362208 1003190 362516 1003246
rect 362572 1003190 362577 1003246
rect 362208 1003188 362577 1003190
rect 359055 1003185 359121 1003188
rect 362511 1003185 362577 1003188
rect 361263 1002656 361329 1002659
rect 361056 1002654 361329 1002656
rect 361056 1002598 361268 1002654
rect 361324 1002598 361329 1002654
rect 361056 1002596 361329 1002598
rect 361263 1002593 361329 1002596
rect 361839 1002508 361905 1002511
rect 361632 1002506 361905 1002508
rect 361632 1002450 361844 1002506
rect 361900 1002450 361905 1002506
rect 361632 1002448 361905 1002450
rect 361839 1002445 361905 1002448
rect 362895 1002360 362961 1002363
rect 363471 1002360 363537 1002363
rect 362688 1002358 362961 1002360
rect 362688 1002302 362900 1002358
rect 362956 1002302 362961 1002358
rect 362688 1002300 362961 1002302
rect 363264 1002358 363537 1002360
rect 363264 1002302 363476 1002358
rect 363532 1002302 363537 1002358
rect 363264 1002300 363537 1002302
rect 362895 1002297 362961 1002300
rect 363471 1002297 363537 1002300
rect 356367 1000880 356433 1000883
rect 360207 1000880 360273 1000883
rect 356160 1000878 356433 1000880
rect 356160 1000822 356372 1000878
rect 356428 1000822 356433 1000878
rect 356160 1000820 356433 1000822
rect 360000 1000878 360273 1000880
rect 360000 1000822 360212 1000878
rect 360268 1000822 360273 1000878
rect 360000 1000820 360273 1000822
rect 356367 1000817 356433 1000820
rect 360207 1000817 360273 1000820
rect 357039 999400 357105 999403
rect 356736 999398 357105 999400
rect 356736 999342 357044 999398
rect 357100 999342 357105 999398
rect 356736 999340 357105 999342
rect 357039 999337 357105 999340
rect 364527 999252 364593 999255
rect 364320 999250 364593 999252
rect 364320 999194 364532 999250
rect 364588 999194 364593 999250
rect 364320 999192 364593 999194
rect 364527 999189 364593 999192
rect 365199 997772 365265 997775
rect 365199 997770 365472 997772
rect 365199 997714 365204 997770
rect 365260 997714 365472 997770
rect 365199 997712 365472 997714
rect 365199 997709 365265 997712
rect 377196 997605 377796 1022158
rect 378530 1022096 379130 1031376
rect 378530 997619 379130 1021496
rect 380080 1021254 380680 1031106
rect 327774 996990 328374 996991
rect 276374 996952 276974 996953
rect 274880 996864 275480 996865
rect 329327 996843 329333 997441
rect 329931 996843 329937 997441
rect 330883 996947 330889 997545
rect 331487 996947 331493 997545
rect 332431 997005 332437 997603
rect 333035 997005 333041 997603
rect 377191 997007 377197 997605
rect 377795 997007 377801 997605
rect 378525 997021 378531 997619
rect 379129 997021 379135 997619
rect 380080 997595 380680 1020654
rect 381548 1020680 382148 1031544
rect 381548 997609 382148 1020080
rect 410146 1022632 410746 1030668
rect 378530 997020 379130 997021
rect 377196 997006 377796 997007
rect 332436 997004 333036 997005
rect 380075 996997 380081 997595
rect 380679 996997 380685 997595
rect 381543 997011 381549 997609
rect 382147 997011 382153 997609
rect 410146 997425 410746 1022032
rect 412148 1021702 412748 1030018
rect 381548 997010 382148 997011
rect 380080 996996 380680 996997
rect 330888 996946 331488 996947
rect 329332 996842 329932 996843
rect 410141 996827 410147 997425
rect 410745 996827 410751 997425
rect 412148 997413 412748 1021102
rect 414358 1021156 414958 1030152
rect 414358 997531 414958 1020556
rect 415922 1020566 416522 1030350
rect 415922 997547 416522 1019966
rect 491650 1022572 492250 1031710
rect 421410 1015916 422526 1015976
rect 421410 1015798 421470 1015916
rect 422466 1015798 422526 1015916
rect 435183 1005912 435249 1005915
rect 465711 1005912 465777 1005915
rect 435183 1005910 465777 1005912
rect 435183 1005854 435188 1005910
rect 435244 1005854 465716 1005910
rect 465772 1005854 465777 1005910
rect 435183 1005852 465777 1005854
rect 435183 1005849 435249 1005852
rect 465711 1005849 465777 1005852
rect 435087 1005172 435153 1005175
rect 443535 1005172 443601 1005175
rect 435087 1005170 443601 1005172
rect 435087 1005114 435092 1005170
rect 435148 1005114 443540 1005170
rect 443596 1005114 443601 1005170
rect 435087 1005112 443601 1005114
rect 435087 1005109 435153 1005112
rect 443535 1005109 443601 1005112
rect 426063 1003248 426129 1003251
rect 429231 1003248 429297 1003251
rect 425760 1003246 426129 1003248
rect 425760 1003190 426068 1003246
rect 426124 1003190 426129 1003246
rect 425760 1003188 426129 1003190
rect 429024 1003246 429297 1003248
rect 429024 1003190 429236 1003246
rect 429292 1003190 429297 1003246
rect 429024 1003188 429297 1003190
rect 426063 1003185 426129 1003188
rect 429231 1003185 429297 1003188
rect 425391 1003100 425457 1003103
rect 430287 1003100 430353 1003103
rect 425184 1003098 425457 1003100
rect 425184 1003042 425396 1003098
rect 425452 1003042 425457 1003098
rect 425184 1003040 425457 1003042
rect 430176 1003098 430353 1003100
rect 430176 1003042 430292 1003098
rect 430348 1003042 430353 1003098
rect 430176 1003040 430353 1003042
rect 425391 1003037 425457 1003040
rect 430287 1003037 430353 1003040
rect 424335 1002952 424401 1002955
rect 428751 1002952 428817 1002955
rect 424128 1002950 424401 1002952
rect 424128 1002894 424340 1002950
rect 424396 1002894 424401 1002950
rect 424128 1002892 424401 1002894
rect 428448 1002950 428817 1002952
rect 428448 1002894 428756 1002950
rect 428812 1002894 428817 1002950
rect 428448 1002892 428817 1002894
rect 424335 1002889 424401 1002892
rect 428751 1002889 428817 1002892
rect 423759 1002804 423825 1002807
rect 428271 1002804 428337 1002807
rect 423648 1002802 423825 1002804
rect 423648 1002746 423764 1002802
rect 423820 1002746 423825 1002802
rect 423648 1002744 423825 1002746
rect 427968 1002802 428337 1002804
rect 427968 1002746 428276 1002802
rect 428332 1002746 428337 1002802
rect 427968 1002744 428337 1002746
rect 423759 1002741 423825 1002744
rect 428271 1002741 428337 1002744
rect 424815 1002656 424881 1002659
rect 427695 1002656 427761 1002659
rect 424704 1002654 424881 1002656
rect 424704 1002598 424820 1002654
rect 424876 1002598 424881 1002654
rect 424704 1002596 424881 1002598
rect 427392 1002654 427761 1002656
rect 427392 1002598 427700 1002654
rect 427756 1002598 427761 1002654
rect 427392 1002596 427761 1002598
rect 424815 1002593 424881 1002596
rect 427695 1002593 427761 1002596
rect 426639 1002508 426705 1002511
rect 427119 1002508 427185 1002511
rect 426336 1002506 426705 1002508
rect 426336 1002450 426644 1002506
rect 426700 1002450 426705 1002506
rect 426336 1002448 426705 1002450
rect 426912 1002506 427185 1002508
rect 426912 1002450 427124 1002506
rect 427180 1002450 427185 1002506
rect 426912 1002448 427185 1002450
rect 426639 1002445 426705 1002448
rect 427119 1002445 427185 1002448
rect 431919 1002360 431985 1002363
rect 431712 1002358 431985 1002360
rect 431712 1002302 431924 1002358
rect 431980 1002302 431985 1002358
rect 431712 1002300 431985 1002302
rect 431919 1002297 431985 1002300
rect 429903 1000880 429969 1000883
rect 430959 1000880 431025 1000883
rect 429600 1000878 429969 1000880
rect 429600 1000822 429908 1000878
rect 429964 1000822 429969 1000878
rect 429600 1000820 429969 1000822
rect 430656 1000878 431025 1000880
rect 430656 1000822 430964 1000878
rect 431020 1000822 431025 1000878
rect 430656 1000820 431025 1000822
rect 429903 1000817 429969 1000820
rect 430959 1000817 431025 1000820
rect 410146 996826 410746 996827
rect 412143 996815 412149 997413
rect 412747 996815 412753 997413
rect 414353 996933 414359 997531
rect 414957 996933 414963 997531
rect 415917 996949 415923 997547
rect 416521 996949 416527 997547
rect 491650 997381 492250 1021972
rect 493070 1021882 493670 1031664
rect 493070 997381 493670 1021282
rect 494582 1021166 495182 1031852
rect 494582 997523 495182 1020566
rect 496096 1020550 496696 1031616
rect 496096 997571 496696 1019950
rect 568178 1022764 568778 1029852
rect 499266 1015916 500094 1015976
rect 499266 1015828 499326 1015916
rect 498912 1015768 499326 1015828
rect 500034 999400 500094 1015916
rect 501327 1003100 501393 1003103
rect 502383 1003100 502449 1003103
rect 502959 1003100 503025 1003103
rect 504015 1003100 504081 1003103
rect 501120 1003098 501393 1003100
rect 501120 1003042 501332 1003098
rect 501388 1003042 501393 1003098
rect 501120 1003040 501393 1003042
rect 502176 1003098 502449 1003100
rect 502176 1003042 502388 1003098
rect 502444 1003042 502449 1003098
rect 502176 1003040 502449 1003042
rect 502752 1003098 503025 1003100
rect 502752 1003042 502964 1003098
rect 503020 1003042 503025 1003098
rect 502752 1003040 503025 1003042
rect 503904 1003098 504081 1003100
rect 503904 1003042 504020 1003098
rect 504076 1003042 504081 1003098
rect 503904 1003040 504081 1003042
rect 501327 1003037 501393 1003040
rect 502383 1003037 502449 1003040
rect 502959 1003037 503025 1003040
rect 504015 1003037 504081 1003040
rect 554895 1002952 554961 1002955
rect 554688 1002950 554961 1002952
rect 554688 1002894 554900 1002950
rect 554956 1002894 554961 1002950
rect 554688 1002892 554961 1002894
rect 554895 1002889 554961 1002892
rect 554319 1002804 554385 1002807
rect 554208 1002802 554385 1002804
rect 554208 1002746 554324 1002802
rect 554380 1002746 554385 1002802
rect 554208 1002744 554385 1002746
rect 554319 1002741 554385 1002744
rect 553743 1002656 553809 1002659
rect 553632 1002654 553809 1002656
rect 553632 1002598 553748 1002654
rect 553804 1002598 553809 1002654
rect 553632 1002596 553809 1002598
rect 553743 1002593 553809 1002596
rect 503439 1002360 503505 1002363
rect 553263 1002360 553329 1002363
rect 555375 1002360 555441 1002363
rect 503328 1002358 503505 1002360
rect 503328 1002302 503444 1002358
rect 503500 1002302 503505 1002358
rect 503328 1002300 503505 1002302
rect 553056 1002358 553329 1002360
rect 553056 1002302 553268 1002358
rect 553324 1002302 553329 1002358
rect 553056 1002300 553329 1002302
rect 555264 1002358 555441 1002360
rect 555264 1002302 555380 1002358
rect 555436 1002302 555441 1002358
rect 555264 1002300 555441 1002302
rect 503439 1002297 503505 1002300
rect 553263 1002297 553329 1002300
rect 555375 1002297 555441 1002300
rect 506223 1001472 506289 1001475
rect 506016 1001470 506289 1001472
rect 506016 1001414 506228 1001470
rect 506284 1001414 506289 1001470
rect 506016 1001412 506289 1001414
rect 506223 1001409 506289 1001412
rect 557775 1001324 557841 1001327
rect 557472 1001322 557841 1001324
rect 557472 1001266 557780 1001322
rect 557836 1001266 557841 1001322
rect 557472 1001264 557841 1001266
rect 557775 1001261 557841 1001264
rect 507855 1001028 507921 1001031
rect 507648 1001026 507921 1001028
rect 507648 1000970 507860 1001026
rect 507916 1000970 507921 1001026
rect 507648 1000968 507921 1000970
rect 507855 1000965 507921 1000968
rect 512655 1001028 512721 1001031
rect 523791 1001028 523857 1001031
rect 512655 1001026 523857 1001028
rect 512655 1000970 512660 1001026
rect 512716 1000970 523796 1001026
rect 523852 1000970 523857 1001026
rect 512655 1000968 523857 1000970
rect 512655 1000965 512721 1000968
rect 523791 1000965 523857 1000968
rect 500751 1000880 500817 1000883
rect 500640 1000878 500817 1000880
rect 500640 1000822 500756 1000878
rect 500812 1000822 500817 1000878
rect 500640 1000820 500817 1000822
rect 500751 1000817 500817 1000820
rect 513999 1000880 514065 1000883
rect 523503 1000880 523569 1000883
rect 552303 1000880 552369 1000883
rect 552879 1000880 552945 1000883
rect 513999 1000878 523569 1000880
rect 513999 1000822 514004 1000878
rect 514060 1000822 523508 1000878
rect 523564 1000822 523569 1000878
rect 513999 1000820 523569 1000822
rect 552000 1000878 552369 1000880
rect 552000 1000822 552308 1000878
rect 552364 1000822 552369 1000878
rect 552000 1000820 552369 1000822
rect 552480 1000878 552945 1000880
rect 552480 1000822 552884 1000878
rect 552940 1000822 552945 1000878
rect 552480 1000820 552945 1000822
rect 513999 1000817 514065 1000820
rect 523503 1000817 523569 1000820
rect 552303 1000817 552369 1000820
rect 552879 1000817 552945 1000820
rect 506895 1000732 506961 1000735
rect 506592 1000730 506961 1000732
rect 506592 1000674 506900 1000730
rect 506956 1000674 506961 1000730
rect 506592 1000672 506961 1000674
rect 506895 1000669 506961 1000672
rect 512079 1000732 512145 1000735
rect 523983 1000732 524049 1000735
rect 512079 1000730 524049 1000732
rect 512079 1000674 512084 1000730
rect 512140 1000674 523988 1000730
rect 524044 1000674 524049 1000730
rect 512079 1000672 524049 1000674
rect 512079 1000669 512145 1000672
rect 523983 1000669 524049 1000672
rect 518415 999844 518481 999847
rect 523887 999844 523953 999847
rect 518415 999842 523953 999844
rect 518415 999786 518420 999842
rect 518476 999786 523892 999842
rect 523948 999786 523953 999842
rect 518415 999784 523953 999786
rect 518415 999781 518481 999784
rect 523887 999781 523953 999784
rect 501999 999696 502065 999699
rect 501696 999694 502065 999696
rect 501696 999638 502004 999694
rect 502060 999638 502065 999694
rect 501696 999636 502065 999638
rect 501999 999633 502065 999636
rect 512079 999696 512145 999699
rect 523695 999696 523761 999699
rect 512079 999694 523761 999696
rect 512079 999638 512084 999694
rect 512140 999638 523700 999694
rect 523756 999638 523761 999694
rect 512079 999636 523761 999638
rect 512079 999633 512145 999636
rect 523695 999633 523761 999636
rect 504687 999548 504753 999551
rect 504384 999546 504753 999548
rect 504384 999490 504692 999546
rect 504748 999490 504753 999546
rect 504384 999488 504753 999490
rect 504687 999485 504753 999488
rect 512079 999548 512145 999551
rect 524079 999548 524145 999551
rect 512079 999546 524145 999548
rect 512079 999490 512084 999546
rect 512140 999490 524084 999546
rect 524140 999490 524145 999546
rect 512079 999488 524145 999490
rect 512079 999485 512145 999488
rect 524079 999485 524145 999488
rect 500175 999400 500241 999403
rect 500034 999398 500241 999400
rect 500034 999370 500180 999398
rect 500064 999342 500180 999370
rect 500236 999342 500241 999398
rect 500064 999340 500241 999342
rect 500175 999337 500241 999340
rect 518511 999400 518577 999403
rect 523599 999400 523665 999403
rect 518511 999398 523665 999400
rect 518511 999342 518516 999398
rect 518572 999342 523604 999398
rect 523660 999342 523665 999398
rect 518511 999340 523665 999342
rect 518511 999337 518577 999340
rect 523599 999337 523665 999340
rect 557199 999104 557265 999107
rect 556896 999102 557265 999104
rect 556896 999046 557204 999102
rect 557260 999046 557265 999102
rect 556896 999044 557265 999046
rect 557199 999041 557265 999044
rect 558831 998956 558897 998959
rect 558528 998954 558897 998956
rect 558528 998898 558836 998954
rect 558892 998898 558897 998954
rect 558528 998896 558897 998898
rect 558831 998893 558897 998896
rect 555951 997772 556017 997775
rect 555744 997770 556017 997772
rect 555744 997714 555956 997770
rect 556012 997714 556017 997770
rect 555744 997712 556017 997714
rect 555951 997709 556017 997712
rect 415922 996948 416522 996949
rect 414358 996932 414958 996933
rect 412148 996814 412748 996815
rect 491645 996783 491651 997381
rect 492249 996783 492255 997381
rect 493065 996783 493071 997381
rect 493669 996783 493675 997381
rect 494577 996925 494583 997523
rect 495181 996925 495187 997523
rect 496091 996973 496097 997571
rect 496695 996973 496701 997571
rect 558159 997476 558225 997479
rect 557952 997474 558225 997476
rect 557952 997418 558164 997474
rect 558220 997418 558225 997474
rect 568178 997451 568778 1022164
rect 570328 1022042 570928 1030392
rect 570328 997543 570928 1021442
rect 571834 1021444 572434 1030832
rect 571834 997585 572434 1020844
rect 573446 1020596 574046 1031176
rect 557952 997416 558225 997418
rect 558159 997413 558225 997416
rect 559407 997328 559473 997331
rect 559008 997326 559473 997328
rect 559008 997270 559412 997326
rect 559468 997270 559473 997326
rect 559008 997268 559473 997270
rect 559407 997265 559473 997268
rect 496096 996972 496696 996973
rect 494582 996924 495182 996925
rect 568173 996853 568179 997451
rect 568777 996853 568783 997451
rect 570323 996945 570329 997543
rect 570927 996945 570933 997543
rect 571829 996987 571835 997585
rect 572433 996987 572439 997585
rect 573446 997527 574046 1019996
rect 571834 996986 572434 996987
rect 570328 996944 570928 996945
rect 573441 996929 573447 997527
rect 574045 996929 574051 997527
rect 576108 997132 580206 997948
rect 585714 997132 589812 997914
rect 576108 997072 589812 997132
rect 573446 996928 574046 996929
rect 568178 996852 568778 996853
rect 491650 996782 492250 996783
rect 493070 996782 493670 996783
rect 298120 996745 298240 996766
rect 225484 996706 226084 996707
rect 298120 996675 298159 996745
rect 298229 996675 298240 996745
rect 298120 996664 298240 996675
rect 156015 996588 156081 996591
rect 205263 996588 205329 996591
rect 259983 996588 260049 996591
rect 505647 996588 505713 996591
rect 507279 996588 507345 996591
rect 156015 996586 156288 996588
rect 156015 996530 156020 996586
rect 156076 996530 156288 996586
rect 156015 996528 156288 996530
rect 205263 996586 205536 996588
rect 205263 996530 205268 996586
rect 205324 996530 205536 996586
rect 205263 996528 205536 996530
rect 259983 996586 260160 996588
rect 259983 996530 259988 996586
rect 260044 996530 260160 996586
rect 259983 996528 260160 996530
rect 505440 996586 505713 996588
rect 505440 996530 505652 996586
rect 505708 996530 505713 996586
rect 505440 996528 505713 996530
rect 507168 996586 507345 996588
rect 507168 996530 507284 996586
rect 507340 996530 507345 996586
rect 507168 996528 507345 996530
rect 156015 996525 156081 996528
rect 205263 996525 205329 996528
rect 259983 996525 260049 996528
rect 505647 996525 505713 996528
rect 507279 996525 507345 996528
rect 262095 996292 262161 996295
rect 432591 996292 432657 996295
rect 508335 996292 508401 996295
rect 262095 996290 262368 996292
rect 262095 996234 262100 996290
rect 262156 996234 262368 996290
rect 262095 996232 262368 996234
rect 432591 996290 432864 996292
rect 432591 996234 432596 996290
rect 432652 996234 432864 996290
rect 432591 996232 432864 996234
rect 508224 996290 508401 996292
rect 508224 996234 508340 996290
rect 508396 996234 508401 996290
rect 508224 996232 508401 996234
rect 262095 996229 262161 996232
rect 432591 996229 432657 996232
rect 508335 996229 508401 996232
rect 159183 996144 159249 996147
rect 159759 996144 159825 996147
rect 158976 996142 159249 996144
rect 158976 996086 159188 996142
rect 159244 996086 159249 996142
rect 158976 996084 159249 996086
rect 159552 996142 159825 996144
rect 159552 996086 159764 996142
rect 159820 996086 159825 996142
rect 159552 996084 159825 996086
rect 159183 996081 159249 996084
rect 159759 996081 159825 996084
rect 204015 996144 204081 996147
rect 210159 996144 210225 996147
rect 261999 996144 262065 996147
rect 263055 996144 263121 996147
rect 204015 996142 204384 996144
rect 204015 996086 204020 996142
rect 204076 996086 204384 996142
rect 204015 996084 204384 996086
rect 210159 996142 210432 996144
rect 210159 996086 210164 996142
rect 210220 996086 210432 996142
rect 210159 996084 210432 996086
rect 261792 996142 262065 996144
rect 261792 996086 262004 996142
rect 262060 996086 262065 996142
rect 261792 996084 262065 996086
rect 262944 996142 263121 996144
rect 262944 996086 263060 996142
rect 263116 996086 263121 996142
rect 262944 996084 263121 996086
rect 204015 996081 204081 996084
rect 210159 996081 210225 996084
rect 261999 996081 262065 996084
rect 263055 996081 263121 996084
rect 313167 996144 313233 996147
rect 314799 996144 314865 996147
rect 432495 996144 432561 996147
rect 313167 996142 313440 996144
rect 313167 996086 313172 996142
rect 313228 996086 313440 996142
rect 313167 996084 313440 996086
rect 314799 996142 314976 996144
rect 314799 996086 314804 996142
rect 314860 996086 314976 996142
rect 314799 996084 314976 996086
rect 432288 996142 432561 996144
rect 432288 996086 432500 996142
rect 432556 996086 432561 996142
rect 432288 996084 432561 996086
rect 313167 996081 313233 996084
rect 314799 996081 314865 996084
rect 432495 996081 432561 996084
rect 463695 996144 463761 996147
rect 476602 996144 476608 996146
rect 463695 996142 476608 996144
rect 463695 996086 463700 996142
rect 463756 996086 476608 996142
rect 463695 996084 476608 996086
rect 463695 996081 463761 996084
rect 476602 996082 476608 996084
rect 476672 996082 476678 996146
rect 508527 996144 508593 996147
rect 509583 996144 509649 996147
rect 561039 996144 561105 996147
rect 508527 996142 508704 996144
rect 508527 996086 508532 996142
rect 508588 996086 508704 996142
rect 508527 996084 508704 996086
rect 509583 996142 509856 996144
rect 509583 996086 509588 996142
rect 509644 996086 509856 996142
rect 509583 996084 509856 996086
rect 561039 996142 561216 996144
rect 561039 996086 561044 996142
rect 561100 996086 561216 996142
rect 561039 996084 561216 996086
rect 508527 996081 508593 996084
rect 509583 996081 509649 996084
rect 561039 996081 561105 996084
rect 576108 996004 580256 997072
rect 585666 996004 589812 997072
rect 576108 996002 589812 996004
rect 99567 995996 99633 995999
rect 102927 995996 102993 995999
rect 108975 995996 109041 995999
rect 99567 995994 99936 995996
rect 99567 995938 99572 995994
rect 99628 995938 99936 995994
rect 99567 995936 99936 995938
rect 102927 995994 103200 995996
rect 102927 995938 102932 995994
rect 102988 995938 103200 995994
rect 102927 995936 103200 995938
rect 108672 995994 109041 995996
rect 108672 995938 108980 995994
rect 109036 995938 109041 995994
rect 108672 995936 109041 995938
rect 99567 995933 99633 995936
rect 102927 995933 102993 995936
rect 108975 995933 109041 995936
rect 109551 995996 109617 995999
rect 152079 995996 152145 995999
rect 160431 995996 160497 995999
rect 198639 995996 198705 995999
rect 109551 995994 109728 995996
rect 109551 995938 109556 995994
rect 109612 995938 109728 995994
rect 109551 995936 109728 995938
rect 150018 995936 150240 995996
rect 152079 995994 152448 995996
rect 152079 995938 152084 995994
rect 152140 995938 152448 995994
rect 152079 995936 152448 995938
rect 160431 995994 160608 995996
rect 160431 995938 160436 995994
rect 160492 995938 160608 995994
rect 160431 995936 160608 995938
rect 189186 995994 198705 995996
rect 189186 995938 198644 995994
rect 198700 995938 198705 995994
rect 189186 995936 198705 995938
rect 109551 995933 109617 995936
rect 102447 995848 102513 995851
rect 104463 995848 104529 995851
rect 107919 995848 107985 995851
rect 126639 995848 126705 995851
rect 134319 995848 134385 995851
rect 97935 995846 98430 995848
rect 81039 995788 95025 995790
rect 81039 995785 81105 995788
rect 94959 995785 95025 995788
rect 85935 995700 86001 995703
rect 97794 995700 97854 995818
rect 97935 995790 97940 995846
rect 97996 995818 98430 995846
rect 97996 995790 98400 995818
rect 97935 995788 98400 995790
rect 97935 995785 98001 995788
rect 98850 995700 98910 995818
rect 85935 995698 94014 995700
rect 85935 995642 85940 995698
rect 85996 995642 94014 995698
rect 85935 995640 94014 995642
rect 97794 995640 98910 995700
rect 98991 995700 99057 995703
rect 100482 995700 100542 995818
rect 98991 995698 100542 995700
rect 98991 995642 98996 995698
rect 99052 995642 100542 995698
rect 98991 995640 100542 995642
rect 85935 995637 86001 995640
rect 85359 995404 85425 995407
rect 93807 995404 93873 995407
rect 85359 995402 93873 995404
rect 85359 995346 85364 995402
rect 85420 995346 93812 995402
rect 93868 995346 93873 995402
rect 85359 995344 93873 995346
rect 93954 995404 94014 995640
rect 98991 995637 99057 995640
rect 97839 995552 97905 995555
rect 101058 995552 101118 995818
rect 97839 995550 101118 995552
rect 97839 995494 97844 995550
rect 97900 995494 101118 995550
rect 97839 995492 101118 995494
rect 101442 995788 101664 995848
rect 102447 995846 102720 995848
rect 97839 995489 97905 995492
rect 101442 995404 101502 995788
rect 93954 995344 101502 995404
rect 85359 995341 85425 995344
rect 93807 995341 93873 995344
rect 86415 995256 86481 995259
rect 99567 995256 99633 995259
rect 86415 995254 99633 995256
rect 86415 995198 86420 995254
rect 86476 995198 99572 995254
rect 99628 995198 99633 995254
rect 86415 995196 99633 995198
rect 86415 995193 86481 995196
rect 99567 995193 99633 995196
rect 87759 995108 87825 995111
rect 102114 995108 102174 995818
rect 102447 995790 102452 995846
rect 102508 995790 102720 995846
rect 104463 995846 104928 995848
rect 102447 995788 102720 995790
rect 102447 995785 102513 995788
rect 87759 995106 102174 995108
rect 87759 995050 87764 995106
rect 87820 995050 102174 995106
rect 87759 995048 102174 995050
rect 87759 995045 87825 995048
rect 97839 994960 97905 994963
rect 103746 994960 103806 995818
rect 104463 995790 104468 995846
rect 104524 995790 104928 995846
rect 107919 995846 108192 995848
rect 104463 995788 104928 995790
rect 104463 995785 104529 995788
rect 105378 995259 105438 995818
rect 105954 995407 106014 995818
rect 105903 995402 106014 995407
rect 105903 995346 105908 995402
rect 105964 995346 106014 995402
rect 105903 995344 106014 995346
rect 105903 995341 105969 995344
rect 107010 995259 107070 995818
rect 107586 995555 107646 995818
rect 107919 995790 107924 995846
rect 107980 995790 108192 995846
rect 126639 995846 134385 995848
rect 107919 995788 108192 995790
rect 107919 995785 107985 995788
rect 109218 995555 109278 995818
rect 107535 995550 107646 995555
rect 107535 995494 107540 995550
rect 107596 995494 107646 995550
rect 107535 995492 107646 995494
rect 109167 995550 109278 995555
rect 109167 995494 109172 995550
rect 109228 995494 109278 995550
rect 109167 995492 109278 995494
rect 107535 995489 107601 995492
rect 109167 995489 109233 995492
rect 110274 995259 110334 995818
rect 105327 995254 105438 995259
rect 105327 995198 105332 995254
rect 105388 995198 105438 995254
rect 105327 995196 105438 995198
rect 106959 995254 107070 995259
rect 106959 995198 106964 995254
rect 107020 995198 107070 995254
rect 106959 995196 107070 995198
rect 110223 995254 110334 995259
rect 110223 995198 110228 995254
rect 110284 995198 110334 995254
rect 110223 995196 110334 995198
rect 105327 995193 105393 995196
rect 106959 995193 107025 995196
rect 110223 995193 110289 995196
rect 109359 995108 109425 995111
rect 110850 995108 110910 995818
rect 126639 995790 126644 995846
rect 126700 995790 134324 995846
rect 134380 995790 134385 995846
rect 126639 995788 134385 995790
rect 126639 995785 126705 995788
rect 134319 995785 134385 995788
rect 136143 995848 136209 995851
rect 144111 995848 144177 995851
rect 136143 995846 144177 995848
rect 136143 995790 136148 995846
rect 136204 995790 144116 995846
rect 144172 995790 144177 995846
rect 136143 995788 144177 995790
rect 136143 995785 136209 995788
rect 144111 995785 144177 995788
rect 149154 995700 149214 995818
rect 150018 995700 150078 995936
rect 152079 995933 152145 995936
rect 160431 995933 160497 995936
rect 151695 995848 151761 995851
rect 154863 995848 154929 995851
rect 158223 995848 158289 995851
rect 161487 995848 161553 995851
rect 188751 995848 188817 995851
rect 189186 995848 189246 995936
rect 198639 995933 198705 995936
rect 207375 995996 207441 995999
rect 210639 995996 210705 995999
rect 211791 995996 211857 995999
rect 219087 995996 219153 995999
rect 246927 995996 246993 995999
rect 207375 995994 207648 995996
rect 207375 995938 207380 995994
rect 207436 995938 207648 995994
rect 207375 995936 207648 995938
rect 210639 995994 210912 995996
rect 210639 995938 210644 995994
rect 210700 995938 210912 995994
rect 210639 995936 210912 995938
rect 211791 995994 212064 995996
rect 211791 995938 211796 995994
rect 211852 995938 212064 995994
rect 211791 995936 212064 995938
rect 212640 995936 212862 995996
rect 213696 995994 219153 995996
rect 213696 995938 219092 995994
rect 219148 995938 219153 995994
rect 213696 995936 219153 995938
rect 207375 995933 207441 995936
rect 210639 995933 210705 995936
rect 211791 995933 211857 995936
rect 151695 995846 151968 995848
rect 151695 995790 151700 995846
rect 151756 995790 151968 995846
rect 151695 995788 151968 995790
rect 153504 995788 153726 995848
rect 154863 995846 155232 995848
rect 151695 995785 151761 995788
rect 153666 995700 153726 995788
rect 149154 995640 150078 995700
rect 153474 995640 153726 995700
rect 139215 995552 139281 995555
rect 153474 995552 153534 995640
rect 139215 995550 153534 995552
rect 139215 995494 139220 995550
rect 139276 995494 153534 995550
rect 139215 995492 153534 995494
rect 139215 995489 139281 995492
rect 144687 995404 144753 995407
rect 154050 995404 154110 995818
rect 144687 995402 154110 995404
rect 144687 995346 144692 995402
rect 144748 995346 154110 995402
rect 144687 995344 154110 995346
rect 144687 995341 144753 995344
rect 149679 995256 149745 995259
rect 154626 995256 154686 995818
rect 154863 995790 154868 995846
rect 154924 995790 155232 995846
rect 154863 995788 155232 995790
rect 156768 995788 156990 995848
rect 158223 995846 158496 995848
rect 154863 995785 154929 995788
rect 156930 995700 156990 995788
rect 156738 995640 156990 995700
rect 154767 995404 154833 995407
rect 156738 995404 156798 995640
rect 154767 995402 156798 995404
rect 154767 995346 154772 995402
rect 154828 995346 156798 995402
rect 154767 995344 156798 995346
rect 154767 995341 154833 995344
rect 157314 995259 157374 995818
rect 158223 995790 158228 995846
rect 158284 995790 158496 995846
rect 158223 995788 158496 995790
rect 161487 995846 161760 995848
rect 161487 995790 161492 995846
rect 161548 995790 161760 995846
rect 188751 995846 189246 995848
rect 161487 995788 161760 995790
rect 158223 995785 158289 995788
rect 161487 995785 161553 995788
rect 149679 995254 154686 995256
rect 149679 995198 149684 995254
rect 149740 995198 154686 995254
rect 149679 995196 154686 995198
rect 157263 995254 157374 995259
rect 157263 995198 157268 995254
rect 157324 995198 157374 995254
rect 157263 995196 157374 995198
rect 161679 995256 161745 995259
rect 162210 995256 162270 995818
rect 188751 995790 188756 995846
rect 188812 995790 189246 995846
rect 188751 995788 189246 995790
rect 189423 995848 189489 995851
rect 198639 995848 198705 995851
rect 202479 995848 202545 995851
rect 202959 995848 203025 995851
rect 205647 995848 205713 995851
rect 189423 995846 198705 995848
rect 189423 995790 189428 995846
rect 189484 995790 198644 995846
rect 198700 995790 198705 995846
rect 189423 995788 198705 995790
rect 201120 995788 201534 995848
rect 202479 995846 202848 995848
rect 188751 995785 188817 995788
rect 189423 995785 189489 995788
rect 198639 995785 198705 995788
rect 197199 995700 197265 995703
rect 201474 995700 201534 995788
rect 202242 995700 202302 995818
rect 202479 995790 202484 995846
rect 202540 995790 202848 995846
rect 202479 995788 202848 995790
rect 202959 995846 203328 995848
rect 202959 995790 202964 995846
rect 203020 995790 203328 995846
rect 205647 995846 206112 995848
rect 202959 995788 203328 995790
rect 202479 995785 202545 995788
rect 202959 995785 203025 995788
rect 197199 995698 202302 995700
rect 197199 995642 197204 995698
rect 197260 995642 202302 995698
rect 197199 995640 202302 995642
rect 197199 995637 197265 995640
rect 188079 995552 188145 995555
rect 198447 995552 198513 995555
rect 188079 995550 198513 995552
rect 188079 995494 188084 995550
rect 188140 995494 198452 995550
rect 198508 995494 198513 995550
rect 188079 995492 198513 995494
rect 188079 995489 188145 995492
rect 198447 995489 198513 995492
rect 198639 995552 198705 995555
rect 203874 995552 203934 995818
rect 198639 995550 203934 995552
rect 198639 995494 198644 995550
rect 198700 995494 203934 995550
rect 198639 995492 203934 995494
rect 198639 995489 198705 995492
rect 190575 995404 190641 995407
rect 204930 995404 204990 995818
rect 205647 995790 205652 995846
rect 205708 995790 206112 995846
rect 205647 995788 206112 995790
rect 205647 995785 205713 995788
rect 190575 995402 204990 995404
rect 190575 995346 190580 995402
rect 190636 995346 204990 995402
rect 190575 995344 204990 995346
rect 190575 995341 190641 995344
rect 161679 995254 162270 995256
rect 161679 995198 161684 995254
rect 161740 995198 162270 995254
rect 161679 995196 162270 995198
rect 198639 995256 198705 995259
rect 206562 995256 206622 995818
rect 208194 995259 208254 995818
rect 208770 995259 208830 995818
rect 209826 995259 209886 995818
rect 212802 995700 212862 995936
rect 219087 995933 219153 995936
rect 243330 995994 246993 995996
rect 243330 995938 246932 995994
rect 246988 995938 246993 995994
rect 243330 995936 246993 995938
rect 213327 995848 213393 995851
rect 213120 995846 213393 995848
rect 213120 995790 213332 995846
rect 213388 995790 213393 995846
rect 213120 995788 213393 995790
rect 213327 995785 213393 995788
rect 243183 995848 243249 995851
rect 243330 995848 243390 995936
rect 246927 995933 246993 995936
rect 254511 995996 254577 995999
rect 257679 995996 257745 995999
rect 263247 995996 263313 995999
rect 303951 995996 304017 995999
rect 254511 995994 254688 995996
rect 254511 995938 254516 995994
rect 254572 995938 254688 995994
rect 254511 995936 254688 995938
rect 257679 995994 257952 995996
rect 257679 995938 257684 995994
rect 257740 995938 257952 995994
rect 257679 995936 257952 995938
rect 263247 995994 263424 995996
rect 263247 995938 263252 995994
rect 263308 995938 263424 995994
rect 263247 995936 263424 995938
rect 303648 995994 304017 995996
rect 303648 995938 303956 995994
rect 304012 995938 304017 995994
rect 303648 995936 304017 995938
rect 254511 995933 254577 995936
rect 257679 995933 257745 995936
rect 263247 995933 263313 995936
rect 303951 995933 304017 995936
rect 304335 995996 304401 995999
rect 311535 995996 311601 995999
rect 319599 995996 319665 995999
rect 363951 995996 364017 995999
rect 304335 995994 304704 995996
rect 304335 995938 304340 995994
rect 304396 995938 304704 995994
rect 304335 995936 304704 995938
rect 311535 995994 311712 995996
rect 311535 995938 311540 995994
rect 311596 995938 311712 995994
rect 311535 995936 311712 995938
rect 316704 995994 319665 995996
rect 316704 995938 319604 995994
rect 319660 995938 319665 995994
rect 316704 995936 319665 995938
rect 363744 995994 364017 995996
rect 363744 995938 363956 995994
rect 364012 995938 364017 995994
rect 363744 995936 364017 995938
rect 304335 995933 304401 995936
rect 311535 995933 311601 995936
rect 319599 995933 319665 995936
rect 363951 995933 364017 995936
rect 430959 995996 431025 995999
rect 437871 995996 437937 995999
rect 430959 995994 431232 995996
rect 430959 995938 430964 995994
rect 431020 995938 431232 995994
rect 430959 995936 431232 995938
rect 434496 995994 437937 995996
rect 434496 995938 437876 995994
rect 437932 995938 437937 995994
rect 434496 995936 437937 995938
rect 430959 995933 431025 995936
rect 437871 995933 437937 995936
rect 467823 995996 467889 995999
rect 510543 995996 510609 995999
rect 515535 995996 515601 995999
rect 561903 995996 561969 995999
rect 467823 995994 481662 995996
rect 467823 995938 467828 995994
rect 467884 995938 481662 995994
rect 467823 995936 481662 995938
rect 510432 995994 510609 995996
rect 510432 995938 510548 995994
rect 510604 995938 510609 995994
rect 510432 995936 510609 995938
rect 511488 995994 515601 995996
rect 511488 995938 515540 995994
rect 515596 995938 515601 995994
rect 511488 995936 515601 995938
rect 561792 995994 561969 995996
rect 561792 995938 561908 995994
rect 561964 995938 561969 995994
rect 579686 995980 589812 996002
rect 585714 995968 589812 995980
rect 561792 995936 561969 995938
rect 467823 995933 467889 995936
rect 243183 995846 243390 995848
rect 243183 995790 243188 995846
rect 243244 995790 243390 995846
rect 243183 995788 243390 995790
rect 243951 995848 244017 995851
rect 246831 995848 246897 995851
rect 243951 995846 246897 995848
rect 243951 995790 243956 995846
rect 244012 995790 246836 995846
rect 246892 995790 246897 995846
rect 256143 995848 256209 995851
rect 259407 995848 259473 995851
rect 270735 995848 270801 995851
rect 256143 995846 256416 995848
rect 243951 995788 246897 995790
rect 243183 995785 243249 995788
rect 243951 995785 244017 995788
rect 246831 995785 246897 995788
rect 216015 995700 216081 995703
rect 212802 995698 216081 995700
rect 212802 995642 216020 995698
rect 216076 995642 216081 995698
rect 212802 995640 216081 995642
rect 216015 995637 216081 995640
rect 241839 995700 241905 995703
rect 247599 995700 247665 995703
rect 241839 995698 247665 995700
rect 241839 995642 241844 995698
rect 241900 995642 247604 995698
rect 247660 995642 247665 995698
rect 241839 995640 247665 995642
rect 241839 995637 241905 995640
rect 247599 995637 247665 995640
rect 247791 995700 247857 995703
rect 252546 995700 252606 995818
rect 253602 995700 253662 995818
rect 247791 995698 253662 995700
rect 247791 995642 247796 995698
rect 247852 995642 253662 995698
rect 247791 995640 253662 995642
rect 247791 995637 247857 995640
rect 236463 995552 236529 995555
rect 255234 995552 255294 995818
rect 256143 995790 256148 995846
rect 256204 995790 256416 995846
rect 259407 995846 259680 995848
rect 256143 995788 256416 995790
rect 256143 995785 256209 995788
rect 236463 995550 255294 995552
rect 236463 995494 236468 995550
rect 236524 995494 255294 995550
rect 236463 995492 255294 995494
rect 236463 995489 236529 995492
rect 238959 995404 239025 995407
rect 247023 995404 247089 995407
rect 238959 995402 247089 995404
rect 238959 995346 238964 995402
rect 239020 995346 247028 995402
rect 247084 995346 247089 995402
rect 238959 995344 247089 995346
rect 238959 995341 239025 995344
rect 247023 995341 247089 995344
rect 247599 995404 247665 995407
rect 256866 995404 256926 995818
rect 247599 995402 256926 995404
rect 247599 995346 247604 995402
rect 247660 995346 256926 995402
rect 247599 995344 256926 995346
rect 247599 995341 247665 995344
rect 198639 995254 206622 995256
rect 198639 995198 198644 995254
rect 198700 995198 206622 995254
rect 198639 995196 206622 995198
rect 208143 995254 208254 995259
rect 208143 995198 208148 995254
rect 208204 995198 208254 995254
rect 208143 995196 208254 995198
rect 208719 995254 208830 995259
rect 208719 995198 208724 995254
rect 208780 995198 208830 995254
rect 208719 995196 208830 995198
rect 209775 995254 209886 995259
rect 209775 995198 209780 995254
rect 209836 995198 209886 995254
rect 209775 995196 209886 995198
rect 250479 995256 250545 995259
rect 257442 995256 257502 995818
rect 259407 995790 259412 995846
rect 259468 995790 259680 995846
rect 259407 995788 259680 995790
rect 261216 995788 261438 995848
rect 259407 995785 259473 995788
rect 261378 995700 261438 995788
rect 250479 995254 257502 995256
rect 250479 995198 250484 995254
rect 250540 995198 257502 995254
rect 250479 995196 257502 995198
rect 261186 995640 261438 995700
rect 149679 995193 149745 995196
rect 157263 995193 157329 995196
rect 161679 995193 161745 995196
rect 198639 995193 198705 995196
rect 208143 995193 208209 995196
rect 208719 995193 208785 995196
rect 209775 995193 209841 995196
rect 250479 995193 250545 995196
rect 109359 995106 110910 995108
rect 109359 995050 109364 995106
rect 109420 995050 110910 995106
rect 109359 995048 110910 995050
rect 109359 995045 109425 995048
rect 97839 994958 103806 994960
rect 97839 994902 97844 994958
rect 97900 994902 103806 994958
rect 97839 994900 103806 994902
rect 97839 994897 97905 994900
rect 133647 994516 133713 994519
rect 146799 994516 146865 994519
rect 133647 994514 146865 994516
rect 133647 994458 133652 994514
rect 133708 994458 146804 994514
rect 146860 994458 146865 994514
rect 133647 994456 146865 994458
rect 133647 994453 133713 994456
rect 146799 994453 146865 994456
rect 132783 994368 132849 994371
rect 144687 994368 144753 994371
rect 132783 994366 144753 994368
rect 132783 994310 132788 994366
rect 132844 994310 144692 994366
rect 144748 994310 144753 994366
rect 132783 994308 144753 994310
rect 132783 994305 132849 994308
rect 144687 994305 144753 994308
rect 146895 994368 146961 994371
rect 185775 994368 185841 994371
rect 187311 994368 187377 994371
rect 207375 994368 207441 994371
rect 146895 994366 185982 994368
rect 146895 994310 146900 994366
rect 146956 994310 185780 994366
rect 185836 994310 185982 994366
rect 146895 994308 185982 994310
rect 146895 994305 146961 994308
rect 185775 994305 185841 994308
rect 131823 994220 131889 994223
rect 154767 994220 154833 994223
rect 131823 994218 154833 994220
rect 131823 994162 131828 994218
rect 131884 994162 154772 994218
rect 154828 994162 154833 994218
rect 131823 994160 154833 994162
rect 185922 994220 185982 994308
rect 187311 994366 207441 994368
rect 187311 994310 187316 994366
rect 187372 994310 207380 994366
rect 207436 994310 207441 994366
rect 187311 994308 207441 994310
rect 187311 994305 187377 994308
rect 207375 994305 207441 994308
rect 232527 994368 232593 994371
rect 261186 994368 261246 995640
rect 263970 995552 264030 995818
rect 264480 995788 264702 995848
rect 265056 995846 270801 995848
rect 265056 995790 270740 995846
rect 270796 995790 270801 995846
rect 265056 995788 270801 995790
rect 264642 995700 264702 995788
rect 270735 995785 270801 995788
rect 290511 995848 290577 995851
rect 298383 995848 298449 995851
rect 290511 995846 298449 995848
rect 290511 995790 290516 995846
rect 290572 995790 298388 995846
rect 298444 995790 298449 995846
rect 306063 995848 306129 995851
rect 306543 995848 306609 995851
rect 358095 995848 358161 995851
rect 366159 995848 366225 995851
rect 366735 995848 366801 995851
rect 371535 995848 371601 995851
rect 306063 995846 306336 995848
rect 290511 995788 298449 995790
rect 290511 995785 290577 995788
rect 298383 995785 298449 995788
rect 267951 995700 268017 995703
rect 264642 995698 268017 995700
rect 264642 995642 267956 995698
rect 268012 995642 268017 995698
rect 264642 995640 268017 995642
rect 267951 995637 268017 995640
rect 292527 995700 292593 995703
rect 305730 995700 305790 995818
rect 306063 995790 306068 995846
rect 306124 995790 306336 995846
rect 306063 995788 306336 995790
rect 306543 995846 306912 995848
rect 306543 995790 306548 995846
rect 306604 995790 306912 995846
rect 306543 995788 306912 995790
rect 306063 995785 306129 995788
rect 306543 995785 306609 995788
rect 292527 995698 305790 995700
rect 292527 995642 292532 995698
rect 292588 995642 305790 995698
rect 292527 995640 305790 995642
rect 306447 995700 306513 995703
rect 307362 995700 307422 995818
rect 306447 995698 307422 995700
rect 306447 995642 306452 995698
rect 306508 995642 307422 995698
rect 306447 995640 307422 995642
rect 292527 995637 292593 995640
rect 306447 995637 306513 995640
rect 267855 995552 267921 995555
rect 263970 995550 267921 995552
rect 263970 995494 267860 995550
rect 267916 995494 267921 995550
rect 263970 995492 267921 995494
rect 267855 995489 267921 995492
rect 293583 995552 293649 995555
rect 307938 995552 307998 995818
rect 293583 995550 307998 995552
rect 293583 995494 293588 995550
rect 293644 995494 307998 995550
rect 293583 995492 307998 995494
rect 293583 995489 293649 995492
rect 288015 994664 288081 994667
rect 288975 994664 289041 994667
rect 308079 994664 308145 994667
rect 288015 994662 308145 994664
rect 288015 994606 288020 994662
rect 288076 994606 288980 994662
rect 289036 994606 308084 994662
rect 308140 994606 308145 994662
rect 288015 994604 308145 994606
rect 288015 994601 288081 994604
rect 288975 994601 289041 994604
rect 308079 994601 308145 994604
rect 285999 994516 286065 994519
rect 311202 994516 311262 995818
rect 312834 995407 312894 995818
rect 315522 995700 315582 995818
rect 353952 995788 354366 995848
rect 319695 995700 319761 995703
rect 315522 995698 319761 995700
rect 315522 995642 319700 995698
rect 319756 995642 319761 995698
rect 315522 995640 319761 995642
rect 354306 995700 354366 995788
rect 355074 995700 355134 995818
rect 357216 995788 357630 995848
rect 357792 995846 358161 995848
rect 357792 995790 358100 995846
rect 358156 995790 358161 995846
rect 357792 995788 358161 995790
rect 354306 995640 355134 995700
rect 357570 995700 357630 995788
rect 358095 995785 358161 995788
rect 358191 995700 358257 995703
rect 357570 995698 358257 995700
rect 357570 995642 358196 995698
rect 358252 995642 358257 995698
rect 357570 995640 358257 995642
rect 319695 995637 319761 995640
rect 358191 995637 358257 995640
rect 312783 995402 312894 995407
rect 312783 995346 312788 995402
rect 312844 995346 312894 995402
rect 312783 995344 312894 995346
rect 312783 995341 312849 995344
rect 358338 994664 358398 995818
rect 359394 994960 359454 995818
rect 360480 995788 360702 995848
rect 365952 995846 366225 995848
rect 360642 995552 360702 995788
rect 364866 995700 364926 995818
rect 365952 995790 366164 995846
rect 366220 995790 366225 995846
rect 365952 995788 366225 995790
rect 366528 995846 366801 995848
rect 366528 995790 366740 995846
rect 366796 995790 366801 995846
rect 366528 995788 366801 995790
rect 367008 995846 371601 995848
rect 367008 995790 371540 995846
rect 371596 995790 371601 995846
rect 367008 995788 371601 995790
rect 366159 995785 366225 995788
rect 366735 995785 366801 995788
rect 371535 995785 371601 995788
rect 383055 995848 383121 995851
rect 393711 995848 393777 995851
rect 422127 995848 422193 995851
rect 472239 995848 472305 995851
rect 476463 995848 476529 995851
rect 383055 995846 393777 995848
rect 383055 995790 383060 995846
rect 383116 995790 393716 995846
rect 393772 995790 393777 995846
rect 383055 995788 393777 995790
rect 421920 995846 422334 995848
rect 421920 995790 422132 995846
rect 422188 995790 422334 995846
rect 421920 995788 422334 995790
rect 383055 995785 383121 995788
rect 393711 995785 393777 995788
rect 422127 995785 422193 995788
rect 368655 995700 368721 995703
rect 364866 995698 368721 995700
rect 364866 995642 368660 995698
rect 368716 995642 368721 995698
rect 364866 995640 368721 995642
rect 368655 995637 368721 995640
rect 377199 995700 377265 995703
rect 387471 995700 387537 995703
rect 377199 995698 387537 995700
rect 377199 995642 377204 995698
rect 377260 995642 387476 995698
rect 387532 995642 387537 995698
rect 377199 995640 387537 995642
rect 422274 995700 422334 995788
rect 423042 995700 423102 995818
rect 422274 995640 423102 995700
rect 433218 995788 433440 995848
rect 433218 995700 433278 995788
rect 433890 995700 433950 995818
rect 439170 995788 459198 995848
rect 437775 995700 437841 995703
rect 433218 995640 433470 995700
rect 433890 995698 437841 995700
rect 433890 995642 437780 995698
rect 437836 995642 437841 995698
rect 433890 995640 437841 995642
rect 377199 995637 377265 995640
rect 387471 995637 387537 995640
rect 365775 995552 365841 995555
rect 360642 995550 365841 995552
rect 360642 995494 365780 995550
rect 365836 995494 365841 995550
rect 360642 995492 365841 995494
rect 433410 995552 433470 995640
rect 437775 995637 437841 995640
rect 437967 995552 438033 995555
rect 433410 995550 438033 995552
rect 433410 995494 437972 995550
rect 438028 995494 438033 995550
rect 433410 995492 438033 995494
rect 365775 995489 365841 995492
rect 437967 995489 438033 995492
rect 391119 995404 391185 995407
rect 439170 995404 439230 995788
rect 391119 995402 439230 995404
rect 391119 995346 391124 995402
rect 391180 995346 439230 995402
rect 391119 995344 439230 995346
rect 391119 995341 391185 995344
rect 459138 995256 459198 995788
rect 472239 995846 476529 995848
rect 472239 995790 472244 995846
rect 472300 995790 476468 995846
rect 476524 995790 476529 995846
rect 472239 995788 476529 995790
rect 472239 995785 472305 995788
rect 476463 995785 476529 995788
rect 476602 995786 476608 995850
rect 476672 995848 476678 995850
rect 481455 995848 481521 995851
rect 476672 995846 481521 995848
rect 476672 995790 481460 995846
rect 481516 995790 481521 995846
rect 476672 995788 481521 995790
rect 481602 995848 481662 995936
rect 510543 995933 510609 995936
rect 515535 995933 515601 995936
rect 561903 995933 561969 995936
rect 482031 995848 482097 995851
rect 511119 995848 511185 995851
rect 481602 995846 482097 995848
rect 481602 995790 482036 995846
rect 482092 995790 482097 995846
rect 510912 995846 511185 995848
rect 481602 995788 482097 995790
rect 476672 995786 476678 995788
rect 481455 995785 481521 995788
rect 482031 995785 482097 995788
rect 463791 995700 463857 995703
rect 477711 995700 477777 995703
rect 482703 995700 482769 995703
rect 463791 995698 477777 995700
rect 463791 995642 463796 995698
rect 463852 995642 477716 995698
rect 477772 995642 477777 995698
rect 463791 995640 477777 995642
rect 463791 995637 463857 995640
rect 477711 995637 477777 995640
rect 477954 995698 482769 995700
rect 477954 995642 482708 995698
rect 482764 995642 482769 995698
rect 477954 995640 482769 995642
rect 498402 995700 498462 995818
rect 499458 995700 499518 995818
rect 498402 995640 499518 995700
rect 465327 995552 465393 995555
rect 477954 995552 478014 995640
rect 482703 995637 482769 995640
rect 465327 995550 478014 995552
rect 465327 995494 465332 995550
rect 465388 995494 478014 995550
rect 465327 995492 478014 995494
rect 504930 995552 504990 995818
rect 509250 995700 509310 995818
rect 510912 995790 511124 995846
rect 511180 995790 511185 995846
rect 510912 995788 511185 995790
rect 511119 995785 511185 995788
rect 521199 995848 521265 995851
rect 532239 995848 532305 995851
rect 521199 995846 532305 995848
rect 521199 995790 521204 995846
rect 521260 995790 532244 995846
rect 532300 995790 532305 995846
rect 550479 995848 550545 995851
rect 559791 995848 559857 995851
rect 569871 995848 569937 995851
rect 550479 995846 550944 995848
rect 521199 995788 532305 995790
rect 521199 995785 521265 995788
rect 532239 995785 532305 995788
rect 518415 995700 518481 995703
rect 509250 995698 518481 995700
rect 509250 995642 518420 995698
rect 518476 995642 518481 995698
rect 509250 995640 518481 995642
rect 518415 995637 518481 995640
rect 523503 995700 523569 995703
rect 529071 995700 529137 995703
rect 523503 995698 529137 995700
rect 523503 995642 523508 995698
rect 523564 995642 529076 995698
rect 529132 995642 529137 995698
rect 523503 995640 529137 995642
rect 523503 995637 523569 995640
rect 529071 995637 529137 995640
rect 521295 995552 521361 995555
rect 504930 995550 521361 995552
rect 504930 995494 521300 995550
rect 521356 995494 521361 995550
rect 504930 995492 521361 995494
rect 549762 995552 549822 995818
rect 550338 995700 550398 995818
rect 550479 995790 550484 995846
rect 550540 995790 550944 995846
rect 559584 995846 559857 995848
rect 550479 995788 550944 995790
rect 550479 995785 550545 995788
rect 551394 995700 551454 995818
rect 555375 995700 555441 995703
rect 550338 995698 555441 995700
rect 550338 995642 555380 995698
rect 555436 995642 555441 995698
rect 550338 995640 555441 995642
rect 555375 995637 555441 995640
rect 550479 995552 550545 995555
rect 549762 995550 550545 995552
rect 549762 995494 550484 995550
rect 550540 995494 550545 995550
rect 549762 995492 550545 995494
rect 465327 995489 465393 995492
rect 521295 995489 521361 995492
rect 550479 995489 550545 995492
rect 556290 995404 556350 995818
rect 559584 995790 559796 995846
rect 559852 995790 559857 995846
rect 559584 995788 559857 995790
rect 559791 995785 559857 995788
rect 560130 995703 560190 995818
rect 560514 995788 560736 995848
rect 562272 995788 562686 995848
rect 562848 995846 569937 995848
rect 562848 995790 569876 995846
rect 569932 995790 569937 995846
rect 562848 995788 569937 995790
rect 560130 995698 560241 995703
rect 560130 995642 560180 995698
rect 560236 995642 560241 995698
rect 560130 995640 560241 995642
rect 560514 995700 560574 995788
rect 562626 995700 562686 995788
rect 569871 995785 569937 995788
rect 569679 995700 569745 995703
rect 560514 995640 560766 995700
rect 562626 995698 569745 995700
rect 562626 995642 569684 995698
rect 569740 995642 569745 995698
rect 562626 995640 569745 995642
rect 560175 995637 560241 995640
rect 560706 995552 560766 995640
rect 569679 995637 569745 995640
rect 573807 995700 573873 995703
rect 633999 995700 634065 995703
rect 573807 995698 634065 995700
rect 573807 995642 573812 995698
rect 573868 995642 634004 995698
rect 634060 995642 634065 995698
rect 573807 995640 634065 995642
rect 573807 995637 573873 995640
rect 633999 995637 634065 995640
rect 565839 995552 565905 995555
rect 560706 995550 565905 995552
rect 560706 995494 565844 995550
rect 565900 995494 565905 995550
rect 560706 995492 565905 995494
rect 565839 995489 565905 995492
rect 573039 995552 573105 995555
rect 630927 995552 630993 995555
rect 573039 995550 630993 995552
rect 573039 995494 573044 995550
rect 573100 995494 630932 995550
rect 630988 995494 630993 995550
rect 573039 995492 630993 995494
rect 573039 995489 573105 995492
rect 630927 995489 630993 995492
rect 561615 995404 561681 995407
rect 556290 995402 561681 995404
rect 556290 995346 561620 995402
rect 561676 995346 561681 995402
rect 556290 995344 561681 995346
rect 561615 995341 561681 995344
rect 575151 995404 575217 995407
rect 634575 995404 634641 995407
rect 575151 995402 634641 995404
rect 575151 995346 575156 995402
rect 575212 995346 634580 995402
rect 634636 995346 634641 995402
rect 575151 995344 634641 995346
rect 575151 995341 575217 995344
rect 634575 995341 634641 995344
rect 478095 995256 478161 995259
rect 459138 995254 478161 995256
rect 459138 995198 478100 995254
rect 478156 995198 478161 995254
rect 459138 995196 478161 995198
rect 478095 995193 478161 995196
rect 573231 995256 573297 995259
rect 636111 995256 636177 995259
rect 573231 995254 636177 995256
rect 573231 995198 573236 995254
rect 573292 995198 636116 995254
rect 636172 995198 636177 995254
rect 573231 995196 636177 995198
rect 573231 995193 573297 995196
rect 636111 995193 636177 995196
rect 377103 995108 377169 995111
rect 396975 995108 397041 995111
rect 377103 995106 397041 995108
rect 377103 995050 377108 995106
rect 377164 995050 396980 995106
rect 397036 995050 397041 995106
rect 377103 995048 397041 995050
rect 377103 995045 377169 995048
rect 396975 995045 397041 995048
rect 472143 995108 472209 995111
rect 481071 995108 481137 995111
rect 472143 995106 481137 995108
rect 472143 995050 472148 995106
rect 472204 995050 481076 995106
rect 481132 995050 481137 995106
rect 472143 995048 481137 995050
rect 472143 995045 472209 995048
rect 481071 995045 481137 995048
rect 573519 995108 573585 995111
rect 639183 995108 639249 995111
rect 573519 995106 639249 995108
rect 573519 995050 573524 995106
rect 573580 995050 639188 995106
rect 639244 995050 639249 995106
rect 573519 995048 639249 995050
rect 573519 995045 573585 995048
rect 639183 995045 639249 995048
rect 388335 994960 388401 994963
rect 359394 994958 388401 994960
rect 359394 994902 388340 994958
rect 388396 994902 388401 994958
rect 359394 994900 388401 994902
rect 388335 994897 388401 994900
rect 467055 994960 467121 994963
rect 484143 994960 484209 994963
rect 467055 994958 484209 994960
rect 467055 994902 467060 994958
rect 467116 994902 484148 994958
rect 484204 994902 484209 994958
rect 467055 994900 484209 994902
rect 467055 994897 467121 994900
rect 484143 994897 484209 994900
rect 572943 994960 573009 994963
rect 635247 994960 635313 994963
rect 572943 994958 635313 994960
rect 572943 994902 572948 994958
rect 573004 994902 635252 994958
rect 635308 994902 635313 994958
rect 572943 994900 635313 994902
rect 572943 994897 573009 994900
rect 635247 994897 635313 994900
rect 358479 994812 358545 994815
rect 389391 994812 389457 994815
rect 358479 994810 389457 994812
rect 358479 994754 358484 994810
rect 358540 994754 389396 994810
rect 389452 994754 389457 994810
rect 358479 994752 389457 994754
rect 358479 994749 358545 994752
rect 389391 994749 389457 994752
rect 464751 994812 464817 994815
rect 485967 994812 486033 994815
rect 464751 994810 486033 994812
rect 464751 994754 464756 994810
rect 464812 994754 485972 994810
rect 486028 994754 486033 994810
rect 464751 994752 486033 994754
rect 464751 994749 464817 994752
rect 485967 994749 486033 994752
rect 572847 994812 572913 994815
rect 637359 994812 637425 994815
rect 572847 994810 637425 994812
rect 572847 994754 572852 994810
rect 572908 994754 637364 994810
rect 637420 994754 637425 994810
rect 572847 994752 637425 994754
rect 572847 994749 572913 994752
rect 637359 994749 637425 994752
rect 395151 994664 395217 994667
rect 358338 994662 395217 994664
rect 358338 994606 395156 994662
rect 395212 994606 395217 994662
rect 358338 994604 395217 994606
rect 395151 994601 395217 994604
rect 478095 994664 478161 994667
rect 479823 994664 479889 994667
rect 524079 994664 524145 994667
rect 478095 994662 524145 994664
rect 478095 994606 478100 994662
rect 478156 994606 479828 994662
rect 479884 994606 524084 994662
rect 524140 994606 524145 994662
rect 478095 994604 524145 994606
rect 478095 994601 478161 994604
rect 479823 994601 479889 994604
rect 524079 994601 524145 994604
rect 536751 994664 536817 994667
rect 634287 994664 634353 994667
rect 536751 994662 634353 994664
rect 536751 994606 536756 994662
rect 536812 994606 634292 994662
rect 634348 994606 634353 994662
rect 536751 994604 634353 994606
rect 536751 994601 536817 994604
rect 634287 994601 634353 994604
rect 285999 994514 311262 994516
rect 285999 994458 286004 994514
rect 286060 994458 311262 994514
rect 285999 994456 311262 994458
rect 358095 994516 358161 994519
rect 393039 994516 393105 994519
rect 358095 994514 393105 994516
rect 358095 994458 358100 994514
rect 358156 994458 393044 994514
rect 393100 994458 393105 994514
rect 358095 994456 393105 994458
rect 285999 994453 286065 994456
rect 358095 994453 358161 994456
rect 393039 994453 393105 994456
rect 485583 994516 485649 994519
rect 650031 994516 650097 994519
rect 485583 994514 650097 994516
rect 485583 994458 485588 994514
rect 485644 994458 650036 994514
rect 650092 994458 650097 994514
rect 485583 994456 650097 994458
rect 485583 994453 485649 994456
rect 650031 994453 650097 994456
rect 232527 994366 261246 994368
rect 232527 994310 232532 994366
rect 232588 994310 261246 994366
rect 232527 994308 261246 994310
rect 308079 994368 308145 994371
rect 390831 994368 390897 994371
rect 308079 994366 390897 994368
rect 308079 994310 308084 994366
rect 308140 994310 390836 994366
rect 390892 994310 390897 994366
rect 308079 994308 390897 994310
rect 232527 994305 232593 994308
rect 308079 994305 308145 994308
rect 390831 994305 390897 994308
rect 396303 994368 396369 994371
rect 604623 994368 604689 994371
rect 396303 994366 604689 994368
rect 396303 994310 396308 994366
rect 396364 994310 604628 994366
rect 604684 994310 604689 994366
rect 396303 994308 604689 994310
rect 396303 994305 396369 994308
rect 604623 994305 604689 994308
rect 237519 994220 237585 994223
rect 288015 994220 288081 994223
rect 185922 994218 288081 994220
rect 185922 994162 237524 994218
rect 237580 994162 288020 994218
rect 288076 994162 288081 994218
rect 185922 994160 288081 994162
rect 131823 994157 131889 994160
rect 154767 994157 154833 994160
rect 237519 994157 237585 994160
rect 288015 994157 288081 994160
rect 294543 994220 294609 994223
rect 649743 994220 649809 994223
rect 294543 994218 649809 994220
rect 294543 994162 294548 994218
rect 294604 994162 649748 994218
rect 649804 994162 649809 994218
rect 294543 994160 649809 994162
rect 294543 994157 294609 994160
rect 649743 994157 649809 994160
rect 135183 994072 135249 994075
rect 146895 994072 146961 994075
rect 135183 994070 146961 994072
rect 135183 994014 135188 994070
rect 135244 994014 146900 994070
rect 146956 994014 146961 994070
rect 135183 994012 146961 994014
rect 135183 994009 135249 994012
rect 146895 994009 146961 994012
rect 191535 994072 191601 994075
rect 649647 994072 649713 994075
rect 191535 994070 649713 994072
rect 191535 994014 191540 994070
rect 191596 994014 649652 994070
rect 649708 994014 649713 994070
rect 191535 994012 649713 994014
rect 191535 994009 191601 994012
rect 649647 994009 649713 994012
rect 88719 993924 88785 993927
rect 576303 993924 576369 993927
rect 88719 993922 576369 993924
rect 88719 993866 88724 993922
rect 88780 993866 576308 993922
rect 576364 993866 576369 993922
rect 88719 993864 576369 993866
rect 88719 993861 88785 993864
rect 576303 993861 576369 993864
rect 638511 993924 638577 993927
rect 642255 993924 642321 993927
rect 638511 993922 642321 993924
rect 638511 993866 638516 993922
rect 638572 993866 642260 993922
rect 642316 993866 642321 993922
rect 638511 993864 642321 993866
rect 638511 993861 638577 993864
rect 642255 993861 642321 993864
rect 84495 993776 84561 993779
rect 104463 993776 104529 993779
rect 84495 993774 104529 993776
rect 84495 993718 84500 993774
rect 84556 993718 104468 993774
rect 104524 993718 104529 993774
rect 84495 993716 104529 993718
rect 84495 993713 84561 993716
rect 104463 993713 104529 993716
rect 140367 993776 140433 993779
rect 641103 993776 641169 993779
rect 140367 993774 641169 993776
rect 140367 993718 140372 993774
rect 140428 993718 641108 993774
rect 641164 993718 641169 993774
rect 140367 993716 641169 993718
rect 140367 993713 140433 993716
rect 641103 993713 641169 993716
rect 423375 993628 423441 993631
rect 443439 993628 443505 993631
rect 423375 993626 443505 993628
rect 423375 993570 423380 993626
rect 423436 993570 443444 993626
rect 443500 993570 443505 993626
rect 423375 993568 443505 993570
rect 423375 993565 423441 993568
rect 443439 993565 443505 993568
rect 362895 993332 362961 993335
rect 382959 993332 383025 993335
rect 362895 993330 383025 993332
rect 362895 993274 362900 993330
rect 362956 993274 382964 993330
rect 383020 993274 383025 993330
rect 362895 993272 383025 993274
rect 362895 993269 362961 993272
rect 382959 993269 383025 993272
rect 30656 988352 31778 988394
rect 30656 984370 30806 988352
rect 31614 988174 31778 988352
rect 31614 988042 42224 988174
rect 31614 984584 41196 988042
rect 42102 984584 42224 988042
rect 31614 984474 42224 984584
rect 31614 984370 31778 984474
rect 30656 984336 31778 984370
rect 655119 976756 655185 976759
rect 650208 976754 655185 976756
rect 650208 976698 655124 976754
rect 655180 976698 655185 976754
rect 650208 976696 655185 976698
rect 655119 976693 655185 976696
rect 59439 975424 59505 975427
rect 59439 975422 64416 975424
rect 59439 975366 59444 975422
rect 59500 975366 64416 975422
rect 59439 975364 64416 975366
rect 59439 975361 59505 975364
rect 42063 968766 42129 968767
rect 42063 968762 42112 968766
rect 42176 968764 42182 968766
rect 42063 968706 42068 968762
rect 42063 968702 42112 968706
rect 42176 968704 42220 968764
rect 42176 968702 42182 968704
rect 42063 968701 42129 968702
rect 674319 967580 674385 967583
rect 674991 967580 675057 967583
rect 674319 967578 675057 967580
rect 674319 967522 674324 967578
rect 674380 967522 674996 967578
rect 675052 967522 675057 967578
rect 674319 967520 675057 967522
rect 674319 967517 674385 967520
rect 674991 967517 675057 967520
rect 674511 967432 674577 967435
rect 675706 967432 675712 967434
rect 674511 967430 675712 967432
rect 674511 967374 674516 967430
rect 674572 967374 675712 967430
rect 674511 967372 675712 967374
rect 674511 967369 674577 967372
rect 675706 967370 675712 967372
rect 675776 967370 675782 967434
rect 41338 967074 41344 967138
rect 41408 967136 41414 967138
rect 41775 967136 41841 967139
rect 41408 967134 41841 967136
rect 41408 967078 41780 967134
rect 41836 967078 41841 967134
rect 41408 967076 41841 967078
rect 41408 967074 41414 967076
rect 41775 967073 41841 967076
rect 675759 965656 675825 965659
rect 676090 965656 676096 965658
rect 675759 965654 676096 965656
rect 675759 965598 675764 965654
rect 675820 965598 676096 965654
rect 675759 965596 676096 965598
rect 675759 965593 675825 965596
rect 676090 965594 676096 965596
rect 676160 965594 676166 965658
rect 42063 965064 42129 965067
rect 42298 965064 42304 965066
rect 42063 965062 42304 965064
rect 42063 965006 42068 965062
rect 42124 965006 42304 965062
rect 42063 965004 42304 965006
rect 42063 965001 42129 965004
rect 42298 965002 42304 965004
rect 42368 965002 42374 965066
rect 655215 965064 655281 965067
rect 650208 965062 655281 965064
rect 650208 965006 655220 965062
rect 655276 965006 655281 965062
rect 650208 965004 655281 965006
rect 655215 965001 655281 965004
rect 674362 965002 674368 965066
rect 674432 965064 674438 965066
rect 675279 965064 675345 965067
rect 674432 965062 675345 965064
rect 674432 965006 675284 965062
rect 675340 965006 675345 965062
rect 674432 965004 675345 965006
rect 674432 965002 674438 965004
rect 675279 965001 675345 965004
rect 675183 964918 675249 964919
rect 675130 964916 675136 964918
rect 675092 964856 675136 964916
rect 675200 964914 675249 964918
rect 675244 964858 675249 964914
rect 675130 964854 675136 964856
rect 675200 964854 675249 964858
rect 675183 964853 675249 964854
rect 40954 963966 40960 964030
rect 41024 964028 41030 964030
rect 41775 964028 41841 964031
rect 41024 964026 41841 964028
rect 41024 963970 41780 964026
rect 41836 963970 41841 964026
rect 41024 963968 41841 963970
rect 41024 963966 41030 963968
rect 41775 963965 41841 963968
rect 41146 963226 41152 963290
rect 41216 963288 41222 963290
rect 41775 963288 41841 963291
rect 41216 963286 41841 963288
rect 41216 963230 41780 963286
rect 41836 963230 41841 963286
rect 41216 963228 41841 963230
rect 41216 963226 41222 963228
rect 41775 963225 41841 963228
rect 42831 963288 42897 963291
rect 62031 963288 62097 963291
rect 42831 963286 62097 963288
rect 42831 963230 42836 963286
rect 42892 963230 62036 963286
rect 62092 963230 62097 963286
rect 42831 963228 62097 963230
rect 42831 963225 42897 963228
rect 62031 963225 62097 963228
rect 674938 962782 674944 962846
rect 675008 962844 675014 962846
rect 675087 962844 675153 962847
rect 675008 962842 675153 962844
rect 675008 962786 675092 962842
rect 675148 962786 675153 962842
rect 675008 962784 675153 962786
rect 675008 962782 675014 962784
rect 675087 962781 675153 962784
rect 40762 962634 40768 962698
rect 40832 962696 40838 962698
rect 41775 962696 41841 962699
rect 40832 962694 41841 962696
rect 40832 962638 41780 962694
rect 41836 962638 41841 962694
rect 40832 962636 41841 962638
rect 40832 962634 40838 962636
rect 41775 962633 41841 962636
rect 674554 962486 674560 962550
rect 674624 962548 674630 962550
rect 675183 962548 675249 962551
rect 674624 962546 675249 962548
rect 674624 962490 675188 962546
rect 675244 962490 675249 962546
rect 674624 962488 675249 962490
rect 674624 962486 674630 962488
rect 675183 962485 675249 962488
rect 675759 962252 675825 962255
rect 676282 962252 676288 962254
rect 675759 962250 676288 962252
rect 675759 962194 675764 962250
rect 675820 962194 676288 962250
rect 675759 962192 676288 962194
rect 675759 962189 675825 962192
rect 676282 962190 676288 962192
rect 676352 962190 676358 962254
rect 40378 962042 40384 962106
rect 40448 962104 40454 962106
rect 41871 962104 41937 962107
rect 40448 962102 41937 962104
rect 40448 962046 41876 962102
rect 41932 962046 41937 962102
rect 40448 962044 41937 962046
rect 40448 962042 40454 962044
rect 41871 962041 41937 962044
rect 42682 961894 42688 961958
rect 42752 961956 42758 961958
rect 61839 961956 61905 961959
rect 42752 961954 61905 961956
rect 42752 961898 61844 961954
rect 61900 961898 61905 961954
rect 42752 961896 61905 961898
rect 42752 961894 42758 961896
rect 61839 961893 61905 961896
rect 674746 961450 674752 961514
rect 674816 961512 674822 961514
rect 675375 961512 675441 961515
rect 674816 961510 675441 961512
rect 674816 961454 675380 961510
rect 675436 961454 675441 961510
rect 674816 961452 675441 961454
rect 674816 961450 674822 961452
rect 675375 961449 675441 961452
rect 675663 961070 675729 961071
rect 675663 961068 675712 961070
rect 675620 961066 675712 961068
rect 675620 961010 675668 961066
rect 675620 961008 675712 961010
rect 675663 961006 675712 961008
rect 675776 961006 675782 961070
rect 675663 961005 675729 961006
rect 59535 960920 59601 960923
rect 59535 960918 64416 960920
rect 59535 960862 59540 960918
rect 59596 960862 64416 960918
rect 59535 960860 64416 960862
rect 59535 960857 59601 960860
rect 42159 960476 42225 960479
rect 42682 960476 42688 960478
rect 42159 960474 42688 960476
rect 42159 960418 42164 960474
rect 42220 960418 42688 960474
rect 42159 960416 42688 960418
rect 42159 960413 42225 960416
rect 42682 960414 42688 960416
rect 42752 960414 42758 960478
rect 675759 960180 675825 960183
rect 675898 960180 675904 960182
rect 675759 960178 675904 960180
rect 675759 960122 675764 960178
rect 675820 960122 675904 960178
rect 675759 960120 675904 960122
rect 675759 960117 675825 960120
rect 675898 960118 675904 960120
rect 675968 960118 675974 960182
rect 41530 959674 41536 959738
rect 41600 959736 41606 959738
rect 41775 959736 41841 959739
rect 41600 959734 41841 959736
rect 41600 959678 41780 959734
rect 41836 959678 41841 959734
rect 41600 959676 41841 959678
rect 41600 959674 41606 959676
rect 41775 959673 41841 959676
rect 41775 959146 41841 959147
rect 41722 959144 41728 959146
rect 41684 959084 41728 959144
rect 41792 959142 41841 959146
rect 41836 959086 41841 959142
rect 41722 959082 41728 959084
rect 41792 959082 41841 959086
rect 675322 959082 675328 959146
rect 675392 959144 675398 959146
rect 675471 959144 675537 959147
rect 675392 959142 675537 959144
rect 675392 959086 675476 959142
rect 675532 959086 675537 959142
rect 675392 959084 675537 959086
rect 675392 959082 675398 959084
rect 41775 959081 41841 959082
rect 675471 959081 675537 959084
rect 40570 958490 40576 958554
rect 40640 958552 40646 958554
rect 41775 958552 41841 958555
rect 40640 958550 41841 958552
rect 40640 958494 41780 958550
rect 41836 958494 41841 958550
rect 40640 958492 41841 958494
rect 40640 958490 40646 958492
rect 41775 958489 41841 958492
rect 41871 957814 41937 957815
rect 41871 957810 41920 957814
rect 41984 957812 41990 957814
rect 41871 957754 41876 957810
rect 41871 957750 41920 957754
rect 41984 957752 42028 957812
rect 41984 957750 41990 957752
rect 41871 957749 41937 957750
rect 675471 957666 675537 957667
rect 675471 957662 675520 957666
rect 675584 957664 675590 957666
rect 675471 957606 675476 957662
rect 675471 957602 675520 957606
rect 675584 957604 675628 957664
rect 675584 957602 675590 957604
rect 675471 957601 675537 957602
rect 673978 955974 673984 956038
rect 674048 956036 674054 956038
rect 675471 956036 675537 956039
rect 674048 956034 675537 956036
rect 674048 955978 675476 956034
rect 675532 955978 675537 956034
rect 674048 955976 675537 955978
rect 674048 955974 674054 955976
rect 675471 955973 675537 955976
rect 42159 955888 42225 955891
rect 42490 955888 42496 955890
rect 42159 955886 42496 955888
rect 42159 955830 42164 955886
rect 42220 955830 42496 955886
rect 42159 955828 42496 955830
rect 42159 955825 42225 955828
rect 42490 955826 42496 955828
rect 42560 955826 42566 955890
rect 675087 953520 675153 953523
rect 677050 953520 677056 953522
rect 675087 953518 677056 953520
rect 675087 953462 675092 953518
rect 675148 953462 677056 953518
rect 675087 953460 677056 953462
rect 675087 953457 675153 953460
rect 677050 953458 677056 953460
rect 677120 953458 677126 953522
rect 655311 953372 655377 953375
rect 650208 953370 655377 953372
rect 650208 953314 655316 953370
rect 655372 953314 655377 953370
rect 650208 953312 655377 953314
rect 655311 953309 655377 953312
rect 675183 953372 675249 953375
rect 676858 953372 676864 953374
rect 675183 953370 676864 953372
rect 675183 953314 675188 953370
rect 675244 953314 676864 953370
rect 675183 953312 676864 953314
rect 675183 953309 675249 953312
rect 676858 953310 676864 953312
rect 676928 953310 676934 953374
rect 6594 952032 8752 952832
rect 9552 952831 50926 952832
rect 9552 952033 50127 952831
rect 50925 952033 50931 952831
rect 9552 952032 50926 952033
rect 6562 950306 16320 951106
rect 17120 951105 52718 951106
rect 17120 950307 51919 951105
rect 52717 950307 52723 951105
rect 671682 950872 699411 950873
rect 17120 950306 52718 950307
rect 42429 950151 42499 950153
rect 42429 950150 42515 950151
rect 42829 950150 42899 950155
rect 42429 950148 42834 950150
rect 42429 950088 42434 950148
rect 42494 950090 42834 950148
rect 42894 950090 42899 950150
rect 42494 950088 42515 950090
rect 42429 950083 42515 950088
rect 42829 950085 42899 950090
rect 42445 950081 42515 950083
rect 671677 949780 671683 950872
rect 672775 949780 699411 950872
rect 671682 949779 699411 949780
rect 700505 949779 710805 950873
rect 666066 949401 709356 949402
rect 6276 948482 7286 949282
rect 8086 949281 54502 949282
rect 8086 948483 53703 949281
rect 54501 948483 54507 949281
rect 8086 948482 54502 948483
rect 666061 948219 666067 949401
rect 667249 948219 709356 949401
rect 666066 948218 709356 948219
rect 710540 948218 710676 949402
rect 6468 946946 17618 947746
rect 18418 947745 56068 947746
rect 18418 946947 55269 947745
rect 56067 946947 56073 947745
rect 662178 947415 700802 947416
rect 18418 946946 56068 946947
rect 59535 946712 59601 946715
rect 59535 946710 64416 946712
rect 59535 946654 59540 946710
rect 59596 946654 64416 946710
rect 59535 946652 64416 946654
rect 59535 946649 59601 946652
rect 662173 946233 662179 947415
rect 663361 946233 700802 947415
rect 662178 946232 700802 946233
rect 701986 946232 710734 947416
rect 42298 945614 42304 945678
rect 42368 945676 42374 945678
rect 42874 945676 42880 945678
rect 42368 945616 42880 945676
rect 42368 945614 42374 945616
rect 42874 945614 42880 945616
rect 42944 945614 42950 945678
rect 659368 945491 708038 945492
rect 42639 944936 42705 944939
rect 42528 944934 42705 944936
rect 42528 944878 42644 944934
rect 42700 944878 42705 944934
rect 42528 944876 42705 944878
rect 42639 944873 42705 944876
rect 42639 944344 42705 944347
rect 42528 944342 42705 944344
rect 42528 944286 42644 944342
rect 42700 944286 42705 944342
rect 659363 944309 659369 945491
rect 660551 944309 708038 945491
rect 659368 944308 708038 944309
rect 709222 944308 710908 945492
rect 42528 944284 42705 944286
rect 42639 944281 42705 944284
rect 42735 943826 42801 943829
rect 42528 943824 42801 943826
rect 42528 943768 42740 943824
rect 42796 943768 42801 943824
rect 42528 943766 42801 943768
rect 42735 943763 42801 943766
rect 40386 943015 40446 943278
rect 40335 943010 40446 943015
rect 40335 942954 40340 943010
rect 40396 942954 40446 943010
rect 40335 942952 40446 942954
rect 40335 942949 40401 942952
rect 42639 942716 42705 942719
rect 42528 942714 42705 942716
rect 42528 942658 42644 942714
rect 42700 942658 42705 942714
rect 42528 942656 42705 942658
rect 42639 942653 42705 942656
rect 42639 942198 42705 942201
rect 42528 942196 42705 942198
rect 42528 942140 42644 942196
rect 42700 942140 42705 942196
rect 42528 942138 42705 942140
rect 42639 942135 42705 942138
rect 649647 941828 649713 941831
rect 649602 941826 649713 941828
rect 649602 941770 649652 941826
rect 649708 941770 649713 941826
rect 649602 941765 649713 941770
rect 47439 941680 47505 941683
rect 40224 941678 47505 941680
rect 40224 941650 47444 941678
rect 40194 941622 47444 941650
rect 47500 941622 47505 941678
rect 40194 941620 47505 941622
rect 40194 941386 40254 941620
rect 47439 941617 47505 941620
rect 649602 941502 649662 941765
rect 40186 941322 40192 941386
rect 40256 941322 40262 941386
rect 42490 941322 42496 941386
rect 42560 941322 42566 941386
rect 42498 941058 42558 941322
rect 676866 940943 676926 941280
rect 41338 940878 41344 940942
rect 41408 940878 41414 940942
rect 676815 940938 676926 940943
rect 676815 940882 676820 940938
rect 676876 940882 676926 940938
rect 676815 940880 676926 940882
rect 41346 940540 41406 940878
rect 676815 940877 676881 940880
rect 676866 940499 676926 940762
rect 676866 940494 676977 940499
rect 676866 940438 676916 940494
rect 676972 940438 676977 940494
rect 676866 940436 676977 940438
rect 676911 940433 676977 940436
rect 42351 940348 42417 940351
rect 42306 940346 42417 940348
rect 42306 940290 42356 940346
rect 42412 940290 42417 940346
rect 42306 940285 42417 940290
rect 42306 940022 42366 940285
rect 674607 939904 674673 939907
rect 674754 939904 674814 940170
rect 674607 939902 674814 939904
rect 674607 939846 674612 939902
rect 674668 939846 674814 939902
rect 674607 939844 674814 939846
rect 674607 939841 674673 939844
rect 41914 939694 41920 939758
rect 41984 939694 41990 939758
rect 41922 939430 41982 939694
rect 674415 939608 674481 939611
rect 674415 939606 674784 939608
rect 674415 939550 674420 939606
rect 674476 939550 674784 939606
rect 674415 939548 674784 939550
rect 674415 939545 674481 939548
rect 40378 939102 40384 939166
rect 40448 939102 40454 939166
rect 673839 939164 673905 939167
rect 673839 939162 674784 939164
rect 673839 939106 673844 939162
rect 673900 939106 674784 939162
rect 673839 939104 674784 939106
rect 40386 938912 40446 939102
rect 673839 939101 673905 939104
rect 42106 938658 42112 938722
rect 42176 938658 42182 938722
rect 42114 938394 42174 938658
rect 676866 938279 676926 938542
rect 676815 938274 676926 938279
rect 676815 938218 676820 938274
rect 676876 938218 676926 938274
rect 676815 938216 676926 938218
rect 676815 938213 676881 938216
rect 42159 938128 42225 938131
rect 42114 938126 42225 938128
rect 42114 938070 42164 938126
rect 42220 938070 42225 938126
rect 42114 938065 42225 938070
rect 42114 937802 42174 938065
rect 674415 937980 674481 937983
rect 674415 937978 674784 937980
rect 674415 937922 674420 937978
rect 674476 937922 674784 937978
rect 674415 937920 674784 937922
rect 674415 937917 674481 937920
rect 40570 937622 40576 937686
rect 40640 937622 40646 937686
rect 40578 937284 40638 937622
rect 674362 937474 674368 937538
rect 674432 937536 674438 937538
rect 674432 937476 674784 937536
rect 674432 937474 674438 937476
rect 41722 937030 41728 937094
rect 41792 937030 41798 937094
rect 41730 936766 41790 937030
rect 674127 936944 674193 936947
rect 674127 936942 674784 936944
rect 674127 936886 674132 936942
rect 674188 936886 674784 936942
rect 674127 936884 674784 936886
rect 674127 936881 674193 936884
rect 675130 936586 675136 936650
rect 675200 936586 675206 936650
rect 675138 936322 675198 936586
rect 42874 936204 42880 936206
rect 42528 936144 42880 936204
rect 42874 936142 42880 936144
rect 42944 936142 42950 936206
rect 674938 935994 674944 936058
rect 675008 935994 675014 936058
rect 41146 935846 41152 935910
rect 41216 935846 41222 935910
rect 674946 935878 675006 935994
rect 41154 935656 41214 935846
rect 675322 935550 675328 935614
rect 675392 935550 675398 935614
rect 41530 935402 41536 935466
rect 41600 935402 41606 935466
rect 41538 935138 41598 935402
rect 675330 935286 675390 935550
rect 40762 934810 40768 934874
rect 40832 934810 40838 934874
rect 40770 934546 40830 934810
rect 674031 934724 674097 934727
rect 674031 934722 674784 934724
rect 674031 934666 674036 934722
rect 674092 934666 674784 934722
rect 674031 934664 674784 934666
rect 674031 934661 674097 934664
rect 676090 934514 676096 934578
rect 676160 934514 676166 934578
rect 40954 934366 40960 934430
rect 41024 934366 41030 934430
rect 40962 933954 41022 934366
rect 676098 934250 676158 934514
rect 674554 933922 674560 933986
rect 674624 933984 674630 933986
rect 674624 933924 674814 933984
rect 674624 933922 674630 933924
rect 674754 933658 674814 933924
rect 42498 933244 42558 933510
rect 676282 933330 676288 933394
rect 676352 933330 676358 933394
rect 42498 933184 42750 933244
rect 35202 932655 35262 932918
rect 42690 932800 42750 933184
rect 676290 933066 676350 933330
rect 35151 932650 35262 932655
rect 35151 932594 35156 932650
rect 35212 932594 35262 932650
rect 35151 932592 35262 932594
rect 42498 932740 42750 932800
rect 35151 932589 35217 932592
rect 35151 932208 35217 932211
rect 42498 932208 42558 932740
rect 673978 932590 673984 932654
rect 674048 932652 674054 932654
rect 674048 932592 674784 932652
rect 674048 932590 674054 932592
rect 675514 932294 675520 932358
rect 675584 932294 675590 932358
rect 42639 932208 42705 932211
rect 35151 932206 35262 932208
rect 35151 932150 35156 932206
rect 35212 932150 35262 932206
rect 35151 932145 35262 932150
rect 42498 932206 42705 932208
rect 42498 932150 42644 932206
rect 42700 932150 42705 932206
rect 42498 932148 42705 932150
rect 42639 932145 42705 932148
rect 59535 932208 59601 932211
rect 59535 932206 64416 932208
rect 59535 932150 59540 932206
rect 59596 932150 64416 932206
rect 59535 932148 64416 932150
rect 59535 932145 59601 932148
rect 35202 931882 35262 932145
rect 675522 932030 675582 932294
rect 674746 931702 674752 931766
rect 674816 931702 674822 931766
rect 674754 931438 674814 931702
rect 677050 931258 677056 931322
rect 677120 931258 677126 931322
rect 677058 930920 677118 931258
rect 676858 930666 676864 930730
rect 676928 930666 676934 930730
rect 676866 930402 676926 930666
rect 654447 929840 654513 929843
rect 650208 929838 654513 929840
rect 650208 929782 654452 929838
rect 654508 929782 654513 929838
rect 650208 929780 654513 929782
rect 654447 929777 654513 929780
rect 677058 929547 677118 929810
rect 677007 929542 677118 929547
rect 677007 929486 677012 929542
rect 677068 929486 677118 929542
rect 677007 929484 677118 929486
rect 677007 929481 677073 929484
rect 676866 928955 676926 929292
rect 676815 928950 676926 928955
rect 676815 928894 676820 928950
rect 676876 928894 676926 928950
rect 676815 928892 676926 928894
rect 676815 928889 676881 928892
rect 677058 928511 677118 928774
rect 676815 928508 676881 928511
rect 676815 928506 676926 928508
rect 676815 928450 676820 928506
rect 676876 928450 676926 928506
rect 676815 928445 676926 928450
rect 677007 928506 677118 928511
rect 677007 928450 677012 928506
rect 677068 928450 677118 928506
rect 677007 928448 677118 928450
rect 677007 928445 677073 928448
rect 676866 928182 676926 928445
rect 40143 927324 40209 927327
rect 40143 927322 40254 927324
rect 40143 927266 40148 927322
rect 40204 927266 40254 927322
rect 40143 927261 40254 927266
rect 39855 927176 39921 927179
rect 40194 927176 40254 927261
rect 39855 927174 40254 927176
rect 39855 927118 39860 927174
rect 39916 927118 40254 927174
rect 39855 927116 40254 927118
rect 39855 927113 39921 927116
rect 38546 922378 45882 926250
rect 38546 922334 43192 922378
rect 42960 916604 43192 922334
rect 44420 916604 45882 922378
rect 671748 921504 679012 921540
rect 653967 918148 654033 918151
rect 650208 918146 654033 918148
rect 650208 918090 653972 918146
rect 654028 918090 654033 918146
rect 650208 918088 654033 918090
rect 653967 918085 654033 918088
rect 671698 918086 679012 921504
rect 59535 917852 59601 917855
rect 59535 917850 64416 917852
rect 59535 917794 59540 917850
rect 59596 917794 64416 917850
rect 59535 917792 64416 917794
rect 671698 917844 675116 918086
rect 59535 917789 59601 917792
rect 42960 916534 45882 916604
rect 38842 912792 45882 916534
rect 671698 912320 671794 917844
rect 674916 912320 675116 917844
rect 671698 912256 675116 912320
rect 671698 908802 678962 912256
rect 654447 906456 654513 906459
rect 650208 906454 654513 906456
rect 650208 906398 654452 906454
rect 654508 906398 654513 906454
rect 650208 906396 654513 906398
rect 654447 906393 654513 906396
rect 59535 903496 59601 903499
rect 59535 903494 64416 903496
rect 59535 903438 59540 903494
rect 59596 903438 64416 903494
rect 59535 903436 64416 903438
rect 59535 903433 59601 903436
rect 650127 895208 650193 895211
rect 650127 895206 650238 895208
rect 650127 895150 650132 895206
rect 650188 895150 650238 895206
rect 650127 895145 650238 895150
rect 650178 894586 650238 895145
rect 59535 889140 59601 889143
rect 59535 889138 64416 889140
rect 59535 889082 59540 889138
rect 59596 889082 64416 889138
rect 59535 889080 64416 889082
rect 59535 889077 59601 889080
rect 653967 882924 654033 882927
rect 650208 882922 654033 882924
rect 650208 882866 653972 882922
rect 654028 882866 654033 882922
rect 650208 882864 654033 882866
rect 653967 882861 654033 882864
rect 674746 876942 674752 877006
rect 674816 877004 674822 877006
rect 675375 877004 675441 877007
rect 674816 877002 675441 877004
rect 674816 876946 675380 877002
rect 675436 876946 675441 877002
rect 674816 876944 675441 876946
rect 674816 876942 674822 876944
rect 675375 876941 675441 876944
rect 673978 876498 673984 876562
rect 674048 876560 674054 876562
rect 675375 876560 675441 876563
rect 674048 876558 675441 876560
rect 674048 876502 675380 876558
rect 675436 876502 675441 876558
rect 674048 876500 675441 876502
rect 674048 876498 674054 876500
rect 675375 876497 675441 876500
rect 675279 875968 675345 875971
rect 675706 875968 675712 875970
rect 675279 875966 675712 875968
rect 675279 875910 675284 875966
rect 675340 875910 675712 875966
rect 675279 875908 675712 875910
rect 675279 875905 675345 875908
rect 675706 875906 675712 875908
rect 675776 875906 675782 875970
rect 674554 875758 674560 875822
rect 674624 875820 674630 875822
rect 675375 875820 675441 875823
rect 674624 875818 675441 875820
rect 674624 875762 675380 875818
rect 675436 875762 675441 875818
rect 674624 875760 675441 875762
rect 674624 875758 674630 875760
rect 675375 875757 675441 875760
rect 675087 875672 675153 875675
rect 675898 875672 675904 875674
rect 675087 875670 675904 875672
rect 675087 875614 675092 875670
rect 675148 875614 675904 875670
rect 675087 875612 675904 875614
rect 675087 875609 675153 875612
rect 675898 875610 675904 875612
rect 675968 875610 675974 875674
rect 59535 874784 59601 874787
rect 59535 874782 64416 874784
rect 59535 874726 59540 874782
rect 59596 874726 64416 874782
rect 59535 874724 64416 874726
rect 59535 874721 59601 874724
rect 674170 874130 674176 874194
rect 674240 874192 674246 874194
rect 675471 874192 675537 874195
rect 674240 874190 675537 874192
rect 674240 874134 675476 874190
rect 675532 874134 675537 874190
rect 674240 874132 675537 874134
rect 674240 874130 674246 874132
rect 675471 874129 675537 874132
rect 674938 873390 674944 873454
rect 675008 873452 675014 873454
rect 675375 873452 675441 873455
rect 675008 873450 675441 873452
rect 675008 873394 675380 873450
rect 675436 873394 675441 873450
rect 675008 873392 675441 873394
rect 675008 873390 675014 873392
rect 675375 873389 675441 873392
rect 674362 872798 674368 872862
rect 674432 872860 674438 872862
rect 675375 872860 675441 872863
rect 674432 872858 675441 872860
rect 674432 872802 675380 872858
rect 675436 872802 675441 872858
rect 674432 872800 675441 872802
rect 674432 872798 674438 872800
rect 675375 872797 675441 872800
rect 654447 871232 654513 871235
rect 650208 871230 654513 871232
rect 650208 871174 654452 871230
rect 654508 871174 654513 871230
rect 650208 871172 654513 871174
rect 654447 871169 654513 871172
rect 675130 869838 675136 869902
rect 675200 869900 675206 869902
rect 675375 869900 675441 869903
rect 675200 869898 675441 869900
rect 675200 869842 675380 869898
rect 675436 869842 675441 869898
rect 675200 869840 675441 869842
rect 675200 869838 675206 869840
rect 675375 869837 675441 869840
rect 675375 864722 675441 864723
rect 675322 864720 675328 864722
rect 675284 864660 675328 864720
rect 675392 864718 675441 864722
rect 675436 864662 675441 864718
rect 675322 864658 675328 864660
rect 675392 864658 675441 864662
rect 675375 864657 675441 864658
rect 674895 862204 674961 862207
rect 675183 862204 675249 862207
rect 674895 862202 675249 862204
rect 674895 862146 674900 862202
rect 674956 862146 675188 862202
rect 675244 862146 675249 862202
rect 674895 862144 675249 862146
rect 674895 862141 674961 862144
rect 675183 862141 675249 862144
rect 58575 860428 58641 860431
rect 58575 860426 64416 860428
rect 58575 860370 58580 860426
rect 58636 860370 64416 860426
rect 58575 860368 64416 860370
rect 58575 860365 58641 860368
rect 654159 859540 654225 859543
rect 650208 859538 654225 859540
rect 650208 859482 654164 859538
rect 654220 859482 654225 859538
rect 650208 859480 654225 859482
rect 654159 859477 654225 859480
rect 649743 848292 649809 848295
rect 649743 848290 649854 848292
rect 649743 848234 649748 848290
rect 649804 848234 649854 848290
rect 649743 848229 649854 848234
rect 649794 847670 649854 848229
rect 59535 846072 59601 846075
rect 59535 846070 64416 846072
rect 59535 846014 59540 846070
rect 59596 846014 64416 846070
rect 59535 846012 64416 846014
rect 59535 846009 59601 846012
rect 38170 841394 45946 841526
rect 38170 837942 44902 841394
rect 43396 832312 44902 837942
rect 38826 828278 44902 832312
rect 45730 828278 45946 841394
rect 653967 836008 654033 836011
rect 650208 836006 654033 836008
rect 650208 835950 653972 836006
rect 654028 835950 654033 836006
rect 650208 835948 654033 835950
rect 653967 835945 654033 835948
rect 668662 832500 673560 832542
rect 668662 832382 679954 832500
rect 59535 831716 59601 831719
rect 59535 831714 64416 831716
rect 59535 831658 59540 831714
rect 59596 831658 64416 831714
rect 59535 831656 64416 831658
rect 59535 831653 59601 831656
rect 38826 828272 45946 828278
rect 6142 825720 8804 826520
rect 9604 826519 50926 826520
rect 9604 825721 50127 826519
rect 50925 825721 50931 826519
rect 9604 825720 50926 825721
rect 5860 824258 16354 825058
rect 17154 825057 52718 825058
rect 17154 824259 51919 825057
rect 52717 824259 52723 825057
rect 653967 824316 654033 824319
rect 650208 824314 654033 824316
rect 17154 824258 52718 824259
rect 650208 824258 653972 824314
rect 654028 824258 654033 824314
rect 650208 824256 654033 824258
rect 653967 824253 654033 824256
rect 6474 822700 7284 823500
rect 8084 823499 54502 823500
rect 8084 822701 53703 823499
rect 54501 822701 54507 823499
rect 8084 822700 54502 822701
rect 6804 821426 17446 822226
rect 18246 822225 56068 822226
rect 18246 821427 55269 822225
rect 56067 821427 56073 822225
rect 18246 821426 56068 821427
rect 668662 819526 668858 832382
rect 670730 828600 679954 832382
rect 670730 822546 673560 828600
rect 670730 819526 679356 822546
rect 668662 819350 679356 819526
rect 668662 819328 673560 819350
rect 42639 819136 42705 819139
rect 42528 819134 42705 819136
rect 42528 819078 42644 819134
rect 42700 819078 42705 819134
rect 42528 819076 42705 819078
rect 42639 819073 42705 819076
rect 41679 818840 41745 818843
rect 41679 818838 41790 818840
rect 41679 818782 41684 818838
rect 41740 818782 41790 818838
rect 41679 818777 41790 818782
rect 41730 818514 41790 818777
rect 42639 818100 42705 818103
rect 42498 818098 42705 818100
rect 42498 818042 42644 818098
rect 42700 818042 42705 818098
rect 42498 818040 42705 818042
rect 42498 817922 42558 818040
rect 42639 818037 42705 818040
rect 43215 817508 43281 817511
rect 42528 817506 43281 817508
rect 42528 817450 43220 817506
rect 43276 817450 43281 817506
rect 42528 817448 43281 817450
rect 43215 817445 43281 817448
rect 59535 817360 59601 817363
rect 59535 817358 64416 817360
rect 59535 817302 59540 817358
rect 59596 817302 64416 817358
rect 59535 817300 64416 817302
rect 59535 817297 59601 817300
rect 40335 817212 40401 817215
rect 40335 817210 40446 817212
rect 40335 817154 40340 817210
rect 40396 817154 40446 817210
rect 40335 817149 40446 817154
rect 40386 816886 40446 817149
rect 40239 816768 40305 816771
rect 40194 816766 40305 816768
rect 40194 816710 40244 816766
rect 40300 816710 40305 816766
rect 40194 816705 40305 816710
rect 40194 816294 40254 816705
rect 40378 815966 40384 816030
rect 40448 815966 40454 816030
rect 40386 815850 40446 815966
rect 41730 814995 41790 815258
rect 41730 814990 41841 814995
rect 41730 814934 41780 814990
rect 41836 814934 41841 814990
rect 41730 814932 41841 814934
rect 41775 814929 41841 814932
rect 42498 814400 42558 814666
rect 42639 814400 42705 814403
rect 42498 814398 42705 814400
rect 42498 814342 42644 814398
rect 42700 814342 42705 814398
rect 42498 814340 42705 814342
rect 42639 814337 42705 814340
rect 40578 813958 40638 814222
rect 40570 813894 40576 813958
rect 40640 813894 40646 813958
rect 41730 813367 41790 813630
rect 41679 813362 41790 813367
rect 41679 813306 41684 813362
rect 41740 813306 41790 813362
rect 41679 813304 41790 813306
rect 41679 813301 41745 813304
rect 41922 812775 41982 813038
rect 41922 812770 42033 812775
rect 41922 812714 41972 812770
rect 42028 812714 42033 812770
rect 41922 812712 42033 812714
rect 41967 812709 42033 812712
rect 654447 812624 654513 812627
rect 650208 812622 654513 812624
rect 41922 812331 41982 812594
rect 650208 812566 654452 812622
rect 654508 812566 654513 812622
rect 650208 812564 654513 812566
rect 654447 812561 654513 812564
rect 41871 812326 41982 812331
rect 41871 812270 41876 812326
rect 41932 812270 41982 812326
rect 41871 812268 41982 812270
rect 41871 812265 41937 812268
rect 40770 811738 40830 812002
rect 40762 811674 40768 811738
rect 40832 811674 40838 811738
rect 42114 811147 42174 811410
rect 42063 811142 42174 811147
rect 42063 811086 42068 811142
rect 42124 811086 42174 811142
rect 42063 811084 42174 811086
rect 42063 811081 42129 811084
rect 42114 810555 42174 810966
rect 42114 810550 42225 810555
rect 42114 810494 42164 810550
rect 42220 810494 42225 810550
rect 42114 810492 42225 810494
rect 42159 810489 42225 810492
rect 43023 810404 43089 810407
rect 42528 810402 43089 810404
rect 42528 810346 43028 810402
rect 43084 810346 43089 810402
rect 42528 810344 43089 810346
rect 43023 810341 43089 810344
rect 42306 809519 42366 809782
rect 42306 809514 42417 809519
rect 42306 809458 42356 809514
rect 42412 809458 42417 809514
rect 42306 809456 42417 809458
rect 42351 809453 42417 809456
rect 42735 809294 42801 809297
rect 42528 809292 42801 809294
rect 42528 809236 42740 809292
rect 42796 809236 42801 809292
rect 42528 809234 42801 809236
rect 42735 809231 42801 809234
rect 43119 808776 43185 808779
rect 42528 808774 43185 808776
rect 42528 808718 43124 808774
rect 43180 808718 43185 808774
rect 42528 808716 43185 808718
rect 43119 808713 43185 808716
rect 42831 808184 42897 808187
rect 42528 808182 42897 808184
rect 42528 808126 42836 808182
rect 42892 808126 42897 808182
rect 42528 808124 42897 808126
rect 42831 808121 42897 808124
rect 42498 807296 42558 807636
rect 42498 807236 42750 807296
rect 35202 806855 35262 807118
rect 35151 806850 35262 806855
rect 42690 806852 42750 807236
rect 35151 806794 35156 806850
rect 35212 806794 35262 806850
rect 35151 806792 35262 806794
rect 42498 806792 42750 806852
rect 35151 806789 35217 806792
rect 42498 806556 42558 806792
rect 44559 806556 44625 806559
rect 42498 806554 44625 806556
rect 42498 806526 44564 806554
rect 42528 806498 44564 806526
rect 44620 806498 44625 806554
rect 42528 806496 44625 806498
rect 44559 806493 44625 806496
rect 35151 806408 35217 806411
rect 35151 806406 35262 806408
rect 35151 806350 35156 806406
rect 35212 806350 35262 806406
rect 35151 806345 35262 806350
rect 35202 806008 35262 806345
rect 59535 802856 59601 802859
rect 59535 802854 64416 802856
rect 59535 802798 59540 802854
rect 59596 802798 64416 802854
rect 59535 802796 64416 802798
rect 59535 802793 59601 802796
rect 37359 802116 37425 802119
rect 40954 802116 40960 802118
rect 37359 802114 40960 802116
rect 37359 802058 37364 802114
rect 37420 802058 40960 802114
rect 37359 802056 40960 802058
rect 37359 802053 37425 802056
rect 40954 802054 40960 802056
rect 41024 802054 41030 802118
rect 650223 801376 650289 801379
rect 650178 801374 650289 801376
rect 650178 801318 650228 801374
rect 650284 801318 650289 801374
rect 650178 801313 650289 801318
rect 650178 800754 650238 801313
rect 41914 800426 41920 800490
rect 41984 800488 41990 800490
rect 42063 800488 42129 800491
rect 41984 800486 42129 800488
rect 41984 800430 42068 800486
rect 42124 800430 42129 800486
rect 41984 800428 42129 800430
rect 41984 800426 41990 800428
rect 42063 800425 42129 800428
rect 41967 800340 42033 800343
rect 42298 800340 42304 800342
rect 41967 800338 42304 800340
rect 41967 800282 41972 800338
rect 42028 800282 42304 800338
rect 41967 800280 42304 800282
rect 41967 800277 42033 800280
rect 42298 800278 42304 800280
rect 42368 800278 42374 800342
rect 42351 799748 42417 799751
rect 42490 799748 42496 799750
rect 42351 799746 42496 799748
rect 42351 799690 42356 799746
rect 42412 799690 42496 799746
rect 42351 799688 42496 799690
rect 42351 799685 42417 799688
rect 42490 799686 42496 799688
rect 42560 799686 42566 799750
rect 42106 797614 42112 797678
rect 42176 797676 42182 797678
rect 42447 797676 42513 797679
rect 42176 797674 42513 797676
rect 42176 797618 42452 797674
rect 42508 797618 42513 797674
rect 42176 797616 42513 797618
rect 42176 797614 42182 797616
rect 42447 797613 42513 797616
rect 42447 797530 42513 797531
rect 42447 797528 42496 797530
rect 42404 797526 42496 797528
rect 42404 797470 42452 797526
rect 42404 797468 42496 797470
rect 42447 797466 42496 797468
rect 42560 797466 42566 797530
rect 42447 797465 42513 797466
rect 42298 797022 42304 797086
rect 42368 797084 42374 797086
rect 42543 797084 42609 797087
rect 42368 797082 42609 797084
rect 42368 797026 42548 797082
rect 42604 797026 42609 797082
rect 42368 797024 42609 797026
rect 42368 797022 42374 797024
rect 42543 797021 42609 797024
rect 41914 792582 41920 792646
rect 41984 792644 41990 792646
rect 42543 792644 42609 792647
rect 41984 792642 42609 792644
rect 41984 792586 42548 792642
rect 42604 792586 42609 792642
rect 41984 792584 42609 792586
rect 41984 792582 41990 792584
rect 42543 792581 42609 792584
rect 40762 791842 40768 791906
rect 40832 791904 40838 791906
rect 42351 791904 42417 791907
rect 40832 791902 42417 791904
rect 40832 791846 42356 791902
rect 42412 791846 42417 791902
rect 40832 791844 42417 791846
rect 40832 791842 40838 791844
rect 42351 791841 42417 791844
rect 40570 791694 40576 791758
rect 40640 791756 40646 791758
rect 42447 791756 42513 791759
rect 40640 791754 42513 791756
rect 40640 791698 42452 791754
rect 42508 791698 42513 791754
rect 40640 791696 42513 791698
rect 40640 791694 40646 791696
rect 42447 791693 42513 791696
rect 42063 791314 42129 791315
rect 42063 791312 42112 791314
rect 42020 791310 42112 791312
rect 42020 791254 42068 791310
rect 42020 791252 42112 791254
rect 42063 791250 42112 791252
rect 42176 791250 42182 791314
rect 42063 791249 42129 791250
rect 41722 791102 41728 791166
rect 41792 791164 41798 791166
rect 42159 791164 42225 791167
rect 42682 791164 42688 791166
rect 41792 791162 42688 791164
rect 41792 791106 42164 791162
rect 42220 791106 42688 791162
rect 41792 791104 42688 791106
rect 41792 791102 41798 791104
rect 42159 791101 42225 791104
rect 42682 791102 42688 791104
rect 42752 791102 42758 791166
rect 654063 789092 654129 789095
rect 650208 789090 654129 789092
rect 650208 789034 654068 789090
rect 654124 789034 654129 789090
rect 650208 789032 654129 789034
rect 654063 789029 654129 789032
rect 59535 788648 59601 788651
rect 59535 788646 64416 788648
rect 59535 788590 59540 788646
rect 59596 788590 64416 788646
rect 59535 788588 64416 788590
rect 59535 788585 59601 788588
rect 675759 788056 675825 788059
rect 675898 788056 675904 788058
rect 675759 788054 675904 788056
rect 675759 787998 675764 788054
rect 675820 787998 675904 788054
rect 675759 787996 675904 787998
rect 675759 787993 675825 787996
rect 675898 787994 675904 787996
rect 675968 787994 675974 788058
rect 675471 787170 675537 787171
rect 675471 787166 675520 787170
rect 675584 787168 675590 787170
rect 675471 787110 675476 787166
rect 675471 787106 675520 787110
rect 675584 787108 675628 787168
rect 675584 787106 675590 787108
rect 675471 787105 675537 787106
rect 675759 786724 675825 786727
rect 676090 786724 676096 786726
rect 675759 786722 676096 786724
rect 675759 786666 675764 786722
rect 675820 786666 676096 786722
rect 675759 786664 676096 786666
rect 675759 786661 675825 786664
rect 676090 786662 676096 786664
rect 676160 786662 676166 786726
rect 675759 784948 675825 784951
rect 676282 784948 676288 784950
rect 675759 784946 676288 784948
rect 675759 784890 675764 784946
rect 675820 784890 676288 784946
rect 675759 784888 676288 784890
rect 675759 784885 675825 784888
rect 676282 784886 676288 784888
rect 676352 784886 676358 784950
rect 675663 784210 675729 784211
rect 675663 784206 675712 784210
rect 675776 784208 675782 784210
rect 675663 784150 675668 784206
rect 675663 784146 675712 784150
rect 675776 784148 675820 784208
rect 675776 784146 675782 784148
rect 675663 784145 675729 784146
rect 7168 782976 8578 783776
rect 9378 783775 50926 783776
rect 9378 782977 50127 783775
rect 50925 782977 50931 783775
rect 9378 782976 50926 782977
rect 6604 781848 16310 782648
rect 17110 782647 52718 782648
rect 17110 781849 51919 782647
rect 52717 781849 52723 782647
rect 675759 781988 675825 781991
rect 676666 781988 676672 781990
rect 675759 781986 676672 781988
rect 675759 781930 675764 781986
rect 675820 781930 676672 781986
rect 675759 781928 676672 781930
rect 675759 781925 675825 781928
rect 676666 781926 676672 781928
rect 676736 781926 676742 781990
rect 17110 781848 52718 781849
rect 6042 780440 7234 781240
rect 8034 781239 54502 781240
rect 8034 780441 53703 781239
rect 54501 780441 54507 781239
rect 675759 780656 675825 780659
rect 676474 780656 676480 780658
rect 675759 780654 676480 780656
rect 675759 780598 675764 780654
rect 675820 780598 676480 780654
rect 675759 780596 676480 780598
rect 675759 780593 675825 780596
rect 676474 780594 676480 780596
rect 676544 780594 676550 780658
rect 8034 780440 54502 780441
rect 5712 778984 17582 779784
rect 18382 779783 56068 779784
rect 18382 778985 55269 779783
rect 56067 778985 56073 779783
rect 18382 778984 56068 778985
rect 674511 777548 674577 777551
rect 677050 777548 677056 777550
rect 674511 777546 677056 777548
rect 674511 777490 674516 777546
rect 674572 777490 677056 777546
rect 674511 777488 677056 777490
rect 674511 777485 674577 777488
rect 677050 777486 677056 777488
rect 677120 777486 677126 777550
rect 654063 777400 654129 777403
rect 650208 777398 654129 777400
rect 650208 777342 654068 777398
rect 654124 777342 654129 777398
rect 650208 777340 654129 777342
rect 654063 777337 654129 777340
rect 674607 776956 674673 776959
rect 677050 776956 677056 776958
rect 674607 776954 677056 776956
rect 674607 776898 674612 776954
rect 674668 776898 677056 776954
rect 674607 776896 677056 776898
rect 674607 776893 674673 776896
rect 677050 776894 677056 776896
rect 677120 776894 677126 776958
rect 674895 776216 674961 776219
rect 677050 776216 677056 776218
rect 674895 776214 677056 776216
rect 674895 776158 674900 776214
rect 674956 776158 677056 776214
rect 674895 776156 677056 776158
rect 674895 776153 674961 776156
rect 677050 776154 677056 776156
rect 677120 776154 677126 776218
rect 42447 776068 42513 776071
rect 42447 776066 42558 776068
rect 42447 776010 42452 776066
rect 42508 776010 42558 776066
rect 42447 776005 42558 776010
rect 42498 775890 42558 776005
rect 42831 775328 42897 775331
rect 42528 775326 42897 775328
rect 42528 775270 42836 775326
rect 42892 775270 42897 775326
rect 42528 775268 42897 775270
rect 42831 775265 42897 775268
rect 674895 774884 674961 774887
rect 676858 774884 676864 774886
rect 674895 774882 676864 774884
rect 674895 774826 674900 774882
rect 674956 774826 676864 774882
rect 674895 774824 676864 774826
rect 674895 774821 674961 774824
rect 676858 774822 676864 774824
rect 676928 774822 676934 774886
rect 42831 774810 42897 774813
rect 42528 774808 42897 774810
rect 42528 774752 42836 774808
rect 42892 774752 42897 774808
rect 42528 774750 42897 774752
rect 42831 774747 42897 774750
rect 43407 774292 43473 774295
rect 42528 774290 43473 774292
rect 42528 774234 43412 774290
rect 43468 774234 43473 774290
rect 42528 774232 43473 774234
rect 43407 774229 43473 774232
rect 59535 774144 59601 774147
rect 59535 774142 64416 774144
rect 59535 774086 59540 774142
rect 59596 774086 64416 774142
rect 59535 774084 64416 774086
rect 59535 774081 59601 774084
rect 43215 773700 43281 773703
rect 42528 773698 43281 773700
rect 42528 773642 43220 773698
rect 43276 773642 43281 773698
rect 42528 773640 43281 773642
rect 43215 773637 43281 773640
rect 40954 773342 40960 773406
rect 41024 773342 41030 773406
rect 40962 773182 41022 773342
rect 40416 773152 41022 773182
rect 40386 773122 40992 773152
rect 40386 772814 40446 773122
rect 674319 773108 674385 773111
rect 677626 773108 677632 773110
rect 674319 773106 677632 773108
rect 674319 773050 674324 773106
rect 674380 773050 677632 773106
rect 674319 773048 677632 773050
rect 674319 773045 674385 773048
rect 677626 773046 677632 773048
rect 677696 773046 677702 773110
rect 40378 772750 40384 772814
rect 40448 772750 40454 772814
rect 40578 772370 40638 772634
rect 40570 772306 40576 772370
rect 40640 772306 40646 772370
rect 43023 772072 43089 772075
rect 42528 772070 43089 772072
rect 42528 772014 43028 772070
rect 43084 772014 43089 772070
rect 42528 772012 43089 772014
rect 43023 772009 43089 772012
rect 671682 771920 699229 771921
rect 42114 771187 42174 771524
rect 42063 771182 42174 771187
rect 42063 771126 42068 771182
rect 42124 771126 42174 771182
rect 42063 771124 42174 771126
rect 42063 771121 42129 771124
rect 40194 770743 40254 771006
rect 671677 770828 671683 771920
rect 672775 770828 699229 771920
rect 671682 770827 699229 770828
rect 700323 770827 711635 771921
rect 40194 770738 40305 770743
rect 40194 770682 40244 770738
rect 40300 770682 40305 770738
rect 40194 770680 40305 770682
rect 40239 770677 40305 770680
rect 666066 770527 709390 770528
rect 42831 770444 42897 770447
rect 42528 770442 42897 770444
rect 42528 770386 42836 770442
rect 42892 770386 42897 770442
rect 42528 770384 42897 770386
rect 42831 770381 42897 770384
rect 41730 769559 41790 769896
rect 41679 769554 41790 769559
rect 41679 769498 41684 769554
rect 41740 769498 41790 769554
rect 41679 769496 41790 769498
rect 41679 769493 41745 769496
rect 42306 769115 42366 769378
rect 666061 769345 666067 770527
rect 667249 769345 709390 770527
rect 666066 769344 709390 769345
rect 710574 769344 711450 770528
rect 42306 769110 42417 769115
rect 42306 769054 42356 769110
rect 42412 769054 42417 769110
rect 42306 769052 42417 769054
rect 42351 769049 42417 769052
rect 41346 768670 41406 768786
rect 41338 768606 41344 768670
rect 41408 768606 41414 768670
rect 662178 768629 700828 768630
rect 42114 767931 42174 768194
rect 42114 767926 42225 767931
rect 42114 767870 42164 767926
rect 42220 767870 42225 767926
rect 42114 767868 42225 767870
rect 42159 767865 42225 767868
rect 42927 767780 42993 767783
rect 42528 767778 42993 767780
rect 42528 767722 42932 767778
rect 42988 767722 42993 767778
rect 42528 767720 42993 767722
rect 42927 767717 42993 767720
rect 662173 767447 662179 768629
rect 663361 767447 700828 768629
rect 662178 767446 700828 767447
rect 702012 767446 711624 768630
rect 43119 767188 43185 767191
rect 42528 767186 43185 767188
rect 42528 767130 43124 767186
rect 43180 767130 43185 767186
rect 42528 767128 43185 767130
rect 43119 767125 43185 767128
rect 659368 766959 707978 766960
rect 41922 766303 41982 766566
rect 41871 766298 41982 766303
rect 41871 766242 41876 766298
rect 41932 766242 41982 766298
rect 41871 766240 41982 766242
rect 41871 766237 41937 766240
rect 41730 765859 41790 766122
rect 41730 765854 41841 765859
rect 41730 765798 41780 765854
rect 41836 765798 41841 765854
rect 41730 765796 41841 765798
rect 41775 765793 41841 765796
rect 659363 765777 659369 766959
rect 660551 765777 707978 766959
rect 659368 765776 707978 765777
rect 709162 765776 711336 766960
rect 653967 765560 654033 765563
rect 650208 765558 654033 765560
rect 42306 765266 42366 765530
rect 650208 765502 653972 765558
rect 654028 765502 654033 765558
rect 650208 765500 654033 765502
rect 653967 765497 654033 765500
rect 42298 765202 42304 765266
rect 42368 765202 42374 765266
rect 41538 764823 41598 764938
rect 41538 764818 41649 764823
rect 41538 764762 41588 764818
rect 41644 764762 41649 764818
rect 41538 764760 41649 764762
rect 41583 764757 41649 764760
rect 42498 764080 42558 764494
rect 42498 764020 42750 764080
rect 35202 763639 35262 763902
rect 35151 763634 35262 763639
rect 42690 763636 42750 764020
rect 35151 763578 35156 763634
rect 35212 763578 35262 763634
rect 35151 763576 35262 763578
rect 42306 763576 42750 763636
rect 35151 763573 35217 763576
rect 42306 763340 42366 763576
rect 53295 763340 53361 763343
rect 42306 763310 42528 763340
rect 42690 763338 53361 763340
rect 42336 763280 42558 763310
rect 35151 763192 35217 763195
rect 42498 763192 42558 763280
rect 42690 763282 53300 763338
rect 53356 763282 53361 763338
rect 42690 763280 53361 763282
rect 42690 763192 42750 763280
rect 53295 763277 53361 763280
rect 35151 763190 35262 763192
rect 35151 763134 35156 763190
rect 35212 763134 35262 763190
rect 35151 763129 35262 763134
rect 42498 763132 42750 763192
rect 35202 762866 35262 763129
rect 674319 762896 674385 762899
rect 674319 762894 674784 762896
rect 674319 762838 674324 762894
rect 674380 762838 674784 762894
rect 674319 762836 674784 762838
rect 674319 762833 674385 762836
rect 674319 762304 674385 762307
rect 674319 762302 674784 762304
rect 674319 762246 674324 762302
rect 674380 762246 674784 762302
rect 674319 762244 674784 762246
rect 674319 762241 674385 762244
rect 674607 762008 674673 762011
rect 674607 762006 674814 762008
rect 674607 761950 674612 762006
rect 674668 761950 674814 762006
rect 674607 761948 674814 761950
rect 674607 761945 674673 761948
rect 674754 761830 674814 761948
rect 673839 761268 673905 761271
rect 673839 761266 674784 761268
rect 673839 761210 673844 761266
rect 673900 761210 674784 761266
rect 673839 761208 674784 761210
rect 673839 761205 673905 761208
rect 673839 760676 673905 760679
rect 673839 760674 674784 760676
rect 673839 760618 673844 760674
rect 673900 760618 674784 760674
rect 673839 760616 674784 760618
rect 673839 760613 673905 760616
rect 677050 760318 677056 760382
rect 677120 760380 677126 760382
rect 677871 760380 677937 760383
rect 677120 760378 677937 760380
rect 677120 760322 677876 760378
rect 677932 760322 677937 760378
rect 677120 760320 677937 760322
rect 677120 760318 677126 760320
rect 677871 760317 677937 760320
rect 40239 760232 40305 760235
rect 40762 760232 40768 760234
rect 40239 760230 40768 760232
rect 40239 760174 40244 760230
rect 40300 760174 40768 760230
rect 40239 760172 40768 760174
rect 40239 760169 40305 760172
rect 40762 760170 40768 760172
rect 40832 760170 40838 760234
rect 42063 760232 42129 760235
rect 42490 760232 42496 760234
rect 42063 760230 42496 760232
rect 42063 760174 42068 760230
rect 42124 760174 42496 760230
rect 42063 760172 42496 760174
rect 42063 760169 42129 760172
rect 42490 760170 42496 760172
rect 42560 760170 42566 760234
rect 676866 759791 676926 760202
rect 677871 759938 677937 759939
rect 677818 759874 677824 759938
rect 677888 759936 677937 759938
rect 677888 759934 677980 759936
rect 677932 759878 677980 759934
rect 677888 759876 677980 759878
rect 677888 759874 677937 759876
rect 677871 759873 677937 759874
rect 59535 759788 59601 759791
rect 59535 759786 64416 759788
rect 59535 759730 59540 759786
rect 59596 759730 64416 759786
rect 59535 759728 64416 759730
rect 676866 759786 676977 759791
rect 676866 759730 676916 759786
rect 676972 759730 676977 759786
rect 676866 759728 676977 759730
rect 59535 759725 59601 759728
rect 676911 759725 676977 759728
rect 677634 759347 677694 759610
rect 674554 759282 674560 759346
rect 674624 759344 674630 759346
rect 674624 759284 674814 759344
rect 674624 759282 674630 759284
rect 42831 759196 42897 759199
rect 43066 759196 43072 759198
rect 42831 759194 43072 759196
rect 42831 759138 42836 759194
rect 42892 759138 43072 759194
rect 42831 759136 43072 759138
rect 42831 759133 42897 759136
rect 43066 759134 43072 759136
rect 43136 759134 43142 759198
rect 674754 759018 674814 759284
rect 677583 759342 677694 759347
rect 677583 759286 677588 759342
rect 677644 759286 677694 759342
rect 677583 759284 677694 759286
rect 677583 759281 677649 759284
rect 675322 758838 675328 758902
rect 675392 758838 675398 758902
rect 675330 758574 675390 758838
rect 674746 758246 674752 758310
rect 674816 758246 674822 758310
rect 674754 757982 674814 758246
rect 41583 757422 41649 757423
rect 41530 757420 41536 757422
rect 41492 757360 41536 757420
rect 41600 757418 41649 757422
rect 41644 757362 41649 757418
rect 41530 757358 41536 757360
rect 41600 757358 41649 757362
rect 674170 757358 674176 757422
rect 674240 757420 674246 757422
rect 674240 757360 674784 757420
rect 674240 757358 674246 757360
rect 41583 757357 41649 757358
rect 675130 757210 675136 757274
rect 675200 757210 675206 757274
rect 41871 757126 41937 757127
rect 41871 757122 41920 757126
rect 41984 757124 41990 757126
rect 42159 757124 42225 757127
rect 42682 757124 42688 757126
rect 41871 757066 41876 757122
rect 41871 757062 41920 757066
rect 41984 757064 42028 757124
rect 42159 757122 42688 757124
rect 42159 757066 42164 757122
rect 42220 757066 42688 757122
rect 42159 757064 42688 757066
rect 41984 757062 41990 757064
rect 41871 757061 41937 757062
rect 42159 757061 42225 757064
rect 42682 757062 42688 757064
rect 42752 757062 42758 757126
rect 675138 756872 675198 757210
rect 676858 756618 676864 756682
rect 676928 756618 676934 756682
rect 676866 756354 676926 756618
rect 676911 756090 676977 756091
rect 676858 756088 676864 756090
rect 676820 756028 676864 756088
rect 676928 756086 676977 756090
rect 676972 756030 676977 756086
rect 676858 756026 676864 756028
rect 676928 756026 676977 756030
rect 676911 756025 676977 756026
rect 673978 755730 673984 755794
rect 674048 755792 674054 755794
rect 674048 755732 674784 755792
rect 674048 755730 674054 755732
rect 674938 755582 674944 755646
rect 675008 755582 675014 755646
rect 674946 755244 675006 755582
rect 42063 754904 42129 754907
rect 42490 754904 42496 754906
rect 42063 754902 42496 754904
rect 42063 754846 42068 754902
rect 42124 754846 42496 754902
rect 42063 754844 42496 754846
rect 42063 754841 42129 754844
rect 42490 754842 42496 754844
rect 42560 754842 42566 754906
rect 674362 754694 674368 754758
rect 674432 754756 674438 754758
rect 674432 754696 674784 754756
rect 674432 754694 674438 754696
rect 650031 754460 650097 754463
rect 649986 754458 650097 754460
rect 649986 754402 650036 754458
rect 650092 754402 650097 754458
rect 649986 754397 650097 754402
rect 677434 754398 677440 754462
rect 677504 754398 677510 754462
rect 649986 753838 650046 754397
rect 677442 754134 677502 754398
rect 677626 753954 677632 754018
rect 677696 753954 677702 754018
rect 677634 753616 677694 753954
rect 677583 753426 677649 753427
rect 677242 753362 677248 753426
rect 677312 753362 677318 753426
rect 677583 753422 677632 753426
rect 677696 753424 677702 753426
rect 677583 753366 677588 753422
rect 677583 753362 677632 753366
rect 677696 753364 677740 753424
rect 677696 753362 677702 753364
rect 677250 753098 677310 753362
rect 677583 753361 677649 753362
rect 677818 752770 677824 752834
rect 677888 752770 677894 752834
rect 677826 752506 677886 752770
rect 673359 752092 673425 752095
rect 673359 752090 674814 752092
rect 673359 752034 673364 752090
rect 673420 752034 674814 752090
rect 673359 752032 674814 752034
rect 673359 752029 673425 752032
rect 674754 751988 674814 752032
rect 42874 751882 42880 751946
rect 42944 751944 42950 751946
rect 43023 751944 43089 751947
rect 42944 751942 43089 751944
rect 42944 751886 43028 751942
rect 43084 751886 43089 751942
rect 42944 751884 43089 751886
rect 42944 751882 42950 751884
rect 43023 751881 43089 751884
rect 41530 751734 41536 751798
rect 41600 751796 41606 751798
rect 42063 751796 42129 751799
rect 41600 751794 42129 751796
rect 41600 751738 42068 751794
rect 42124 751738 42129 751794
rect 41600 751736 42129 751738
rect 41600 751734 41606 751736
rect 42063 751733 42129 751736
rect 42735 751650 42801 751651
rect 42682 751586 42688 751650
rect 42752 751648 42801 751650
rect 42752 751646 42844 751648
rect 42796 751590 42844 751646
rect 42752 751588 42844 751590
rect 42752 751586 42801 751588
rect 42735 751585 42801 751586
rect 677058 751207 677118 751470
rect 677007 751202 677118 751207
rect 677007 751146 677012 751202
rect 677068 751146 677118 751202
rect 677007 751144 677118 751146
rect 677007 751141 677073 751144
rect 41871 751058 41937 751059
rect 41871 751054 41920 751058
rect 41984 751056 41990 751058
rect 41871 750998 41876 751054
rect 41871 750994 41920 750998
rect 41984 750996 42028 751056
rect 41984 750994 41990 750996
rect 41871 750993 41937 750994
rect 676866 750615 676926 750878
rect 42159 750612 42225 750615
rect 42298 750612 42304 750614
rect 42159 750610 42304 750612
rect 42159 750554 42164 750610
rect 42220 750554 42304 750610
rect 42159 750552 42304 750554
rect 42159 750549 42225 750552
rect 42298 750550 42304 750552
rect 42368 750550 42374 750614
rect 676815 750610 676926 750615
rect 676815 750554 676820 750610
rect 676876 750554 676926 750610
rect 676815 750552 676926 750554
rect 677007 750612 677073 750615
rect 677007 750610 677118 750612
rect 677007 750554 677012 750610
rect 677068 750554 677118 750610
rect 676815 750549 676881 750552
rect 677007 750549 677118 750554
rect 677058 750360 677118 750549
rect 43023 750318 43089 750319
rect 43023 750316 43072 750318
rect 42980 750314 43072 750316
rect 42980 750258 43028 750314
rect 42980 750256 43072 750258
rect 43023 750254 43072 750256
rect 43136 750254 43142 750318
rect 43023 750253 43089 750254
rect 676815 750168 676881 750171
rect 676815 750166 676926 750168
rect 676815 750110 676820 750166
rect 676876 750110 676926 750166
rect 676815 750105 676926 750110
rect 676866 749842 676926 750105
rect 42831 749726 42897 749727
rect 42831 749724 42880 749726
rect 42788 749722 42880 749724
rect 42788 749666 42836 749722
rect 42788 749664 42880 749666
rect 42831 749662 42880 749664
rect 42944 749662 42950 749726
rect 42831 749661 42897 749662
rect 41967 748690 42033 748691
rect 41914 748626 41920 748690
rect 41984 748688 42033 748690
rect 41984 748686 42076 748688
rect 42028 748630 42076 748686
rect 41984 748628 42076 748630
rect 41984 748626 42033 748628
rect 41967 748625 42033 748626
rect 41530 747146 41536 747210
rect 41600 747208 41606 747210
rect 41775 747208 41841 747211
rect 41600 747206 41841 747208
rect 41600 747150 41780 747206
rect 41836 747150 41841 747206
rect 41600 747148 41841 747150
rect 41600 747146 41606 747148
rect 41775 747145 41841 747148
rect 40762 746850 40768 746914
rect 40832 746912 40838 746914
rect 43119 746912 43185 746915
rect 40832 746910 43185 746912
rect 40832 746854 43124 746910
rect 43180 746854 43185 746910
rect 40832 746852 43185 746854
rect 40832 746850 40838 746852
rect 43119 746849 43185 746852
rect 41338 746110 41344 746174
rect 41408 746172 41414 746174
rect 42735 746172 42801 746175
rect 41408 746170 42801 746172
rect 41408 746114 42740 746170
rect 42796 746114 42801 746170
rect 41408 746112 42801 746114
rect 41408 746110 41414 746112
rect 42735 746109 42801 746112
rect 59535 745580 59601 745583
rect 59535 745578 64416 745580
rect 59535 745522 59540 745578
rect 59596 745522 64416 745578
rect 59535 745520 64416 745522
rect 59535 745517 59601 745520
rect 676858 744482 676864 744546
rect 676928 744544 676934 744546
rect 677242 744544 677248 744546
rect 676928 744484 677248 744544
rect 676928 744482 676934 744484
rect 677242 744482 677248 744484
rect 677312 744482 677318 744546
rect 676858 744334 676864 744398
rect 676928 744396 676934 744398
rect 677626 744396 677632 744398
rect 676928 744336 677632 744396
rect 676928 744334 676934 744336
rect 677626 744334 677632 744336
rect 677696 744334 677702 744398
rect 674170 743150 674176 743214
rect 674240 743212 674246 743214
rect 675375 743212 675441 743215
rect 674240 743210 675441 743212
rect 674240 743154 675380 743210
rect 675436 743154 675441 743210
rect 674240 743152 675441 743154
rect 674240 743150 674246 743152
rect 675375 743149 675441 743152
rect 673978 742410 673984 742474
rect 674048 742472 674054 742474
rect 675471 742472 675537 742475
rect 674048 742470 675537 742472
rect 674048 742414 675476 742470
rect 675532 742414 675537 742470
rect 674048 742412 675537 742414
rect 674048 742410 674054 742412
rect 675471 742409 675537 742412
rect 653967 742176 654033 742179
rect 650208 742174 654033 742176
rect 650208 742118 653972 742174
rect 654028 742118 654033 742174
rect 650208 742116 654033 742118
rect 653967 742113 654033 742116
rect 674362 741670 674368 741734
rect 674432 741732 674438 741734
rect 675471 741732 675537 741735
rect 674432 741730 675537 741732
rect 674432 741674 675476 741730
rect 675532 741674 675537 741730
rect 674432 741672 675537 741674
rect 674432 741670 674438 741672
rect 675471 741669 675537 741672
rect 6206 739788 8760 740588
rect 9560 740587 50926 740588
rect 9560 739789 50127 740587
rect 50925 739789 50931 740587
rect 675183 740400 675249 740403
rect 676666 740400 676672 740402
rect 675183 740398 676672 740400
rect 675183 740342 675188 740398
rect 675244 740342 676672 740398
rect 675183 740340 676672 740342
rect 675183 740337 675249 740340
rect 676666 740338 676672 740340
rect 676736 740338 676742 740402
rect 675130 740042 675136 740106
rect 675200 740104 675206 740106
rect 675375 740104 675441 740107
rect 675200 740102 675441 740104
rect 675200 740046 675380 740102
rect 675436 740046 675441 740102
rect 675200 740044 675441 740046
rect 675200 740042 675206 740044
rect 675375 740041 675441 740044
rect 9560 739788 50926 739789
rect 6206 738434 16424 739234
rect 17224 739233 52718 739234
rect 17224 738435 51919 739233
rect 52717 738435 52723 739233
rect 674938 739154 674944 739218
rect 675008 739216 675014 739218
rect 675471 739216 675537 739219
rect 675008 739214 675537 739216
rect 675008 739158 675476 739214
rect 675532 739158 675537 739214
rect 675008 739156 675537 739158
rect 675008 739154 675014 739156
rect 675471 739153 675537 739156
rect 674746 738562 674752 738626
rect 674816 738624 674822 738626
rect 675375 738624 675441 738627
rect 674816 738622 675441 738624
rect 674816 738566 675380 738622
rect 675436 738566 675441 738622
rect 674816 738564 675441 738566
rect 674816 738562 674822 738564
rect 675375 738561 675441 738564
rect 17224 738434 52718 738435
rect 5926 737032 7422 737832
rect 8222 737831 54502 737832
rect 8222 737033 53703 737831
rect 54501 737033 54507 737831
rect 8222 737032 54502 737033
rect 6160 735350 17528 736150
rect 18328 736149 56068 736150
rect 18328 735351 55269 736149
rect 56067 735351 56073 736149
rect 18328 735350 56068 735351
rect 675375 734482 675441 734483
rect 675322 734480 675328 734482
rect 675284 734420 675328 734480
rect 675392 734478 675441 734482
rect 675436 734422 675441 734478
rect 675322 734418 675328 734420
rect 675392 734418 675441 734422
rect 675375 734417 675441 734418
rect 42735 732704 42801 732707
rect 42528 732702 42801 732704
rect 42528 732646 42740 732702
rect 42796 732646 42801 732702
rect 42528 732644 42801 732646
rect 42735 732641 42801 732644
rect 42735 732112 42801 732115
rect 42528 732110 42801 732112
rect 42528 732054 42740 732110
rect 42796 732054 42801 732110
rect 42528 732052 42801 732054
rect 42735 732049 42801 732052
rect 42351 731816 42417 731819
rect 42306 731814 42417 731816
rect 42306 731758 42356 731814
rect 42412 731758 42417 731814
rect 42306 731753 42417 731758
rect 42306 731638 42366 731753
rect 43695 731076 43761 731079
rect 42528 731074 43761 731076
rect 42528 731018 43700 731074
rect 43756 731018 43761 731074
rect 42528 731016 43761 731018
rect 43695 731013 43761 731016
rect 59535 731076 59601 731079
rect 59535 731074 64416 731076
rect 59535 731018 59540 731074
rect 59596 731018 64416 731074
rect 59535 731016 64416 731018
rect 59535 731013 59601 731016
rect 43407 730484 43473 730487
rect 655215 730484 655281 730487
rect 42528 730482 43473 730484
rect 42528 730426 43412 730482
rect 43468 730426 43473 730482
rect 42528 730424 43473 730426
rect 650208 730482 655281 730484
rect 650208 730426 655220 730482
rect 655276 730426 655281 730482
rect 650208 730424 655281 730426
rect 43407 730421 43473 730424
rect 655215 730421 655281 730424
rect 40578 729598 40638 729936
rect 40570 729534 40576 729598
rect 40640 729534 40646 729598
rect 41154 729154 41214 729418
rect 41146 729090 41152 729154
rect 41216 729090 41222 729154
rect 41538 728711 41598 728826
rect 41538 728706 41649 728711
rect 41538 728650 41588 728706
rect 41644 728650 41649 728706
rect 41538 728648 41649 728650
rect 41583 728645 41649 728648
rect 41922 727971 41982 728308
rect 674511 728116 674577 728119
rect 677242 728116 677248 728118
rect 674511 728114 677248 728116
rect 674511 728058 674516 728114
rect 674572 728058 677248 728114
rect 674511 728056 677248 728058
rect 674511 728053 674577 728056
rect 677242 728054 677248 728056
rect 677312 728054 677318 728118
rect 41871 727966 41982 727971
rect 41871 727910 41876 727966
rect 41932 727910 41982 727966
rect 41871 727908 41982 727910
rect 41871 727905 41937 727908
rect 41346 727526 41406 727790
rect 671682 727724 699315 727725
rect 41338 727462 41344 727526
rect 41408 727462 41414 727526
rect 41730 726935 41790 727198
rect 41679 726930 41790 726935
rect 41679 726874 41684 726930
rect 41740 726874 41790 726930
rect 41679 726872 41790 726874
rect 41679 726869 41745 726872
rect 41730 726343 41790 726680
rect 671677 726632 671683 727724
rect 672775 726632 699315 727724
rect 671682 726631 699315 726632
rect 700409 726631 711179 727725
rect 41730 726338 41841 726343
rect 41730 726282 41780 726338
rect 41836 726282 41841 726338
rect 41730 726280 41841 726282
rect 41775 726277 41841 726280
rect 42306 725899 42366 726162
rect 676666 725982 676672 726046
rect 676736 726044 676742 726046
rect 676736 725984 677502 726044
rect 676736 725982 676742 725984
rect 42306 725894 42417 725899
rect 677442 725898 677502 725984
rect 42306 725838 42356 725894
rect 42412 725838 42417 725894
rect 42306 725836 42417 725838
rect 42351 725833 42417 725836
rect 677434 725834 677440 725898
rect 677504 725834 677510 725898
rect 40962 725306 41022 725570
rect 666066 725405 709350 725406
rect 40954 725242 40960 725306
rect 41024 725242 41030 725306
rect 42874 725082 42880 725084
rect 42528 725022 42880 725082
rect 42874 725020 42880 725022
rect 42944 725020 42950 725084
rect 40770 724271 40830 724534
rect 40719 724266 40830 724271
rect 40719 724210 40724 724266
rect 40780 724210 40830 724266
rect 666061 724223 666067 725405
rect 667249 724223 709350 725405
rect 666066 724222 709350 724223
rect 710534 724222 710694 725406
rect 40719 724208 40830 724210
rect 40719 724205 40785 724208
rect 42114 723679 42174 723942
rect 42114 723674 42225 723679
rect 42114 723618 42164 723674
rect 42220 723618 42225 723674
rect 42114 723616 42225 723618
rect 42159 723613 42225 723616
rect 41538 723087 41598 723424
rect 662178 723371 700686 723372
rect 41487 723082 41598 723087
rect 41487 723026 41492 723082
rect 41548 723026 41598 723082
rect 41487 723024 41598 723026
rect 41487 723021 41553 723024
rect 43023 722936 43089 722939
rect 42528 722934 43089 722936
rect 42528 722878 43028 722934
rect 43084 722878 43089 722934
rect 42528 722876 43089 722878
rect 43023 722873 43089 722876
rect 41730 722050 41790 722314
rect 662173 722189 662179 723371
rect 663361 722189 700686 723371
rect 662178 722188 700686 722189
rect 701870 722188 710750 723372
rect 41722 721986 41728 722050
rect 41792 721986 41798 722050
rect 42735 721826 42801 721829
rect 42528 721824 42801 721826
rect 42528 721768 42740 721824
rect 42796 721768 42801 721824
rect 42528 721766 42801 721768
rect 42735 721763 42801 721766
rect 659368 721281 708076 721282
rect 42498 721012 42558 721278
rect 42498 720952 42750 721012
rect 35202 720423 35262 720686
rect 42690 720568 42750 720952
rect 35151 720418 35262 720423
rect 35151 720362 35156 720418
rect 35212 720362 35262 720418
rect 35151 720360 35262 720362
rect 42498 720508 42750 720568
rect 35151 720357 35217 720360
rect 42498 720124 42558 720508
rect 53391 720124 53457 720127
rect 42498 720122 53457 720124
rect 42498 720066 53396 720122
rect 53452 720066 53457 720122
rect 659363 720099 659369 721281
rect 660551 720099 708076 721281
rect 659368 720098 708076 720099
rect 709260 720098 710694 721282
rect 42498 720064 53457 720066
rect 53391 720061 53457 720064
rect 35151 719976 35217 719979
rect 35151 719974 35262 719976
rect 35151 719918 35156 719974
rect 35212 719918 35262 719974
rect 35151 719913 35262 719918
rect 35202 719650 35262 719913
rect 654255 718644 654321 718647
rect 650208 718642 654321 718644
rect 650208 718586 654260 718642
rect 654316 718586 654321 718642
rect 650208 718584 654321 718586
rect 654255 718581 654321 718584
rect 674415 717904 674481 717907
rect 674415 717902 674784 717904
rect 674415 717846 674420 717902
rect 674476 717846 674784 717902
rect 674415 717844 674784 717846
rect 674415 717841 674481 717844
rect 674415 717312 674481 717315
rect 674415 717310 674784 717312
rect 674415 717254 674420 717310
rect 674476 717254 674784 717310
rect 674415 717252 674784 717254
rect 674415 717249 674481 717252
rect 674415 716868 674481 716871
rect 674415 716866 674784 716868
rect 674415 716810 674420 716866
rect 674476 716810 674784 716866
rect 674415 716808 674784 716810
rect 674415 716805 674481 716808
rect 59535 716720 59601 716723
rect 59535 716718 64416 716720
rect 59535 716662 59540 716718
rect 59596 716662 64416 716718
rect 59535 716660 64416 716662
rect 59535 716657 59601 716660
rect 674415 716276 674481 716279
rect 674415 716274 674784 716276
rect 674415 716218 674420 716274
rect 674476 716218 674784 716274
rect 674415 716216 674784 716218
rect 674415 716213 674481 716216
rect 43244 715834 43342 715848
rect 41914 715770 41920 715834
rect 41984 715832 41990 715834
rect 43244 715832 43270 715834
rect 41984 715772 43270 715832
rect 41984 715770 41990 715772
rect 43244 715770 43270 715772
rect 43334 715770 43342 715834
rect 43244 715748 43342 715770
rect 41530 715622 41536 715686
rect 41600 715684 41606 715686
rect 42490 715684 42496 715686
rect 41600 715624 42496 715684
rect 41600 715622 41606 715624
rect 42490 715622 42496 715624
rect 42560 715622 42566 715686
rect 673743 715684 673809 715687
rect 673743 715682 674784 715684
rect 673743 715626 673748 715682
rect 673804 715626 674784 715682
rect 673743 715624 674784 715626
rect 673743 715621 673809 715624
rect 676858 715474 676864 715538
rect 676928 715536 676934 715538
rect 676928 715476 677502 715536
rect 676928 715474 676934 715476
rect 677442 714946 677502 715476
rect 677434 714882 677440 714946
rect 677504 714882 677510 714946
rect 677626 714882 677632 714946
rect 677696 714882 677702 714946
rect 677634 714648 677694 714882
rect 677088 714618 677694 714648
rect 677058 714588 677664 714618
rect 41583 714352 41649 714355
rect 677058 714354 677118 714588
rect 43066 714352 43072 714354
rect 41583 714350 43072 714352
rect 41583 714294 41588 714350
rect 41644 714294 43072 714350
rect 41583 714292 43072 714294
rect 41583 714289 41649 714292
rect 43066 714290 43072 714292
rect 43136 714290 43142 714354
rect 676090 714290 676096 714354
rect 676160 714290 676166 714354
rect 677050 714290 677056 714354
rect 677120 714290 677126 714354
rect 40719 714206 40785 714207
rect 40719 714202 40768 714206
rect 40832 714204 40838 714206
rect 41487 714204 41553 714207
rect 41722 714204 41728 714206
rect 40719 714146 40724 714202
rect 40719 714142 40768 714146
rect 40832 714144 40876 714204
rect 41487 714202 41728 714204
rect 41487 714146 41492 714202
rect 41548 714146 41728 714202
rect 41487 714144 41728 714146
rect 40832 714142 40838 714144
rect 40719 714141 40785 714142
rect 41487 714141 41553 714144
rect 41722 714142 41728 714144
rect 41792 714142 41798 714206
rect 676098 714026 676158 714290
rect 41871 713910 41937 713911
rect 42159 713910 42225 713911
rect 41871 713908 41920 713910
rect 41828 713906 41920 713908
rect 41828 713850 41876 713906
rect 41828 713848 41920 713850
rect 41871 713846 41920 713848
rect 41984 713846 41990 713910
rect 42106 713908 42112 713910
rect 42068 713848 42112 713908
rect 42176 713906 42225 713910
rect 42220 713850 42225 713906
rect 42106 713846 42112 713848
rect 42176 713846 42225 713850
rect 41871 713845 41937 713846
rect 42159 713845 42225 713846
rect 674127 713612 674193 713615
rect 674127 713610 674814 713612
rect 674127 713554 674132 713610
rect 674188 713554 674814 713610
rect 674127 713552 674814 713554
rect 674127 713549 674193 713552
rect 674754 713508 674814 713552
rect 675898 713254 675904 713318
rect 675968 713254 675974 713318
rect 675906 712990 675966 713254
rect 676282 712662 676288 712726
rect 676352 712662 676358 712726
rect 676290 712398 676350 712662
rect 676474 712218 676480 712282
rect 676544 712218 676550 712282
rect 676482 711880 676542 712218
rect 41914 711626 41920 711690
rect 41984 711688 41990 711690
rect 42063 711688 42129 711691
rect 41984 711686 42129 711688
rect 41984 711630 42068 711686
rect 42124 711630 42129 711686
rect 41984 711628 42129 711630
rect 41984 711626 41990 711628
rect 42063 711625 42129 711628
rect 42298 711626 42304 711690
rect 42368 711688 42374 711690
rect 43023 711688 43089 711691
rect 42368 711686 43089 711688
rect 42368 711630 43028 711686
rect 43084 711630 43089 711686
rect 42368 711628 43089 711630
rect 42368 711626 42374 711628
rect 43023 711625 43089 711628
rect 677242 711626 677248 711690
rect 677312 711626 677318 711690
rect 42735 711540 42801 711543
rect 42735 711538 43134 711540
rect 42735 711482 42740 711538
rect 42796 711482 43134 711538
rect 42735 711480 43134 711482
rect 42735 711477 42801 711480
rect 43074 711392 43134 711480
rect 43215 711392 43281 711395
rect 43074 711390 43281 711392
rect 43074 711334 43220 711390
rect 43276 711334 43281 711390
rect 677250 711362 677310 711626
rect 43074 711332 43281 711334
rect 43215 711329 43281 711332
rect 41722 711182 41728 711246
rect 41792 711244 41798 711246
rect 42447 711244 42513 711247
rect 41792 711242 42513 711244
rect 41792 711186 42452 711242
rect 42508 711186 42513 711242
rect 41792 711184 42513 711186
rect 41792 711182 41798 711184
rect 42447 711181 42513 711184
rect 41722 711034 41728 711098
rect 41792 711096 41798 711098
rect 42490 711096 42496 711098
rect 41792 711036 42496 711096
rect 41792 711034 41798 711036
rect 42490 711034 42496 711036
rect 42560 711034 42566 711098
rect 675514 711034 675520 711098
rect 675584 711034 675590 711098
rect 42298 710886 42304 710950
rect 42368 710948 42374 710950
rect 43023 710948 43089 710951
rect 42368 710946 43089 710948
rect 42368 710890 43028 710946
rect 43084 710890 43089 710946
rect 42368 710888 43089 710890
rect 42368 710886 42374 710888
rect 43023 710885 43089 710888
rect 675522 710770 675582 711034
rect 675706 710590 675712 710654
rect 675776 710590 675782 710654
rect 675714 710252 675774 710590
rect 42159 709914 42225 709915
rect 42106 709912 42112 709914
rect 42068 709852 42112 709912
rect 42176 709910 42225 709914
rect 42220 709854 42225 709910
rect 42106 709850 42112 709852
rect 42176 709850 42225 709854
rect 42159 709849 42225 709850
rect 674415 709764 674481 709767
rect 674415 709762 674784 709764
rect 674415 709706 674420 709762
rect 674476 709706 674784 709762
rect 674415 709704 674784 709706
rect 674415 709701 674481 709704
rect 674415 709172 674481 709175
rect 674415 709170 674784 709172
rect 674415 709114 674420 709170
rect 674476 709114 674784 709170
rect 674415 709112 674784 709114
rect 674415 709109 674481 709112
rect 674415 708654 674481 708657
rect 674415 708652 674784 708654
rect 674415 708596 674420 708652
rect 674476 708596 674784 708652
rect 674415 708594 674784 708596
rect 674415 708591 674481 708594
rect 673263 708136 673329 708139
rect 673263 708134 674784 708136
rect 673263 708078 673268 708134
rect 673324 708078 674784 708134
rect 673263 708076 674784 708078
rect 673263 708073 673329 708076
rect 649839 707544 649905 707547
rect 649794 707542 649905 707544
rect 649794 707486 649844 707542
rect 649900 707486 649905 707542
rect 649794 707481 649905 707486
rect 673071 707544 673137 707547
rect 673071 707542 674784 707544
rect 673071 707486 673076 707542
rect 673132 707486 674784 707542
rect 673071 707484 674784 707486
rect 673071 707481 673137 707484
rect 41530 707334 41536 707398
rect 41600 707396 41606 707398
rect 41775 707396 41841 707399
rect 41600 707394 41841 707396
rect 41600 707338 41780 707394
rect 41836 707338 41841 707394
rect 41600 707336 41841 707338
rect 41600 707334 41606 707336
rect 41775 707333 41841 707336
rect 40762 707186 40768 707250
rect 40832 707248 40838 707250
rect 42447 707248 42513 707251
rect 40832 707246 42513 707248
rect 40832 707190 42452 707246
rect 42508 707190 42513 707246
rect 40832 707188 42513 707190
rect 40832 707186 40838 707188
rect 42447 707185 42513 707188
rect 42682 706890 42688 706954
rect 42752 706952 42758 706954
rect 43258 706952 43268 706954
rect 42752 706892 43268 706952
rect 42752 706890 42758 706892
rect 43258 706890 43268 706892
rect 43332 706890 43338 706954
rect 649794 706922 649854 707481
rect 673167 707100 673233 707103
rect 673167 707098 674814 707100
rect 673167 707042 673172 707098
rect 673228 707042 674814 707098
rect 673167 707040 674814 707042
rect 673167 707037 673233 707040
rect 674754 706996 674814 707040
rect 42874 706446 42880 706510
rect 42944 706508 42950 706510
rect 43119 706508 43185 706511
rect 42944 706506 43185 706508
rect 42944 706450 43124 706506
rect 43180 706450 43185 706506
rect 42944 706448 43185 706450
rect 42944 706446 42950 706448
rect 43119 706445 43185 706448
rect 677058 706215 677118 706478
rect 677007 706210 677118 706215
rect 677007 706154 677012 706210
rect 677068 706154 677118 706210
rect 677007 706152 677118 706154
rect 677007 706149 677073 706152
rect 676866 705623 676926 705886
rect 676815 705618 676926 705623
rect 676815 705562 676820 705618
rect 676876 705562 676926 705618
rect 676815 705560 676926 705562
rect 677007 705620 677073 705623
rect 677007 705618 677118 705620
rect 677007 705562 677012 705618
rect 677068 705562 677118 705618
rect 676815 705557 676881 705560
rect 677007 705557 677118 705562
rect 677058 705368 677118 705557
rect 41338 705114 41344 705178
rect 41408 705176 41414 705178
rect 42351 705176 42417 705179
rect 41408 705174 42417 705176
rect 41408 705118 42356 705174
rect 42412 705118 42417 705174
rect 41408 705116 42417 705118
rect 41408 705114 41414 705116
rect 42351 705113 42417 705116
rect 676815 705176 676881 705179
rect 676815 705174 676926 705176
rect 676815 705118 676820 705174
rect 676876 705118 676926 705174
rect 676815 705113 676926 705118
rect 676866 704850 676926 705113
rect 42159 704584 42225 704587
rect 42490 704584 42496 704586
rect 42159 704582 42496 704584
rect 42159 704526 42164 704582
rect 42220 704526 42496 704582
rect 42159 704524 42496 704526
rect 42159 704521 42225 704524
rect 42490 704522 42496 704524
rect 42560 704522 42566 704586
rect 41775 704142 41841 704143
rect 41722 704078 41728 704142
rect 41792 704140 41841 704142
rect 41792 704138 41884 704140
rect 41836 704082 41884 704138
rect 41792 704080 41884 704082
rect 41792 704078 41841 704080
rect 41775 704077 41841 704078
rect 40954 703338 40960 703402
rect 41024 703400 41030 703402
rect 42447 703400 42513 703403
rect 41024 703398 42513 703400
rect 41024 703342 42452 703398
rect 42508 703342 42513 703398
rect 41024 703340 42513 703342
rect 41024 703338 41030 703340
rect 42447 703337 42513 703340
rect 59535 702364 59601 702367
rect 59535 702362 64416 702364
rect 59535 702306 59540 702362
rect 59596 702306 64416 702362
rect 59535 702304 64416 702306
rect 59535 702301 59601 702304
rect 42063 700588 42129 700591
rect 43066 700588 43072 700590
rect 42063 700586 43072 700588
rect 42063 700530 42068 700586
rect 42124 700530 43072 700586
rect 42063 700528 43072 700530
rect 42063 700525 42129 700528
rect 43066 700526 43072 700528
rect 43136 700526 43142 700590
rect 675471 697926 675537 697927
rect 675471 697922 675520 697926
rect 675584 697924 675590 697926
rect 675471 697866 675476 697922
rect 675471 697862 675520 697866
rect 675584 697864 675628 697924
rect 675584 697862 675590 697864
rect 675471 697861 675537 697862
rect 675759 697332 675825 697335
rect 676666 697332 676672 697334
rect 675759 697330 676672 697332
rect 675759 697274 675764 697330
rect 675820 697274 676672 697330
rect 675759 697272 676672 697274
rect 675759 697269 675825 697272
rect 676666 697270 676672 697272
rect 676736 697270 676742 697334
rect 6412 696342 8706 697142
rect 9506 697141 50926 697142
rect 9506 696343 50127 697141
rect 50925 696343 50931 697141
rect 675322 696974 675328 697038
rect 675392 697036 675398 697038
rect 676282 697036 676288 697038
rect 675392 696976 676288 697036
rect 675392 696974 675398 696976
rect 676282 696974 676288 696976
rect 676352 696974 676358 697038
rect 675375 696890 675441 696891
rect 675322 696888 675328 696890
rect 675284 696828 675328 696888
rect 675392 696886 675441 696890
rect 675436 696830 675441 696886
rect 675322 696826 675328 696828
rect 675392 696826 675441 696830
rect 675375 696825 675441 696826
rect 9506 696342 50926 696343
rect 6252 695068 16332 695868
rect 17132 695867 52718 695868
rect 17132 695069 51919 695867
rect 52717 695069 52723 695867
rect 654447 695260 654513 695263
rect 650208 695258 654513 695260
rect 650208 695202 654452 695258
rect 654508 695202 654513 695258
rect 650208 695200 654513 695202
rect 654447 695197 654513 695200
rect 17132 695068 52718 695069
rect 675663 694818 675729 694819
rect 675663 694814 675712 694818
rect 675776 694816 675782 694818
rect 675663 694758 675668 694814
rect 675663 694754 675712 694758
rect 675776 694756 675820 694816
rect 675776 694754 675782 694756
rect 6160 693954 7212 694754
rect 8012 694753 54502 694754
rect 675663 694753 675729 694754
rect 8012 693955 53703 694753
rect 54501 693955 54507 694753
rect 674554 694310 674560 694374
rect 674624 694372 674630 694374
rect 675471 694372 675537 694375
rect 674624 694370 675537 694372
rect 674624 694314 675476 694370
rect 675532 694314 675537 694370
rect 674624 694312 675537 694314
rect 674624 694310 674630 694312
rect 675471 694309 675537 694312
rect 8012 693954 54502 693955
rect 6066 692284 17798 693084
rect 18598 693083 56068 693084
rect 18598 692285 55269 693083
rect 56067 692285 56073 693083
rect 18598 692284 56068 692285
rect 675759 692004 675825 692007
rect 676474 692004 676480 692006
rect 675759 692002 676480 692004
rect 675759 691946 675764 692002
rect 675820 691946 676480 692002
rect 675759 691944 676480 691946
rect 675759 691941 675825 691944
rect 676474 691942 676480 691944
rect 676544 691942 676550 692006
rect 43215 689488 43281 689491
rect 42528 689486 43281 689488
rect 42528 689430 43220 689486
rect 43276 689430 43281 689486
rect 42528 689428 43281 689430
rect 43215 689425 43281 689428
rect 675759 689192 675825 689195
rect 675898 689192 675904 689194
rect 675759 689190 675904 689192
rect 675759 689134 675764 689190
rect 675820 689134 675904 689190
rect 675759 689132 675904 689134
rect 675759 689129 675825 689132
rect 675898 689130 675904 689132
rect 675968 689130 675974 689194
rect 43119 689044 43185 689047
rect 42498 689042 43185 689044
rect 42498 688986 43124 689042
rect 43180 688986 43185 689042
rect 42498 688984 43185 688986
rect 42498 688866 42558 688984
rect 43119 688981 43185 688984
rect 42831 688452 42897 688455
rect 42528 688450 42897 688452
rect 42528 688394 42836 688450
rect 42892 688394 42897 688450
rect 42528 688392 42897 688394
rect 42831 688389 42897 688392
rect 675087 688304 675153 688307
rect 676090 688304 676096 688306
rect 675087 688302 676096 688304
rect 675087 688246 675092 688302
rect 675148 688246 676096 688302
rect 675087 688244 676096 688246
rect 675087 688241 675153 688244
rect 676090 688242 676096 688244
rect 676160 688242 676166 688306
rect 59535 688008 59601 688011
rect 59535 688006 64416 688008
rect 59535 687950 59540 688006
rect 59596 687950 64416 688006
rect 59535 687948 64416 687950
rect 59535 687945 59601 687948
rect 43407 687860 43473 687863
rect 42528 687858 43473 687860
rect 42528 687802 43412 687858
rect 43468 687802 43473 687858
rect 42528 687800 43473 687802
rect 43407 687797 43473 687800
rect 43503 687712 43569 687715
rect 42498 687710 43569 687712
rect 42498 687654 43508 687710
rect 43564 687654 43569 687710
rect 42498 687652 43569 687654
rect 42498 687238 42558 687652
rect 43503 687649 43569 687652
rect 40570 686910 40576 686974
rect 40640 686910 40646 686974
rect 40578 686824 40638 686910
rect 40578 686794 42144 686824
rect 40608 686764 42174 686794
rect 42114 686530 42174 686764
rect 42106 686466 42112 686530
rect 42176 686466 42182 686530
rect 40386 685938 40446 686202
rect 40378 685874 40384 685938
rect 40448 685936 40454 685938
rect 41146 685936 41152 685938
rect 40448 685876 41152 685936
rect 40448 685874 40454 685876
rect 41146 685874 41152 685876
rect 41216 685874 41222 685938
rect 42114 685495 42174 685610
rect 42063 685490 42174 685495
rect 42063 685434 42068 685490
rect 42124 685434 42174 685490
rect 42063 685432 42174 685434
rect 42063 685429 42129 685432
rect 41922 684903 41982 685166
rect 41871 684898 41982 684903
rect 41871 684842 41876 684898
rect 41932 684842 41982 684898
rect 41871 684840 41982 684842
rect 41871 684837 41937 684840
rect 40578 684310 40638 684574
rect 40570 684246 40576 684310
rect 40640 684246 40646 684310
rect 42498 683716 42558 683982
rect 43695 683716 43761 683719
rect 42498 683714 43761 683716
rect 42498 683658 43700 683714
rect 43756 683658 43761 683714
rect 42498 683656 43761 683658
rect 43695 683653 43761 683656
rect 655119 683568 655185 683571
rect 650208 683566 655185 683568
rect 42498 683124 42558 683538
rect 650208 683510 655124 683566
rect 655180 683510 655185 683566
rect 650208 683508 655185 683510
rect 655119 683505 655185 683508
rect 43066 683124 43072 683126
rect 42498 683064 43072 683124
rect 43066 683062 43072 683064
rect 43136 683062 43142 683126
rect 42306 682683 42366 682946
rect 42306 682678 42417 682683
rect 42306 682622 42356 682678
rect 42412 682622 42417 682678
rect 42306 682620 42417 682622
rect 42351 682617 42417 682620
rect 40770 682090 40830 682354
rect 671682 682316 699121 682317
rect 40762 682026 40768 682090
rect 40832 682026 40838 682090
rect 40962 681499 41022 681910
rect 40962 681494 41073 681499
rect 40962 681438 41012 681494
rect 41068 681438 41073 681494
rect 40962 681436 41073 681438
rect 41007 681433 41073 681436
rect 43215 681348 43281 681351
rect 42528 681346 43281 681348
rect 42528 681290 43220 681346
rect 43276 681290 43281 681346
rect 42528 681288 43281 681290
rect 43215 681285 43281 681288
rect 671677 681224 671683 682316
rect 672775 681224 699121 682316
rect 671682 681223 699121 681224
rect 700215 681223 711345 682317
rect 666066 680803 709418 680804
rect 42114 680463 42174 680726
rect 42114 680458 42225 680463
rect 42114 680402 42164 680458
rect 42220 680402 42225 680458
rect 42114 680400 42225 680402
rect 42159 680397 42225 680400
rect 41967 679868 42033 679871
rect 41922 679866 42033 679868
rect 41922 679810 41972 679866
rect 42028 679810 42033 679866
rect 41922 679805 42033 679810
rect 42498 679868 42558 680208
rect 43119 679868 43185 679871
rect 42498 679866 43185 679868
rect 42498 679810 43124 679866
rect 43180 679810 43185 679866
rect 42498 679808 43185 679810
rect 43119 679805 43185 679808
rect 41922 679690 41982 679805
rect 666061 679621 666067 680803
rect 667249 679621 709418 680803
rect 666066 679620 709418 679621
rect 710602 679620 711056 680804
rect 41730 678835 41790 679098
rect 662178 678967 700498 678968
rect 41730 678830 41841 678835
rect 41730 678774 41780 678830
rect 41836 678774 41841 678830
rect 41730 678772 41841 678774
rect 41775 678769 41841 678772
rect 41538 678242 41598 678580
rect 41530 678178 41536 678242
rect 41600 678178 41606 678242
rect 42498 677796 42558 678062
rect 42498 677736 42750 677796
rect 662173 677785 662179 678967
rect 663361 677785 700498 678967
rect 662178 677784 700498 677785
rect 701682 677784 711334 678968
rect 35202 677207 35262 677470
rect 42690 677352 42750 677736
rect 35151 677202 35262 677207
rect 35151 677146 35156 677202
rect 35212 677146 35262 677202
rect 35151 677144 35262 677146
rect 42498 677292 42750 677352
rect 35151 677141 35217 677144
rect 42498 676908 42558 677292
rect 659368 677243 708330 677244
rect 53583 676908 53649 676911
rect 42498 676906 53649 676908
rect 42498 676850 53588 676906
rect 53644 676850 53649 676906
rect 42498 676848 53649 676850
rect 53583 676845 53649 676848
rect 35151 676760 35217 676763
rect 35151 676758 35262 676760
rect 35151 676702 35156 676758
rect 35212 676702 35262 676758
rect 35151 676697 35262 676702
rect 35202 676434 35262 676697
rect 659363 676061 659369 677243
rect 660551 676061 708330 677243
rect 659368 676060 708330 676061
rect 709514 676060 711000 677244
rect 41679 675578 41745 675579
rect 41679 675574 41728 675578
rect 41792 675576 41798 675578
rect 41679 675518 41684 675574
rect 41679 675514 41728 675518
rect 41792 675516 41836 675576
rect 41792 675514 41798 675516
rect 41679 675513 41745 675514
rect 59535 673652 59601 673655
rect 59535 673650 64416 673652
rect 59535 673594 59540 673650
rect 59596 673594 64416 673650
rect 59535 673592 64416 673594
rect 59535 673589 59601 673592
rect 674415 672690 674481 672693
rect 674415 672688 674784 672690
rect 674415 672632 674420 672688
rect 674476 672632 674784 672688
rect 674415 672630 674784 672632
rect 674415 672627 674481 672630
rect 674415 672172 674481 672175
rect 674415 672170 674784 672172
rect 674415 672114 674420 672170
rect 674476 672114 674784 672170
rect 674415 672112 674784 672114
rect 674415 672109 674481 672112
rect 654447 671728 654513 671731
rect 650208 671726 654513 671728
rect 650208 671670 654452 671726
rect 654508 671670 654513 671726
rect 650208 671668 654513 671670
rect 654447 671665 654513 671668
rect 674415 671580 674481 671583
rect 674415 671578 674784 671580
rect 674415 671522 674420 671578
rect 674476 671522 674784 671578
rect 674415 671520 674784 671522
rect 674415 671517 674481 671520
rect 673743 671136 673809 671139
rect 673743 671134 674814 671136
rect 673743 671078 673748 671134
rect 673804 671078 674814 671134
rect 673743 671076 674814 671078
rect 673743 671073 673809 671076
rect 674754 671032 674814 671076
rect 41007 670988 41073 670991
rect 41338 670988 41344 670990
rect 41007 670986 41344 670988
rect 41007 670930 41012 670986
rect 41068 670930 41344 670986
rect 41007 670928 41344 670930
rect 41007 670925 41073 670928
rect 41338 670926 41344 670928
rect 41408 670926 41414 670990
rect 41679 670986 41745 670991
rect 41679 670930 41684 670986
rect 41740 670930 41745 670986
rect 41679 670925 41745 670930
rect 42298 670926 42304 670990
rect 42368 670988 42374 670990
rect 42927 670988 42993 670991
rect 42368 670986 42993 670988
rect 42368 670930 42932 670986
rect 42988 670930 42993 670986
rect 42368 670928 42993 670930
rect 42368 670926 42374 670928
rect 42927 670925 42993 670928
rect 41682 670544 41742 670925
rect 42063 670692 42129 670695
rect 43023 670694 43089 670695
rect 42490 670692 42496 670694
rect 42063 670690 42496 670692
rect 42063 670634 42068 670690
rect 42124 670634 42496 670690
rect 42063 670632 42496 670634
rect 42063 670629 42129 670632
rect 42490 670630 42496 670632
rect 42560 670630 42566 670694
rect 43023 670692 43072 670694
rect 42980 670690 43072 670692
rect 42980 670634 43028 670690
rect 42980 670632 43072 670634
rect 43023 670630 43072 670632
rect 43136 670630 43142 670694
rect 43023 670629 43089 670630
rect 41914 670544 41920 670546
rect 41682 670484 41920 670544
rect 41914 670482 41920 670484
rect 41984 670482 41990 670546
rect 677250 670250 677310 670514
rect 677242 670186 677248 670250
rect 677312 670186 677318 670250
rect 677434 670186 677440 670250
rect 677504 670186 677510 670250
rect 677442 669922 677502 670186
rect 677050 669594 677056 669658
rect 677120 669594 677126 669658
rect 677058 669404 677118 669594
rect 674362 668854 674368 668918
rect 674432 668916 674438 668918
rect 674432 668856 674784 668916
rect 674432 668854 674438 668856
rect 674607 668620 674673 668623
rect 674607 668618 674814 668620
rect 674607 668562 674612 668618
rect 674668 668562 674814 668618
rect 674607 668560 674814 668562
rect 674607 668557 674673 668560
rect 674754 668294 674814 668560
rect 674170 667744 674176 667808
rect 674240 667806 674246 667808
rect 674240 667746 674784 667806
rect 674240 667744 674246 667746
rect 675130 667522 675136 667586
rect 675200 667522 675206 667586
rect 675138 667258 675198 667522
rect 674223 666696 674289 666699
rect 674223 666694 674784 666696
rect 674223 666638 674228 666694
rect 674284 666638 674784 666694
rect 674223 666636 674784 666638
rect 674223 666633 674289 666636
rect 674511 666400 674577 666403
rect 674511 666398 674814 666400
rect 674511 666342 674516 666398
rect 674572 666342 674814 666398
rect 674511 666340 674814 666342
rect 674511 666337 674577 666340
rect 674754 666148 674814 666340
rect 673978 665598 673984 665662
rect 674048 665660 674054 665662
rect 674048 665600 674784 665660
rect 674048 665598 674054 665600
rect 41530 665302 41536 665366
rect 41600 665364 41606 665366
rect 42159 665364 42225 665367
rect 41600 665362 42225 665364
rect 41600 665306 42164 665362
rect 42220 665306 42225 665362
rect 41600 665304 42225 665306
rect 41600 665302 41606 665304
rect 42159 665301 42225 665304
rect 674938 665302 674944 665366
rect 675008 665302 675014 665366
rect 674946 665038 675006 665302
rect 674746 664858 674752 664922
rect 674816 664858 674822 664922
rect 42159 664772 42225 664775
rect 42298 664772 42304 664774
rect 42159 664770 42304 664772
rect 42159 664714 42164 664770
rect 42220 664714 42304 664770
rect 42159 664712 42304 664714
rect 42159 664709 42225 664712
rect 42298 664710 42304 664712
rect 42368 664710 42374 664774
rect 674754 664520 674814 664858
rect 674895 664180 674961 664183
rect 674895 664178 675006 664180
rect 674895 664122 674900 664178
rect 674956 664122 675006 664178
rect 674895 664117 675006 664122
rect 41338 663970 41344 664034
rect 41408 664032 41414 664034
rect 42639 664032 42705 664035
rect 41408 664030 42705 664032
rect 41408 663974 42644 664030
rect 42700 663974 42705 664030
rect 674946 664002 675006 664117
rect 41408 663972 42705 663974
rect 41408 663970 41414 663972
rect 42639 663969 42705 663972
rect 676282 663674 676288 663738
rect 676352 663674 676358 663738
rect 676290 663410 676350 663674
rect 42351 662848 42417 662851
rect 42490 662848 42496 662850
rect 42351 662846 42496 662848
rect 42351 662790 42356 662846
rect 42412 662790 42496 662846
rect 42351 662788 42496 662790
rect 42351 662785 42417 662788
rect 42490 662786 42496 662788
rect 42560 662786 42566 662850
rect 673839 662848 673905 662851
rect 673839 662846 674784 662848
rect 673839 662790 673844 662846
rect 673900 662790 674784 662846
rect 673839 662788 674784 662790
rect 673839 662785 673905 662788
rect 40762 662342 40768 662406
rect 40832 662404 40838 662406
rect 43023 662404 43089 662407
rect 40832 662402 43089 662404
rect 40832 662346 43028 662402
rect 43084 662346 43089 662402
rect 40832 662344 43089 662346
rect 40832 662342 40838 662344
rect 43023 662341 43089 662344
rect 673359 662404 673425 662407
rect 673359 662402 674784 662404
rect 673359 662346 673364 662402
rect 673420 662346 674784 662402
rect 673359 662344 674784 662346
rect 673359 662341 673425 662344
rect 41722 662194 41728 662258
rect 41792 662256 41798 662258
rect 42063 662256 42129 662259
rect 42682 662256 42688 662258
rect 41792 662254 42688 662256
rect 41792 662198 42068 662254
rect 42124 662198 42688 662254
rect 41792 662196 42688 662198
rect 41792 662194 41798 662196
rect 42063 662193 42129 662196
rect 42682 662194 42688 662196
rect 42752 662194 42758 662258
rect 673839 661812 673905 661815
rect 673839 661810 674784 661812
rect 673839 661754 673844 661810
rect 673900 661754 674784 661810
rect 673839 661752 674784 661754
rect 673839 661749 673905 661752
rect 41871 661074 41937 661075
rect 41871 661072 41920 661074
rect 41828 661070 41920 661072
rect 41828 661014 41876 661070
rect 41828 661012 41920 661014
rect 41871 661010 41920 661012
rect 41984 661010 41990 661074
rect 41871 661009 41937 661010
rect 674946 660927 675006 661190
rect 40570 660862 40576 660926
rect 40640 660924 40646 660926
rect 43119 660924 43185 660927
rect 40640 660922 43185 660924
rect 40640 660866 43124 660922
rect 43180 660866 43185 660922
rect 40640 660864 43185 660866
rect 40640 660862 40646 660864
rect 43119 660861 43185 660864
rect 674895 660922 675006 660927
rect 674895 660866 674900 660922
rect 674956 660866 675006 660922
rect 674895 660864 675006 660866
rect 674895 660861 674961 660864
rect 650319 660628 650385 660631
rect 650178 660626 650385 660628
rect 650178 660570 650324 660626
rect 650380 660570 650385 660626
rect 650178 660568 650385 660570
rect 650178 660006 650238 660568
rect 650319 660565 650385 660568
rect 675138 660483 675198 660746
rect 674895 660480 674961 660483
rect 674895 660478 675006 660480
rect 674895 660422 674900 660478
rect 674956 660422 675006 660478
rect 674895 660417 675006 660422
rect 675087 660478 675198 660483
rect 675087 660422 675092 660478
rect 675148 660422 675198 660478
rect 675087 660420 675198 660422
rect 675087 660417 675153 660420
rect 674946 660154 675006 660417
rect 675087 659888 675153 659891
rect 675087 659886 675198 659888
rect 675087 659830 675092 659886
rect 675148 659830 675198 659886
rect 675087 659825 675198 659830
rect 675138 659562 675198 659825
rect 59535 659296 59601 659299
rect 59535 659294 64416 659296
rect 59535 659238 59540 659294
rect 59596 659238 64416 659294
rect 59535 659236 64416 659238
rect 59535 659233 59601 659236
rect 6860 653016 8566 653816
rect 9366 653815 50926 653816
rect 9366 653017 50127 653815
rect 50925 653017 50931 653815
rect 675087 653672 675153 653675
rect 676474 653672 676480 653674
rect 675087 653670 676480 653672
rect 675087 653614 675092 653670
rect 675148 653614 676480 653670
rect 675087 653612 676480 653614
rect 675087 653609 675153 653612
rect 676474 653610 676480 653612
rect 676544 653610 676550 653674
rect 9366 653016 50926 653017
rect 6674 651820 16290 652620
rect 17090 652619 52718 652620
rect 17090 651821 51919 652619
rect 52717 651821 52723 652619
rect 674746 652574 674752 652638
rect 674816 652636 674822 652638
rect 675375 652636 675441 652639
rect 674816 652634 675441 652636
rect 674816 652578 675380 652634
rect 675436 652578 675441 652634
rect 674816 652576 675441 652578
rect 674816 652574 674822 652576
rect 675375 652573 675441 652576
rect 674170 652130 674176 652194
rect 674240 652192 674246 652194
rect 675471 652192 675537 652195
rect 674240 652190 675537 652192
rect 674240 652134 675476 652190
rect 675532 652134 675537 652190
rect 674240 652132 675537 652134
rect 674240 652130 674246 652132
rect 675471 652129 675537 652132
rect 17090 651820 52718 651821
rect 6674 650716 7184 651516
rect 7984 651515 54502 651516
rect 7984 650717 53703 651515
rect 54501 650717 54507 651515
rect 675130 651390 675136 651454
rect 675200 651452 675206 651454
rect 675471 651452 675537 651455
rect 675200 651450 675537 651452
rect 675200 651394 675476 651450
rect 675532 651394 675537 651450
rect 675200 651392 675537 651394
rect 675200 651390 675206 651392
rect 675471 651389 675537 651392
rect 7984 650716 54502 650717
rect 6122 649150 17672 649950
rect 18472 649949 56068 649950
rect 18472 649151 55269 649949
rect 56067 649151 56073 649949
rect 673978 649762 673984 649826
rect 674048 649824 674054 649826
rect 674746 649824 674752 649826
rect 674048 649764 674752 649824
rect 674048 649762 674054 649764
rect 674746 649762 674752 649764
rect 674816 649762 674822 649826
rect 674746 649614 674752 649678
rect 674816 649676 674822 649678
rect 675375 649676 675441 649679
rect 674816 649674 675441 649676
rect 674816 649618 675380 649674
rect 675436 649618 675441 649674
rect 674816 649616 675441 649618
rect 674816 649614 674822 649616
rect 675375 649613 675441 649616
rect 18472 649150 56068 649151
rect 674362 648874 674368 648938
rect 674432 648936 674438 648938
rect 675471 648936 675537 648939
rect 674432 648934 675537 648936
rect 674432 648878 675476 648934
rect 675532 648878 675537 648934
rect 674432 648876 675537 648878
rect 674432 648874 674438 648876
rect 675471 648873 675537 648876
rect 654255 648344 654321 648347
rect 650208 648342 654321 648344
rect 650208 648286 654260 648342
rect 654316 648286 654321 648342
rect 650208 648284 654321 648286
rect 654255 648281 654321 648284
rect 42106 647098 42112 647162
rect 42176 647160 42182 647162
rect 43791 647160 43857 647163
rect 42176 647158 43857 647160
rect 42176 647102 43796 647158
rect 43852 647102 43857 647158
rect 42176 647100 43857 647102
rect 42176 647098 42182 647100
rect 43791 647097 43857 647100
rect 40378 646950 40384 647014
rect 40448 647012 40454 647014
rect 43599 647012 43665 647015
rect 40448 647010 43665 647012
rect 40448 646954 43604 647010
rect 43660 646954 43665 647010
rect 40448 646952 43665 646954
rect 40448 646950 40454 646952
rect 43599 646949 43665 646952
rect 42927 646272 42993 646275
rect 42528 646270 42993 646272
rect 42528 646214 42932 646270
rect 42988 646214 42993 646270
rect 42528 646212 42993 646214
rect 42927 646209 42993 646212
rect 42306 645535 42366 645724
rect 42306 645530 42417 645535
rect 42306 645474 42356 645530
rect 42412 645474 42417 645530
rect 42306 645472 42417 645474
rect 42351 645469 42417 645472
rect 675759 645384 675825 645387
rect 676282 645384 676288 645386
rect 675759 645382 676288 645384
rect 675759 645326 675764 645382
rect 675820 645326 676288 645382
rect 675759 645324 676288 645326
rect 675759 645321 675825 645324
rect 676282 645322 676288 645324
rect 676352 645322 676358 645386
rect 43215 645236 43281 645239
rect 42528 645234 43281 645236
rect 42528 645178 43220 645234
rect 43276 645178 43281 645234
rect 42528 645176 43281 645178
rect 43215 645173 43281 645176
rect 59535 644940 59601 644943
rect 59535 644938 64416 644940
rect 59535 644882 59540 644938
rect 59596 644882 64416 644938
rect 59535 644880 64416 644882
rect 59535 644877 59601 644880
rect 43983 644644 44049 644647
rect 42528 644642 44049 644644
rect 42528 644586 43988 644642
rect 44044 644586 44049 644642
rect 42528 644584 44049 644586
rect 43983 644581 44049 644584
rect 43311 644496 43377 644499
rect 42498 644494 43377 644496
rect 42498 644438 43316 644494
rect 43372 644438 43377 644494
rect 42498 644436 43377 644438
rect 42498 644096 42558 644436
rect 43311 644433 43377 644436
rect 43791 643608 43857 643611
rect 42528 643606 43857 643608
rect 42528 643550 43796 643606
rect 43852 643550 43857 643606
rect 42528 643548 43857 643550
rect 43791 643545 43857 643548
rect 43599 643016 43665 643019
rect 42528 643014 43665 643016
rect 42528 642958 43604 643014
rect 43660 642958 43665 643014
rect 42528 642956 43665 642958
rect 43599 642953 43665 642956
rect 42498 642128 42558 642468
rect 43503 642128 43569 642131
rect 42498 642126 43569 642128
rect 42498 642070 43508 642126
rect 43564 642070 43569 642126
rect 42498 642068 43569 642070
rect 43503 642065 43569 642068
rect 41730 641687 41790 641950
rect 41730 641682 41841 641687
rect 41730 641626 41780 641682
rect 41836 641626 41841 641682
rect 41730 641624 41841 641626
rect 41775 641621 41841 641624
rect 40962 641094 41022 641358
rect 40954 641030 40960 641094
rect 41024 641030 41030 641094
rect 40962 640503 41022 640840
rect 40962 640498 41073 640503
rect 40962 640442 41012 640498
rect 41068 640442 41073 640498
rect 40962 640440 41073 640442
rect 41007 640437 41073 640440
rect 41538 640059 41598 640322
rect 673978 640290 673984 640354
rect 674048 640352 674054 640354
rect 675375 640352 675441 640355
rect 674048 640350 675441 640352
rect 674048 640294 675380 640350
rect 675436 640294 675441 640350
rect 674048 640292 675441 640294
rect 674048 640290 674054 640292
rect 675375 640289 675441 640292
rect 41538 640054 41649 640059
rect 41538 639998 41588 640054
rect 41644 639998 41649 640054
rect 41538 639996 41649 639998
rect 41583 639993 41649 639996
rect 41922 639467 41982 639730
rect 41871 639462 41982 639467
rect 41871 639406 41876 639462
rect 41932 639406 41982 639462
rect 41871 639404 41982 639406
rect 41871 639401 41937 639404
rect 40578 638874 40638 639138
rect 40570 638810 40576 638874
rect 40640 638810 40646 638874
rect 41538 638431 41598 638694
rect 675759 638576 675825 638579
rect 676474 638576 676480 638578
rect 675759 638574 676480 638576
rect 675759 638518 675764 638574
rect 675820 638518 676480 638574
rect 675759 638516 676480 638518
rect 675759 638513 675825 638516
rect 676474 638514 676480 638516
rect 676544 638514 676550 638578
rect 41487 638426 41598 638431
rect 41487 638370 41492 638426
rect 41548 638370 41598 638426
rect 41487 638368 41598 638370
rect 41487 638365 41553 638368
rect 41922 637839 41982 638102
rect 41922 637834 42033 637839
rect 41922 637778 41972 637834
rect 42028 637778 42033 637834
rect 41922 637776 42033 637778
rect 41967 637773 42033 637776
rect 42498 637244 42558 637510
rect 43215 637244 43281 637247
rect 42498 637242 43281 637244
rect 42498 637186 43220 637242
rect 43276 637186 43281 637242
rect 42498 637184 43281 637186
rect 43215 637181 43281 637184
rect 42114 636803 42174 637066
rect 671682 636972 699309 636973
rect 42114 636798 42225 636803
rect 42114 636742 42164 636798
rect 42220 636742 42225 636798
rect 42114 636740 42225 636742
rect 42159 636737 42225 636740
rect 655311 636652 655377 636655
rect 650208 636650 655377 636652
rect 650208 636594 655316 636650
rect 655372 636594 655377 636650
rect 650208 636592 655377 636594
rect 655311 636589 655377 636592
rect 42114 636211 42174 636474
rect 42063 636206 42174 636211
rect 42063 636150 42068 636206
rect 42124 636150 42174 636206
rect 42063 636148 42174 636150
rect 42063 636145 42129 636148
rect 42498 635616 42558 635882
rect 671677 635880 671683 636972
rect 672775 635880 699309 636972
rect 671682 635879 699309 635880
rect 700403 635879 712145 636973
rect 43311 635616 43377 635619
rect 42498 635614 43377 635616
rect 42498 635558 43316 635614
rect 43372 635558 43377 635614
rect 42498 635556 43377 635558
rect 43311 635553 43377 635556
rect 666066 635485 709374 635486
rect 42306 635175 42366 635438
rect 42306 635170 42417 635175
rect 42306 635114 42356 635170
rect 42412 635114 42417 635170
rect 42306 635112 42417 635114
rect 42351 635109 42417 635112
rect 42498 634580 42558 634846
rect 42498 634520 42750 634580
rect 35202 633991 35262 634254
rect 42690 634136 42750 634520
rect 666061 634303 666067 635485
rect 667249 634303 709374 635485
rect 666066 634302 709374 634303
rect 710558 634302 711918 635486
rect 35151 633986 35262 633991
rect 35151 633930 35156 633986
rect 35212 633930 35262 633986
rect 35151 633928 35262 633930
rect 42498 634076 42750 634136
rect 42498 633988 42558 634076
rect 56079 633988 56145 633991
rect 42498 633986 56145 633988
rect 42498 633930 56084 633986
rect 56140 633930 56145 633986
rect 42498 633928 56145 633930
rect 35151 633925 35217 633928
rect 42498 633810 42558 633928
rect 56079 633925 56145 633928
rect 662178 633625 700650 633626
rect 35151 633544 35217 633547
rect 35151 633542 35262 633544
rect 35151 633486 35156 633542
rect 35212 633486 35262 633542
rect 35151 633481 35262 633486
rect 35202 633218 35262 633481
rect 662173 632443 662179 633625
rect 663361 632443 700650 633625
rect 662178 632442 700650 632443
rect 701834 632442 711808 633626
rect 673786 630818 673792 630882
rect 673856 630880 673862 630882
rect 674938 630880 674944 630882
rect 673856 630820 674944 630880
rect 673856 630818 673862 630820
rect 674938 630818 674944 630820
rect 675008 630818 675014 630882
rect 674127 630732 674193 630735
rect 674362 630732 674368 630734
rect 674127 630730 674368 630732
rect 674127 630674 674132 630730
rect 674188 630674 674368 630730
rect 674127 630672 674368 630674
rect 674127 630669 674193 630672
rect 674362 630670 674368 630672
rect 674432 630670 674438 630734
rect 674991 630732 675057 630735
rect 675130 630732 675136 630734
rect 674991 630730 675136 630732
rect 674991 630674 674996 630730
rect 675052 630674 675136 630730
rect 674991 630672 675136 630674
rect 674991 630669 675057 630672
rect 675130 630670 675136 630672
rect 675200 630670 675206 630734
rect 59535 630584 59601 630587
rect 59535 630582 64416 630584
rect 59535 630526 59540 630582
rect 59596 630526 64416 630582
rect 59535 630524 64416 630526
rect 59535 630521 59601 630524
rect 659368 630015 708128 630016
rect 659363 628833 659369 630015
rect 660551 628833 708128 630015
rect 659368 628832 708128 628833
rect 709312 628832 711140 630016
rect 42159 628216 42225 628219
rect 42639 628216 42705 628219
rect 42159 628214 42705 628216
rect 42159 628158 42164 628214
rect 42220 628158 42644 628214
rect 42700 628158 42705 628214
rect 42159 628156 42705 628158
rect 42159 628153 42225 628156
rect 42639 628153 42705 628156
rect 41487 627774 41553 627775
rect 41487 627772 41536 627774
rect 41444 627770 41536 627772
rect 41444 627714 41492 627770
rect 41444 627712 41536 627714
rect 41487 627710 41536 627712
rect 41600 627710 41606 627774
rect 673839 627772 673905 627775
rect 673839 627770 674814 627772
rect 673839 627714 673844 627770
rect 673900 627714 674814 627770
rect 673839 627712 674814 627714
rect 41487 627709 41553 627710
rect 673839 627709 673905 627712
rect 674754 627668 674814 627712
rect 42063 627626 42129 627627
rect 42063 627624 42112 627626
rect 42020 627622 42112 627624
rect 42020 627566 42068 627622
rect 42020 627564 42112 627566
rect 42063 627562 42112 627564
rect 42176 627562 42182 627626
rect 42063 627561 42129 627562
rect 41967 627476 42033 627479
rect 42298 627476 42304 627478
rect 41967 627474 42304 627476
rect 41967 627418 41972 627474
rect 42028 627418 42304 627474
rect 41967 627416 42304 627418
rect 41967 627413 42033 627416
rect 42298 627414 42304 627416
rect 42368 627414 42374 627478
rect 674607 627328 674673 627331
rect 674607 627326 674814 627328
rect 674607 627270 674612 627326
rect 674668 627270 674814 627326
rect 674607 627268 674814 627270
rect 674607 627265 674673 627268
rect 674754 627150 674814 627268
rect 42351 627032 42417 627035
rect 42490 627032 42496 627034
rect 42351 627030 42496 627032
rect 42351 626974 42356 627030
rect 42412 626974 42496 627030
rect 42351 626972 42496 626974
rect 42351 626969 42417 626972
rect 42490 626970 42496 626972
rect 42560 626970 42566 627034
rect 674607 626884 674673 626887
rect 674607 626882 674814 626884
rect 674607 626826 674612 626882
rect 674668 626826 674814 626882
rect 674607 626824 674814 626826
rect 674607 626821 674673 626824
rect 674754 626558 674814 626824
rect 677242 626378 677248 626442
rect 677312 626378 677318 626442
rect 677250 626040 677310 626378
rect 674607 625256 674673 625259
rect 674754 625256 674814 625522
rect 674607 625254 674814 625256
rect 674607 625198 674612 625254
rect 674668 625198 674814 625254
rect 674607 625196 674814 625198
rect 674607 625193 674673 625196
rect 677434 625157 677440 625221
rect 677504 625157 677510 625221
rect 654063 624812 654129 624815
rect 650208 624810 654129 624812
rect 650208 624754 654068 624810
rect 654124 624754 654129 624810
rect 650208 624752 654129 624754
rect 654063 624749 654129 624752
rect 677050 624602 677056 624666
rect 677120 624602 677126 624666
rect 677199 624664 677265 624667
rect 677442 624664 677502 625157
rect 677199 624662 677502 624664
rect 677199 624606 677204 624662
rect 677260 624606 677502 624662
rect 677199 624604 677502 624606
rect 42447 624518 42513 624519
rect 42447 624516 42496 624518
rect 42404 624514 42496 624516
rect 42404 624458 42452 624514
rect 42404 624456 42496 624458
rect 42447 624454 42496 624456
rect 42560 624454 42566 624518
rect 42447 624453 42513 624454
rect 675322 624158 675328 624222
rect 675392 624158 675398 624222
rect 675330 623894 675390 624158
rect 676815 624072 676881 624075
rect 677058 624072 677118 624602
rect 677199 624601 677265 624604
rect 676815 624070 677118 624072
rect 676815 624014 676820 624070
rect 676876 624014 677118 624070
rect 676815 624012 677118 624014
rect 676815 624009 676881 624012
rect 674319 623332 674385 623335
rect 674319 623330 674784 623332
rect 674319 623274 674324 623330
rect 674380 623274 674784 623330
rect 674319 623272 674784 623274
rect 674319 623269 674385 623272
rect 675514 623122 675520 623186
rect 675584 623122 675590 623186
rect 675522 622784 675582 623122
rect 675706 622530 675712 622594
rect 675776 622530 675782 622594
rect 675714 622266 675774 622530
rect 42298 622086 42304 622150
rect 42368 622148 42374 622150
rect 42447 622148 42513 622151
rect 42368 622146 42513 622148
rect 42368 622090 42452 622146
rect 42508 622090 42513 622146
rect 42368 622088 42513 622090
rect 42368 622086 42374 622088
rect 42447 622085 42513 622088
rect 674895 622000 674961 622003
rect 674895 621998 675006 622000
rect 674895 621942 674900 621998
rect 674956 621942 675006 621998
rect 674895 621937 675006 621942
rect 674946 621674 675006 621937
rect 42106 621494 42112 621558
rect 42176 621556 42182 621558
rect 42639 621556 42705 621559
rect 42176 621554 42705 621556
rect 42176 621498 42644 621554
rect 42700 621498 42705 621554
rect 42176 621496 42705 621498
rect 42176 621494 42182 621496
rect 42639 621493 42705 621496
rect 674415 621112 674481 621115
rect 674415 621110 674784 621112
rect 674415 621054 674420 621110
rect 674476 621054 674784 621110
rect 674415 621052 674784 621054
rect 674415 621049 674481 621052
rect 676666 620902 676672 620966
rect 676736 620902 676742 620966
rect 674991 620818 675057 620819
rect 674938 620816 674944 620818
rect 674900 620756 674944 620816
rect 675008 620814 675057 620818
rect 675052 620758 675057 620814
rect 674938 620754 674944 620756
rect 675008 620754 675057 620758
rect 674991 620753 675057 620754
rect 676674 620638 676734 620902
rect 674554 620310 674560 620374
rect 674624 620372 674630 620374
rect 674624 620312 674814 620372
rect 674624 620310 674630 620312
rect 674754 620046 674814 620312
rect 674127 619928 674193 619931
rect 674554 619928 674560 619930
rect 674127 619926 674560 619928
rect 674127 619870 674132 619926
rect 674188 619870 674560 619926
rect 674127 619868 674560 619870
rect 674127 619865 674193 619868
rect 674554 619866 674560 619868
rect 674624 619866 674630 619930
rect 676090 619866 676096 619930
rect 676160 619866 676166 619930
rect 41530 619570 41536 619634
rect 41600 619632 41606 619634
rect 42351 619632 42417 619635
rect 41600 619630 42417 619632
rect 41600 619574 42356 619630
rect 42412 619574 42417 619630
rect 41600 619572 42417 619574
rect 41600 619570 41606 619572
rect 42351 619569 42417 619572
rect 676098 619454 676158 619866
rect 674895 619188 674961 619191
rect 674895 619186 675006 619188
rect 674895 619130 674900 619186
rect 674956 619130 675006 619186
rect 674895 619125 675006 619130
rect 674946 619010 675006 619125
rect 675898 618682 675904 618746
rect 675968 618682 675974 618746
rect 675906 618418 675966 618682
rect 41722 618238 41728 618302
rect 41792 618300 41798 618302
rect 42159 618300 42225 618303
rect 42298 618300 42304 618302
rect 41792 618298 42304 618300
rect 41792 618242 42164 618298
rect 42220 618242 42304 618298
rect 41792 618240 42304 618242
rect 41792 618238 41798 618240
rect 42159 618237 42225 618240
rect 42298 618238 42304 618240
rect 42368 618238 42374 618302
rect 673839 617856 673905 617859
rect 673839 617854 674784 617856
rect 673839 617798 673844 617854
rect 673900 617798 674784 617854
rect 673839 617796 674784 617798
rect 673839 617793 673905 617796
rect 41967 617710 42033 617711
rect 41914 617708 41920 617710
rect 41840 617648 41920 617708
rect 41984 617708 42033 617710
rect 42490 617708 42496 617710
rect 41984 617706 42496 617708
rect 42028 617650 42496 617706
rect 41914 617646 41920 617648
rect 41984 617648 42496 617650
rect 41984 617646 42033 617648
rect 42490 617646 42496 617648
rect 42560 617646 42566 617710
rect 41967 617645 42033 617646
rect 673263 617412 673329 617415
rect 673263 617410 674784 617412
rect 673263 617354 673268 617410
rect 673324 617354 674784 617410
rect 673263 617352 674784 617354
rect 673263 617349 673329 617352
rect 40954 617202 40960 617266
rect 41024 617264 41030 617266
rect 42447 617264 42513 617267
rect 41024 617262 42513 617264
rect 41024 617206 42452 617262
rect 42508 617206 42513 617262
rect 41024 617204 42513 617206
rect 41024 617202 41030 617204
rect 42447 617201 42513 617204
rect 673071 616820 673137 616823
rect 673071 616818 674784 616820
rect 673071 616762 673076 616818
rect 673132 616762 674784 616818
rect 673071 616760 674784 616762
rect 673071 616757 673137 616760
rect 40570 616462 40576 616526
rect 40640 616524 40646 616526
rect 42351 616524 42417 616527
rect 40640 616522 42417 616524
rect 40640 616466 42356 616522
rect 42412 616466 42417 616522
rect 40640 616464 42417 616466
rect 40640 616462 40646 616464
rect 42351 616461 42417 616464
rect 59535 616228 59601 616231
rect 59535 616226 64416 616228
rect 59535 616170 59540 616226
rect 59596 616170 64416 616226
rect 59535 616168 64416 616170
rect 59535 616165 59601 616168
rect 677058 615935 677118 616198
rect 677058 615930 677169 615935
rect 677058 615874 677108 615930
rect 677164 615874 677169 615930
rect 677058 615872 677169 615874
rect 677103 615869 677169 615872
rect 676866 615343 676926 615754
rect 676866 615338 676977 615343
rect 677103 615340 677169 615343
rect 676866 615282 676916 615338
rect 676972 615282 676977 615338
rect 676866 615280 676977 615282
rect 676911 615277 676977 615280
rect 677058 615338 677169 615340
rect 677058 615282 677108 615338
rect 677164 615282 677169 615338
rect 677058 615277 677169 615282
rect 677058 615162 677118 615277
rect 676911 614896 676977 614899
rect 676866 614894 676977 614896
rect 676866 614838 676916 614894
rect 676972 614838 676977 614894
rect 676866 614833 676977 614838
rect 676866 614570 676926 614833
rect 674746 613798 674752 613862
rect 674816 613860 674822 613862
rect 676090 613860 676096 613862
rect 674816 613800 676096 613860
rect 674816 613798 674822 613800
rect 676090 613798 676096 613800
rect 676160 613798 676166 613862
rect 673978 613650 673984 613714
rect 674048 613712 674054 613714
rect 675514 613712 675520 613714
rect 674048 613652 675520 613712
rect 674048 613650 674054 613652
rect 675514 613650 675520 613652
rect 675584 613650 675590 613714
rect 654351 613120 654417 613123
rect 650208 613118 654417 613120
rect 650208 613062 654356 613118
rect 654412 613062 654417 613118
rect 650208 613060 654417 613062
rect 654351 613057 654417 613060
rect 6648 609926 8736 610726
rect 9536 610725 50926 610726
rect 9536 609927 50127 610725
rect 50925 609927 50931 610725
rect 9536 609926 50926 609927
rect 6648 608646 16282 609446
rect 17082 609445 52718 609446
rect 17082 608647 51919 609445
rect 52717 608647 52723 609445
rect 17082 608646 52718 608647
rect 6192 607092 7318 607892
rect 8118 607891 54502 607892
rect 8118 607093 53703 607891
rect 54501 607093 54507 607891
rect 673978 607730 673984 607794
rect 674048 607792 674054 607794
rect 675375 607792 675441 607795
rect 674048 607790 675441 607792
rect 674048 607734 675380 607790
rect 675436 607734 675441 607790
rect 674048 607732 675441 607734
rect 674048 607730 674054 607732
rect 675375 607729 675441 607732
rect 675130 607138 675136 607202
rect 675200 607200 675206 607202
rect 675471 607200 675537 607203
rect 675200 607198 675537 607200
rect 675200 607142 675476 607198
rect 675532 607142 675537 607198
rect 675200 607140 675537 607142
rect 675200 607138 675206 607140
rect 675471 607137 675537 607140
rect 8118 607092 54502 607093
rect 675322 606546 675328 606610
rect 675392 606608 675398 606610
rect 675898 606608 675904 606610
rect 675392 606548 675904 606608
rect 675392 606546 675398 606548
rect 675898 606546 675904 606548
rect 675968 606546 675974 606610
rect 675322 606398 675328 606462
rect 675392 606460 675398 606462
rect 675471 606460 675537 606463
rect 675392 606458 675537 606460
rect 675392 606402 675476 606458
rect 675532 606402 675537 606458
rect 675392 606400 675537 606402
rect 675392 606398 675398 606400
rect 675471 606397 675537 606400
rect 6282 605356 17654 606156
rect 18454 606155 56068 606156
rect 18454 605357 55269 606155
rect 56067 605357 56073 606155
rect 18454 605356 56068 605357
rect 42298 605066 42304 605130
rect 42368 605066 42374 605130
rect 42490 605066 42496 605130
rect 42560 605066 42566 605130
rect 42306 604982 42366 605066
rect 42498 604982 42558 605066
rect 42298 604918 42304 604982
rect 42368 604918 42374 604982
rect 42490 604918 42496 604982
rect 42560 604918 42566 604982
rect 674362 604770 674368 604834
rect 674432 604832 674438 604834
rect 675375 604832 675441 604835
rect 674432 604830 675441 604832
rect 674432 604774 675380 604830
rect 675436 604774 675441 604830
rect 674432 604772 675441 604774
rect 674432 604770 674438 604772
rect 675375 604769 675441 604772
rect 42498 602911 42558 603026
rect 42447 602906 42558 602911
rect 42447 602850 42452 602906
rect 42508 602850 42558 602906
rect 42447 602848 42558 602850
rect 42447 602845 42513 602848
rect 42498 602464 42558 602582
rect 43215 602464 43281 602467
rect 42498 602462 43281 602464
rect 42498 602406 43220 602462
rect 43276 602406 43281 602462
rect 42498 602404 43281 602406
rect 43215 602401 43281 602404
rect 42351 602168 42417 602171
rect 42306 602166 42417 602168
rect 42306 602110 42356 602166
rect 42412 602110 42417 602166
rect 42306 602105 42417 602110
rect 42306 601990 42366 602105
rect 59535 601872 59601 601875
rect 59535 601870 64416 601872
rect 59535 601814 59540 601870
rect 59596 601814 64416 601870
rect 59535 601812 64416 601814
rect 59535 601809 59601 601812
rect 43215 601428 43281 601431
rect 654447 601428 654513 601431
rect 42528 601426 43281 601428
rect 42528 601370 43220 601426
rect 43276 601370 43281 601426
rect 42528 601368 43281 601370
rect 650208 601426 654513 601428
rect 650208 601370 654452 601426
rect 654508 601370 654513 601426
rect 650208 601368 654513 601370
rect 43215 601365 43281 601368
rect 654447 601365 654513 601368
rect 43983 601280 44049 601283
rect 42498 601278 44049 601280
rect 42498 601222 43988 601278
rect 44044 601222 44049 601278
rect 42498 601220 44049 601222
rect 42498 600880 42558 601220
rect 43983 601217 44049 601220
rect 675514 600478 675520 600542
rect 675584 600540 675590 600542
rect 676666 600540 676672 600542
rect 675584 600480 676672 600540
rect 675584 600478 675590 600480
rect 676666 600478 676672 600480
rect 676736 600478 676742 600542
rect 43791 600392 43857 600395
rect 42528 600390 43857 600392
rect 42528 600334 43796 600390
rect 43852 600334 43857 600390
rect 42528 600332 43857 600334
rect 43791 600329 43857 600332
rect 43407 600096 43473 600099
rect 43599 600096 43665 600099
rect 42498 600094 43665 600096
rect 42498 600038 43412 600094
rect 43468 600038 43604 600094
rect 43660 600038 43665 600094
rect 42498 600036 43665 600038
rect 42498 599770 42558 600036
rect 43407 600033 43473 600036
rect 43599 600033 43665 600036
rect 42874 599282 42880 599284
rect 42528 599222 42880 599282
rect 42874 599220 42880 599222
rect 42944 599220 42950 599284
rect 43119 598764 43185 598767
rect 42528 598762 43185 598764
rect 42528 598706 43124 598762
rect 43180 598706 43185 598762
rect 42528 598704 43185 598706
rect 43119 598701 43185 598704
rect 40386 597878 40446 598142
rect 40378 597814 40384 597878
rect 40448 597814 40454 597878
rect 41538 597287 41598 597624
rect 41538 597282 41649 597287
rect 41538 597226 41588 597282
rect 41644 597226 41649 597282
rect 41538 597224 41649 597226
rect 41583 597221 41649 597224
rect 41730 596843 41790 597106
rect 41730 596838 41841 596843
rect 41730 596782 41780 596838
rect 41836 596782 41841 596838
rect 41730 596780 41841 596782
rect 41775 596777 41841 596780
rect 41922 596251 41982 596514
rect 41871 596246 41982 596251
rect 41871 596190 41876 596246
rect 41932 596190 41982 596246
rect 41871 596188 41982 596190
rect 41871 596185 41937 596188
rect 40578 595658 40638 595996
rect 40570 595594 40576 595658
rect 40640 595594 40646 595658
rect 675087 595508 675153 595511
rect 676090 595508 676096 595510
rect 675087 595506 676096 595508
rect 41922 595215 41982 595478
rect 675087 595450 675092 595506
rect 675148 595450 676096 595506
rect 675087 595448 676096 595450
rect 675087 595445 675153 595448
rect 676090 595446 676096 595448
rect 676160 595446 676166 595510
rect 675759 595360 675825 595363
rect 676090 595360 676096 595362
rect 675759 595358 676096 595360
rect 675759 595302 675764 595358
rect 675820 595302 676096 595358
rect 675759 595300 676096 595302
rect 675759 595297 675825 595300
rect 676090 595298 676096 595300
rect 676160 595298 676166 595362
rect 41922 595210 42033 595215
rect 41922 595154 41972 595210
rect 42028 595154 42033 595210
rect 41922 595152 42033 595154
rect 41967 595149 42033 595152
rect 41730 594623 41790 594886
rect 674746 594706 674752 594770
rect 674816 594768 674822 594770
rect 675898 594768 675904 594770
rect 674816 594708 675904 594768
rect 674816 594706 674822 594708
rect 675898 594706 675904 594708
rect 675968 594706 675974 594770
rect 41679 594618 41790 594623
rect 41679 594562 41684 594618
rect 41740 594562 41790 594618
rect 41679 594560 41790 594562
rect 41679 594557 41745 594560
rect 42927 594398 42993 594401
rect 42528 594396 42993 594398
rect 42528 594340 42932 594396
rect 42988 594340 42993 594396
rect 42528 594338 42993 594340
rect 42927 594335 42993 594338
rect 42114 593587 42174 593850
rect 42063 593582 42174 593587
rect 42063 593526 42068 593582
rect 42124 593526 42174 593582
rect 42063 593524 42174 593526
rect 42063 593521 42129 593524
rect 675759 593436 675825 593439
rect 675898 593436 675904 593438
rect 675759 593434 675904 593436
rect 675759 593378 675764 593434
rect 675820 593378 675904 593434
rect 675759 593376 675904 593378
rect 675759 593373 675825 593376
rect 675898 593374 675904 593376
rect 675968 593374 675974 593438
rect 42114 592994 42174 593258
rect 42106 592930 42112 592994
rect 42176 592930 42182 592994
rect 43023 592770 43089 592773
rect 42528 592768 43089 592770
rect 42528 592712 43028 592768
rect 43084 592712 43089 592768
rect 42528 592710 43089 592712
rect 43023 592707 43089 592710
rect 671682 592642 699395 592643
rect 42498 591958 42558 592222
rect 42490 591894 42496 591958
rect 42560 591894 42566 591958
rect 42498 591364 42558 591630
rect 671677 591550 671683 592642
rect 672775 591550 699395 592642
rect 671682 591549 699395 591550
rect 700489 591549 711191 592643
rect 42498 591304 42750 591364
rect 30594 590774 30654 591112
rect 42690 590920 42750 591304
rect 42498 590860 42750 590920
rect 30586 590710 30592 590774
rect 30656 590710 30662 590774
rect 42498 590624 42558 590860
rect 674938 590858 674944 590922
rect 675008 590920 675014 590922
rect 676666 590920 676672 590922
rect 675008 590860 676672 590920
rect 675008 590858 675014 590860
rect 676666 590858 676672 590860
rect 676736 590858 676742 590922
rect 53775 590624 53841 590627
rect 42498 590622 53841 590624
rect 42498 590594 53780 590622
rect 42528 590566 53780 590594
rect 53836 590566 53841 590622
rect 42528 590564 53841 590566
rect 53775 590561 53841 590564
rect 674554 590562 674560 590626
rect 674624 590624 674630 590626
rect 674895 590624 674961 590627
rect 674624 590622 674961 590624
rect 674624 590566 674900 590622
rect 674956 590566 674961 590622
rect 674624 590564 674961 590566
rect 674624 590562 674630 590564
rect 674895 590561 674961 590564
rect 674607 590476 674673 590479
rect 675706 590476 675712 590478
rect 674607 590474 675712 590476
rect 674607 590418 674612 590474
rect 674668 590418 675712 590474
rect 674607 590416 675712 590418
rect 674607 590413 674673 590416
rect 675706 590414 675712 590416
rect 675776 590414 675782 590478
rect 675471 590330 675537 590331
rect 30586 590266 30592 590330
rect 30656 590328 30662 590330
rect 30656 590268 30846 590328
rect 30656 590266 30662 590268
rect 30786 590002 30846 590268
rect 674554 590266 674560 590330
rect 674624 590328 674630 590330
rect 675130 590328 675136 590330
rect 674624 590268 675136 590328
rect 674624 590266 674630 590268
rect 675130 590266 675136 590268
rect 675200 590266 675206 590330
rect 675471 590328 675520 590330
rect 675428 590326 675520 590328
rect 675428 590270 675476 590326
rect 675428 590268 675520 590270
rect 675471 590266 675520 590268
rect 675584 590266 675590 590330
rect 675471 590265 675537 590266
rect 674746 590118 674752 590182
rect 674816 590180 674822 590182
rect 674895 590180 674961 590183
rect 674816 590178 674961 590180
rect 674816 590122 674900 590178
rect 674956 590122 674961 590178
rect 674816 590120 674961 590122
rect 674816 590118 674822 590120
rect 674895 590117 674961 590120
rect 675130 589970 675136 590034
rect 675200 590032 675206 590034
rect 676474 590032 676480 590034
rect 675200 589972 676480 590032
rect 675200 589970 675206 589972
rect 676474 589970 676480 589972
rect 676544 589970 676550 590034
rect 676474 589822 676480 589886
rect 676544 589884 676550 589886
rect 676858 589884 676864 589886
rect 676544 589824 676864 589884
rect 676544 589822 676550 589824
rect 676858 589822 676864 589824
rect 676928 589822 676934 589886
rect 654447 589588 654513 589591
rect 650208 589586 654513 589588
rect 650208 589530 654452 589586
rect 654508 589530 654513 589586
rect 650208 589528 654513 589530
rect 654447 589525 654513 589528
rect 666066 589137 709314 589138
rect 41914 588934 41920 588998
rect 41984 588996 41990 588998
rect 42682 588996 42688 588998
rect 41984 588936 42688 588996
rect 41984 588934 41990 588936
rect 42682 588934 42688 588936
rect 42752 588934 42758 588998
rect 666061 587955 666067 589137
rect 667249 587955 709314 589137
rect 666066 587954 709314 587955
rect 710498 587954 710528 589138
rect 58767 587516 58833 587519
rect 58767 587514 64416 587516
rect 58767 587458 58772 587514
rect 58828 587458 64416 587514
rect 58767 587456 64416 587458
rect 58767 587453 58833 587456
rect 662178 587355 700810 587356
rect 662173 586173 662179 587355
rect 663361 586173 700810 587355
rect 662178 586172 700810 586173
rect 701994 586172 710096 587356
rect 659368 585085 708068 585086
rect 41967 584260 42033 584263
rect 42298 584260 42304 584262
rect 41967 584258 42304 584260
rect 41967 584202 41972 584258
rect 42028 584202 42304 584258
rect 41967 584200 42304 584202
rect 41967 584197 42033 584200
rect 42298 584198 42304 584200
rect 42368 584198 42374 584262
rect 659363 583903 659369 585085
rect 660551 583903 708068 585085
rect 659368 583902 708068 583903
rect 709252 583902 709934 585086
rect 674607 582188 674673 582191
rect 674754 582188 674814 582454
rect 674607 582186 674814 582188
rect 674607 582130 674612 582186
rect 674668 582130 674814 582186
rect 674607 582128 674814 582130
rect 674607 582125 674673 582128
rect 674415 581966 674481 581969
rect 674415 581964 674784 581966
rect 674415 581908 674420 581964
rect 674476 581908 674784 581964
rect 674415 581906 674784 581908
rect 674415 581903 674481 581906
rect 674607 581596 674673 581599
rect 674607 581594 674814 581596
rect 674607 581538 674612 581594
rect 674668 581538 674814 581594
rect 674607 581536 674814 581538
rect 674607 581533 674673 581536
rect 674754 581418 674814 581536
rect 42298 581238 42304 581302
rect 42368 581300 42374 581302
rect 42447 581300 42513 581303
rect 42368 581298 42513 581300
rect 42368 581242 42452 581298
rect 42508 581242 42513 581298
rect 42368 581240 42513 581242
rect 42368 581238 42374 581240
rect 42447 581237 42513 581240
rect 674415 580856 674481 580859
rect 674415 580854 674784 580856
rect 674415 580798 674420 580854
rect 674476 580798 674784 580854
rect 674415 580796 674784 580798
rect 674415 580793 674481 580796
rect 674607 580116 674673 580119
rect 674754 580116 674814 580234
rect 674607 580114 674814 580116
rect 674607 580058 674612 580114
rect 674668 580058 674814 580114
rect 674607 580056 674814 580058
rect 676911 580116 676977 580119
rect 676911 580114 677310 580116
rect 676911 580058 676916 580114
rect 676972 580058 677310 580114
rect 676911 580056 677310 580058
rect 674607 580053 674673 580056
rect 676911 580053 676977 580056
rect 676815 579524 676881 579527
rect 677250 579526 677310 580056
rect 676815 579522 677118 579524
rect 676815 579466 676820 579522
rect 676876 579466 677118 579522
rect 676815 579464 677118 579466
rect 676815 579461 676881 579464
rect 41722 579166 41728 579230
rect 41792 579228 41798 579230
rect 41914 579228 41920 579230
rect 41792 579168 41920 579228
rect 41792 579166 41798 579168
rect 41914 579166 41920 579168
rect 41984 579166 41990 579230
rect 677058 579082 677118 579464
rect 677242 579462 677248 579526
rect 677312 579462 677318 579526
rect 41530 579018 41536 579082
rect 41600 579080 41606 579082
rect 41600 579020 41838 579080
rect 41600 579018 41606 579020
rect 41778 578932 41838 579020
rect 42106 579018 42112 579082
rect 42176 579080 42182 579082
rect 42298 579080 42304 579082
rect 42176 579020 42304 579080
rect 42176 579018 42182 579020
rect 42298 579018 42304 579020
rect 42368 579018 42374 579082
rect 677050 579018 677056 579082
rect 677120 579018 677126 579082
rect 41914 578932 41920 578934
rect 41778 578872 41920 578932
rect 41914 578870 41920 578872
rect 41984 578870 41990 578934
rect 42159 578932 42225 578935
rect 42682 578932 42688 578934
rect 42159 578930 42688 578932
rect 42159 578874 42164 578930
rect 42220 578874 42688 578930
rect 42159 578872 42688 578874
rect 42159 578869 42225 578872
rect 42682 578870 42688 578872
rect 42752 578870 42758 578934
rect 676666 578870 676672 578934
rect 676736 578870 676742 578934
rect 676674 578606 676734 578870
rect 676474 578426 676480 578490
rect 676544 578426 676550 578490
rect 676482 578162 676542 578426
rect 654447 577896 654513 577899
rect 650208 577894 654513 577896
rect 650208 577838 654452 577894
rect 654508 577838 654513 577894
rect 650208 577836 654513 577838
rect 654447 577833 654513 577836
rect 674938 577834 674944 577898
rect 675008 577834 675014 577898
rect 674946 577570 675006 577834
rect 675514 577242 675520 577306
rect 675584 577242 675590 577306
rect 42927 577010 42993 577011
rect 42874 576946 42880 577010
rect 42944 577008 42993 577010
rect 42944 577006 43036 577008
rect 42988 576950 43036 577006
rect 675522 576978 675582 577242
rect 42944 576948 43036 576950
rect 42944 576946 42993 576948
rect 42927 576945 42993 576946
rect 676282 576798 676288 576862
rect 676352 576798 676358 576862
rect 676290 576534 676350 576798
rect 675130 576206 675136 576270
rect 675200 576206 675206 576270
rect 41967 575974 42033 575975
rect 41914 575910 41920 575974
rect 41984 575972 42033 575974
rect 41984 575970 42076 575972
rect 42028 575914 42076 575970
rect 675138 575942 675198 576206
rect 41984 575912 42076 575914
rect 41984 575910 42033 575912
rect 41967 575909 42033 575910
rect 674170 575318 674176 575382
rect 674240 575380 674246 575382
rect 674240 575320 674784 575380
rect 674240 575318 674246 575320
rect 674746 575170 674752 575234
rect 674816 575170 674822 575234
rect 674754 574906 674814 575170
rect 42063 574642 42129 574643
rect 42063 574640 42112 574642
rect 42020 574638 42112 574640
rect 42020 574582 42068 574638
rect 42020 574580 42112 574582
rect 42063 574578 42112 574580
rect 42176 574578 42182 574642
rect 42063 574577 42129 574578
rect 41775 574494 41841 574495
rect 41722 574430 41728 574494
rect 41792 574492 41841 574494
rect 674607 574492 674673 574495
rect 41792 574490 41884 574492
rect 41836 574434 41884 574490
rect 41792 574432 41884 574434
rect 674607 574490 674814 574492
rect 674607 574434 674612 574490
rect 674668 574434 674814 574490
rect 674607 574432 674814 574434
rect 41792 574430 41841 574432
rect 41775 574429 41841 574430
rect 674607 574429 674673 574432
rect 674754 574314 674814 574432
rect 40378 573838 40384 573902
rect 40448 573900 40454 573902
rect 43119 573900 43185 573903
rect 40448 573898 43185 573900
rect 40448 573842 43124 573898
rect 43180 573842 43185 573898
rect 40448 573840 43185 573842
rect 40448 573838 40454 573840
rect 43119 573837 43185 573840
rect 673359 573752 673425 573755
rect 673359 573750 674784 573752
rect 673359 573694 673364 573750
rect 673420 573694 674784 573750
rect 673359 573692 674784 573694
rect 673359 573689 673425 573692
rect 674607 573456 674673 573459
rect 674607 573454 674814 573456
rect 674607 573398 674612 573454
rect 674668 573398 674814 573454
rect 674607 573396 674814 573398
rect 674607 573393 674673 573396
rect 674754 573278 674814 573396
rect 40570 573098 40576 573162
rect 40640 573160 40646 573162
rect 42447 573160 42513 573163
rect 40640 573158 42513 573160
rect 40640 573102 42452 573158
rect 42508 573102 42513 573158
rect 40640 573100 42513 573102
rect 40640 573098 40646 573100
rect 42447 573097 42513 573100
rect 59535 573012 59601 573015
rect 59535 573010 64416 573012
rect 59535 572954 59540 573010
rect 59596 572954 64416 573010
rect 59535 572952 64416 572954
rect 59535 572949 59601 572952
rect 674607 572864 674673 572867
rect 674607 572862 674814 572864
rect 674607 572806 674612 572862
rect 674668 572806 674814 572862
rect 674607 572804 674814 572806
rect 674607 572801 674673 572804
rect 674754 572686 674814 572804
rect 673743 572124 673809 572127
rect 673743 572122 674784 572124
rect 673743 572066 673748 572122
rect 673804 572066 674784 572122
rect 673743 572064 674784 572066
rect 673743 572061 673809 572064
rect 674607 571828 674673 571831
rect 674607 571826 674814 571828
rect 674607 571770 674612 571826
rect 674668 571770 674814 571826
rect 674607 571768 674814 571770
rect 674607 571765 674673 571768
rect 674754 571576 674814 571768
rect 677058 570795 677118 571058
rect 677007 570790 677118 570795
rect 677007 570734 677012 570790
rect 677068 570734 677118 570790
rect 677007 570732 677118 570734
rect 677007 570729 677073 570732
rect 43791 570348 43857 570351
rect 43791 570346 43902 570348
rect 43791 570290 43796 570346
rect 43852 570290 43902 570346
rect 43791 570285 43902 570290
rect 43842 570203 43902 570285
rect 676866 570203 676926 570466
rect 43791 570198 43902 570203
rect 43791 570142 43796 570198
rect 43852 570142 43902 570198
rect 43791 570140 43902 570142
rect 676815 570198 676926 570203
rect 676815 570142 676820 570198
rect 676876 570142 676926 570198
rect 676815 570140 676926 570142
rect 677007 570200 677073 570203
rect 677007 570198 677118 570200
rect 677007 570142 677012 570198
rect 677068 570142 677118 570198
rect 43791 570137 43857 570140
rect 676815 570137 676881 570140
rect 677007 570137 677118 570142
rect 677058 569948 677118 570137
rect 676815 569756 676881 569759
rect 676815 569754 676926 569756
rect 676815 569698 676820 569754
rect 676876 569698 676926 569754
rect 676815 569693 676926 569698
rect 676866 569430 676926 569693
rect 7652 566846 8620 567646
rect 9420 567645 50926 567646
rect 9420 566847 50127 567645
rect 50925 566847 50931 567645
rect 9420 566846 50926 566847
rect 7108 565744 16256 566544
rect 17056 566543 52718 566544
rect 17056 565745 51919 566543
rect 52717 565745 52723 566543
rect 654447 566204 654513 566207
rect 650208 566202 654513 566204
rect 650208 566146 654452 566202
rect 654508 566146 654513 566202
rect 650208 566144 654513 566146
rect 654447 566141 654513 566144
rect 17056 565744 52718 565745
rect 6836 564474 7348 565274
rect 8148 565273 54502 565274
rect 8148 564475 53703 565273
rect 54501 564475 54507 565273
rect 8148 564474 54502 564475
rect 6564 563022 17620 563822
rect 18420 563821 56068 563822
rect 18420 563023 55269 563821
rect 56067 563023 56073 563821
rect 18420 563022 56068 563023
rect 674938 562442 674944 562506
rect 675008 562504 675014 562506
rect 675471 562504 675537 562507
rect 675008 562502 675537 562504
rect 675008 562446 675476 562502
rect 675532 562446 675537 562502
rect 675008 562444 675537 562446
rect 675008 562442 675014 562444
rect 675471 562441 675537 562444
rect 674170 561998 674176 562062
rect 674240 562060 674246 562062
rect 675471 562060 675537 562063
rect 674240 562058 675537 562060
rect 674240 562002 675476 562058
rect 675532 562002 675537 562058
rect 674240 562000 675537 562002
rect 674240 561998 674246 562000
rect 675471 561997 675537 562000
rect 41914 561554 41920 561618
rect 41984 561616 41990 561618
rect 42490 561616 42496 561618
rect 41984 561556 42496 561616
rect 41984 561554 41990 561556
rect 42490 561554 42496 561556
rect 42560 561554 42566 561618
rect 675130 561406 675136 561470
rect 675200 561468 675206 561470
rect 675375 561468 675441 561471
rect 675200 561466 675441 561468
rect 675200 561410 675380 561466
rect 675436 561410 675441 561466
rect 675200 561408 675441 561410
rect 675200 561406 675206 561408
rect 675375 561405 675441 561408
rect 40186 560518 40192 560582
rect 40256 560580 40262 560582
rect 43503 560580 43569 560583
rect 40256 560578 43569 560580
rect 40256 560522 43508 560578
rect 43564 560522 43569 560578
rect 40256 560520 43569 560522
rect 40256 560518 40262 560520
rect 43503 560517 43569 560520
rect 42498 559547 42558 559810
rect 42498 559542 42609 559547
rect 42498 559486 42548 559542
rect 42604 559486 42609 559542
rect 42498 559484 42609 559486
rect 42543 559481 42609 559484
rect 42498 559103 42558 559366
rect 42447 559098 42558 559103
rect 42447 559042 42452 559098
rect 42508 559042 42558 559098
rect 42447 559040 42558 559042
rect 42447 559037 42513 559040
rect 59535 558952 59601 558955
rect 59535 558950 64416 558952
rect 59535 558894 59540 558950
rect 59596 558894 64416 558950
rect 59535 558892 64416 558894
rect 59535 558889 59601 558892
rect 674746 558890 674752 558954
rect 674816 558952 674822 558954
rect 675471 558952 675537 558955
rect 674816 558950 675537 558952
rect 674816 558894 675476 558950
rect 675532 558894 675537 558950
rect 674816 558892 675537 558894
rect 674816 558890 674822 558892
rect 675471 558889 675537 558892
rect 42927 558804 42993 558807
rect 42528 558802 42993 558804
rect 42528 558746 42932 558802
rect 42988 558746 42993 558802
rect 42528 558744 42993 558746
rect 42927 558741 42993 558744
rect 43407 558508 43473 558511
rect 42306 558506 43473 558508
rect 42306 558450 43412 558506
rect 43468 558450 43473 558506
rect 42306 558448 43473 558450
rect 42306 558182 42366 558448
rect 43407 558445 43473 558448
rect 43215 558064 43281 558067
rect 42498 558062 43281 558064
rect 42498 558006 43220 558062
rect 43276 558006 43281 558062
rect 42498 558004 43281 558006
rect 42498 557738 42558 558004
rect 43215 558001 43281 558004
rect 40186 556818 40192 556882
rect 40256 556818 40262 556882
rect 42498 556880 42558 557146
rect 43599 556880 43665 556883
rect 42498 556878 43665 556880
rect 42498 556822 43604 556878
rect 43660 556822 43665 556878
rect 42498 556820 43665 556822
rect 40194 556554 40254 556818
rect 43599 556817 43665 556820
rect 41730 555847 41790 556110
rect 41679 555842 41790 555847
rect 41679 555786 41684 555842
rect 41740 555786 41790 555842
rect 41679 555784 41790 555786
rect 41679 555781 41745 555784
rect 41922 555255 41982 555518
rect 41922 555250 42033 555255
rect 41922 555194 41972 555250
rect 42028 555194 42033 555250
rect 41922 555192 42033 555194
rect 41967 555189 42033 555192
rect 40386 554662 40446 554926
rect 40378 554598 40384 554662
rect 40448 554598 40454 554662
rect 654447 554512 654513 554515
rect 650208 554510 654513 554512
rect 41730 554071 41790 554482
rect 650208 554454 654452 554510
rect 654508 554454 654513 554510
rect 650208 554452 654513 554454
rect 654447 554449 654513 554452
rect 675759 554512 675825 554515
rect 676858 554512 676864 554514
rect 675759 554510 676864 554512
rect 675759 554454 675764 554510
rect 675820 554454 676864 554510
rect 675759 554452 676864 554454
rect 675759 554449 675825 554452
rect 676858 554450 676864 554452
rect 676928 554450 676934 554514
rect 41730 554066 41841 554071
rect 41730 554010 41780 554066
rect 41836 554010 41841 554066
rect 41730 554008 41841 554010
rect 41775 554005 41841 554008
rect 42927 553920 42993 553923
rect 42528 553918 42993 553920
rect 42528 553862 42932 553918
rect 42988 553862 42993 553918
rect 42528 553860 42993 553862
rect 42927 553857 42993 553860
rect 42498 553035 42558 553298
rect 42447 553030 42558 553035
rect 42447 552974 42452 553030
rect 42508 552974 42558 553030
rect 42447 552972 42558 552974
rect 42447 552969 42513 552972
rect 40578 552442 40638 552854
rect 40570 552378 40576 552442
rect 40640 552378 40646 552442
rect 42114 551999 42174 552262
rect 42063 551994 42174 551999
rect 42063 551938 42068 551994
rect 42124 551938 42174 551994
rect 42063 551936 42174 551938
rect 42063 551933 42129 551936
rect 41922 551407 41982 551670
rect 41871 551402 41982 551407
rect 41871 551346 41876 551402
rect 41932 551346 41982 551402
rect 41871 551344 41982 551346
rect 41871 551341 41937 551344
rect 43023 551182 43089 551185
rect 42528 551180 43089 551182
rect 42528 551124 43028 551180
rect 43084 551124 43089 551180
rect 42528 551122 43089 551124
rect 43023 551119 43089 551122
rect 42114 550371 42174 550634
rect 42114 550366 42225 550371
rect 42114 550310 42164 550366
rect 42220 550310 42225 550366
rect 42114 550308 42225 550310
rect 42159 550305 42225 550308
rect 41730 549779 41790 550042
rect 41730 549774 41841 549779
rect 41730 549718 41780 549774
rect 41836 549718 41841 549774
rect 41730 549716 41841 549718
rect 41775 549713 41841 549716
rect 42831 549554 42897 549557
rect 42528 549552 42897 549554
rect 42528 549496 42836 549552
rect 42892 549496 42897 549552
rect 42528 549494 42897 549496
rect 42831 549491 42897 549494
rect 43023 549036 43089 549039
rect 42528 549034 43089 549036
rect 42528 548978 43028 549034
rect 43084 548978 43089 549034
rect 42528 548976 43089 548978
rect 43023 548973 43089 548976
rect 42498 548148 42558 548414
rect 42498 548088 42750 548148
rect 35202 547559 35262 547896
rect 42690 547704 42750 548088
rect 35151 547554 35262 547559
rect 35151 547498 35156 547554
rect 35212 547498 35262 547554
rect 35151 547496 35262 547498
rect 42498 547644 42750 547704
rect 35151 547493 35217 547496
rect 42498 547408 42558 547644
rect 44847 547408 44913 547411
rect 42498 547406 44913 547408
rect 42498 547378 44852 547406
rect 42528 547350 44852 547378
rect 44908 547350 44913 547406
rect 42528 547348 44913 547350
rect 44847 547345 44913 547348
rect 671682 547150 699205 547151
rect 35151 547112 35217 547115
rect 35151 547110 35262 547112
rect 35151 547054 35156 547110
rect 35212 547054 35262 547110
rect 35151 547049 35262 547054
rect 35202 546786 35262 547049
rect 671677 546058 671683 547150
rect 672775 546058 699205 547150
rect 671682 546057 699205 546058
rect 700299 546057 710823 547151
rect 666066 545495 709418 545496
rect 59535 544448 59601 544451
rect 59535 544446 64416 544448
rect 59535 544390 59540 544446
rect 59596 544390 64416 544446
rect 59535 544388 64416 544390
rect 59535 544385 59601 544388
rect 666061 544313 666067 545495
rect 667249 544313 709418 545495
rect 666066 544312 709418 544313
rect 710602 544312 711294 545496
rect 662178 543901 700596 543902
rect 662173 542719 662179 543901
rect 663361 542719 700596 543901
rect 662178 542718 700596 542719
rect 701780 542718 711028 543902
rect 654447 542672 654513 542675
rect 650208 542670 654513 542672
rect 650208 542614 654452 542670
rect 654508 542614 654513 542670
rect 650208 542612 654513 542614
rect 654447 542609 654513 542612
rect 659368 541881 707930 541882
rect 42927 541638 42993 541639
rect 42874 541636 42880 541638
rect 42836 541576 42880 541636
rect 42944 541634 42993 541638
rect 42988 541578 42993 541634
rect 42874 541574 42880 541576
rect 42944 541574 42993 541578
rect 42927 541573 42993 541574
rect 41679 541340 41745 541343
rect 42682 541340 42688 541342
rect 41679 541338 42688 541340
rect 41679 541282 41684 541338
rect 41740 541282 42688 541338
rect 41679 541280 42688 541282
rect 41679 541277 41745 541280
rect 42682 541278 42688 541280
rect 42752 541278 42758 541342
rect 41775 541192 41841 541195
rect 42298 541192 42304 541194
rect 41775 541190 42304 541192
rect 41775 541134 41780 541190
rect 41836 541134 42304 541190
rect 41775 541132 42304 541134
rect 41775 541129 41841 541132
rect 42298 541130 42304 541132
rect 42368 541130 42374 541194
rect 41871 541046 41937 541047
rect 41871 541044 41920 541046
rect 41828 541042 41920 541044
rect 41828 540986 41876 541042
rect 41828 540984 41920 540986
rect 41871 540982 41920 540984
rect 41984 540982 41990 541046
rect 41871 540981 41937 540982
rect 42159 540748 42225 540751
rect 42447 540748 42513 540751
rect 42159 540746 42513 540748
rect 42159 540690 42164 540746
rect 42220 540690 42452 540746
rect 42508 540690 42513 540746
rect 659363 540699 659369 541881
rect 660551 540699 707930 541881
rect 659368 540698 707930 540699
rect 709114 540698 711506 541882
rect 42159 540688 42513 540690
rect 42159 540685 42225 540688
rect 42447 540685 42513 540688
rect 676866 537199 676926 537462
rect 676815 537194 676926 537199
rect 676815 537138 676820 537194
rect 676876 537138 676926 537194
rect 676815 537136 676926 537138
rect 676815 537133 676881 537136
rect 41914 536838 41920 536902
rect 41984 536900 41990 536902
rect 42447 536900 42513 536903
rect 41984 536898 42513 536900
rect 41984 536842 42452 536898
rect 42508 536842 42513 536898
rect 41984 536840 42513 536842
rect 41984 536838 41990 536840
rect 42447 536837 42513 536840
rect 673743 536900 673809 536903
rect 673743 536898 674784 536900
rect 673743 536842 673748 536898
rect 673804 536842 674784 536898
rect 673743 536840 674784 536842
rect 673743 536837 673809 536840
rect 674607 536604 674673 536607
rect 674607 536602 674814 536604
rect 674607 536546 674612 536602
rect 674668 536546 674814 536602
rect 674607 536544 674814 536546
rect 674607 536541 674673 536544
rect 674754 536426 674814 536544
rect 673743 535864 673809 535867
rect 673743 535862 674784 535864
rect 673743 535806 673748 535862
rect 673804 535806 674784 535862
rect 673743 535804 674784 535806
rect 673743 535801 673809 535804
rect 42874 535654 42880 535718
rect 42944 535716 42950 535718
rect 43023 535716 43089 535719
rect 42944 535714 43089 535716
rect 42944 535658 43028 535714
rect 43084 535658 43089 535714
rect 42944 535656 43089 535658
rect 42944 535654 42950 535656
rect 43023 535653 43089 535656
rect 677242 535062 677248 535126
rect 677312 535062 677318 535126
rect 677250 534535 677310 535062
rect 677442 534979 677502 535242
rect 677391 534974 677502 534979
rect 677391 534918 677396 534974
rect 677452 534918 677502 534974
rect 677391 534916 677502 534918
rect 677391 534913 677457 534916
rect 677050 534470 677056 534534
rect 677120 534470 677126 534534
rect 677199 534530 677310 534535
rect 677199 534474 677204 534530
rect 677260 534474 677310 534530
rect 677199 534472 677310 534474
rect 42682 534322 42688 534386
rect 42752 534384 42758 534386
rect 42927 534384 42993 534387
rect 42752 534382 42993 534384
rect 42752 534326 42932 534382
rect 42988 534326 42993 534382
rect 42752 534324 42993 534326
rect 42752 534322 42758 534324
rect 42927 534321 42993 534324
rect 677058 533943 677118 534470
rect 677199 534469 677265 534472
rect 675322 533878 675328 533942
rect 675392 533878 675398 533942
rect 677007 533938 677118 533943
rect 677007 533882 677012 533938
rect 677068 533882 677118 533938
rect 677007 533880 677118 533882
rect 675330 533614 675390 533878
rect 677007 533877 677073 533880
rect 676090 533434 676096 533498
rect 676160 533434 676166 533498
rect 42351 533350 42417 533351
rect 42298 533286 42304 533350
rect 42368 533348 42417 533350
rect 42368 533346 42460 533348
rect 42412 533290 42460 533346
rect 42368 533288 42460 533290
rect 42368 533286 42417 533288
rect 42351 533285 42417 533286
rect 676098 533170 676158 533434
rect 42159 532756 42225 532759
rect 42490 532756 42496 532758
rect 42159 532754 42496 532756
rect 42159 532698 42164 532754
rect 42220 532698 42496 532754
rect 42159 532696 42496 532698
rect 42159 532693 42225 532696
rect 42490 532694 42496 532696
rect 42560 532694 42566 532758
rect 673978 532546 673984 532610
rect 674048 532608 674054 532610
rect 674048 532548 674784 532608
rect 674048 532546 674054 532548
rect 674362 531954 674368 532018
rect 674432 532016 674438 532018
rect 674432 531956 674784 532016
rect 674432 531954 674438 531956
rect 41914 531806 41920 531870
rect 41984 531868 41990 531870
rect 42159 531868 42225 531871
rect 41984 531866 42225 531868
rect 41984 531810 42164 531866
rect 42220 531810 42225 531866
rect 41984 531808 42225 531810
rect 41984 531806 41990 531808
rect 42159 531805 42225 531808
rect 675706 531806 675712 531870
rect 675776 531806 675782 531870
rect 41775 531722 41841 531723
rect 41722 531658 41728 531722
rect 41792 531720 41841 531722
rect 41792 531718 41884 531720
rect 41836 531662 41884 531718
rect 41792 531660 41884 531662
rect 41792 531658 41841 531660
rect 41775 531657 41841 531658
rect 675714 531542 675774 531806
rect 40570 531214 40576 531278
rect 40640 531276 40646 531278
rect 42351 531276 42417 531279
rect 40640 531274 42417 531276
rect 40640 531218 42356 531274
rect 42412 531218 42417 531274
rect 40640 531216 42417 531218
rect 40640 531214 40646 531216
rect 42351 531213 42417 531216
rect 675898 531214 675904 531278
rect 675968 531214 675974 531278
rect 654063 530980 654129 530983
rect 650208 530978 654129 530980
rect 650208 530922 654068 530978
rect 654124 530922 654129 530978
rect 675906 530950 675966 531214
rect 650208 530920 654129 530922
rect 654063 530917 654129 530920
rect 40378 530622 40384 530686
rect 40448 530684 40454 530686
rect 42927 530684 42993 530687
rect 40448 530682 42993 530684
rect 40448 530626 42932 530682
rect 42988 530626 42993 530682
rect 40448 530624 42993 530626
rect 40448 530622 40454 530624
rect 42927 530621 42993 530624
rect 674554 530622 674560 530686
rect 674624 530684 674630 530686
rect 674624 530624 674814 530684
rect 674624 530622 674630 530624
rect 674754 530358 674814 530624
rect 59535 530092 59601 530095
rect 59535 530090 64416 530092
rect 59535 530034 59540 530090
rect 59596 530034 64416 530090
rect 59535 530032 64416 530034
rect 59535 530029 59601 530032
rect 673743 529944 673809 529947
rect 673743 529942 674814 529944
rect 673743 529886 673748 529942
rect 673804 529886 674814 529942
rect 673743 529884 674814 529886
rect 673743 529881 673809 529884
rect 674754 529840 674814 529884
rect 674895 529500 674961 529503
rect 674895 529498 675006 529500
rect 674895 529442 674900 529498
rect 674956 529442 675006 529498
rect 674895 529437 675006 529442
rect 674946 529322 675006 529437
rect 673743 528760 673809 528763
rect 673743 528758 674784 528760
rect 673743 528702 673748 528758
rect 673804 528702 674784 528758
rect 673743 528700 674784 528702
rect 673743 528697 673809 528700
rect 673743 528316 673809 528319
rect 673743 528314 674814 528316
rect 673743 528258 673748 528314
rect 673804 528258 674814 528314
rect 673743 528256 674814 528258
rect 673743 528253 673809 528256
rect 674754 528212 674814 528256
rect 673263 527724 673329 527727
rect 673263 527722 674784 527724
rect 673263 527666 673268 527722
rect 673324 527666 674784 527722
rect 673263 527664 674784 527666
rect 673263 527661 673329 527664
rect 673071 527132 673137 527135
rect 673071 527130 674784 527132
rect 673071 527074 673076 527130
rect 673132 527074 674784 527130
rect 673071 527072 674784 527074
rect 673071 527069 673137 527072
rect 672975 526688 673041 526691
rect 672975 526686 674814 526688
rect 672975 526630 672980 526686
rect 673036 526630 674814 526686
rect 672975 526628 674814 526630
rect 672975 526625 673041 526628
rect 674754 526584 674814 526628
rect 677058 525803 677118 526066
rect 677058 525798 677169 525803
rect 677058 525742 677108 525798
rect 677164 525742 677169 525798
rect 677058 525740 677169 525742
rect 677103 525737 677169 525740
rect 676866 525211 676926 525474
rect 676815 525206 676926 525211
rect 677103 525208 677169 525211
rect 676815 525150 676820 525206
rect 676876 525150 676926 525206
rect 676815 525148 676926 525150
rect 677058 525206 677169 525208
rect 677058 525150 677108 525206
rect 677164 525150 677169 525206
rect 676815 525145 676881 525148
rect 677058 525145 677169 525150
rect 677058 524956 677118 525145
rect 676815 524764 676881 524767
rect 676815 524762 676926 524764
rect 676815 524706 676820 524762
rect 676876 524706 676926 524762
rect 676815 524701 676926 524706
rect 676866 524438 676926 524701
rect 654447 519288 654513 519291
rect 650208 519286 654513 519288
rect 650208 519230 654452 519286
rect 654508 519230 654513 519286
rect 650208 519228 654513 519230
rect 654447 519225 654513 519228
rect 669318 518470 677862 518476
rect 669304 518424 677862 518470
rect 669304 518422 669372 518424
rect 59535 515736 59601 515739
rect 59535 515734 64416 515736
rect 59535 515678 59540 515734
rect 59596 515678 64416 515734
rect 59535 515676 64416 515678
rect 59535 515673 59601 515676
rect 669304 514106 669368 518422
rect 654447 507448 654513 507451
rect 650208 507446 654513 507448
rect 650208 507390 654452 507446
rect 654508 507390 654513 507446
rect 650208 507388 654513 507390
rect 654447 507385 654513 507388
rect 669304 504232 669372 514106
rect 670344 514050 677862 518424
rect 670344 508556 670422 514050
rect 670344 508462 677998 508556
rect 670350 504232 677998 508462
rect 669304 504156 677998 504232
rect 669304 504066 670422 504156
rect 674895 504044 674961 504047
rect 675087 504044 675153 504047
rect 674895 504042 675153 504044
rect 674895 503986 674900 504042
rect 674956 503986 675092 504042
rect 675148 503986 675153 504042
rect 674895 503984 675153 503986
rect 674895 503981 674961 503984
rect 675087 503981 675153 503984
rect 671682 503088 699153 503089
rect 671677 501996 671683 503088
rect 672775 501996 699153 503088
rect 671682 501995 699153 501996
rect 700247 501995 711355 503089
rect 666066 501273 709152 501274
rect 59535 501232 59601 501235
rect 59535 501230 64416 501232
rect 59535 501174 59540 501230
rect 59596 501174 64416 501230
rect 59535 501172 64416 501174
rect 59535 501169 59601 501172
rect 666061 500091 666067 501273
rect 667249 500091 709152 501273
rect 666066 500090 709152 500091
rect 710336 500090 711188 501274
rect 662178 499413 700596 499414
rect 662173 498231 662179 499413
rect 663361 498231 700596 499413
rect 662178 498230 700596 498231
rect 701780 498230 710816 499414
rect 659368 497499 708036 497500
rect 42530 497306 47070 497352
rect 38434 497304 47070 497306
rect 38434 493252 45974 497304
rect 42530 487666 45974 493252
rect 38012 483786 45974 487666
rect 46716 483786 47070 497304
rect 659363 496317 659369 497499
rect 660551 496317 708036 497499
rect 659368 496316 708036 496317
rect 709220 496316 710444 497500
rect 654351 495756 654417 495759
rect 650208 495754 654417 495756
rect 650208 495698 654356 495754
rect 654412 495698 654417 495754
rect 650208 495696 654417 495698
rect 654351 495693 654417 495696
rect 674607 493240 674673 493243
rect 674754 493240 674814 493506
rect 674607 493238 674814 493240
rect 674607 493182 674612 493238
rect 674668 493182 674814 493238
rect 674607 493180 674814 493182
rect 674607 493177 674673 493180
rect 674319 492944 674385 492947
rect 674319 492942 674784 492944
rect 674319 492886 674324 492942
rect 674380 492886 674784 492942
rect 674319 492884 674784 492886
rect 674319 492881 674385 492884
rect 673839 492352 673905 492355
rect 673839 492350 674784 492352
rect 673839 492294 673844 492350
rect 673900 492294 674784 492350
rect 673839 492292 674784 492294
rect 673839 492289 673905 492292
rect 677391 492204 677457 492207
rect 677391 492202 677502 492204
rect 677391 492146 677396 492202
rect 677452 492146 677502 492202
rect 677391 492141 677502 492146
rect 677442 491878 677502 492141
rect 677199 491168 677265 491171
rect 677199 491166 677694 491168
rect 677199 491110 677204 491166
rect 677260 491110 677694 491166
rect 677199 491108 677694 491110
rect 677199 491105 677265 491108
rect 676815 490576 676881 490579
rect 677634 490578 677694 491108
rect 677826 491022 677886 491286
rect 677818 490958 677824 491022
rect 677888 490958 677894 491022
rect 676815 490574 676926 490576
rect 676815 490518 676820 490574
rect 676876 490518 676926 490574
rect 676815 490513 676926 490518
rect 677626 490514 677632 490578
rect 677696 490514 677702 490578
rect 676866 490280 676926 490513
rect 676866 490250 677472 490280
rect 676896 490220 677502 490250
rect 677442 489986 677502 490220
rect 675130 489922 675136 489986
rect 675200 489922 675206 489986
rect 677434 489922 677440 489986
rect 677504 489922 677510 489986
rect 675138 489658 675198 489922
rect 674511 489392 674577 489395
rect 674511 489390 674814 489392
rect 674511 489334 674516 489390
rect 674572 489334 674814 489390
rect 674511 489332 674814 489334
rect 674511 489329 674577 489332
rect 674754 489066 674814 489332
rect 674938 488886 674944 488950
rect 675008 488886 675014 488950
rect 674946 488622 675006 488886
rect 675375 488356 675441 488359
rect 675330 488354 675441 488356
rect 675330 488298 675380 488354
rect 675436 488298 675441 488354
rect 675330 488293 675441 488298
rect 675330 488030 675390 488293
rect 674415 487468 674481 487471
rect 674415 487466 674784 487468
rect 674415 487410 674420 487466
rect 674476 487410 674784 487466
rect 674415 487408 674784 487410
rect 674415 487405 674481 487408
rect 674991 487172 675057 487175
rect 674946 487170 675057 487172
rect 674946 487114 674996 487170
rect 675052 487114 675057 487170
rect 674946 487109 675057 487114
rect 674946 486994 675006 487109
rect 58575 486876 58641 486879
rect 58575 486874 64416 486876
rect 58575 486818 58580 486874
rect 58636 486818 64416 486874
rect 58575 486816 64416 486818
rect 58575 486813 58641 486816
rect 674170 486370 674176 486434
rect 674240 486432 674246 486434
rect 674240 486372 674784 486432
rect 674240 486370 674246 486372
rect 674746 486074 674752 486138
rect 674816 486074 674822 486138
rect 674754 485810 674814 486074
rect 674895 485544 674961 485547
rect 674895 485542 675006 485544
rect 674895 485486 674900 485542
rect 674956 485486 675006 485542
rect 674895 485481 675006 485486
rect 674946 485366 675006 485481
rect 674223 484804 674289 484807
rect 674223 484802 674784 484804
rect 674223 484746 674228 484802
rect 674284 484746 674784 484802
rect 674223 484744 674784 484746
rect 674223 484741 674289 484744
rect 673167 484212 673233 484215
rect 673167 484210 674784 484212
rect 673167 484154 673172 484210
rect 673228 484154 674784 484210
rect 673167 484152 674784 484154
rect 673167 484149 673233 484152
rect 654255 484064 654321 484067
rect 650208 484062 654321 484064
rect 650208 484006 654260 484062
rect 654316 484006 654321 484062
rect 650208 484004 654321 484006
rect 654255 484001 654321 484004
rect 38012 483668 47070 483786
rect 673455 483768 673521 483771
rect 673455 483766 674814 483768
rect 673455 483710 673460 483766
rect 673516 483710 674814 483766
rect 673455 483708 674814 483710
rect 673455 483705 673521 483708
rect 674754 483664 674814 483708
rect 676858 483410 676864 483474
rect 676928 483410 676934 483474
rect 676866 483146 676926 483410
rect 673359 482584 673425 482587
rect 673359 482582 674784 482584
rect 673359 482526 673364 482582
rect 673420 482526 674784 482582
rect 673359 482524 674784 482526
rect 673359 482521 673425 482524
rect 677058 481699 677118 482036
rect 677007 481694 677118 481699
rect 677007 481638 677012 481694
rect 677068 481638 677118 481694
rect 677007 481636 677118 481638
rect 677007 481633 677073 481636
rect 676866 481255 676926 481518
rect 676815 481250 676926 481255
rect 676815 481194 676820 481250
rect 676876 481194 676926 481250
rect 676815 481192 676926 481194
rect 677007 481252 677073 481255
rect 677007 481250 677118 481252
rect 677007 481194 677012 481250
rect 677068 481194 677118 481250
rect 676815 481189 676881 481192
rect 677007 481189 677118 481194
rect 677058 480926 677118 481189
rect 676815 480808 676881 480811
rect 676815 480806 676926 480808
rect 676815 480750 676820 480806
rect 676876 480750 676926 480806
rect 676815 480745 676926 480750
rect 676866 480408 676926 480745
rect 674338 474082 680474 474094
rect 674110 474078 680474 474082
rect 659822 473848 680474 474078
rect 59535 472520 59601 472523
rect 59535 472518 64416 472520
rect 59535 472462 59540 472518
rect 59596 472462 64416 472518
rect 59535 472460 64416 472462
rect 59535 472457 59601 472460
rect 654447 472224 654513 472227
rect 650208 472222 654513 472224
rect 650208 472166 654452 472222
rect 654508 472166 654513 472222
rect 650208 472164 654513 472166
rect 654447 472161 654513 472164
rect 654447 460532 654513 460535
rect 650208 460530 654513 460532
rect 650208 460474 654452 460530
rect 654508 460474 654513 460530
rect 650208 460472 654513 460474
rect 654447 460469 654513 460472
rect 659822 460522 665144 473848
rect 668046 470186 680474 473848
rect 668046 464288 676620 470186
rect 668046 460522 681110 464288
rect 659822 460394 681110 460522
rect 659822 460256 676620 460394
rect 59535 458164 59601 458167
rect 59535 458162 64416 458164
rect 59535 458106 59540 458162
rect 59596 458106 64416 458162
rect 59535 458104 64416 458106
rect 59535 458101 59601 458104
rect 37822 454820 44492 454846
rect 47144 454820 49272 454828
rect 37822 454744 49272 454820
rect 37822 451458 47166 454744
rect 42366 445418 47166 451458
rect 36928 441662 47166 445418
rect 49188 441662 49272 454744
rect 654351 448840 654417 448843
rect 650208 448838 654417 448840
rect 650208 448782 654356 448838
rect 654412 448782 654417 448838
rect 650208 448780 654417 448782
rect 654351 448777 654417 448780
rect 59535 443808 59601 443811
rect 59535 443806 64416 443808
rect 59535 443750 59540 443806
rect 59596 443750 64416 443806
rect 59535 443748 64416 443750
rect 59535 443745 59601 443748
rect 36928 441608 49272 441662
rect 36928 441582 44730 441608
rect 47144 441602 49272 441608
rect 6098 439190 8774 439990
rect 9574 439989 50926 439990
rect 9574 439191 50127 439989
rect 50925 439191 50931 439989
rect 9574 439190 50926 439191
rect 6648 437824 16250 438624
rect 17050 438623 52718 438624
rect 17050 437825 51919 438623
rect 52717 437825 52723 438623
rect 17050 437824 52718 437825
rect 6918 436296 7356 437096
rect 8156 437095 54502 437096
rect 8156 436297 53703 437095
rect 54501 436297 54507 437095
rect 654447 437000 654513 437003
rect 650208 436998 654513 437000
rect 650208 436942 654452 436998
rect 654508 436942 654513 436998
rect 650208 436940 654513 436942
rect 654447 436937 654513 436940
rect 8156 436296 54502 436297
rect 6378 434948 17690 435748
rect 18490 435747 56068 435748
rect 18490 434949 55269 435747
rect 56067 434949 56073 435747
rect 18490 434948 56068 434949
rect 42831 432264 42897 432267
rect 42528 432262 42897 432264
rect 42528 432206 42836 432262
rect 42892 432206 42897 432262
rect 42528 432204 42897 432206
rect 42831 432201 42897 432204
rect 42831 431746 42897 431749
rect 42528 431744 42897 431746
rect 42528 431688 42836 431744
rect 42892 431688 42897 431744
rect 42528 431686 42897 431688
rect 42831 431683 42897 431686
rect 42351 431376 42417 431379
rect 42306 431374 42417 431376
rect 42306 431318 42356 431374
rect 42412 431318 42417 431374
rect 42306 431313 42417 431318
rect 42306 431198 42366 431313
rect 43215 430636 43281 430639
rect 42528 430634 43281 430636
rect 42528 430578 43220 430634
rect 43276 430578 43281 430634
rect 42528 430576 43281 430578
rect 43215 430573 43281 430576
rect 43407 430192 43473 430195
rect 42498 430190 43473 430192
rect 42498 430134 43412 430190
rect 43468 430134 43473 430190
rect 42498 430132 43473 430134
rect 42498 430088 42558 430132
rect 43407 430129 43473 430132
rect 42831 429600 42897 429603
rect 40416 429598 42897 429600
rect 40416 429570 42836 429598
rect 40386 429542 42836 429570
rect 42892 429542 42897 429598
rect 40386 429540 42897 429542
rect 40386 429306 40446 429540
rect 42831 429537 42897 429540
rect 59535 429452 59601 429455
rect 59535 429450 64416 429452
rect 59535 429394 59540 429450
rect 59596 429394 64416 429450
rect 59535 429392 64416 429394
rect 59535 429389 59601 429392
rect 40378 429242 40384 429306
rect 40448 429242 40454 429306
rect 43503 429008 43569 429011
rect 40608 429006 43569 429008
rect 40608 428978 43508 429006
rect 40578 428950 43508 428978
rect 43564 428950 43569 429006
rect 40578 428948 43569 428950
rect 40578 428714 40638 428948
rect 43503 428945 43569 428948
rect 40570 428650 40576 428714
rect 40640 428650 40646 428714
rect 40962 428122 41022 428460
rect 40954 428058 40960 428122
rect 41024 428058 41030 428122
rect 42831 427972 42897 427975
rect 42528 427970 42897 427972
rect 42528 427914 42836 427970
rect 42892 427914 42897 427970
rect 42528 427912 42897 427914
rect 42831 427909 42897 427912
rect 40770 427086 40830 427350
rect 40762 427022 40768 427086
rect 40832 427022 40838 427086
rect 41346 426494 41406 426832
rect 41338 426430 41344 426494
rect 41408 426430 41414 426494
rect 41538 426050 41598 426314
rect 41530 425986 41536 426050
rect 41600 425986 41606 426050
rect 41922 425459 41982 425722
rect 41871 425454 41982 425459
rect 654447 425456 654513 425459
rect 41871 425398 41876 425454
rect 41932 425398 41982 425454
rect 41871 425396 41982 425398
rect 650208 425454 654513 425456
rect 650208 425398 654452 425454
rect 654508 425398 654513 425454
rect 650208 425396 654513 425398
rect 41871 425393 41937 425396
rect 654447 425393 654513 425396
rect 41154 424866 41214 425204
rect 41146 424802 41152 424866
rect 41216 424802 41222 424866
rect 42114 424422 42174 424686
rect 42106 424358 42112 424422
rect 42176 424358 42182 424422
rect 42306 423978 42366 424094
rect 42298 423914 42304 423978
rect 42368 423914 42374 423978
rect 40194 423387 40254 423576
rect 40194 423382 40305 423387
rect 40194 423326 40244 423382
rect 40300 423326 40305 423382
rect 40194 423324 40305 423326
rect 40239 423321 40305 423324
rect 40002 422795 40062 423058
rect 39951 422790 40062 422795
rect 39951 422734 39956 422790
rect 40012 422734 40062 422790
rect 39951 422732 40062 422734
rect 39951 422729 40017 422732
rect 40002 422203 40062 422466
rect 40002 422198 40113 422203
rect 40002 422142 40052 422198
rect 40108 422142 40113 422198
rect 40002 422140 40113 422142
rect 40047 422137 40113 422140
rect 40194 421611 40254 421874
rect 40143 421606 40254 421611
rect 40143 421550 40148 421606
rect 40204 421550 40254 421606
rect 40143 421548 40254 421550
rect 40143 421545 40209 421548
rect 42927 421460 42993 421463
rect 42528 421458 42993 421460
rect 42528 421402 42932 421458
rect 42988 421402 42993 421458
rect 42528 421400 42993 421402
rect 42927 421397 42993 421400
rect 42306 420575 42366 420838
rect 42306 420570 42417 420575
rect 42306 420514 42356 420570
rect 42412 420514 42417 420570
rect 42306 420512 42417 420514
rect 42351 420509 42417 420512
rect 35202 419983 35262 420246
rect 35151 419978 35262 419983
rect 35151 419922 35156 419978
rect 35212 419922 35262 419978
rect 35151 419920 35262 419922
rect 35151 419917 35217 419920
rect 42306 419539 42366 419802
rect 35151 419536 35217 419539
rect 35151 419534 35262 419536
rect 35151 419478 35156 419534
rect 35212 419478 35262 419534
rect 35151 419473 35262 419478
rect 42306 419534 42417 419539
rect 42306 419478 42356 419534
rect 42412 419478 42417 419534
rect 42306 419476 42417 419478
rect 42351 419473 42417 419476
rect 35202 419210 35262 419473
rect 58383 415096 58449 415099
rect 58383 415094 64416 415096
rect 58383 415038 58388 415094
rect 58444 415038 64416 415094
rect 58383 415036 64416 415038
rect 58383 415033 58449 415036
rect 671682 414948 699209 414949
rect 671677 413856 671683 414948
rect 672775 413856 699209 414948
rect 671682 413855 699209 413856
rect 700303 413855 711689 414949
rect 653871 413616 653937 413619
rect 650208 413614 653937 413616
rect 650208 413558 653876 413614
rect 653932 413558 653937 413614
rect 650208 413556 653937 413558
rect 653871 413553 653937 413556
rect 666066 412999 709366 413000
rect 666061 411817 666067 412999
rect 667249 411817 709366 412999
rect 666066 411816 709366 411817
rect 710550 411816 711682 413000
rect 662178 411215 700720 411216
rect 662173 410033 662179 411215
rect 663361 410033 700720 411215
rect 662178 410032 700720 410033
rect 701904 410032 711578 411216
rect 659368 409431 708100 409432
rect 659363 408249 659369 409431
rect 660551 408249 708100 409431
rect 659368 408248 708100 408249
rect 709284 408248 711786 409432
rect 41530 406006 41536 406070
rect 41600 406068 41606 406070
rect 41775 406068 41841 406071
rect 41600 406066 41841 406068
rect 41600 406010 41780 406066
rect 41836 406010 41841 406066
rect 41600 406008 41841 406010
rect 41600 406006 41606 406008
rect 41775 406005 41841 406008
rect 674703 405476 674769 405479
rect 674703 405474 674814 405476
rect 674703 405418 674708 405474
rect 674764 405418 674814 405474
rect 674703 405413 674814 405418
rect 674754 405298 674814 405413
rect 41871 405182 41937 405183
rect 41871 405180 41920 405182
rect 41828 405178 41920 405180
rect 41828 405122 41876 405178
rect 41828 405120 41920 405122
rect 41871 405118 41920 405120
rect 41984 405118 41990 405182
rect 41871 405117 41937 405118
rect 674415 404736 674481 404739
rect 674415 404734 674784 404736
rect 674415 404678 674420 404734
rect 674476 404678 674784 404734
rect 674415 404676 674784 404678
rect 674415 404673 674481 404676
rect 41775 404442 41841 404443
rect 41722 404378 41728 404442
rect 41792 404440 41841 404442
rect 674703 404440 674769 404443
rect 41792 404438 41884 404440
rect 41836 404382 41884 404438
rect 41792 404380 41884 404382
rect 674703 404438 674814 404440
rect 674703 404382 674708 404438
rect 674764 404382 674814 404438
rect 41792 404378 41841 404380
rect 41775 404377 41841 404378
rect 674703 404377 674814 404382
rect 674754 404188 674814 404377
rect 677818 403934 677824 403998
rect 677888 403934 677894 403998
rect 677826 403670 677886 403934
rect 42159 403108 42225 403111
rect 42298 403108 42304 403110
rect 42159 403106 42304 403108
rect 42159 403050 42164 403106
rect 42220 403050 42304 403106
rect 42159 403048 42304 403050
rect 42159 403045 42225 403048
rect 42298 403046 42304 403048
rect 42368 403046 42374 403110
rect 673647 403108 673713 403111
rect 673647 403106 674784 403108
rect 673647 403050 673652 403106
rect 673708 403050 674784 403106
rect 673647 403048 674784 403050
rect 673647 403045 673713 403048
rect 677626 402750 677632 402814
rect 677696 402750 677702 402814
rect 42159 402666 42225 402667
rect 42106 402664 42112 402666
rect 42068 402604 42112 402664
rect 42176 402662 42225 402666
rect 42220 402606 42225 402662
rect 42106 402602 42112 402604
rect 42176 402602 42225 402606
rect 42159 402601 42225 402602
rect 677295 402368 677361 402371
rect 677634 402368 677694 402750
rect 677295 402366 677694 402368
rect 677295 402310 677300 402366
rect 677356 402310 677694 402366
rect 677295 402308 677694 402310
rect 677295 402305 677361 402308
rect 677434 402158 677440 402222
rect 677504 402158 677510 402222
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 654447 401776 654513 401779
rect 650208 401774 654513 401776
rect 650208 401718 654452 401774
rect 654508 401718 654513 401774
rect 650208 401716 654513 401718
rect 654447 401713 654513 401716
rect 677103 401776 677169 401779
rect 677442 401776 677502 402158
rect 677103 401774 677502 401776
rect 677103 401718 677108 401774
rect 677164 401718 677502 401774
rect 677103 401716 677502 401718
rect 677103 401713 677169 401716
rect 674946 401335 675006 401450
rect 674895 401330 675006 401335
rect 674895 401274 674900 401330
rect 674956 401274 675006 401330
rect 674895 401272 675006 401274
rect 674895 401269 674961 401272
rect 58383 400740 58449 400743
rect 58383 400738 64416 400740
rect 58383 400682 58388 400738
rect 58444 400682 64416 400738
rect 58383 400680 64416 400682
rect 58383 400677 58449 400680
rect 674554 400530 674560 400594
rect 674624 400592 674630 400594
rect 674754 400592 674814 400858
rect 674624 400532 674814 400592
rect 674624 400530 674630 400532
rect 674946 400151 675006 400414
rect 40954 400086 40960 400150
rect 41024 400148 41030 400150
rect 41775 400148 41841 400151
rect 41024 400146 41841 400148
rect 41024 400090 41780 400146
rect 41836 400090 41841 400146
rect 41024 400088 41841 400090
rect 674946 400146 675057 400151
rect 674946 400090 674996 400146
rect 675052 400090 675057 400146
rect 674946 400088 675057 400090
rect 41024 400086 41030 400088
rect 41775 400085 41841 400088
rect 674991 400085 675057 400088
rect 674511 399704 674577 399707
rect 674754 399704 674814 399822
rect 674511 399702 674814 399704
rect 674511 399646 674516 399702
rect 674572 399646 674814 399702
rect 674511 399644 674814 399646
rect 674511 399641 674577 399644
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 674362 399198 674368 399262
rect 674432 399260 674438 399262
rect 674432 399200 674784 399260
rect 674432 399198 674438 399200
rect 40762 398754 40768 398818
rect 40832 398816 40838 398818
rect 41775 398816 41841 398819
rect 40832 398814 41841 398816
rect 40832 398758 41780 398814
rect 41836 398758 41841 398814
rect 40832 398756 41841 398758
rect 40832 398754 40838 398756
rect 41775 398753 41841 398756
rect 674170 398754 674176 398818
rect 674240 398816 674246 398818
rect 674240 398756 674784 398816
rect 674240 398754 674246 398756
rect 675138 397931 675198 398194
rect 675138 397926 675249 397931
rect 675138 397870 675188 397926
rect 675244 397870 675249 397926
rect 675138 397868 675249 397870
rect 675183 397865 675249 397868
rect 674415 397632 674481 397635
rect 674415 397630 674784 397632
rect 674415 397574 674420 397630
rect 674476 397574 674784 397630
rect 674415 397572 674784 397574
rect 674415 397569 674481 397572
rect 675138 396895 675198 397158
rect 675087 396890 675198 396895
rect 6846 396038 8624 396838
rect 9424 396837 50926 396838
rect 9424 396039 50127 396837
rect 50925 396039 50931 396837
rect 675087 396834 675092 396890
rect 675148 396834 675198 396890
rect 675087 396832 675198 396834
rect 675087 396829 675153 396832
rect 673935 396596 674001 396599
rect 673935 396594 674784 396596
rect 673935 396538 673940 396594
rect 673996 396538 674784 396594
rect 673935 396536 674784 396538
rect 673935 396533 674001 396536
rect 9424 396038 50926 396039
rect 674607 395856 674673 395859
rect 674754 395856 674814 395974
rect 674607 395854 674814 395856
rect 674607 395798 674612 395854
rect 674668 395798 674814 395854
rect 674607 395796 674814 395798
rect 674607 395793 674673 395796
rect 6400 394606 16362 395406
rect 17162 395405 52718 395406
rect 17162 394607 51919 395405
rect 52717 394607 52723 395405
rect 674754 395119 674814 395530
rect 674703 395114 674814 395119
rect 674703 395058 674708 395114
rect 674764 395058 674814 395114
rect 674703 395056 674814 395058
rect 674703 395053 674769 395056
rect 674754 394675 674814 394938
rect 674754 394670 674865 394675
rect 674754 394614 674804 394670
rect 674860 394614 674865 394670
rect 674754 394612 674865 394614
rect 674799 394609 674865 394612
rect 17162 394606 52718 394607
rect 674223 394376 674289 394379
rect 674223 394374 674784 394376
rect 674223 394318 674228 394374
rect 674284 394318 674784 394374
rect 674223 394316 674784 394318
rect 674223 394313 674289 394316
rect 6042 393086 7322 393886
rect 8122 393885 54502 393886
rect 8122 393087 53703 393885
rect 54501 393087 54507 393885
rect 677058 393491 677118 393902
rect 677058 393486 677169 393491
rect 677058 393430 677108 393486
rect 677164 393430 677169 393486
rect 677058 393428 677169 393430
rect 677103 393425 677169 393428
rect 8122 393086 54502 393087
rect 676866 393047 676926 393310
rect 676866 393042 676977 393047
rect 677103 393044 677169 393047
rect 676866 392986 676916 393042
rect 676972 392986 676977 393042
rect 676866 392984 676977 392986
rect 676911 392981 676977 392984
rect 677058 393042 677169 393044
rect 677058 392986 677108 393042
rect 677164 392986 677169 393042
rect 677058 392981 677169 392986
rect 677058 392718 677118 392981
rect 676911 392600 676977 392603
rect 676866 392598 676977 392600
rect 676866 392542 676916 392598
rect 676972 392542 676977 392598
rect 676866 392537 676977 392542
rect 6132 391566 17528 392366
rect 18328 392365 56068 392366
rect 18328 391567 55269 392365
rect 56067 391567 56073 392365
rect 676866 392200 676926 392537
rect 18328 391566 56068 391567
rect 654447 390084 654513 390087
rect 650208 390082 654513 390084
rect 650208 390026 654452 390082
rect 654508 390026 654513 390082
rect 650208 390024 654513 390026
rect 654447 390021 654513 390024
rect 42351 389344 42417 389347
rect 42306 389342 42417 389344
rect 42306 389286 42356 389342
rect 42412 389286 42417 389342
rect 42306 389281 42417 389286
rect 42306 389018 42366 389281
rect 42351 388752 42417 388755
rect 42306 388750 42417 388752
rect 42306 388694 42356 388750
rect 42412 388694 42417 388750
rect 42306 388689 42417 388694
rect 42306 388574 42366 388689
rect 42735 388012 42801 388015
rect 42528 388010 42801 388012
rect 42528 387954 42740 388010
rect 42796 387954 42801 388010
rect 42528 387952 42801 387954
rect 42735 387949 42801 387952
rect 42498 387272 42558 387390
rect 43311 387272 43377 387275
rect 42498 387270 43377 387272
rect 42498 387214 43316 387270
rect 43372 387214 43377 387270
rect 42498 387212 43377 387214
rect 43311 387209 43377 387212
rect 43215 387124 43281 387127
rect 42498 387122 43281 387124
rect 42498 387066 43220 387122
rect 43276 387066 43281 387122
rect 42498 387064 43281 387066
rect 42498 386946 42558 387064
rect 43215 387061 43281 387064
rect 59247 386384 59313 386387
rect 59247 386382 64416 386384
rect 40386 386090 40446 386354
rect 59247 386326 59252 386382
rect 59308 386326 64416 386382
rect 59247 386324 64416 386326
rect 59247 386321 59313 386324
rect 40378 386026 40384 386090
rect 40448 386026 40454 386090
rect 40570 386026 40576 386090
rect 40640 386026 40646 386090
rect 40578 385762 40638 386026
rect 40962 384906 41022 385318
rect 40954 384842 40960 384906
rect 41024 384842 41030 384906
rect 42114 384463 42174 384726
rect 42114 384458 42225 384463
rect 42114 384402 42164 384458
rect 42220 384402 42225 384458
rect 42114 384400 42225 384402
rect 42159 384397 42225 384400
rect 40770 383870 40830 384134
rect 40762 383806 40768 383870
rect 40832 383806 40838 383870
rect 41346 383278 41406 383616
rect 41338 383214 41344 383278
rect 41408 383214 41414 383278
rect 41538 382834 41598 383098
rect 41530 382770 41536 382834
rect 41600 382770 41606 382834
rect 42306 382243 42366 382506
rect 42306 382238 42417 382243
rect 42306 382182 42356 382238
rect 42412 382182 42417 382238
rect 42306 382180 42417 382182
rect 42351 382177 42417 382180
rect 41154 381650 41214 381988
rect 41146 381586 41152 381650
rect 41216 381586 41222 381650
rect 40002 381207 40062 381470
rect 40002 381202 40113 381207
rect 40002 381146 40052 381202
rect 40108 381146 40113 381202
rect 40002 381144 40113 381146
rect 40047 381141 40113 381144
rect 40194 380615 40254 380878
rect 40143 380610 40254 380615
rect 40143 380554 40148 380610
rect 40204 380554 40254 380610
rect 40143 380552 40254 380554
rect 40143 380549 40209 380552
rect 40002 380171 40062 380360
rect 39951 380166 40062 380171
rect 39951 380110 39956 380166
rect 40012 380110 40062 380166
rect 39951 380108 40062 380110
rect 39951 380105 40017 380108
rect 42498 379579 42558 379842
rect 42498 379574 42609 379579
rect 42498 379518 42548 379574
rect 42604 379518 42609 379574
rect 42498 379516 42609 379518
rect 42543 379513 42609 379516
rect 39810 378987 39870 379250
rect 39810 378982 39921 378987
rect 39810 378926 39860 378982
rect 39916 378926 39921 378982
rect 39810 378924 39921 378926
rect 39855 378921 39921 378924
rect 674362 378774 674368 378838
rect 674432 378836 674438 378838
rect 675471 378836 675537 378839
rect 674432 378834 675537 378836
rect 674432 378778 675476 378834
rect 675532 378778 675537 378834
rect 674432 378776 675537 378778
rect 674432 378774 674438 378776
rect 675471 378773 675537 378776
rect 40194 378395 40254 378732
rect 654447 378540 654513 378543
rect 650208 378538 654513 378540
rect 650208 378482 654452 378538
rect 654508 378482 654513 378538
rect 650208 378480 654513 378482
rect 654447 378477 654513 378480
rect 40194 378390 40305 378395
rect 40194 378334 40244 378390
rect 40300 378334 40305 378390
rect 40194 378332 40305 378334
rect 40239 378329 40305 378332
rect 43119 378244 43185 378247
rect 42528 378242 43185 378244
rect 42528 378186 43124 378242
rect 43180 378186 43185 378242
rect 42528 378184 43185 378186
rect 43119 378181 43185 378184
rect 42639 377652 42705 377655
rect 42528 377650 42705 377652
rect 42528 377594 42644 377650
rect 42700 377594 42705 377650
rect 42528 377592 42705 377594
rect 42639 377589 42705 377592
rect 35202 376767 35262 377104
rect 35151 376762 35262 376767
rect 35151 376706 35156 376762
rect 35212 376706 35262 376762
rect 35151 376704 35262 376706
rect 35151 376701 35217 376704
rect 42639 376616 42705 376619
rect 42528 376614 42705 376616
rect 42528 376558 42644 376614
rect 42700 376558 42705 376614
rect 42528 376556 42705 376558
rect 42639 376553 42705 376556
rect 35151 376320 35217 376323
rect 35151 376318 35262 376320
rect 35151 376262 35156 376318
rect 35212 376262 35262 376318
rect 35151 376257 35262 376262
rect 35202 375994 35262 376257
rect 40047 375136 40113 375139
rect 42106 375136 42112 375138
rect 40047 375134 42112 375136
rect 40047 375078 40052 375134
rect 40108 375078 42112 375134
rect 40047 375076 42112 375078
rect 40047 375073 40113 375076
rect 42106 375074 42112 375076
rect 42176 375074 42182 375138
rect 675087 374544 675153 374547
rect 675322 374544 675328 374546
rect 675087 374542 675328 374544
rect 675087 374486 675092 374542
rect 675148 374486 675328 374542
rect 675087 374484 675328 374486
rect 675087 374481 675153 374484
rect 675322 374482 675328 374484
rect 675392 374482 675398 374546
rect 673359 374396 673425 374399
rect 677050 374396 677056 374398
rect 673359 374394 677056 374396
rect 673359 374338 673364 374394
rect 673420 374338 677056 374394
rect 673359 374336 677056 374338
rect 673359 374333 673425 374336
rect 677050 374334 677056 374336
rect 677120 374334 677126 374398
rect 675183 374100 675249 374103
rect 675514 374100 675520 374102
rect 675183 374098 675520 374100
rect 675183 374042 675188 374098
rect 675244 374042 675520 374098
rect 675183 374040 675520 374042
rect 675183 374037 675249 374040
rect 675514 374038 675520 374040
rect 675584 374038 675590 374102
rect 674554 373890 674560 373954
rect 674624 373952 674630 373954
rect 675471 373952 675537 373955
rect 674624 373950 675537 373952
rect 674624 373894 675476 373950
rect 675532 373894 675537 373950
rect 674624 373892 675537 373894
rect 674624 373890 674630 373892
rect 675471 373889 675537 373892
rect 673455 373064 673521 373067
rect 677050 373064 677056 373066
rect 673455 373062 677056 373064
rect 673455 373006 673460 373062
rect 673516 373006 677056 373062
rect 673455 373004 677056 373006
rect 673455 373001 673521 373004
rect 677050 373002 677056 373004
rect 677120 373002 677126 373066
rect 40143 372916 40209 372919
rect 42298 372916 42304 372918
rect 40143 372914 42304 372916
rect 40143 372858 40148 372914
rect 40204 372858 42304 372914
rect 40143 372856 42304 372858
rect 40143 372853 40209 372856
rect 42298 372854 42304 372856
rect 42368 372854 42374 372918
rect 674170 371966 674176 372030
rect 674240 372028 674246 372030
rect 675375 372028 675441 372031
rect 674240 372026 675441 372028
rect 674240 371970 675380 372026
rect 675436 371970 675441 372026
rect 674240 371968 675441 371970
rect 674240 371966 674246 371968
rect 675375 371965 675441 371968
rect 59535 371880 59601 371883
rect 59535 371878 64416 371880
rect 59535 371822 59540 371878
rect 59596 371822 64416 371878
rect 59535 371820 64416 371822
rect 59535 371817 59601 371820
rect 671682 369980 699307 369981
rect 671677 368888 671683 369980
rect 672775 368888 699307 369980
rect 671682 368887 699307 368888
rect 700401 368887 711389 369981
rect 666066 367915 709268 367916
rect 666061 366733 666067 367915
rect 667249 366733 709268 367915
rect 666066 366732 709268 366733
rect 710452 366732 711590 367916
rect 654447 366552 654513 366555
rect 650208 366550 654513 366552
rect 650208 366494 654452 366550
rect 654508 366494 654513 366550
rect 650208 366492 654513 366494
rect 654447 366489 654513 366492
rect 662178 366061 700568 366062
rect 662173 364879 662179 366061
rect 663361 364879 700568 366061
rect 662178 364878 700568 364879
rect 701752 364878 711486 366062
rect 659368 364311 707888 364312
rect 659363 363129 659369 364311
rect 660551 363129 707888 364311
rect 659368 363128 707888 363129
rect 709072 363128 711640 364312
rect 41530 362790 41536 362854
rect 41600 362852 41606 362854
rect 41775 362852 41841 362855
rect 41600 362850 41841 362852
rect 41600 362794 41780 362850
rect 41836 362794 41841 362850
rect 41600 362792 41841 362794
rect 41600 362790 41606 362792
rect 41775 362789 41841 362792
rect 41914 360866 41920 360930
rect 41984 360928 41990 360930
rect 42063 360928 42129 360931
rect 42490 360928 42496 360930
rect 41984 360926 42496 360928
rect 41984 360870 42068 360926
rect 42124 360870 42496 360926
rect 41984 360868 42496 360870
rect 41984 360866 41990 360868
rect 42063 360865 42129 360868
rect 42490 360866 42496 360868
rect 42560 360866 42566 360930
rect 41722 360570 41728 360634
rect 41792 360632 41798 360634
rect 41967 360632 42033 360635
rect 42682 360632 42688 360634
rect 41792 360630 42688 360632
rect 41792 360574 41972 360630
rect 42028 360574 42688 360630
rect 41792 360572 42688 360574
rect 41792 360570 41798 360572
rect 41967 360569 42033 360572
rect 42682 360570 42688 360572
rect 42752 360570 42758 360634
rect 674415 360040 674481 360043
rect 674415 360038 674784 360040
rect 674415 359982 674420 360038
rect 674476 359982 674784 360038
rect 674415 359980 674784 359982
rect 674415 359977 674481 359980
rect 42159 359892 42225 359895
rect 42298 359892 42304 359894
rect 42159 359890 42304 359892
rect 42159 359834 42164 359890
rect 42220 359834 42304 359890
rect 42159 359832 42304 359834
rect 42159 359829 42225 359832
rect 42298 359830 42304 359832
rect 42368 359830 42374 359894
rect 674703 359744 674769 359747
rect 674703 359742 674814 359744
rect 674703 359686 674708 359742
rect 674764 359686 674814 359742
rect 674703 359681 674814 359686
rect 674754 359566 674814 359681
rect 42063 359450 42129 359451
rect 42063 359446 42112 359450
rect 42176 359448 42182 359450
rect 42063 359390 42068 359446
rect 42063 359386 42112 359390
rect 42176 359388 42220 359448
rect 42176 359386 42182 359388
rect 42063 359385 42129 359386
rect 674415 359004 674481 359007
rect 674415 359002 674784 359004
rect 674415 358946 674420 359002
rect 674476 358946 674784 359002
rect 674415 358944 674784 358946
rect 674415 358941 674481 358944
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 673839 358412 673905 358415
rect 673839 358410 674784 358412
rect 673839 358354 673844 358410
rect 673900 358354 674784 358410
rect 673839 358352 674784 358354
rect 673839 358349 673905 358352
rect 59535 357672 59601 357675
rect 676866 357674 676926 357938
rect 59535 357670 64416 357672
rect 59535 357614 59540 357670
rect 59596 357614 64416 357670
rect 59535 357612 64416 357614
rect 59535 357609 59601 357612
rect 676858 357610 676864 357674
rect 676928 357610 676934 357674
rect 677050 357610 677056 357674
rect 677120 357610 677126 357674
rect 677058 357346 677118 357610
rect 40954 356870 40960 356934
rect 41024 356932 41030 356934
rect 41775 356932 41841 356935
rect 41024 356930 41841 356932
rect 41024 356874 41780 356930
rect 41836 356874 41841 356930
rect 41024 356872 41841 356874
rect 41024 356870 41030 356872
rect 41775 356869 41841 356872
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 677442 356490 677502 356754
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 677434 356426 677440 356490
rect 677504 356426 677510 356490
rect 674415 356340 674481 356343
rect 674415 356338 674784 356340
rect 674415 356282 674420 356338
rect 674476 356282 674784 356338
rect 674415 356280 674784 356282
rect 674415 356277 674481 356280
rect 673978 355686 673984 355750
rect 674048 355748 674054 355750
rect 674048 355688 674784 355748
rect 674048 355686 674054 355688
rect 40762 355538 40768 355602
rect 40832 355600 40838 355602
rect 41775 355600 41841 355603
rect 40832 355598 41841 355600
rect 40832 355542 41780 355598
rect 41836 355542 41841 355598
rect 40832 355540 41841 355542
rect 40832 355538 40838 355540
rect 41775 355537 41841 355540
rect 674754 355011 674814 355126
rect 674754 355006 674865 355011
rect 674754 354950 674804 355006
rect 674860 354950 674865 355006
rect 674754 354948 674865 354950
rect 674799 354945 674865 354948
rect 655215 354860 655281 354863
rect 650208 354858 655281 354860
rect 650208 354802 655220 354858
rect 655276 354802 655281 354858
rect 650208 354800 655281 354802
rect 655215 354797 655281 354800
rect 674607 354416 674673 354419
rect 674754 354416 674814 354682
rect 674607 354414 674814 354416
rect 674607 354358 674612 354414
rect 674668 354358 674814 354414
rect 674607 354356 674814 354358
rect 674607 354353 674673 354356
rect 673935 354120 674001 354123
rect 673935 354118 674784 354120
rect 673935 354062 673940 354118
rect 673996 354062 674784 354118
rect 673935 354060 674784 354062
rect 673935 354057 674001 354060
rect 677058 353235 677118 353498
rect 677007 353230 677118 353235
rect 677007 353174 677012 353230
rect 677068 353174 677118 353230
rect 677007 353172 677118 353174
rect 677007 353169 677073 353172
rect 6168 352300 8636 353100
rect 9436 353099 50926 353100
rect 9436 352301 50127 353099
rect 50925 352301 50931 353099
rect 674946 352791 675006 353054
rect 674895 352786 675006 352791
rect 674895 352730 674900 352786
rect 674956 352730 675006 352786
rect 674895 352728 675006 352730
rect 674895 352725 674961 352728
rect 9436 352300 50926 352301
rect 674511 352196 674577 352199
rect 674754 352196 674814 352462
rect 674511 352194 674814 352196
rect 674511 352138 674516 352194
rect 674572 352138 674814 352194
rect 674511 352136 674814 352138
rect 674511 352133 674577 352136
rect 5372 351238 16348 352038
rect 17148 352037 52718 352038
rect 17148 351239 51919 352037
rect 52717 351239 52723 352037
rect 674946 351755 675006 351870
rect 674946 351750 675057 351755
rect 674946 351694 674996 351750
rect 675052 351694 675057 351750
rect 674946 351692 675057 351694
rect 674991 351689 675057 351692
rect 17148 351238 52718 351239
rect 676866 351163 676926 351352
rect 676815 351158 676926 351163
rect 676815 351102 676820 351158
rect 676876 351102 676926 351158
rect 676815 351100 676926 351102
rect 676815 351097 676881 351100
rect 5814 350088 7236 350888
rect 8036 350887 54502 350888
rect 8036 350089 53703 350887
rect 54501 350089 54507 350887
rect 674319 350864 674385 350867
rect 674319 350862 674784 350864
rect 674319 350806 674324 350862
rect 674380 350806 674784 350862
rect 674319 350804 674784 350806
rect 674319 350801 674385 350804
rect 674754 350127 674814 350242
rect 674703 350122 674814 350127
rect 8036 350088 54502 350089
rect 674703 350066 674708 350122
rect 674764 350066 674814 350122
rect 674703 350064 674814 350066
rect 674703 350061 674769 350064
rect 674223 349754 674289 349757
rect 674223 349752 674784 349754
rect 674223 349696 674228 349752
rect 674284 349696 674784 349752
rect 674223 349694 674784 349696
rect 674223 349691 674289 349694
rect 5636 348586 17548 349386
rect 18348 349385 56068 349386
rect 18348 348587 55269 349385
rect 56067 348587 56073 349385
rect 674031 349236 674097 349239
rect 674031 349234 674784 349236
rect 674031 349178 674036 349234
rect 674092 349178 674784 349234
rect 674031 349176 674784 349178
rect 674031 349173 674097 349176
rect 18348 348586 56068 348587
rect 677058 348351 677118 348614
rect 677058 348346 677169 348351
rect 677058 348290 677108 348346
rect 677164 348290 677169 348346
rect 677058 348288 677169 348290
rect 677103 348285 677169 348288
rect 676866 347759 676926 348096
rect 676866 347754 676977 347759
rect 677103 347756 677169 347759
rect 676866 347698 676916 347754
rect 676972 347698 676977 347754
rect 676866 347696 676977 347698
rect 676911 347693 676977 347696
rect 677058 347754 677169 347756
rect 677058 347698 677108 347754
rect 677164 347698 677169 347754
rect 677058 347693 677169 347698
rect 677058 347578 677118 347693
rect 676911 347312 676977 347315
rect 676866 347310 676977 347312
rect 676866 347254 676916 347310
rect 676972 347254 676977 347310
rect 676866 347249 676977 347254
rect 676866 346986 676926 347249
rect 42447 346128 42513 346131
rect 42447 346126 42558 346128
rect 42447 346070 42452 346126
rect 42508 346070 42558 346126
rect 42447 346065 42558 346070
rect 42498 345876 42558 346065
rect 42447 345536 42513 345539
rect 42447 345534 42558 345536
rect 42447 345478 42452 345534
rect 42508 345478 42558 345534
rect 42447 345473 42558 345478
rect 676474 345474 676480 345538
rect 676544 345536 676550 345538
rect 676815 345536 676881 345539
rect 676544 345534 676881 345536
rect 676544 345478 676820 345534
rect 676876 345478 676881 345534
rect 676544 345476 676881 345478
rect 676544 345474 676550 345476
rect 676815 345473 676881 345476
rect 42498 345358 42558 345473
rect 676666 345326 676672 345390
rect 676736 345388 676742 345390
rect 677007 345388 677073 345391
rect 676736 345386 677073 345388
rect 676736 345330 677012 345386
rect 677068 345330 677073 345386
rect 676736 345328 677073 345330
rect 676736 345326 676742 345328
rect 677007 345325 677073 345328
rect 42927 344796 42993 344799
rect 42528 344794 42993 344796
rect 42528 344738 42932 344794
rect 42988 344738 42993 344794
rect 42528 344736 42993 344738
rect 42927 344733 42993 344736
rect 42498 344056 42558 344248
rect 43119 344056 43185 344059
rect 42498 344054 43185 344056
rect 42498 343998 43124 344054
rect 43180 343998 43185 344054
rect 42498 343996 43185 343998
rect 43119 343993 43185 343996
rect 43215 343760 43281 343763
rect 42528 343758 43281 343760
rect 42528 343702 43220 343758
rect 43276 343702 43281 343758
rect 42528 343700 43281 343702
rect 43215 343697 43281 343700
rect 58383 343168 58449 343171
rect 654447 343168 654513 343171
rect 58383 343166 64416 343168
rect 40386 343022 40446 343138
rect 58383 343110 58388 343166
rect 58444 343110 64416 343166
rect 58383 343108 64416 343110
rect 650208 343166 654513 343168
rect 650208 343110 654452 343166
rect 654508 343110 654513 343166
rect 650208 343108 654513 343110
rect 58383 343105 58449 343108
rect 654447 343105 654513 343108
rect 40378 342958 40384 343022
rect 40448 342958 40454 343022
rect 40570 342810 40576 342874
rect 40640 342810 40646 342874
rect 40578 342546 40638 342810
rect 40770 341838 40830 342102
rect 40762 341774 40768 341838
rect 40832 341774 40838 341838
rect 42927 341540 42993 341543
rect 42528 341538 42993 341540
rect 42528 341482 42932 341538
rect 42988 341482 42993 341538
rect 42528 341480 42993 341482
rect 42927 341477 42993 341480
rect 40962 340654 41022 340918
rect 40954 340590 40960 340654
rect 41024 340590 41030 340654
rect 41346 340210 41406 340474
rect 41338 340146 41344 340210
rect 41408 340146 41414 340210
rect 41538 339618 41598 339882
rect 41530 339554 41536 339618
rect 41600 339554 41606 339618
rect 41922 339027 41982 339290
rect 41871 339022 41982 339027
rect 41871 338966 41876 339022
rect 41932 338966 41982 339022
rect 41871 338964 41982 338966
rect 41871 338961 41937 338964
rect 42490 338962 42496 339026
rect 42560 339024 42566 339026
rect 42874 339024 42880 339026
rect 42560 338964 42880 339024
rect 42560 338962 42566 338964
rect 42874 338962 42880 338964
rect 42944 338962 42950 339026
rect 41154 338582 41214 338846
rect 41146 338518 41152 338582
rect 41216 338518 41222 338582
rect 43066 338284 43072 338286
rect 42528 338224 43072 338284
rect 43066 338222 43072 338224
rect 43136 338222 43142 338286
rect 40194 337399 40254 337662
rect 40143 337394 40254 337399
rect 40143 337338 40148 337394
rect 40204 337338 40254 337394
rect 40143 337336 40254 337338
rect 40143 337333 40209 337336
rect 40002 336955 40062 337218
rect 39951 336950 40062 336955
rect 39951 336894 39956 336950
rect 40012 336894 40062 336950
rect 39951 336892 40062 336894
rect 39951 336889 40017 336892
rect 40002 336363 40062 336626
rect 40002 336358 40113 336363
rect 40002 336302 40052 336358
rect 40108 336302 40113 336358
rect 40002 336300 40113 336302
rect 40047 336297 40113 336300
rect 40194 335771 40254 336034
rect 40194 335766 40305 335771
rect 40194 335710 40244 335766
rect 40300 335710 40305 335766
rect 40194 335708 40305 335710
rect 40239 335705 40305 335708
rect 39810 335179 39870 335590
rect 39810 335174 39921 335179
rect 39810 335118 39860 335174
rect 39916 335118 39921 335174
rect 39810 335116 39921 335118
rect 39855 335113 39921 335116
rect 43023 335028 43089 335031
rect 42528 335026 43089 335028
rect 42528 334970 43028 335026
rect 43084 334970 43089 335026
rect 42528 334968 43089 334970
rect 43023 334965 43089 334968
rect 675279 335030 675345 335031
rect 675279 335026 675328 335030
rect 675392 335028 675398 335030
rect 675279 334970 675284 335026
rect 675279 334966 675328 334970
rect 675392 334968 675436 335028
rect 675392 334966 675398 334968
rect 675279 334965 675345 334966
rect 42498 334140 42558 334406
rect 42498 334080 42750 334140
rect 35202 333551 35262 333888
rect 42690 333696 42750 334080
rect 675471 333846 675537 333847
rect 675471 333844 675520 333846
rect 675428 333842 675520 333844
rect 675428 333786 675476 333842
rect 675428 333784 675520 333786
rect 675471 333782 675520 333784
rect 675584 333782 675590 333846
rect 675471 333781 675537 333782
rect 35151 333546 35262 333551
rect 35151 333490 35156 333546
rect 35212 333490 35262 333546
rect 35151 333488 35262 333490
rect 42498 333636 42750 333696
rect 35151 333485 35217 333488
rect 42498 333400 42558 333636
rect 42831 333400 42897 333403
rect 42498 333398 42897 333400
rect 42498 333370 42836 333398
rect 42528 333342 42836 333370
rect 42892 333342 42897 333398
rect 42528 333340 42897 333342
rect 42831 333337 42897 333340
rect 35151 333104 35217 333107
rect 35151 333102 35262 333104
rect 35151 333046 35156 333102
rect 35212 333046 35262 333102
rect 35151 333041 35262 333046
rect 35202 332778 35262 333041
rect 31956 331648 45488 331678
rect 31956 330486 32020 331648
rect 32604 331636 45488 331648
rect 32604 330504 44906 331636
rect 45450 330504 45488 331636
rect 654447 331624 654513 331627
rect 650208 331622 654513 331624
rect 650208 331566 654452 331622
rect 654508 331566 654513 331622
rect 650208 331564 654513 331566
rect 654447 331561 654513 331564
rect 675759 330588 675825 330591
rect 676474 330588 676480 330590
rect 675759 330586 676480 330588
rect 675759 330530 675764 330586
rect 675820 330530 676480 330586
rect 675759 330528 676480 330530
rect 675759 330525 675825 330528
rect 676474 330526 676480 330528
rect 676544 330526 676550 330590
rect 32604 330486 45488 330504
rect 31956 330458 45488 330486
rect 40143 329848 40209 329851
rect 42298 329848 42304 329850
rect 40143 329846 42304 329848
rect 40143 329790 40148 329846
rect 40204 329790 42304 329846
rect 40143 329788 42304 329790
rect 40143 329785 40209 329788
rect 42298 329786 42304 329788
rect 42368 329786 42374 329850
rect 675183 329552 675249 329555
rect 675322 329552 675328 329554
rect 675183 329550 675328 329552
rect 675183 329494 675188 329550
rect 675244 329494 675328 329550
rect 675183 329492 675328 329494
rect 675183 329489 675249 329492
rect 675322 329490 675328 329492
rect 675392 329490 675398 329554
rect 57807 328812 57873 328815
rect 57807 328810 64416 328812
rect 57807 328754 57812 328810
rect 57868 328754 64416 328810
rect 57807 328752 64416 328754
rect 57807 328749 57873 328752
rect 673978 328306 673984 328370
rect 674048 328368 674054 328370
rect 675375 328368 675441 328371
rect 674048 328366 675441 328368
rect 674048 328310 675380 328366
rect 675436 328310 675441 328366
rect 674048 328308 675441 328310
rect 674048 328306 674054 328308
rect 675375 328305 675441 328308
rect 675759 326888 675825 326891
rect 676666 326888 676672 326890
rect 675759 326886 676672 326888
rect 675759 326830 675764 326886
rect 675820 326830 676672 326886
rect 675759 326828 676672 326830
rect 675759 326825 675825 326828
rect 676666 326826 676672 326828
rect 676736 326826 676742 326890
rect 42351 326592 42417 326595
rect 42490 326592 42496 326594
rect 42351 326590 42496 326592
rect 42351 326534 42356 326590
rect 42412 326534 42496 326590
rect 42351 326532 42496 326534
rect 42351 326529 42417 326532
rect 42490 326530 42496 326532
rect 42560 326530 42566 326594
rect 671682 324236 699295 324237
rect 671677 323144 671683 324236
rect 672775 323144 699295 324236
rect 671682 323143 699295 323144
rect 700389 323143 711573 324237
rect 666066 322605 709502 322606
rect 41914 322534 41920 322598
rect 41984 322596 41990 322598
rect 42874 322596 42880 322598
rect 41984 322536 42880 322596
rect 41984 322534 41990 322536
rect 42874 322534 42880 322536
rect 42944 322534 42950 322598
rect 666061 321423 666067 322605
rect 667249 321423 709502 322605
rect 666066 321422 709502 321423
rect 710686 321422 711466 322606
rect 42447 320970 42513 320971
rect 42447 320968 42496 320970
rect 42404 320966 42496 320968
rect 42404 320910 42452 320966
rect 42404 320908 42496 320910
rect 42447 320906 42496 320908
rect 42560 320906 42566 320970
rect 42447 320905 42513 320906
rect 662178 320471 700628 320472
rect 41530 319722 41536 319786
rect 41600 319784 41606 319786
rect 41775 319784 41841 319787
rect 655119 319784 655185 319787
rect 41600 319782 41841 319784
rect 41600 319726 41780 319782
rect 41836 319726 41841 319782
rect 41600 319724 41841 319726
rect 650208 319782 655185 319784
rect 650208 319726 655124 319782
rect 655180 319726 655185 319782
rect 650208 319724 655185 319726
rect 41600 319722 41606 319724
rect 41775 319721 41841 319724
rect 655119 319721 655185 319724
rect 662173 319289 662179 320471
rect 663361 319289 700628 320471
rect 662178 319288 700628 319289
rect 701812 319288 711110 320472
rect 41967 318750 42033 318751
rect 41914 318686 41920 318750
rect 41984 318748 42033 318750
rect 41984 318746 42076 318748
rect 42028 318690 42076 318746
rect 41984 318688 42076 318690
rect 41984 318686 42033 318688
rect 41967 318685 42033 318686
rect 659368 318185 707920 318186
rect 41967 317862 42033 317863
rect 41914 317798 41920 317862
rect 41984 317860 42033 317862
rect 41984 317858 42076 317860
rect 42028 317802 42076 317858
rect 41984 317800 42076 317802
rect 41984 317798 42033 317800
rect 41967 317797 42033 317798
rect 42106 317058 42112 317122
rect 42176 317120 42182 317122
rect 43066 317120 43072 317122
rect 42176 317060 43072 317120
rect 42176 317058 42182 317060
rect 43066 317058 43072 317060
rect 43136 317058 43142 317122
rect 659363 317003 659369 318185
rect 660551 317003 707920 318185
rect 659368 317002 707920 317003
rect 709104 317002 711668 318186
rect 42063 316676 42129 316679
rect 42298 316676 42304 316678
rect 42063 316674 42304 316676
rect 42063 316618 42068 316674
rect 42124 316618 42304 316674
rect 42063 316616 42304 316618
rect 42063 316613 42129 316616
rect 42298 316614 42304 316616
rect 42368 316614 42374 316678
rect 42063 316086 42129 316087
rect 42063 316082 42112 316086
rect 42176 316084 42182 316086
rect 42063 316026 42068 316082
rect 42063 316022 42112 316026
rect 42176 316024 42220 316084
rect 42176 316022 42182 316024
rect 42063 316021 42129 316022
rect 41338 315430 41344 315494
rect 41408 315492 41414 315494
rect 41775 315492 41841 315495
rect 41408 315490 41841 315492
rect 41408 315434 41780 315490
rect 41836 315434 41841 315490
rect 41408 315432 41841 315434
rect 41408 315430 41414 315432
rect 41775 315429 41841 315432
rect 674415 315048 674481 315051
rect 674415 315046 674784 315048
rect 674415 314990 674420 315046
rect 674476 314990 674784 315046
rect 674415 314988 674784 314990
rect 674415 314985 674481 314988
rect 674703 314752 674769 314755
rect 674703 314750 674814 314752
rect 674703 314694 674708 314750
rect 674764 314694 674814 314750
rect 674703 314689 674814 314694
rect 57999 314604 58065 314607
rect 57999 314602 64416 314604
rect 57999 314546 58004 314602
rect 58060 314546 64416 314602
rect 674754 314574 674814 314689
rect 57999 314544 64416 314546
rect 57999 314541 58065 314544
rect 674415 314012 674481 314015
rect 674415 314010 674784 314012
rect 674415 313954 674420 314010
rect 674476 313954 674784 314010
rect 674415 313952 674784 313954
rect 674415 313949 674481 313952
rect 40762 313654 40768 313718
rect 40832 313716 40838 313718
rect 41871 313716 41937 313719
rect 40832 313714 41937 313716
rect 40832 313658 41876 313714
rect 41932 313658 41937 313714
rect 40832 313656 41937 313658
rect 40832 313654 40838 313656
rect 41871 313653 41937 313656
rect 676858 313654 676864 313718
rect 676928 313654 676934 313718
rect 676866 313390 676926 313654
rect 41146 313210 41152 313274
rect 41216 313272 41222 313274
rect 41775 313272 41841 313275
rect 41216 313270 41841 313272
rect 41216 313214 41780 313270
rect 41836 313214 41841 313270
rect 41216 313212 41841 313214
rect 41216 313210 41222 313212
rect 41775 313209 41841 313212
rect 677250 312534 677310 312946
rect 677242 312470 677248 312534
rect 677312 312470 677318 312534
rect 40954 312322 40960 312386
rect 41024 312384 41030 312386
rect 41775 312384 41841 312387
rect 41024 312382 41841 312384
rect 41024 312326 41780 312382
rect 41836 312326 41841 312382
rect 41024 312324 41841 312326
rect 41024 312322 41030 312324
rect 41775 312321 41841 312324
rect 677058 312090 677118 312354
rect 677050 312026 677056 312090
rect 677120 312026 677126 312090
rect 677434 312026 677440 312090
rect 677504 312026 677510 312090
rect 677442 311792 677502 312026
rect 676896 311762 677502 311792
rect 676866 311732 677472 311762
rect 676866 311498 676926 311732
rect 676858 311434 676864 311498
rect 676928 311434 676934 311498
rect 673935 311348 674001 311351
rect 673935 311346 674784 311348
rect 673935 311290 673940 311346
rect 673996 311290 674784 311346
rect 673935 311288 674784 311290
rect 673935 311285 674001 311288
rect 673978 310694 673984 310758
rect 674048 310756 674054 310758
rect 674048 310696 674784 310756
rect 674048 310694 674054 310696
rect 674754 310019 674814 310134
rect 674703 310014 674814 310019
rect 674703 309958 674708 310014
rect 674764 309958 674814 310014
rect 674703 309956 674814 309958
rect 674703 309953 674769 309956
rect 6176 309136 8738 309936
rect 9538 309935 50926 309936
rect 9538 309137 50127 309935
rect 50925 309137 50931 309935
rect 674319 309646 674385 309649
rect 674319 309644 674784 309646
rect 674319 309588 674324 309644
rect 674380 309588 674784 309644
rect 674319 309586 674784 309588
rect 674319 309583 674385 309586
rect 9538 309136 50926 309137
rect 674946 308835 675006 309098
rect 674946 308830 675057 308835
rect 5914 307998 16328 308798
rect 17128 308797 52718 308798
rect 17128 307999 51919 308797
rect 52717 307999 52723 308797
rect 674946 308774 674996 308830
rect 675052 308774 675057 308830
rect 674946 308772 675057 308774
rect 674991 308769 675057 308772
rect 677058 308243 677118 308506
rect 677007 308238 677118 308243
rect 677007 308182 677012 308238
rect 677068 308182 677118 308238
rect 677007 308180 677118 308182
rect 677007 308177 677073 308180
rect 17128 307998 52718 307999
rect 655311 307944 655377 307947
rect 650208 307942 655377 307944
rect 650208 307886 655316 307942
rect 655372 307886 655377 307942
rect 650208 307884 655377 307886
rect 655311 307881 655377 307884
rect 674946 307799 675006 307988
rect 674895 307794 675006 307799
rect 674895 307738 674900 307794
rect 674956 307738 675006 307794
rect 674895 307736 675006 307738
rect 674895 307733 674961 307736
rect 675138 307207 675198 307470
rect 675087 307202 675198 307207
rect 675087 307146 675092 307202
rect 675148 307146 675198 307202
rect 675087 307144 675198 307146
rect 675087 307141 675153 307144
rect 6002 306336 7378 307136
rect 8178 307135 54502 307136
rect 8178 306337 53703 307135
rect 54501 306337 54507 307135
rect 674754 306763 674814 306878
rect 674754 306758 674865 306763
rect 674754 306702 674804 306758
rect 674860 306702 674865 306758
rect 674754 306700 674865 306702
rect 674799 306697 674865 306700
rect 8178 306336 54502 306337
rect 676866 306023 676926 306360
rect 676866 306018 676977 306023
rect 676866 305962 676916 306018
rect 676972 305962 676977 306018
rect 676866 305960 676977 305962
rect 676911 305957 676977 305960
rect 674031 305872 674097 305875
rect 674031 305870 674784 305872
rect 674031 305814 674036 305870
rect 674092 305814 674784 305870
rect 674031 305812 674784 305814
rect 674031 305809 674097 305812
rect 6176 304848 17732 305648
rect 18532 305647 56068 305648
rect 18532 304849 55269 305647
rect 56067 304849 56073 305647
rect 674607 305132 674673 305135
rect 674754 305132 674814 305250
rect 674607 305130 674814 305132
rect 674607 305074 674612 305130
rect 674668 305074 674814 305130
rect 674607 305072 674814 305074
rect 674607 305069 674673 305072
rect 18532 304848 56068 304849
rect 674511 304540 674577 304543
rect 674754 304540 674814 304732
rect 674511 304538 674814 304540
rect 674511 304482 674516 304538
rect 674572 304482 674814 304538
rect 674511 304480 674814 304482
rect 674511 304477 674577 304480
rect 674223 304244 674289 304247
rect 674223 304242 674784 304244
rect 674223 304186 674228 304242
rect 674284 304186 674784 304242
rect 674223 304184 674784 304186
rect 674223 304181 674289 304184
rect 674415 303652 674481 303655
rect 674415 303650 674784 303652
rect 674415 303594 674420 303650
rect 674476 303594 674784 303650
rect 674415 303592 674784 303594
rect 674415 303589 674481 303592
rect 42543 302912 42609 302915
rect 42498 302910 42609 302912
rect 42498 302854 42548 302910
rect 42604 302854 42609 302910
rect 42498 302849 42609 302854
rect 42498 302660 42558 302849
rect 676866 302767 676926 303104
rect 676815 302762 676926 302767
rect 676815 302706 676820 302762
rect 676876 302706 676926 302762
rect 676815 302704 676926 302706
rect 676815 302701 676881 302704
rect 674415 302616 674481 302619
rect 674415 302614 674784 302616
rect 674415 302558 674420 302614
rect 674476 302558 674784 302614
rect 674415 302556 674784 302558
rect 674415 302553 674481 302556
rect 42543 302320 42609 302323
rect 42498 302318 42609 302320
rect 42498 302262 42548 302318
rect 42604 302262 42609 302318
rect 42498 302257 42609 302262
rect 676815 302320 676881 302323
rect 676815 302318 676926 302320
rect 676815 302262 676820 302318
rect 676876 302262 676926 302318
rect 676815 302257 676926 302262
rect 42498 302142 42558 302257
rect 676866 301994 676926 302257
rect 42543 301876 42609 301879
rect 42498 301874 42609 301876
rect 42498 301818 42548 301874
rect 42604 301818 42609 301874
rect 42498 301813 42609 301818
rect 42498 301550 42558 301813
rect 42498 300988 42558 301032
rect 43311 300988 43377 300991
rect 42498 300986 43377 300988
rect 42498 300930 43316 300986
rect 43372 300930 43377 300986
rect 42498 300928 43377 300930
rect 43311 300925 43377 300928
rect 43215 300544 43281 300547
rect 42528 300542 43281 300544
rect 42528 300486 43220 300542
rect 43276 300486 43281 300542
rect 42528 300484 43281 300486
rect 43215 300481 43281 300484
rect 59439 300100 59505 300103
rect 59439 300098 64416 300100
rect 59439 300042 59444 300098
rect 59500 300042 64416 300098
rect 59439 300040 64416 300042
rect 59439 300037 59505 300040
rect 40386 299806 40446 299922
rect 40378 299742 40384 299806
rect 40448 299742 40454 299806
rect 40570 299594 40576 299658
rect 40640 299656 40646 299658
rect 42298 299656 42304 299658
rect 40640 299596 42304 299656
rect 40640 299594 40646 299596
rect 42298 299594 42304 299596
rect 42368 299594 42374 299658
rect 42306 299404 42366 299594
rect 675898 299446 675904 299510
rect 675968 299508 675974 299510
rect 676911 299508 676977 299511
rect 675968 299506 676977 299508
rect 675968 299450 676916 299506
rect 676972 299450 676977 299506
rect 675968 299448 676977 299450
rect 675968 299446 675974 299448
rect 676911 299445 676977 299448
rect 676666 299298 676672 299362
rect 676736 299360 676742 299362
rect 677007 299360 677073 299363
rect 676736 299358 677073 299360
rect 676736 299302 677012 299358
rect 677068 299302 677073 299358
rect 676736 299300 677073 299302
rect 676736 299298 676742 299300
rect 677007 299297 677073 299300
rect 40770 298622 40830 298886
rect 40762 298558 40768 298622
rect 40832 298558 40838 298622
rect 41154 298031 41214 298294
rect 41154 298026 41265 298031
rect 41154 297970 41204 298026
rect 41260 297970 41265 298026
rect 41154 297968 41265 297970
rect 41199 297965 41265 297968
rect 40962 297438 41022 297776
rect 40954 297374 40960 297438
rect 41024 297374 41030 297438
rect 41346 296994 41406 297258
rect 41338 296930 41344 296994
rect 41408 296930 41414 296994
rect 41538 296550 41598 296666
rect 41530 296486 41536 296550
rect 41600 296486 41606 296550
rect 654543 296252 654609 296255
rect 650208 296250 654609 296252
rect 650208 296194 654548 296250
rect 654604 296194 654609 296250
rect 650208 296192 654609 296194
rect 654543 296189 654609 296192
rect 41922 295811 41982 296148
rect 41922 295806 42033 295811
rect 41922 295750 41972 295806
rect 42028 295750 42033 295806
rect 41922 295748 42033 295750
rect 41967 295745 42033 295748
rect 41154 295366 41214 295630
rect 41146 295302 41152 295366
rect 41216 295302 41222 295366
rect 42114 294922 42174 295038
rect 42106 294858 42112 294922
rect 42176 294858 42182 294922
rect 40194 294183 40254 294520
rect 40194 294178 40305 294183
rect 40194 294122 40244 294178
rect 40300 294122 40305 294178
rect 40194 294120 40305 294122
rect 40239 294117 40305 294120
rect 40194 293739 40254 294002
rect 40143 293734 40254 293739
rect 40143 293678 40148 293734
rect 40204 293678 40254 293734
rect 40143 293676 40254 293678
rect 40143 293673 40209 293676
rect 42682 293440 42688 293442
rect 42528 293380 42688 293440
rect 42682 293378 42688 293380
rect 42752 293378 42758 293442
rect 39810 292555 39870 292818
rect 39810 292550 39921 292555
rect 39810 292494 39860 292550
rect 39916 292494 39921 292550
rect 39810 292492 39921 292494
rect 39855 292489 39921 292492
rect 40002 292111 40062 292374
rect 40002 292106 40113 292111
rect 40002 292050 40052 292106
rect 40108 292050 40113 292106
rect 40002 292048 40113 292050
rect 40047 292045 40113 292048
rect 42927 291812 42993 291815
rect 42528 291810 42993 291812
rect 42528 291754 42932 291810
rect 42988 291754 42993 291810
rect 42528 291752 42993 291754
rect 42927 291749 42993 291752
rect 42498 290924 42558 291190
rect 42498 290864 42750 290924
rect 35202 290483 35262 290746
rect 35151 290478 35262 290483
rect 42690 290480 42750 290864
rect 35151 290422 35156 290478
rect 35212 290422 35262 290478
rect 35151 290420 35262 290422
rect 42498 290420 42750 290480
rect 35151 290417 35217 290420
rect 42498 289891 42558 290420
rect 675279 290038 675345 290039
rect 675279 290034 675328 290038
rect 675392 290036 675398 290038
rect 675279 289978 675284 290034
rect 675279 289974 675328 289978
rect 675392 289976 675436 290036
rect 675392 289974 675398 289976
rect 675279 289973 675345 289974
rect 35151 289888 35217 289891
rect 35151 289886 35262 289888
rect 35151 289830 35156 289886
rect 35212 289830 35262 289886
rect 35151 289825 35262 289830
rect 42498 289886 42609 289891
rect 42498 289830 42548 289886
rect 42604 289830 42609 289886
rect 42498 289828 42609 289830
rect 42543 289825 42609 289828
rect 35202 289562 35262 289825
rect 675471 289594 675537 289595
rect 675471 289590 675520 289594
rect 675584 289592 675590 289594
rect 675471 289534 675476 289590
rect 675471 289530 675520 289534
rect 675584 289532 675628 289592
rect 675584 289530 675590 289532
rect 675471 289529 675537 289530
rect 36308 287744 47008 287772
rect 36308 286660 36346 287744
rect 36976 287742 47008 287744
rect 36976 286664 46158 287742
rect 46718 286664 47008 287742
rect 36976 286660 47008 286664
rect 36308 286640 47008 286660
rect 58095 285892 58161 285895
rect 58095 285890 64416 285892
rect 58095 285834 58100 285890
rect 58156 285834 64416 285890
rect 58095 285832 64416 285834
rect 58095 285829 58161 285832
rect 41914 285534 41920 285598
rect 41984 285596 41990 285598
rect 42490 285596 42496 285598
rect 41984 285536 42496 285596
rect 41984 285534 41990 285536
rect 42490 285534 42496 285536
rect 42560 285534 42566 285598
rect 40239 285152 40305 285155
rect 41722 285152 41728 285154
rect 40239 285150 41728 285152
rect 40239 285094 40244 285150
rect 40300 285094 41728 285150
rect 40239 285092 41728 285094
rect 40239 285089 40305 285092
rect 41722 285090 41728 285092
rect 41792 285090 41798 285154
rect 674554 284942 674560 285006
rect 674624 285004 674630 285006
rect 675183 285004 675249 285007
rect 674624 285002 675249 285004
rect 674624 284946 675188 285002
rect 675244 284946 675249 285002
rect 674624 284944 675249 284946
rect 674624 284942 674630 284944
rect 675183 284941 675249 284944
rect 674362 284794 674368 284858
rect 674432 284856 674438 284858
rect 675087 284856 675153 284859
rect 674432 284854 675153 284856
rect 674432 284798 675092 284854
rect 675148 284798 675153 284854
rect 674432 284796 675153 284798
rect 674432 284794 674438 284796
rect 675087 284793 675153 284796
rect 675759 284856 675825 284859
rect 675898 284856 675904 284858
rect 675759 284854 675904 284856
rect 675759 284798 675764 284854
rect 675820 284798 675904 284854
rect 675759 284796 675904 284798
rect 675759 284793 675825 284796
rect 675898 284794 675904 284796
rect 675968 284794 675974 284858
rect 654063 284708 654129 284711
rect 650208 284706 654129 284708
rect 650208 284650 654068 284706
rect 654124 284650 654129 284706
rect 650208 284648 654129 284650
rect 654063 284645 654129 284648
rect 673978 283610 673984 283674
rect 674048 283672 674054 283674
rect 675375 283672 675441 283675
rect 674048 283670 675441 283672
rect 674048 283614 675380 283670
rect 675436 283614 675441 283670
rect 674048 283612 675441 283614
rect 674048 283610 674054 283612
rect 675375 283609 675441 283612
rect 675759 281896 675825 281899
rect 676666 281896 676672 281898
rect 675759 281894 676672 281896
rect 675759 281838 675764 281894
rect 675820 281838 676672 281894
rect 675759 281836 676672 281838
rect 675759 281833 675825 281836
rect 676666 281834 676672 281836
rect 676736 281834 676742 281898
rect 671682 279568 699329 279569
rect 373167 278640 373233 278643
rect 204546 278638 373233 278640
rect 204546 278582 373172 278638
rect 373228 278582 373233 278638
rect 204546 278580 373233 278582
rect 204546 278495 204606 278580
rect 373167 278577 373233 278580
rect 373359 278640 373425 278643
rect 384015 278640 384081 278643
rect 373359 278638 384081 278640
rect 373359 278582 373364 278638
rect 373420 278582 384020 278638
rect 384076 278582 384081 278638
rect 373359 278580 384081 278582
rect 373359 278577 373425 278580
rect 384015 278577 384081 278580
rect 204495 278490 204606 278495
rect 204495 278434 204500 278490
rect 204556 278434 204606 278490
rect 204495 278432 204606 278434
rect 263727 278492 263793 278495
rect 598479 278492 598545 278495
rect 263727 278490 598545 278492
rect 263727 278434 263732 278490
rect 263788 278434 598484 278490
rect 598540 278434 598545 278490
rect 671677 278476 671683 279568
rect 672775 278476 699329 279568
rect 671682 278475 699329 278476
rect 700423 278475 711799 279569
rect 263727 278432 598545 278434
rect 204495 278429 204561 278432
rect 263727 278429 263793 278432
rect 598479 278429 598545 278432
rect 303375 278344 303441 278347
rect 467535 278344 467601 278347
rect 303375 278342 467601 278344
rect 303375 278286 303380 278342
rect 303436 278286 467540 278342
rect 467596 278286 467601 278342
rect 303375 278284 467601 278286
rect 303375 278281 303441 278284
rect 467535 278281 467601 278284
rect 304527 278196 304593 278199
rect 474735 278196 474801 278199
rect 304527 278194 474801 278196
rect 304527 278138 304532 278194
rect 304588 278138 474740 278194
rect 474796 278138 474801 278194
rect 304527 278136 474801 278138
rect 304527 278133 304593 278136
rect 474735 278133 474801 278136
rect 42159 278048 42225 278051
rect 42682 278048 42688 278050
rect 42159 278046 42688 278048
rect 42159 277990 42164 278046
rect 42220 277990 42688 278046
rect 42159 277988 42688 277990
rect 42159 277985 42225 277988
rect 42682 277986 42688 277988
rect 42752 277986 42758 278050
rect 317103 278048 317169 278051
rect 488943 278048 489009 278051
rect 317103 278046 489009 278048
rect 317103 277990 317108 278046
rect 317164 277990 488948 278046
rect 489004 277990 489009 278046
rect 666066 277999 709390 278000
rect 317103 277988 489009 277990
rect 317103 277985 317169 277988
rect 488943 277985 489009 277988
rect 305199 277900 305265 277903
rect 481839 277900 481905 277903
rect 305199 277898 481905 277900
rect 305199 277842 305204 277898
rect 305260 277842 481844 277898
rect 481900 277842 481905 277898
rect 305199 277840 481905 277842
rect 305199 277837 305265 277840
rect 481839 277837 481905 277840
rect 307119 277752 307185 277755
rect 496143 277752 496209 277755
rect 307119 277750 496209 277752
rect 307119 277694 307124 277750
rect 307180 277694 496148 277750
rect 496204 277694 496209 277750
rect 307119 277692 496209 277694
rect 307119 277689 307185 277692
rect 496143 277689 496209 277692
rect 308367 277604 308433 277607
rect 507087 277604 507153 277607
rect 308367 277602 507153 277604
rect 308367 277546 308372 277602
rect 308428 277546 507092 277602
rect 507148 277546 507153 277602
rect 308367 277544 507153 277546
rect 308367 277541 308433 277544
rect 507087 277541 507153 277544
rect 309519 277456 309585 277459
rect 517743 277456 517809 277459
rect 309519 277454 517809 277456
rect 309519 277398 309524 277454
rect 309580 277398 517748 277454
rect 517804 277398 517809 277454
rect 309519 277396 517809 277398
rect 309519 277393 309585 277396
rect 517743 277393 517809 277396
rect 310959 277308 311025 277311
rect 528495 277308 528561 277311
rect 310959 277306 528561 277308
rect 310959 277250 310964 277306
rect 311020 277250 528500 277306
rect 528556 277250 528561 277306
rect 310959 277248 528561 277250
rect 310959 277245 311025 277248
rect 528495 277245 528561 277248
rect 312399 277160 312465 277163
rect 539247 277160 539313 277163
rect 312399 277158 539313 277160
rect 312399 277102 312404 277158
rect 312460 277102 539252 277158
rect 539308 277102 539313 277158
rect 312399 277100 539313 277102
rect 312399 277097 312465 277100
rect 539247 277097 539313 277100
rect 309423 277012 309489 277015
rect 318351 277012 318417 277015
rect 309423 277010 318417 277012
rect 309423 276954 309428 277010
rect 309484 276954 318356 277010
rect 318412 276954 318417 277010
rect 309423 276952 318417 276954
rect 309423 276949 309489 276952
rect 318351 276949 318417 276952
rect 321423 277012 321489 277015
rect 617679 277012 617745 277015
rect 321423 277010 617745 277012
rect 321423 276954 321428 277010
rect 321484 276954 617684 277010
rect 617740 276954 617745 277010
rect 321423 276952 617745 276954
rect 321423 276949 321489 276952
rect 617679 276949 617745 276952
rect 309615 276864 309681 276867
rect 318447 276864 318513 276867
rect 309615 276862 318513 276864
rect 309615 276806 309620 276862
rect 309676 276806 318452 276862
rect 318508 276806 318513 276862
rect 309615 276804 318513 276806
rect 309615 276801 309681 276804
rect 318447 276801 318513 276804
rect 325071 276864 325137 276867
rect 642735 276864 642801 276867
rect 325071 276862 642801 276864
rect 325071 276806 325076 276862
rect 325132 276806 642740 276862
rect 642796 276806 642801 276862
rect 666061 276817 666067 277999
rect 667249 276817 709390 277999
rect 666066 276816 709390 276817
rect 710574 276816 711542 278000
rect 325071 276804 642801 276806
rect 325071 276801 325137 276804
rect 642735 276801 642801 276804
rect 114639 276716 114705 276719
rect 322095 276716 322161 276719
rect 114639 276714 322161 276716
rect 114639 276658 114644 276714
rect 114700 276658 322100 276714
rect 322156 276658 322161 276714
rect 114639 276656 322161 276658
rect 114639 276653 114705 276656
rect 322095 276653 322161 276656
rect 325551 276716 325617 276719
rect 646287 276716 646353 276719
rect 325551 276714 646353 276716
rect 325551 276658 325556 276714
rect 325612 276658 646292 276714
rect 646348 276658 646353 276714
rect 325551 276656 646353 276658
rect 325551 276653 325617 276656
rect 646287 276653 646353 276656
rect 41530 276506 41536 276570
rect 41600 276568 41606 276570
rect 41775 276568 41841 276571
rect 41600 276566 41841 276568
rect 41600 276510 41780 276566
rect 41836 276510 41841 276566
rect 41600 276508 41841 276510
rect 41600 276506 41606 276508
rect 41775 276505 41841 276508
rect 315087 276568 315153 276571
rect 373359 276568 373425 276571
rect 315087 276566 373425 276568
rect 315087 276510 315092 276566
rect 315148 276510 373364 276566
rect 373420 276510 373425 276566
rect 315087 276508 373425 276510
rect 315087 276505 315153 276508
rect 373359 276505 373425 276508
rect 373935 276568 374001 276571
rect 387855 276568 387921 276571
rect 373935 276566 387921 276568
rect 373935 276510 373940 276566
rect 373996 276510 387860 276566
rect 387916 276510 387921 276566
rect 373935 276508 387921 276510
rect 373935 276505 374001 276508
rect 387855 276505 387921 276508
rect 318639 276420 318705 276423
rect 592719 276420 592785 276423
rect 318639 276418 592785 276420
rect 318639 276362 318644 276418
rect 318700 276362 592724 276418
rect 592780 276362 592785 276418
rect 318639 276360 592785 276362
rect 318639 276357 318705 276360
rect 592719 276357 592785 276360
rect 673551 276420 673617 276423
rect 674554 276420 674560 276422
rect 673551 276418 674560 276420
rect 673551 276362 673556 276418
rect 673612 276362 674560 276418
rect 673551 276360 674560 276362
rect 673551 276357 673617 276360
rect 674554 276358 674560 276360
rect 674624 276358 674630 276422
rect 319599 276272 319665 276275
rect 599823 276272 599889 276275
rect 319599 276270 599889 276272
rect 319599 276214 319604 276270
rect 319660 276214 599828 276270
rect 599884 276214 599889 276270
rect 319599 276212 599889 276214
rect 319599 276209 319665 276212
rect 599823 276209 599889 276212
rect 320847 276124 320913 276127
rect 610575 276124 610641 276127
rect 320847 276122 610641 276124
rect 320847 276066 320852 276122
rect 320908 276066 610580 276122
rect 610636 276066 610641 276122
rect 320847 276064 610641 276066
rect 320847 276061 320913 276064
rect 610575 276061 610641 276064
rect 323919 275976 323985 275979
rect 624879 275976 624945 275979
rect 323919 275974 624945 275976
rect 323919 275918 323924 275974
rect 323980 275918 624884 275974
rect 624940 275918 624945 275974
rect 323919 275916 624945 275918
rect 323919 275913 323985 275916
rect 624879 275913 624945 275916
rect 328527 275828 328593 275831
rect 637935 275828 638001 275831
rect 328527 275826 638001 275828
rect 328527 275770 328532 275826
rect 328588 275770 637940 275826
rect 637996 275770 638001 275826
rect 328527 275768 638001 275770
rect 328527 275765 328593 275768
rect 637935 275765 638001 275768
rect 261615 275680 261681 275683
rect 580911 275680 580977 275683
rect 261615 275678 580977 275680
rect 261615 275622 261620 275678
rect 261676 275622 580916 275678
rect 580972 275622 580977 275678
rect 261615 275620 580977 275622
rect 261615 275617 261681 275620
rect 580911 275617 580977 275620
rect 41967 275534 42033 275535
rect 41914 275470 41920 275534
rect 41984 275532 42033 275534
rect 264399 275532 264465 275535
rect 602223 275532 602289 275535
rect 41984 275530 42076 275532
rect 42028 275474 42076 275530
rect 41984 275472 42076 275474
rect 264399 275530 602289 275532
rect 264399 275474 264404 275530
rect 264460 275474 602228 275530
rect 602284 275474 602289 275530
rect 264399 275472 602289 275474
rect 41984 275470 42033 275472
rect 41967 275469 42033 275470
rect 264399 275469 264465 275472
rect 602223 275469 602289 275472
rect 265935 275384 266001 275387
rect 616527 275384 616593 275387
rect 265935 275382 616593 275384
rect 265935 275326 265940 275382
rect 265996 275326 616532 275382
rect 616588 275326 616593 275382
rect 265935 275324 616593 275326
rect 265935 275321 266001 275324
rect 616527 275321 616593 275324
rect 267087 275236 267153 275239
rect 623631 275236 623697 275239
rect 267087 275234 623697 275236
rect 267087 275178 267092 275234
rect 267148 275178 623636 275234
rect 623692 275178 623697 275234
rect 662178 275227 700624 275228
rect 267087 275176 623697 275178
rect 267087 275173 267153 275176
rect 623631 275173 623697 275176
rect 267183 275088 267249 275091
rect 627279 275088 627345 275091
rect 267183 275086 627345 275088
rect 267183 275030 267188 275086
rect 267244 275030 627284 275086
rect 627340 275030 627345 275086
rect 267183 275028 627345 275030
rect 267183 275025 267249 275028
rect 627279 275025 627345 275028
rect 262863 274940 262929 274943
rect 369231 274940 369297 274943
rect 262863 274938 369297 274940
rect 262863 274882 262868 274938
rect 262924 274882 369236 274938
rect 369292 274882 369297 274938
rect 262863 274880 369297 274882
rect 262863 274877 262929 274880
rect 369231 274877 369297 274880
rect 377487 274940 377553 274943
rect 379023 274940 379089 274943
rect 377487 274938 379089 274940
rect 377487 274882 377492 274938
rect 377548 274882 379028 274938
rect 379084 274882 379089 274938
rect 377487 274880 379089 274882
rect 377487 274877 377553 274880
rect 379023 274877 379089 274880
rect 379407 274940 379473 274943
rect 379983 274940 380049 274943
rect 379407 274938 380049 274940
rect 379407 274882 379412 274938
rect 379468 274882 379988 274938
rect 380044 274882 380049 274938
rect 379407 274880 380049 274882
rect 379407 274877 379473 274880
rect 379983 274877 380049 274880
rect 380175 274940 380241 274943
rect 645135 274940 645201 274943
rect 380175 274938 645201 274940
rect 380175 274882 380180 274938
rect 380236 274882 645140 274938
rect 645196 274882 645201 274938
rect 380175 274880 645201 274882
rect 380175 274877 380241 274880
rect 645135 274877 645201 274880
rect 42159 274792 42225 274795
rect 42490 274792 42496 274794
rect 42159 274790 42496 274792
rect 42159 274734 42164 274790
rect 42220 274734 42496 274790
rect 42159 274732 42496 274734
rect 42159 274729 42225 274732
rect 42490 274730 42496 274732
rect 42560 274792 42566 274794
rect 43119 274792 43185 274795
rect 42560 274790 43185 274792
rect 42560 274734 43124 274790
rect 43180 274734 43185 274790
rect 42560 274732 43185 274734
rect 42560 274730 42566 274732
rect 43119 274729 43185 274732
rect 254127 274792 254193 274795
rect 520143 274792 520209 274795
rect 254127 274790 520209 274792
rect 254127 274734 254132 274790
rect 254188 274734 520148 274790
rect 520204 274734 520209 274790
rect 254127 274732 520209 274734
rect 254127 274729 254193 274732
rect 520143 274729 520209 274732
rect 253935 274644 254001 274647
rect 516591 274644 516657 274647
rect 253935 274642 516657 274644
rect 253935 274586 253940 274642
rect 253996 274586 516596 274642
rect 516652 274586 516657 274642
rect 253935 274584 516657 274586
rect 253935 274581 254001 274584
rect 516591 274581 516657 274584
rect 252399 274496 252465 274499
rect 505935 274496 506001 274499
rect 252399 274494 506001 274496
rect 252399 274438 252404 274494
rect 252460 274438 505940 274494
rect 505996 274438 506001 274494
rect 252399 274436 506001 274438
rect 252399 274433 252465 274436
rect 505935 274433 506001 274436
rect 251823 274348 251889 274351
rect 498831 274348 498897 274351
rect 251823 274346 498897 274348
rect 251823 274290 251828 274346
rect 251884 274290 498836 274346
rect 498892 274290 498897 274346
rect 251823 274288 498897 274290
rect 251823 274285 251889 274288
rect 498831 274285 498897 274288
rect 250671 274200 250737 274203
rect 491631 274200 491697 274203
rect 250671 274198 491697 274200
rect 250671 274142 250676 274198
rect 250732 274142 491636 274198
rect 491692 274142 491697 274198
rect 250671 274140 491697 274142
rect 250671 274137 250737 274140
rect 491631 274137 491697 274140
rect 263343 274052 263409 274055
rect 382959 274052 383025 274055
rect 263343 274050 383025 274052
rect 263343 273994 263348 274050
rect 263404 273994 382964 274050
rect 383020 273994 383025 274050
rect 263343 273992 383025 273994
rect 263343 273989 263409 273992
rect 382959 273989 383025 273992
rect 383151 274052 383217 274055
rect 388623 274052 388689 274055
rect 552303 274052 552369 274055
rect 383151 274050 388689 274052
rect 383151 273994 383156 274050
rect 383212 273994 388628 274050
rect 388684 273994 388689 274050
rect 383151 273992 388689 273994
rect 383151 273989 383217 273992
rect 388623 273989 388689 273992
rect 388818 274050 552369 274052
rect 388818 273994 552308 274050
rect 552364 273994 552369 274050
rect 662173 274045 662179 275227
rect 663361 274045 700624 275227
rect 662178 274044 700624 274045
rect 701808 274044 711240 275228
rect 388818 273992 552369 273994
rect 256815 273904 256881 273907
rect 378255 273904 378321 273907
rect 256815 273902 378321 273904
rect 256815 273846 256820 273902
rect 256876 273846 378260 273902
rect 378316 273846 378321 273902
rect 256815 273844 378321 273846
rect 256815 273841 256881 273844
rect 378255 273841 378321 273844
rect 378447 273904 378513 273907
rect 388818 273904 388878 273992
rect 552303 273989 552369 273992
rect 378447 273902 388878 273904
rect 378447 273846 378452 273902
rect 378508 273846 388878 273902
rect 378447 273844 388878 273846
rect 378447 273841 378513 273844
rect 198735 273756 198801 273759
rect 391407 273756 391473 273759
rect 198735 273754 391473 273756
rect 198735 273698 198740 273754
rect 198796 273698 391412 273754
rect 391468 273698 391473 273754
rect 198735 273696 391473 273698
rect 198735 273693 198801 273696
rect 391407 273693 391473 273696
rect 41775 273610 41841 273611
rect 41722 273608 41728 273610
rect 41684 273548 41728 273608
rect 41792 273606 41841 273610
rect 41836 273550 41841 273606
rect 41722 273546 41728 273548
rect 41792 273546 41841 273550
rect 41775 273545 41841 273546
rect 83631 273608 83697 273611
rect 374319 273608 374385 273611
rect 83631 273606 374385 273608
rect 83631 273550 83636 273606
rect 83692 273550 374324 273606
rect 374380 273550 374385 273606
rect 83631 273548 374385 273550
rect 83631 273545 83697 273548
rect 374319 273545 374385 273548
rect 374458 273546 374464 273610
rect 374528 273608 374534 273610
rect 382767 273608 382833 273611
rect 374528 273606 382833 273608
rect 374528 273550 382772 273606
rect 382828 273550 382833 273606
rect 374528 273548 382833 273550
rect 374528 273546 374534 273548
rect 382767 273545 382833 273548
rect 382959 273608 383025 273611
rect 397359 273608 397425 273611
rect 382959 273606 397425 273608
rect 382959 273550 382964 273606
rect 383020 273550 397364 273606
rect 397420 273550 397425 273606
rect 382959 273548 397425 273550
rect 382959 273545 383025 273548
rect 397359 273545 397425 273548
rect 88431 273460 88497 273463
rect 374127 273460 374193 273463
rect 377295 273460 377361 273463
rect 88431 273458 374193 273460
rect 88431 273402 88436 273458
rect 88492 273402 374132 273458
rect 374188 273402 374193 273458
rect 88431 273400 374193 273402
rect 88431 273397 88497 273400
rect 374127 273397 374193 273400
rect 374466 273458 377361 273460
rect 374466 273402 377300 273458
rect 377356 273402 377361 273458
rect 374466 273400 377361 273402
rect 86031 273312 86097 273315
rect 374466 273312 374526 273400
rect 377295 273397 377361 273400
rect 377487 273460 377553 273463
rect 377679 273460 377745 273463
rect 377487 273458 377745 273460
rect 377487 273402 377492 273458
rect 377548 273402 377684 273458
rect 377740 273402 377745 273458
rect 377487 273400 377745 273402
rect 377487 273397 377553 273400
rect 377679 273397 377745 273400
rect 378255 273460 378321 273463
rect 392847 273460 392913 273463
rect 378255 273458 392913 273460
rect 378255 273402 378260 273458
rect 378316 273402 392852 273458
rect 392908 273402 392913 273458
rect 378255 273400 392913 273402
rect 378255 273397 378321 273400
rect 392847 273397 392913 273400
rect 393135 273460 393201 273463
rect 409402 273460 409408 273462
rect 393135 273458 409408 273460
rect 393135 273402 393140 273458
rect 393196 273402 409408 273458
rect 393135 273400 409408 273402
rect 393135 273397 393201 273400
rect 409402 273398 409408 273400
rect 409472 273398 409478 273462
rect 86031 273310 374526 273312
rect 86031 273254 86036 273310
rect 86092 273254 374526 273310
rect 86031 273252 374526 273254
rect 374703 273312 374769 273315
rect 383823 273312 383889 273315
rect 374703 273310 383889 273312
rect 374703 273254 374708 273310
rect 374764 273254 383828 273310
rect 383884 273254 383889 273310
rect 374703 273252 383889 273254
rect 86031 273249 86097 273252
rect 374703 273249 374769 273252
rect 383823 273249 383889 273252
rect 384058 273250 384064 273314
rect 384128 273312 384134 273314
rect 388335 273312 388401 273315
rect 384128 273310 388401 273312
rect 384128 273254 388340 273310
rect 388396 273254 388401 273310
rect 384128 273252 388401 273254
rect 384128 273250 384134 273252
rect 388335 273249 388401 273252
rect 390831 273312 390897 273315
rect 409786 273312 409792 273314
rect 390831 273310 409792 273312
rect 390831 273254 390836 273310
rect 390892 273254 409792 273310
rect 390831 273252 409792 273254
rect 390831 273249 390897 273252
rect 409786 273250 409792 273252
rect 409856 273250 409862 273314
rect 74895 273164 74961 273167
rect 94863 273164 94929 273167
rect 74895 273162 94929 273164
rect 74895 273106 74900 273162
rect 74956 273106 94868 273162
rect 94924 273106 94929 273162
rect 74895 273104 94929 273106
rect 74895 273101 74961 273104
rect 94863 273101 94929 273104
rect 115215 273164 115281 273167
rect 135279 273164 135345 273167
rect 115215 273162 135345 273164
rect 115215 273106 115220 273162
rect 115276 273106 135284 273162
rect 135340 273106 135345 273162
rect 115215 273104 135345 273106
rect 115215 273101 115281 273104
rect 135279 273101 135345 273104
rect 156879 273164 156945 273167
rect 177039 273164 177105 273167
rect 156879 273162 177105 273164
rect 156879 273106 156884 273162
rect 156940 273106 177044 273162
rect 177100 273106 177105 273162
rect 156879 273104 177105 273106
rect 156879 273101 156945 273104
rect 177039 273101 177105 273104
rect 197199 273164 197265 273167
rect 217359 273164 217425 273167
rect 197199 273162 217425 273164
rect 197199 273106 197204 273162
rect 197260 273106 217364 273162
rect 217420 273106 217425 273162
rect 197199 273104 217425 273106
rect 197199 273101 197265 273104
rect 217359 273101 217425 273104
rect 259599 273164 259665 273167
rect 563055 273164 563121 273167
rect 259599 273162 563121 273164
rect 259599 273106 259604 273162
rect 259660 273106 563060 273162
rect 563116 273106 563121 273162
rect 659368 273109 707924 273110
rect 259599 273104 563121 273106
rect 259599 273101 259665 273104
rect 563055 273101 563121 273104
rect 42063 273018 42129 273019
rect 42063 273014 42112 273018
rect 42176 273016 42182 273018
rect 81327 273016 81393 273019
rect 374458 273016 374464 273018
rect 42063 272958 42068 273014
rect 42063 272954 42112 272958
rect 42176 272956 42220 273016
rect 81327 273014 374464 273016
rect 81327 272958 81332 273014
rect 81388 272958 374464 273014
rect 81327 272956 374464 272958
rect 42176 272954 42182 272956
rect 42063 272953 42129 272954
rect 81327 272953 81393 272956
rect 374458 272954 374464 272956
rect 374528 272954 374534 273018
rect 376527 273016 376593 273019
rect 374658 273014 376593 273016
rect 374658 272958 376532 273014
rect 376588 272958 376593 273014
rect 374658 272956 376593 272958
rect 78927 272868 78993 272871
rect 374658 272868 374718 272956
rect 376527 272953 376593 272956
rect 377295 273016 377361 273019
rect 380079 273016 380145 273019
rect 377295 273014 380145 273016
rect 377295 272958 377300 273014
rect 377356 272958 380084 273014
rect 380140 272958 380145 273014
rect 377295 272956 380145 272958
rect 377295 272953 377361 272956
rect 380079 272953 380145 272956
rect 380271 273016 380337 273019
rect 394479 273016 394545 273019
rect 380271 273014 394545 273016
rect 380271 272958 380276 273014
rect 380332 272958 394484 273014
rect 394540 272958 394545 273014
rect 380271 272956 394545 272958
rect 380271 272953 380337 272956
rect 394479 272953 394545 272956
rect 395631 273016 395697 273019
rect 408250 273016 408256 273018
rect 395631 273014 408256 273016
rect 395631 272958 395636 273014
rect 395692 272958 408256 273014
rect 395631 272956 408256 272958
rect 395631 272953 395697 272956
rect 408250 272954 408256 272956
rect 408320 272954 408326 273018
rect 381135 272868 381201 272871
rect 78927 272866 374718 272868
rect 78927 272810 78932 272866
rect 78988 272810 374718 272866
rect 78927 272808 374718 272810
rect 374850 272866 381201 272868
rect 374850 272810 381140 272866
rect 381196 272810 381201 272866
rect 374850 272808 381201 272810
rect 78927 272805 78993 272808
rect 70575 272720 70641 272723
rect 76335 272720 76401 272723
rect 70575 272718 76401 272720
rect 70575 272662 70580 272718
rect 70636 272662 76340 272718
rect 76396 272662 76401 272718
rect 70575 272660 76401 272662
rect 70575 272657 70641 272660
rect 76335 272657 76401 272660
rect 76527 272720 76593 272723
rect 374703 272720 374769 272723
rect 76527 272718 374769 272720
rect 76527 272662 76532 272718
rect 76588 272662 374708 272718
rect 374764 272662 374769 272718
rect 76527 272660 374769 272662
rect 76527 272657 76593 272660
rect 374703 272657 374769 272660
rect 94767 272572 94833 272575
rect 115311 272572 115377 272575
rect 94767 272570 115377 272572
rect 94767 272514 94772 272570
rect 94828 272514 115316 272570
rect 115372 272514 115377 272570
rect 94767 272512 115377 272514
rect 94767 272509 94833 272512
rect 115311 272509 115377 272512
rect 135226 272510 135232 272574
rect 135296 272572 135302 272574
rect 156975 272572 157041 272575
rect 135296 272570 157041 272572
rect 135296 272514 156980 272570
rect 157036 272514 157041 272570
rect 135296 272512 157041 272514
rect 135296 272510 135302 272512
rect 156975 272509 157041 272512
rect 177135 272572 177201 272575
rect 197391 272572 197457 272575
rect 177135 272570 197457 272572
rect 177135 272514 177140 272570
rect 177196 272514 197396 272570
rect 197452 272514 197457 272570
rect 177135 272512 197457 272514
rect 177135 272509 177201 272512
rect 197391 272509 197457 272512
rect 217455 272572 217521 272575
rect 349167 272572 349233 272575
rect 374850 272572 374910 272808
rect 381135 272805 381201 272808
rect 381327 272868 381393 272871
rect 383055 272868 383121 272871
rect 384879 272868 384945 272871
rect 385935 272868 386001 272871
rect 381327 272866 382590 272868
rect 381327 272810 381332 272866
rect 381388 272810 382590 272866
rect 381327 272808 382590 272810
rect 381327 272805 381393 272808
rect 382287 272720 382353 272723
rect 217455 272570 349233 272572
rect 217455 272514 217460 272570
rect 217516 272514 349172 272570
rect 349228 272514 349233 272570
rect 217455 272512 349233 272514
rect 217455 272509 217521 272512
rect 349167 272509 349233 272512
rect 349314 272512 374910 272572
rect 375426 272718 382353 272720
rect 375426 272662 382292 272718
rect 382348 272662 382353 272718
rect 375426 272660 382353 272662
rect 382530 272720 382590 272808
rect 383055 272866 384945 272868
rect 383055 272810 383060 272866
rect 383116 272810 384884 272866
rect 384940 272810 384945 272866
rect 383055 272808 384945 272810
rect 383055 272805 383121 272808
rect 384879 272805 384945 272808
rect 385026 272866 386001 272868
rect 385026 272810 385940 272866
rect 385996 272810 386001 272866
rect 385026 272808 386001 272810
rect 385026 272720 385086 272808
rect 385935 272805 386001 272808
rect 386607 272868 386673 272871
rect 410554 272868 410560 272870
rect 386607 272866 410560 272868
rect 386607 272810 386612 272866
rect 386668 272810 410560 272866
rect 386607 272808 410560 272810
rect 386607 272805 386673 272808
rect 410554 272806 410560 272808
rect 410624 272806 410630 272870
rect 382530 272660 385086 272720
rect 385359 272720 385425 272723
rect 395631 272720 395697 272723
rect 385359 272718 395697 272720
rect 385359 272662 385364 272718
rect 385420 272662 395636 272718
rect 395692 272662 395697 272718
rect 385359 272660 395697 272662
rect 69423 272424 69489 272427
rect 74895 272424 74961 272427
rect 69423 272422 74961 272424
rect 69423 272366 69428 272422
rect 69484 272366 74900 272422
rect 74956 272366 74961 272422
rect 69423 272364 74961 272366
rect 69423 272361 69489 272364
rect 74895 272361 74961 272364
rect 94863 272424 94929 272427
rect 115215 272424 115281 272427
rect 94863 272422 115281 272424
rect 94863 272366 94868 272422
rect 94924 272366 115220 272422
rect 115276 272366 115281 272422
rect 94863 272364 115281 272366
rect 94863 272361 94929 272364
rect 115215 272361 115281 272364
rect 135279 272424 135345 272427
rect 156879 272424 156945 272427
rect 135279 272422 156945 272424
rect 135279 272366 135284 272422
rect 135340 272366 156884 272422
rect 156940 272366 156945 272422
rect 135279 272364 156945 272366
rect 135279 272361 135345 272364
rect 156879 272361 156945 272364
rect 177039 272424 177105 272427
rect 197199 272424 197265 272427
rect 177039 272422 197265 272424
rect 177039 272366 177044 272422
rect 177100 272366 197204 272422
rect 197260 272366 197265 272422
rect 177039 272364 197265 272366
rect 177039 272361 177105 272364
rect 197199 272361 197265 272364
rect 217359 272424 217425 272427
rect 349314 272424 349374 272512
rect 217359 272422 349374 272424
rect 217359 272366 217364 272422
rect 217420 272366 349374 272422
rect 217359 272364 349374 272366
rect 349455 272424 349521 272427
rect 358287 272424 358353 272427
rect 349455 272422 358353 272424
rect 349455 272366 349460 272422
rect 349516 272366 358292 272422
rect 358348 272366 358353 272422
rect 349455 272364 358353 272366
rect 217359 272361 217425 272364
rect 349455 272361 349521 272364
rect 358287 272361 358353 272364
rect 358479 272424 358545 272427
rect 375426 272424 375486 272660
rect 382287 272657 382353 272660
rect 385359 272657 385425 272660
rect 395631 272657 395697 272660
rect 395823 272720 395889 272723
rect 409594 272720 409600 272722
rect 395823 272718 409600 272720
rect 395823 272662 395828 272718
rect 395884 272662 409600 272718
rect 395823 272660 409600 272662
rect 395823 272657 395889 272660
rect 409594 272658 409600 272660
rect 409664 272658 409670 272722
rect 375663 272572 375729 272575
rect 379599 272572 379665 272575
rect 375663 272570 379665 272572
rect 375663 272514 375668 272570
rect 375724 272514 379604 272570
rect 379660 272514 379665 272570
rect 375663 272512 379665 272514
rect 375663 272509 375729 272512
rect 379599 272509 379665 272512
rect 380175 272572 380241 272575
rect 394287 272572 394353 272575
rect 380175 272570 394353 272572
rect 380175 272514 380180 272570
rect 380236 272514 394292 272570
rect 394348 272514 394353 272570
rect 380175 272512 394353 272514
rect 380175 272509 380241 272512
rect 394287 272509 394353 272512
rect 394434 272512 408702 272572
rect 384111 272424 384177 272427
rect 390927 272424 390993 272427
rect 358479 272422 375486 272424
rect 358479 272366 358484 272422
rect 358540 272366 375486 272422
rect 358479 272364 375486 272366
rect 375810 272422 384177 272424
rect 375810 272366 384116 272422
rect 384172 272366 384177 272422
rect 375810 272364 384177 272366
rect 358479 272361 358545 272364
rect 41338 272214 41344 272278
rect 41408 272276 41414 272278
rect 41775 272276 41841 272279
rect 41408 272274 41841 272276
rect 41408 272218 41780 272274
rect 41836 272218 41841 272274
rect 41408 272216 41841 272218
rect 41408 272214 41414 272216
rect 41775 272213 41841 272216
rect 74127 272276 74193 272279
rect 375810 272276 375870 272364
rect 384111 272361 384177 272364
rect 386178 272422 390993 272424
rect 386178 272366 390932 272422
rect 390988 272366 390993 272422
rect 386178 272364 390993 272366
rect 74127 272274 375870 272276
rect 74127 272218 74132 272274
rect 74188 272218 375870 272274
rect 74127 272216 375870 272218
rect 376527 272276 376593 272279
rect 381807 272276 381873 272279
rect 376527 272274 381873 272276
rect 376527 272218 376532 272274
rect 376588 272218 381812 272274
rect 381868 272218 381873 272274
rect 376527 272216 381873 272218
rect 74127 272213 74193 272216
rect 376527 272213 376593 272216
rect 381807 272213 381873 272216
rect 383055 272276 383121 272279
rect 386178 272276 386238 272364
rect 390927 272361 390993 272364
rect 393999 272424 394065 272427
rect 394434 272424 394494 272512
rect 393999 272422 394494 272424
rect 393999 272366 394004 272422
rect 394060 272366 394494 272422
rect 393999 272364 394494 272366
rect 398415 272424 398481 272427
rect 398415 272422 408510 272424
rect 398415 272366 398420 272422
rect 398476 272366 408510 272422
rect 398415 272364 408510 272366
rect 393999 272361 394065 272364
rect 398415 272361 398481 272364
rect 383055 272274 386238 272276
rect 383055 272218 383060 272274
rect 383116 272218 386238 272274
rect 383055 272216 386238 272218
rect 400143 272276 400209 272279
rect 400143 272274 408318 272276
rect 400143 272218 400148 272274
rect 400204 272218 408318 272274
rect 400143 272216 408318 272218
rect 383055 272213 383121 272216
rect 400143 272213 400209 272216
rect 71727 272128 71793 272131
rect 358479 272128 358545 272131
rect 71727 272126 358545 272128
rect 71727 272070 71732 272126
rect 71788 272070 358484 272126
rect 358540 272070 358545 272126
rect 71727 272068 358545 272070
rect 71727 272065 71793 272068
rect 358479 272065 358545 272068
rect 358671 272128 358737 272131
rect 375183 272128 375249 272131
rect 378159 272128 378225 272131
rect 358671 272126 375102 272128
rect 358671 272070 358676 272126
rect 358732 272070 375102 272126
rect 358671 272068 375102 272070
rect 358671 272065 358737 272068
rect 90831 271980 90897 271983
rect 374895 271980 374961 271983
rect 90831 271978 374961 271980
rect 90831 271922 90836 271978
rect 90892 271922 374900 271978
rect 374956 271922 374961 271978
rect 90831 271920 374961 271922
rect 375042 271980 375102 272068
rect 375183 272126 378225 272128
rect 375183 272070 375188 272126
rect 375244 272070 378164 272126
rect 378220 272070 378225 272126
rect 375183 272068 378225 272070
rect 375183 272065 375249 272068
rect 378159 272065 378225 272068
rect 378298 272066 378304 272130
rect 378368 272128 378374 272130
rect 379023 272128 379089 272131
rect 378368 272126 379089 272128
rect 378368 272070 379028 272126
rect 379084 272070 379089 272126
rect 378368 272068 379089 272070
rect 378368 272066 378374 272068
rect 379023 272065 379089 272068
rect 380271 272128 380337 272131
rect 394479 272128 394545 272131
rect 380271 272126 394545 272128
rect 380271 272070 380276 272126
rect 380332 272070 394484 272126
rect 394540 272070 394545 272126
rect 380271 272068 394545 272070
rect 380271 272065 380337 272068
rect 394479 272065 394545 272068
rect 402735 272128 402801 272131
rect 402735 272126 408126 272128
rect 402735 272070 402740 272126
rect 402796 272070 408126 272126
rect 402735 272068 408126 272070
rect 402735 272065 402801 272068
rect 381615 271980 381681 271983
rect 375042 271978 381681 271980
rect 375042 271922 381620 271978
rect 381676 271922 381681 271978
rect 375042 271920 381681 271922
rect 90831 271917 90897 271920
rect 374895 271917 374961 271920
rect 381615 271917 381681 271920
rect 381807 271980 381873 271983
rect 384399 271980 384465 271983
rect 381807 271978 384465 271980
rect 381807 271922 381812 271978
rect 381868 271922 384404 271978
rect 384460 271922 384465 271978
rect 381807 271920 384465 271922
rect 381807 271917 381873 271920
rect 384399 271917 384465 271920
rect 386319 271980 386385 271983
rect 396303 271980 396369 271983
rect 386319 271978 396369 271980
rect 386319 271922 386324 271978
rect 386380 271922 396308 271978
rect 396364 271922 396369 271978
rect 386319 271920 396369 271922
rect 386319 271917 386385 271920
rect 396303 271917 396369 271920
rect 401871 271980 401937 271983
rect 406671 271980 406737 271983
rect 401871 271978 406737 271980
rect 401871 271922 401876 271978
rect 401932 271922 406676 271978
rect 406732 271922 406737 271978
rect 401871 271920 406737 271922
rect 401871 271917 401937 271920
rect 406671 271917 406737 271920
rect 93231 271832 93297 271835
rect 160815 271832 160881 271835
rect 93231 271830 160881 271832
rect 93231 271774 93236 271830
rect 93292 271774 160820 271830
rect 160876 271774 160881 271830
rect 93231 271772 160881 271774
rect 93231 271769 93297 271772
rect 160815 271769 160881 271772
rect 161199 271832 161265 271835
rect 388143 271832 388209 271835
rect 161199 271830 388209 271832
rect 161199 271774 161204 271830
rect 161260 271774 388148 271830
rect 388204 271774 388209 271830
rect 161199 271772 388209 271774
rect 161199 271769 161265 271772
rect 388143 271769 388209 271772
rect 389103 271832 389169 271835
rect 407866 271832 407872 271834
rect 389103 271830 407872 271832
rect 389103 271774 389108 271830
rect 389164 271774 407872 271830
rect 389103 271772 407872 271774
rect 389103 271769 389169 271772
rect 407866 271770 407872 271772
rect 407936 271770 407942 271834
rect 76335 271684 76401 271687
rect 94767 271684 94833 271687
rect 76335 271682 94833 271684
rect 76335 271626 76340 271682
rect 76396 271626 94772 271682
rect 94828 271626 94833 271682
rect 76335 271624 94833 271626
rect 76335 271621 76401 271624
rect 94767 271621 94833 271624
rect 96783 271684 96849 271687
rect 100815 271684 100881 271687
rect 96783 271682 100881 271684
rect 96783 271626 96788 271682
rect 96844 271626 100820 271682
rect 100876 271626 100881 271682
rect 96783 271624 100881 271626
rect 96783 271621 96849 271624
rect 100815 271621 100881 271624
rect 120783 271684 120849 271687
rect 120975 271684 121041 271687
rect 120783 271682 121041 271684
rect 120783 271626 120788 271682
rect 120844 271626 120980 271682
rect 121036 271626 121041 271682
rect 120783 271624 121041 271626
rect 120783 271621 120849 271624
rect 120975 271621 121041 271624
rect 141039 271684 141105 271687
rect 141327 271684 141393 271687
rect 141039 271682 141393 271684
rect 141039 271626 141044 271682
rect 141100 271626 141332 271682
rect 141388 271626 141393 271682
rect 141039 271624 141393 271626
rect 141039 271621 141105 271624
rect 141327 271621 141393 271624
rect 161103 271684 161169 271687
rect 221775 271684 221841 271687
rect 161103 271682 221841 271684
rect 161103 271626 161108 271682
rect 161164 271626 221780 271682
rect 221836 271626 221841 271682
rect 161103 271624 221841 271626
rect 161103 271621 161169 271624
rect 221775 271621 221841 271624
rect 246159 271684 246225 271687
rect 262191 271684 262257 271687
rect 246159 271682 262257 271684
rect 246159 271626 246164 271682
rect 246220 271626 262196 271682
rect 262252 271626 262257 271682
rect 246159 271624 262257 271626
rect 246159 271621 246225 271624
rect 262191 271621 262257 271624
rect 282159 271684 282225 271687
rect 389295 271684 389361 271687
rect 282159 271682 389361 271684
rect 282159 271626 282164 271682
rect 282220 271626 389300 271682
rect 389356 271626 389361 271682
rect 282159 271624 389361 271626
rect 282159 271621 282225 271624
rect 389295 271621 389361 271624
rect 389679 271684 389745 271687
rect 406138 271684 406144 271686
rect 389679 271682 406144 271684
rect 389679 271626 389684 271682
rect 389740 271626 406144 271682
rect 389679 271624 406144 271626
rect 389679 271621 389745 271624
rect 406138 271622 406144 271624
rect 406208 271622 406214 271686
rect 100719 271536 100785 271539
rect 141135 271536 141201 271539
rect 100719 271534 141201 271536
rect 100719 271478 100724 271534
rect 100780 271478 141140 271534
rect 141196 271478 141201 271534
rect 100719 271476 141201 271478
rect 100719 271473 100785 271476
rect 141135 271473 141201 271476
rect 141615 271536 141681 271539
rect 241551 271536 241617 271539
rect 141615 271534 241617 271536
rect 141615 271478 141620 271534
rect 141676 271478 241556 271534
rect 241612 271478 241617 271534
rect 141615 271476 241617 271478
rect 141615 271473 141681 271476
rect 241551 271473 241617 271476
rect 242031 271536 242097 271539
rect 389871 271536 389937 271539
rect 242031 271534 389937 271536
rect 242031 271478 242036 271534
rect 242092 271478 389876 271534
rect 389932 271478 389937 271534
rect 242031 271476 389937 271478
rect 242031 271473 242097 271476
rect 389871 271473 389937 271476
rect 395151 271536 395217 271539
rect 407482 271536 407488 271538
rect 395151 271534 407488 271536
rect 395151 271478 395156 271534
rect 395212 271478 407488 271534
rect 395151 271476 407488 271478
rect 395151 271473 395217 271476
rect 407482 271474 407488 271476
rect 407552 271474 407558 271538
rect 408066 271536 408126 272068
rect 408258 271684 408318 272216
rect 408450 271980 408510 272364
rect 408642 272276 408702 272512
rect 410170 272276 410176 272278
rect 408642 272216 410176 272276
rect 410170 272214 410176 272216
rect 410240 272214 410246 272278
rect 410938 271980 410944 271982
rect 408450 271920 410944 271980
rect 410938 271918 410944 271920
rect 411008 271918 411014 271982
rect 659363 271927 659369 273109
rect 660551 271927 707924 273109
rect 659368 271926 707924 271927
rect 709108 271926 711038 273110
rect 411130 271684 411136 271686
rect 408258 271624 411136 271684
rect 411130 271622 411136 271624
rect 411200 271622 411206 271686
rect 411322 271536 411328 271538
rect 408066 271476 411328 271536
rect 411322 271474 411328 271476
rect 411392 271474 411398 271538
rect 72975 271388 73041 271391
rect 141135 271388 141201 271391
rect 72975 271386 141201 271388
rect 72975 271330 72980 271386
rect 73036 271330 141140 271386
rect 141196 271330 141201 271386
rect 72975 271328 141201 271330
rect 72975 271325 73041 271328
rect 141135 271325 141201 271328
rect 141615 271388 141681 271391
rect 241647 271388 241713 271391
rect 141615 271386 241713 271388
rect 141615 271330 141620 271386
rect 141676 271330 241652 271386
rect 241708 271330 241713 271386
rect 141615 271328 241713 271330
rect 141615 271325 141681 271328
rect 241647 271325 241713 271328
rect 241935 271388 242001 271391
rect 316527 271388 316593 271391
rect 241935 271386 316593 271388
rect 241935 271330 241940 271386
rect 241996 271330 316532 271386
rect 316588 271330 316593 271386
rect 241935 271328 316593 271330
rect 241935 271325 242001 271328
rect 316527 271325 316593 271328
rect 316719 271388 316785 271391
rect 328527 271388 328593 271391
rect 316719 271386 328593 271388
rect 316719 271330 316724 271386
rect 316780 271330 328532 271386
rect 328588 271330 328593 271386
rect 316719 271328 328593 271330
rect 316719 271325 316785 271328
rect 328527 271325 328593 271328
rect 334095 271388 334161 271391
rect 357039 271388 357105 271391
rect 334095 271386 357105 271388
rect 334095 271330 334100 271386
rect 334156 271330 357044 271386
rect 357100 271330 357105 271386
rect 334095 271328 357105 271330
rect 334095 271325 334161 271328
rect 357039 271325 357105 271328
rect 368655 271388 368721 271391
rect 559407 271388 559473 271391
rect 368655 271386 559473 271388
rect 368655 271330 368660 271386
rect 368716 271330 559412 271386
rect 559468 271330 559473 271386
rect 368655 271328 559473 271330
rect 368655 271325 368721 271328
rect 559407 271325 559473 271328
rect 82575 271240 82641 271243
rect 211695 271240 211761 271243
rect 82575 271238 211761 271240
rect 82575 271182 82580 271238
rect 82636 271182 211700 271238
rect 211756 271182 211761 271238
rect 82575 271180 211761 271182
rect 82575 271177 82641 271180
rect 211695 271177 211761 271180
rect 221775 271240 221841 271243
rect 246159 271240 246225 271243
rect 221775 271238 246225 271240
rect 221775 271182 221780 271238
rect 221836 271182 246164 271238
rect 246220 271182 246225 271238
rect 221775 271180 246225 271182
rect 221775 271177 221841 271180
rect 246159 271177 246225 271180
rect 265455 271240 265521 271243
rect 367119 271240 367185 271243
rect 265455 271238 367185 271240
rect 265455 271182 265460 271238
rect 265516 271182 367124 271238
rect 367180 271182 367185 271238
rect 265455 271180 367185 271182
rect 265455 271177 265521 271180
rect 367119 271177 367185 271180
rect 377295 271240 377361 271243
rect 377914 271240 377920 271242
rect 377295 271238 377920 271240
rect 377295 271182 377300 271238
rect 377356 271182 377920 271238
rect 377295 271180 377920 271182
rect 377295 271177 377361 271180
rect 377914 271178 377920 271180
rect 377984 271178 377990 271242
rect 378159 271240 378225 271243
rect 387759 271240 387825 271243
rect 378159 271238 387825 271240
rect 378159 271182 378164 271238
rect 378220 271182 387764 271238
rect 387820 271182 387825 271238
rect 378159 271180 387825 271182
rect 378159 271177 378225 271180
rect 387759 271177 387825 271180
rect 396879 271240 396945 271243
rect 406522 271240 406528 271242
rect 396879 271238 406528 271240
rect 396879 271182 396884 271238
rect 396940 271182 406528 271238
rect 396879 271180 406528 271182
rect 396879 271177 396945 271180
rect 406522 271178 406528 271180
rect 406592 271178 406598 271242
rect 406671 271240 406737 271243
rect 409210 271240 409216 271242
rect 406671 271238 409216 271240
rect 406671 271182 406676 271238
rect 406732 271182 409216 271238
rect 406671 271180 409216 271182
rect 406671 271177 406737 271180
rect 409210 271178 409216 271180
rect 409280 271178 409286 271242
rect 449295 271240 449361 271243
rect 449583 271240 449649 271243
rect 449295 271238 449649 271240
rect 449295 271182 449300 271238
rect 449356 271182 449588 271238
rect 449644 271182 449649 271238
rect 449295 271180 449649 271182
rect 449295 271177 449361 271180
rect 449583 271177 449649 271180
rect 480975 271240 481041 271243
rect 501039 271240 501105 271243
rect 480975 271238 501105 271240
rect 480975 271182 480980 271238
rect 481036 271182 501044 271238
rect 501100 271182 501105 271238
rect 480975 271180 501105 271182
rect 480975 271177 481041 271180
rect 501039 271177 501105 271180
rect 87183 271092 87249 271095
rect 212079 271092 212145 271095
rect 87183 271090 212145 271092
rect 87183 271034 87188 271090
rect 87244 271034 212084 271090
rect 212140 271034 212145 271090
rect 87183 271032 212145 271034
rect 87183 271029 87249 271032
rect 212079 271029 212145 271032
rect 259311 271092 259377 271095
rect 273519 271092 273585 271095
rect 259311 271090 273585 271092
rect 259311 271034 259316 271090
rect 259372 271034 273524 271090
rect 273580 271034 273585 271090
rect 259311 271032 273585 271034
rect 259311 271029 259377 271032
rect 273519 271029 273585 271032
rect 296751 271092 296817 271095
rect 316623 271092 316689 271095
rect 296751 271090 316689 271092
rect 296751 271034 296756 271090
rect 296812 271034 316628 271090
rect 316684 271034 316689 271090
rect 296751 271032 316689 271034
rect 296751 271029 296817 271032
rect 316623 271029 316689 271032
rect 319503 271092 319569 271095
rect 322383 271092 322449 271095
rect 319503 271090 322449 271092
rect 319503 271034 319508 271090
rect 319564 271034 322388 271090
rect 322444 271034 322449 271090
rect 319503 271032 322449 271034
rect 319503 271029 319569 271032
rect 322383 271029 322449 271032
rect 322575 271092 322641 271095
rect 332271 271092 332337 271095
rect 322575 271090 332337 271092
rect 322575 271034 322580 271090
rect 322636 271034 332276 271090
rect 332332 271034 332337 271090
rect 322575 271032 332337 271034
rect 322575 271029 322641 271032
rect 332271 271029 332337 271032
rect 367119 271092 367185 271095
rect 394479 271092 394545 271095
rect 367119 271090 394545 271092
rect 367119 271034 367124 271090
rect 367180 271034 394484 271090
rect 394540 271034 394545 271090
rect 367119 271032 394545 271034
rect 367119 271029 367185 271032
rect 394479 271029 394545 271032
rect 397743 271092 397809 271095
rect 406714 271092 406720 271094
rect 397743 271090 406720 271092
rect 397743 271034 397748 271090
rect 397804 271034 406720 271090
rect 397743 271032 406720 271034
rect 397743 271029 397809 271032
rect 406714 271030 406720 271032
rect 406784 271030 406790 271094
rect 452175 271092 452241 271095
rect 469455 271092 469521 271095
rect 452175 271090 469521 271092
rect 452175 271034 452180 271090
rect 452236 271034 469460 271090
rect 469516 271034 469521 271090
rect 452175 271032 469521 271034
rect 452175 271029 452241 271032
rect 469455 271029 469521 271032
rect 564495 271092 564561 271095
rect 584367 271092 584433 271095
rect 564495 271090 584433 271092
rect 564495 271034 564500 271090
rect 564556 271034 584372 271090
rect 584428 271034 584433 271090
rect 564495 271032 584433 271034
rect 564495 271029 564561 271032
rect 584367 271029 584433 271032
rect 77775 270944 77841 270947
rect 315087 270944 315153 270947
rect 77775 270942 315153 270944
rect 77775 270886 77780 270942
rect 77836 270886 315092 270942
rect 315148 270886 315153 270942
rect 77775 270884 315153 270886
rect 77775 270881 77841 270884
rect 315087 270881 315153 270884
rect 317487 270944 317553 270947
rect 328623 270944 328689 270947
rect 317487 270942 328689 270944
rect 317487 270886 317492 270942
rect 317548 270886 328628 270942
rect 328684 270886 328689 270942
rect 317487 270884 328689 270886
rect 317487 270881 317553 270884
rect 328623 270881 328689 270884
rect 348538 270882 348544 270946
rect 348608 270944 348614 270946
rect 368559 270944 368625 270947
rect 348608 270942 368625 270944
rect 348608 270886 368564 270942
rect 368620 270886 368625 270942
rect 348608 270884 368625 270886
rect 348608 270882 348614 270884
rect 368559 270881 368625 270884
rect 374319 270944 374385 270947
rect 391599 270944 391665 270947
rect 374319 270942 391665 270944
rect 374319 270886 374324 270942
rect 374380 270886 391604 270942
rect 391660 270886 391665 270942
rect 374319 270884 391665 270886
rect 374319 270881 374385 270884
rect 391599 270881 391665 270884
rect 391738 270882 391744 270946
rect 391808 270944 391814 270946
rect 392943 270944 393009 270947
rect 391808 270942 393009 270944
rect 391808 270886 392948 270942
rect 393004 270886 393009 270942
rect 391808 270884 393009 270886
rect 391808 270882 391814 270884
rect 392943 270881 393009 270884
rect 399471 270944 399537 270947
rect 406906 270944 406912 270946
rect 399471 270942 406912 270944
rect 399471 270886 399476 270942
rect 399532 270886 406912 270942
rect 399471 270884 406912 270886
rect 399471 270881 399537 270884
rect 406906 270882 406912 270884
rect 406976 270882 406982 270946
rect 428175 270944 428241 270947
rect 446319 270944 446385 270947
rect 428175 270942 446385 270944
rect 428175 270886 428180 270942
rect 428236 270886 446324 270942
rect 446380 270886 446385 270942
rect 428175 270884 446385 270886
rect 428175 270881 428241 270884
rect 446319 270881 446385 270884
rect 452175 270944 452241 270947
rect 452463 270944 452529 270947
rect 452175 270942 452529 270944
rect 452175 270886 452180 270942
rect 452236 270886 452468 270942
rect 452524 270886 452529 270942
rect 452175 270884 452529 270886
rect 452175 270881 452241 270884
rect 452463 270881 452529 270884
rect 115311 270796 115377 270799
rect 135226 270796 135232 270798
rect 115311 270794 135232 270796
rect 115311 270738 115316 270794
rect 115372 270738 135232 270794
rect 115311 270736 135232 270738
rect 115311 270733 115377 270736
rect 135226 270734 135232 270736
rect 135296 270734 135302 270798
rect 156975 270796 157041 270799
rect 177135 270796 177201 270799
rect 156975 270794 177201 270796
rect 156975 270738 156980 270794
rect 157036 270738 177140 270794
rect 177196 270738 177201 270794
rect 156975 270736 177201 270738
rect 156975 270733 157041 270736
rect 177135 270733 177201 270736
rect 197391 270796 197457 270799
rect 217455 270796 217521 270799
rect 197391 270794 217521 270796
rect 197391 270738 197396 270794
rect 197452 270738 217460 270794
rect 217516 270738 217521 270794
rect 197391 270736 217521 270738
rect 197391 270733 197457 270736
rect 217455 270733 217521 270736
rect 260655 270796 260721 270799
rect 394383 270796 394449 270799
rect 260655 270794 394449 270796
rect 260655 270738 260660 270794
rect 260716 270738 394388 270794
rect 394444 270738 394449 270794
rect 260655 270736 394449 270738
rect 260655 270733 260721 270736
rect 394383 270733 394449 270736
rect 401199 270796 401265 270799
rect 407674 270796 407680 270798
rect 401199 270794 407680 270796
rect 401199 270738 401204 270794
rect 401260 270738 407680 270794
rect 401199 270736 407680 270738
rect 401199 270733 401265 270736
rect 407674 270734 407680 270736
rect 407744 270734 407750 270798
rect 408975 270796 409041 270799
rect 419151 270796 419217 270799
rect 408975 270794 419217 270796
rect 408975 270738 408980 270794
rect 409036 270738 419156 270794
rect 419212 270738 419217 270794
rect 408975 270736 419217 270738
rect 408975 270733 409041 270736
rect 419151 270733 419217 270736
rect 452175 270796 452241 270799
rect 452655 270796 452721 270799
rect 452175 270794 452721 270796
rect 452175 270738 452180 270794
rect 452236 270738 452660 270794
rect 452716 270738 452721 270794
rect 452175 270736 452721 270738
rect 452175 270733 452241 270736
rect 452655 270733 452721 270736
rect 40762 270586 40768 270650
rect 40832 270648 40838 270650
rect 41775 270648 41841 270651
rect 40832 270646 41841 270648
rect 40832 270590 41780 270646
rect 41836 270590 41841 270646
rect 40832 270588 41841 270590
rect 40832 270586 40838 270588
rect 41775 270585 41841 270588
rect 41914 270586 41920 270650
rect 41984 270648 41990 270650
rect 42874 270648 42880 270650
rect 41984 270588 42880 270648
rect 41984 270586 41990 270588
rect 42874 270586 42880 270588
rect 42944 270586 42950 270650
rect 196335 270648 196401 270651
rect 317103 270648 317169 270651
rect 196335 270646 317169 270648
rect 196335 270590 196340 270646
rect 196396 270590 317108 270646
rect 317164 270590 317169 270646
rect 196335 270588 317169 270590
rect 196335 270585 196401 270588
rect 317103 270585 317169 270588
rect 317967 270648 318033 270651
rect 368463 270648 368529 270651
rect 369423 270650 369489 270651
rect 369807 270650 369873 270651
rect 369423 270648 369472 270650
rect 317967 270646 368529 270648
rect 317967 270590 317972 270646
rect 318028 270590 368468 270646
rect 368524 270590 368529 270646
rect 317967 270588 368529 270590
rect 369380 270646 369472 270648
rect 369380 270590 369428 270646
rect 369380 270588 369472 270590
rect 317967 270585 318033 270588
rect 368463 270585 368529 270588
rect 369423 270586 369472 270588
rect 369536 270586 369542 270650
rect 369807 270648 369856 270650
rect 369764 270646 369856 270648
rect 369764 270590 369812 270646
rect 369764 270588 369856 270590
rect 369807 270586 369856 270588
rect 369920 270586 369926 270650
rect 369999 270648 370065 270651
rect 641487 270648 641553 270651
rect 369999 270646 641553 270648
rect 369999 270590 370004 270646
rect 370060 270590 641492 270646
rect 641548 270590 641553 270646
rect 369999 270588 641553 270590
rect 369423 270585 369489 270586
rect 369807 270585 369873 270586
rect 369999 270585 370065 270588
rect 641487 270585 641553 270588
rect 253359 270500 253425 270503
rect 513039 270500 513105 270503
rect 548559 270500 548625 270503
rect 253359 270498 513105 270500
rect 253359 270442 253364 270498
rect 253420 270442 513044 270498
rect 513100 270442 513105 270498
rect 253359 270440 513105 270442
rect 253359 270437 253425 270440
rect 513039 270437 513105 270440
rect 513234 270498 548625 270500
rect 513234 270442 548564 270498
rect 548620 270442 548625 270498
rect 513234 270440 548625 270442
rect 315567 270352 315633 270355
rect 317967 270352 318033 270355
rect 315567 270350 318033 270352
rect 315567 270294 315572 270350
rect 315628 270294 317972 270350
rect 318028 270294 318033 270350
rect 315567 270292 318033 270294
rect 315567 270289 315633 270292
rect 317967 270289 318033 270292
rect 318159 270352 318225 270355
rect 338511 270352 338577 270355
rect 418959 270352 419025 270355
rect 318159 270350 338430 270352
rect 318159 270294 318164 270350
rect 318220 270294 338430 270350
rect 318159 270292 338430 270294
rect 318159 270289 318225 270292
rect 304911 270204 304977 270207
rect 317103 270204 317169 270207
rect 304911 270202 317169 270204
rect 304911 270146 304916 270202
rect 304972 270146 317108 270202
rect 317164 270146 317169 270202
rect 304911 270144 317169 270146
rect 304911 270141 304977 270144
rect 317103 270141 317169 270144
rect 319407 270204 319473 270207
rect 338370 270204 338430 270292
rect 338511 270350 419025 270352
rect 338511 270294 338516 270350
rect 338572 270294 418964 270350
rect 419020 270294 419025 270350
rect 338511 270292 419025 270294
rect 338511 270289 338577 270292
rect 418959 270289 419025 270292
rect 419151 270352 419217 270355
rect 438927 270352 438993 270355
rect 419151 270350 438993 270352
rect 419151 270294 419156 270350
rect 419212 270294 438932 270350
rect 438988 270294 438993 270350
rect 419151 270292 438993 270294
rect 419151 270289 419217 270292
rect 438927 270289 438993 270292
rect 449199 270352 449265 270355
rect 469455 270352 469521 270355
rect 449199 270350 469521 270352
rect 449199 270294 449204 270350
rect 449260 270294 469460 270350
rect 469516 270294 469521 270350
rect 449199 270292 469521 270294
rect 449199 270289 449265 270292
rect 469455 270289 469521 270292
rect 489519 270352 489585 270355
rect 513234 270352 513294 270440
rect 548559 270437 548625 270440
rect 575919 270500 575985 270503
rect 575919 270498 579006 270500
rect 575919 270442 575924 270498
rect 575980 270442 579006 270498
rect 575919 270440 579006 270442
rect 575919 270437 575985 270440
rect 489519 270350 513294 270352
rect 489519 270294 489524 270350
rect 489580 270294 513294 270350
rect 489519 270292 513294 270294
rect 578946 270352 579006 270440
rect 582063 270352 582129 270355
rect 578946 270350 582129 270352
rect 578946 270294 582068 270350
rect 582124 270294 582129 270350
rect 578946 270292 582129 270294
rect 489519 270289 489585 270292
rect 582063 270289 582129 270292
rect 428943 270204 429009 270207
rect 319407 270202 338238 270204
rect 319407 270146 319412 270202
rect 319468 270146 338238 270202
rect 319407 270144 338238 270146
rect 338370 270202 429009 270204
rect 338370 270146 428948 270202
rect 429004 270146 429009 270202
rect 338370 270144 429009 270146
rect 319407 270141 319473 270144
rect 41146 269994 41152 270058
rect 41216 270056 41222 270058
rect 41775 270056 41841 270059
rect 41216 270054 41841 270056
rect 41216 269998 41780 270054
rect 41836 269998 41841 270054
rect 41216 269996 41841 269998
rect 41216 269994 41222 269996
rect 41775 269993 41841 269996
rect 288015 270056 288081 270059
rect 308079 270056 308145 270059
rect 288015 270054 308145 270056
rect 288015 269998 288020 270054
rect 288076 269998 308084 270054
rect 308140 269998 308145 270054
rect 288015 269996 308145 269998
rect 288015 269993 288081 269996
rect 308079 269993 308145 269996
rect 316527 270056 316593 270059
rect 319503 270056 319569 270059
rect 316527 270054 319569 270056
rect 316527 269998 316532 270054
rect 316588 269998 319508 270054
rect 319564 269998 319569 270054
rect 316527 269996 319569 269998
rect 316527 269993 316593 269996
rect 319503 269993 319569 269996
rect 319695 270056 319761 270059
rect 328431 270056 328497 270059
rect 319695 270054 328497 270056
rect 319695 269998 319700 270054
rect 319756 269998 328436 270054
rect 328492 269998 328497 270054
rect 319695 269996 328497 269998
rect 319695 269993 319761 269996
rect 328431 269993 328497 269996
rect 328623 270056 328689 270059
rect 338031 270056 338097 270059
rect 328623 270054 338097 270056
rect 328623 269998 328628 270054
rect 328684 269998 338036 270054
rect 338092 269998 338097 270054
rect 328623 269996 338097 269998
rect 338178 270056 338238 270144
rect 428943 270141 429009 270144
rect 429231 270204 429297 270207
rect 539919 270204 539985 270207
rect 429231 270202 539985 270204
rect 429231 270146 429236 270202
rect 429292 270146 539924 270202
rect 539980 270146 539985 270202
rect 429231 270144 539985 270146
rect 429231 270141 429297 270144
rect 539919 270141 539985 270144
rect 560175 270204 560241 270207
rect 589167 270204 589233 270207
rect 560175 270202 589233 270204
rect 560175 270146 560180 270202
rect 560236 270146 589172 270202
rect 589228 270146 589233 270202
rect 560175 270144 589233 270146
rect 560175 270141 560241 270144
rect 589167 270141 589233 270144
rect 408975 270056 409041 270059
rect 338178 270054 409041 270056
rect 338178 269998 408980 270054
rect 409036 269998 409041 270054
rect 338178 269996 409041 269998
rect 328623 269993 328689 269996
rect 338031 269993 338097 269996
rect 408975 269993 409041 269996
rect 449199 270056 449265 270059
rect 540015 270056 540081 270059
rect 449199 270054 540081 270056
rect 449199 269998 449204 270054
rect 449260 269998 540020 270054
rect 540076 269998 540081 270054
rect 449199 269996 540081 269998
rect 449199 269993 449265 269996
rect 540015 269993 540081 269996
rect 560079 270056 560145 270059
rect 580239 270056 580305 270059
rect 560079 270054 580305 270056
rect 560079 269998 560084 270054
rect 560140 269998 580244 270054
rect 580300 269998 580305 270054
rect 560079 269996 580305 269998
rect 560079 269993 560145 269996
rect 580239 269993 580305 269996
rect 673839 270056 673905 270059
rect 673839 270054 674784 270056
rect 673839 269998 673844 270054
rect 673900 269998 674784 270054
rect 673839 269996 674784 269998
rect 673839 269993 673905 269996
rect 269199 269908 269265 269911
rect 316719 269908 316785 269911
rect 269199 269906 316785 269908
rect 269199 269850 269204 269906
rect 269260 269850 316724 269906
rect 316780 269850 316785 269906
rect 269199 269848 316785 269850
rect 269199 269845 269265 269848
rect 316719 269845 316785 269848
rect 320175 269908 320241 269911
rect 603375 269908 603441 269911
rect 320175 269906 603441 269908
rect 320175 269850 320180 269906
rect 320236 269850 603380 269906
rect 603436 269850 603441 269906
rect 320175 269848 603441 269850
rect 320175 269845 320241 269848
rect 603375 269845 603441 269848
rect 264879 269760 264945 269763
rect 605775 269760 605841 269763
rect 264879 269758 605841 269760
rect 264879 269702 264884 269758
rect 264940 269702 605780 269758
rect 605836 269702 605841 269758
rect 264879 269700 605841 269702
rect 264879 269697 264945 269700
rect 605775 269697 605841 269700
rect 674703 269760 674769 269763
rect 674703 269758 674814 269760
rect 674703 269702 674708 269758
rect 674764 269702 674814 269758
rect 674703 269697 674814 269702
rect 266607 269612 266673 269615
rect 620079 269612 620145 269615
rect 266607 269610 620145 269612
rect 266607 269554 266612 269610
rect 266668 269554 620084 269610
rect 620140 269554 620145 269610
rect 674754 269582 674814 269697
rect 266607 269552 620145 269554
rect 266607 269549 266673 269552
rect 620079 269549 620145 269552
rect 267663 269464 267729 269467
rect 630831 269464 630897 269467
rect 267663 269462 630897 269464
rect 267663 269406 267668 269462
rect 267724 269406 630836 269462
rect 630892 269406 630897 269462
rect 267663 269404 630897 269406
rect 267663 269401 267729 269404
rect 630831 269401 630897 269404
rect 268143 269316 268209 269319
rect 634287 269316 634353 269319
rect 268143 269314 634353 269316
rect 268143 269258 268148 269314
rect 268204 269258 634292 269314
rect 634348 269258 634353 269314
rect 268143 269256 634353 269258
rect 268143 269253 268209 269256
rect 634287 269253 634353 269256
rect 40954 269106 40960 269170
rect 41024 269168 41030 269170
rect 41775 269168 41841 269171
rect 41024 269166 41841 269168
rect 41024 269110 41780 269166
rect 41836 269110 41841 269166
rect 41024 269108 41841 269110
rect 41024 269106 41030 269108
rect 41775 269105 41841 269108
rect 260559 269168 260625 269171
rect 280815 269168 280881 269171
rect 260559 269166 280881 269168
rect 260559 269110 260564 269166
rect 260620 269110 280820 269166
rect 280876 269110 280881 269166
rect 260559 269108 280881 269110
rect 260559 269105 260625 269108
rect 280815 269105 280881 269108
rect 290746 269106 290752 269170
rect 290816 269168 290822 269170
rect 296655 269168 296721 269171
rect 290816 269166 296721 269168
rect 290816 269110 296660 269166
rect 296716 269110 296721 269166
rect 290816 269108 296721 269110
rect 290816 269106 290822 269108
rect 296655 269105 296721 269108
rect 316666 269106 316672 269170
rect 316736 269168 316742 269170
rect 334095 269168 334161 269171
rect 347247 269170 347313 269171
rect 316736 269166 334161 269168
rect 316736 269110 334100 269166
rect 334156 269110 334161 269166
rect 316736 269108 334161 269110
rect 316736 269106 316742 269108
rect 334095 269105 334161 269108
rect 347194 269106 347200 269170
rect 347264 269168 347313 269170
rect 347535 269170 347601 269171
rect 347264 269166 347356 269168
rect 347308 269110 347356 269166
rect 347264 269108 347356 269110
rect 347535 269166 347584 269170
rect 347648 269168 347654 269170
rect 348015 269168 348081 269171
rect 367119 269168 367185 269171
rect 347535 269110 347540 269166
rect 347264 269106 347313 269108
rect 347247 269105 347313 269106
rect 347535 269106 347584 269110
rect 347648 269108 347692 269168
rect 348015 269166 367185 269168
rect 348015 269110 348020 269166
rect 348076 269110 367124 269166
rect 367180 269110 367185 269166
rect 348015 269108 367185 269110
rect 347648 269106 347654 269108
rect 347535 269105 347601 269106
rect 348015 269105 348081 269108
rect 367119 269105 367185 269108
rect 368751 269168 368817 269171
rect 376911 269168 376977 269171
rect 368751 269166 376977 269168
rect 368751 269110 368756 269166
rect 368812 269110 376916 269166
rect 376972 269110 376977 269166
rect 368751 269108 376977 269110
rect 368751 269105 368817 269108
rect 376911 269105 376977 269108
rect 377103 269168 377169 269171
rect 379215 269168 379281 269171
rect 377103 269166 379281 269168
rect 377103 269110 377108 269166
rect 377164 269110 379220 269166
rect 379276 269110 379281 269166
rect 377103 269108 379281 269110
rect 377103 269105 377169 269108
rect 379215 269105 379281 269108
rect 380079 269168 380145 269171
rect 640335 269168 640401 269171
rect 380079 269166 640401 269168
rect 380079 269110 380084 269166
rect 380140 269110 640340 269166
rect 640396 269110 640401 269166
rect 380079 269108 640401 269110
rect 380079 269105 380145 269108
rect 640335 269105 640401 269108
rect 674703 269168 674769 269171
rect 674703 269166 674814 269168
rect 674703 269110 674708 269166
rect 674764 269110 674814 269166
rect 674703 269105 674814 269110
rect 252879 269020 252945 269023
rect 282255 269020 282321 269023
rect 317583 269020 317649 269023
rect 252879 269018 261822 269020
rect 252879 268962 252884 269018
rect 252940 268962 261822 269018
rect 252879 268960 261822 268962
rect 252879 268957 252945 268960
rect 252015 268872 252081 268875
rect 261762 268872 261822 268960
rect 282255 269018 317649 269020
rect 282255 268962 282260 269018
rect 282316 268962 317588 269018
rect 317644 268962 317649 269018
rect 282255 268960 317649 268962
rect 282255 268957 282321 268960
rect 317583 268957 317649 268960
rect 317775 269020 317841 269023
rect 574863 269020 574929 269023
rect 317775 269018 574929 269020
rect 317775 268962 317780 269018
rect 317836 268962 574868 269018
rect 574924 268962 574929 269018
rect 674754 268990 674814 269105
rect 317775 268960 574929 268962
rect 317775 268957 317841 268960
rect 574863 268957 574929 268960
rect 509487 268872 509553 268875
rect 252015 268870 261630 268872
rect 252015 268814 252020 268870
rect 252076 268814 261630 268870
rect 252015 268812 261630 268814
rect 261762 268870 509553 268872
rect 261762 268814 509492 268870
rect 509548 268814 509553 268870
rect 261762 268812 509553 268814
rect 252015 268809 252081 268812
rect 211503 268724 211569 268727
rect 257391 268724 257457 268727
rect 211503 268722 257457 268724
rect 211503 268666 211508 268722
rect 211564 268666 257396 268722
rect 257452 268666 257457 268722
rect 211503 268664 257457 268666
rect 211503 268661 211569 268664
rect 257391 268661 257457 268664
rect 250287 268576 250353 268579
rect 261327 268576 261393 268579
rect 250287 268574 261393 268576
rect 250287 268518 250292 268574
rect 250348 268518 261332 268574
rect 261388 268518 261393 268574
rect 250287 268516 261393 268518
rect 261570 268576 261630 268812
rect 509487 268809 509553 268812
rect 539919 268872 539985 268875
rect 560175 268872 560241 268875
rect 539919 268870 560241 268872
rect 539919 268814 539924 268870
rect 539980 268814 560180 268870
rect 560236 268814 560241 268870
rect 539919 268812 560241 268814
rect 539919 268809 539985 268812
rect 560175 268809 560241 268812
rect 580239 268872 580305 268875
rect 596367 268872 596433 268875
rect 580239 268870 596433 268872
rect 580239 268814 580244 268870
rect 580300 268814 596372 268870
rect 596428 268814 596433 268870
rect 580239 268812 596433 268814
rect 580239 268809 580305 268812
rect 596367 268809 596433 268812
rect 265071 268724 265137 268727
rect 277839 268724 277905 268727
rect 265071 268722 277905 268724
rect 265071 268666 265076 268722
rect 265132 268666 277844 268722
rect 277900 268666 277905 268722
rect 265071 268664 277905 268666
rect 265071 268661 265137 268664
rect 277839 268661 277905 268664
rect 280815 268724 280881 268727
rect 288303 268724 288369 268727
rect 280815 268722 288369 268724
rect 280815 268666 280820 268722
rect 280876 268666 288308 268722
rect 288364 268666 288369 268722
rect 280815 268664 288369 268666
rect 280815 268661 280881 268664
rect 288303 268661 288369 268664
rect 291855 268724 291921 268727
rect 315567 268724 315633 268727
rect 291855 268722 315633 268724
rect 291855 268666 291860 268722
rect 291916 268666 315572 268722
rect 315628 268666 315633 268722
rect 291855 268664 315633 268666
rect 291855 268661 291921 268664
rect 315567 268661 315633 268664
rect 315759 268724 315825 268727
rect 567759 268724 567825 268727
rect 315759 268722 567825 268724
rect 315759 268666 315764 268722
rect 315820 268666 567764 268722
rect 567820 268666 567825 268722
rect 315759 268664 567825 268666
rect 315759 268661 315825 268664
rect 567759 268661 567825 268664
rect 677242 268662 677248 268726
rect 677312 268662 677318 268726
rect 502287 268576 502353 268579
rect 261570 268574 502353 268576
rect 261570 268518 502292 268574
rect 502348 268518 502353 268574
rect 261570 268516 502353 268518
rect 250287 268513 250353 268516
rect 261327 268513 261393 268516
rect 502287 268513 502353 268516
rect 540015 268576 540081 268579
rect 560079 268576 560145 268579
rect 540015 268574 560145 268576
rect 540015 268518 540020 268574
rect 540076 268518 560084 268574
rect 560140 268518 560145 268574
rect 540015 268516 560145 268518
rect 540015 268513 540081 268516
rect 560079 268513 560145 268516
rect 258927 268428 258993 268431
rect 288015 268428 288081 268431
rect 258927 268426 288081 268428
rect 258927 268370 258932 268426
rect 258988 268370 288020 268426
rect 288076 268370 288081 268426
rect 258927 268368 288081 268370
rect 258927 268365 258993 268368
rect 288015 268365 288081 268368
rect 288303 268428 288369 268431
rect 290746 268428 290752 268430
rect 288303 268426 290752 268428
rect 288303 268370 288308 268426
rect 288364 268370 290752 268426
rect 288303 268368 290752 268370
rect 288303 268365 288369 268368
rect 290746 268366 290752 268368
rect 290816 268366 290822 268430
rect 308079 268428 308145 268431
rect 348346 268428 348352 268430
rect 308079 268426 348352 268428
rect 308079 268370 308084 268426
rect 308140 268370 348352 268426
rect 308079 268368 348352 268370
rect 308079 268365 308145 268368
rect 348346 268366 348352 268368
rect 348416 268366 348422 268430
rect 348591 268428 348657 268431
rect 377530 268428 377536 268430
rect 348591 268426 377536 268428
rect 348591 268370 348596 268426
rect 348652 268370 377536 268426
rect 348591 268368 377536 268370
rect 348591 268365 348657 268368
rect 377530 268366 377536 268368
rect 377600 268366 377606 268430
rect 378159 268428 378225 268431
rect 388623 268428 388689 268431
rect 378159 268426 388689 268428
rect 378159 268370 378164 268426
rect 378220 268370 388628 268426
rect 388684 268370 388689 268426
rect 378159 268368 388689 268370
rect 378159 268365 378225 268368
rect 388623 268365 388689 268368
rect 388815 268428 388881 268431
rect 389199 268428 389265 268431
rect 388815 268426 389265 268428
rect 388815 268370 388820 268426
rect 388876 268370 389204 268426
rect 389260 268370 389265 268426
rect 388815 268368 389265 268370
rect 388815 268365 388881 268368
rect 389199 268365 389265 268368
rect 389391 268428 389457 268431
rect 403695 268428 403761 268431
rect 389391 268426 403761 268428
rect 389391 268370 389396 268426
rect 389452 268370 403700 268426
rect 403756 268370 403761 268426
rect 389391 268368 403761 268370
rect 389391 268365 389457 268368
rect 403695 268365 403761 268368
rect 403887 268428 403953 268431
rect 405946 268428 405952 268430
rect 403887 268426 405952 268428
rect 403887 268370 403892 268426
rect 403948 268370 405952 268426
rect 403887 268368 405952 268370
rect 403887 268365 403953 268368
rect 405946 268366 405952 268368
rect 406016 268366 406022 268430
rect 406095 268428 406161 268431
rect 626031 268428 626097 268431
rect 406095 268426 626097 268428
rect 406095 268370 406100 268426
rect 406156 268370 626036 268426
rect 626092 268370 626097 268426
rect 677250 268398 677310 268662
rect 406095 268368 626097 268370
rect 406095 268365 406161 268368
rect 626031 268365 626097 268368
rect 261135 268280 261201 268283
rect 254466 268278 261201 268280
rect 254466 268222 261140 268278
rect 261196 268222 261201 268278
rect 254466 268220 261201 268222
rect 211119 268132 211185 268135
rect 254466 268132 254526 268220
rect 261135 268217 261201 268220
rect 261327 268280 261393 268283
rect 488079 268280 488145 268283
rect 261327 268278 488145 268280
rect 261327 268222 261332 268278
rect 261388 268222 488084 268278
rect 488140 268222 488145 268278
rect 261327 268220 488145 268222
rect 261327 268217 261393 268220
rect 488079 268217 488145 268220
rect 211119 268130 254526 268132
rect 211119 268074 211124 268130
rect 211180 268074 254526 268130
rect 211119 268072 254526 268074
rect 257295 268132 257361 268135
rect 277647 268132 277713 268135
rect 257295 268130 277713 268132
rect 257295 268074 257300 268130
rect 257356 268074 277652 268130
rect 277708 268074 277713 268130
rect 257295 268072 277713 268074
rect 211119 268069 211185 268072
rect 257295 268069 257361 268072
rect 277647 268069 277713 268072
rect 277839 268132 277905 268135
rect 291855 268132 291921 268135
rect 277839 268130 291921 268132
rect 277839 268074 277844 268130
rect 277900 268074 291860 268130
rect 291916 268074 291921 268130
rect 277839 268072 291921 268074
rect 277839 268069 277905 268072
rect 291855 268069 291921 268072
rect 292282 268070 292288 268134
rect 292352 268132 292358 268134
rect 312442 268132 312448 268134
rect 292352 268072 312448 268132
rect 292352 268070 292358 268072
rect 312442 268070 312448 268072
rect 312512 268070 312518 268134
rect 312687 268132 312753 268135
rect 316666 268132 316672 268134
rect 312687 268130 316672 268132
rect 312687 268074 312692 268130
rect 312748 268074 316672 268130
rect 312687 268072 316672 268074
rect 312687 268069 312753 268072
rect 316666 268070 316672 268072
rect 316736 268070 316742 268134
rect 317583 268132 317649 268135
rect 336207 268132 336273 268135
rect 317583 268130 336273 268132
rect 317583 268074 317588 268130
rect 317644 268074 336212 268130
rect 336268 268074 336273 268130
rect 317583 268072 336273 268074
rect 317583 268069 317649 268072
rect 336207 268069 336273 268072
rect 336399 268134 336465 268135
rect 336399 268130 336448 268134
rect 336512 268132 336518 268134
rect 336975 268132 337041 268135
rect 560655 268132 560721 268135
rect 336399 268074 336404 268130
rect 336399 268070 336448 268074
rect 336512 268072 336556 268132
rect 336975 268130 560721 268132
rect 336975 268074 336980 268130
rect 337036 268074 560660 268130
rect 560716 268074 560721 268130
rect 336975 268072 560721 268074
rect 336512 268070 336518 268072
rect 336399 268069 336465 268070
rect 336975 268069 337041 268072
rect 560655 268069 560721 268072
rect 254607 267984 254673 267987
rect 377199 267984 377265 267987
rect 395439 267984 395505 267987
rect 397551 267984 397617 267987
rect 401679 267984 401745 267987
rect 254607 267982 377265 267984
rect 254607 267926 254612 267982
rect 254668 267926 377204 267982
rect 377260 267926 377265 267982
rect 254607 267924 377265 267926
rect 254607 267921 254673 267924
rect 377199 267921 377265 267924
rect 377346 267982 395505 267984
rect 377346 267926 395444 267982
rect 395500 267926 395505 267982
rect 377346 267924 395505 267926
rect 211023 267836 211089 267839
rect 211503 267836 211569 267839
rect 211023 267834 211569 267836
rect 211023 267778 211028 267834
rect 211084 267778 211508 267834
rect 211564 267778 211569 267834
rect 211023 267776 211569 267778
rect 211023 267773 211089 267776
rect 211503 267773 211569 267776
rect 261999 267836 262065 267839
rect 267375 267836 267441 267839
rect 261999 267834 267441 267836
rect 261999 267778 262004 267834
rect 262060 267778 267380 267834
rect 267436 267778 267441 267834
rect 261999 267776 267441 267778
rect 261999 267773 262065 267776
rect 267375 267773 267441 267776
rect 267759 267836 267825 267839
rect 267898 267836 267904 267838
rect 267759 267834 267904 267836
rect 267759 267778 267764 267834
rect 267820 267778 267904 267834
rect 267759 267776 267904 267778
rect 267759 267773 267825 267776
rect 267898 267774 267904 267776
rect 267968 267774 267974 267838
rect 268047 267834 268113 267839
rect 268047 267778 268052 267834
rect 268108 267778 268113 267834
rect 268047 267773 268113 267778
rect 268239 267836 268305 267839
rect 287535 267836 287601 267839
rect 288495 267836 288561 267839
rect 307834 267836 307840 267838
rect 268239 267834 287601 267836
rect 268239 267778 268244 267834
rect 268300 267778 287540 267834
rect 287596 267778 287601 267834
rect 268239 267776 287601 267778
rect 268239 267773 268305 267776
rect 287535 267773 287601 267776
rect 287682 267776 288318 267836
rect 268050 267688 268110 267773
rect 287682 267688 287742 267776
rect 268050 267628 287742 267688
rect 288258 267688 288318 267776
rect 288495 267834 307840 267836
rect 288495 267778 288500 267834
rect 288556 267778 307840 267834
rect 288495 267776 307840 267778
rect 288495 267773 288561 267776
rect 307834 267774 307840 267776
rect 307904 267774 307910 267838
rect 308410 267774 308416 267838
rect 308480 267836 308486 267838
rect 312111 267836 312177 267839
rect 327855 267836 327921 267839
rect 376570 267836 376576 267838
rect 308480 267834 312177 267836
rect 308480 267778 312116 267834
rect 312172 267778 312177 267834
rect 308480 267776 312177 267778
rect 308480 267774 308486 267776
rect 312111 267773 312177 267776
rect 312258 267834 327921 267836
rect 312258 267778 327860 267834
rect 327916 267778 327921 267834
rect 312258 267776 327921 267778
rect 312258 267688 312318 267776
rect 327855 267773 327921 267776
rect 328002 267776 376576 267836
rect 288258 267628 312318 267688
rect 312442 267626 312448 267690
rect 312512 267688 312518 267690
rect 328002 267688 328062 267776
rect 376570 267774 376576 267776
rect 376640 267774 376646 267838
rect 376815 267836 376881 267839
rect 376770 267834 376881 267836
rect 376770 267778 376820 267834
rect 376876 267778 376881 267834
rect 376770 267773 376881 267778
rect 377007 267836 377073 267839
rect 377346 267836 377406 267924
rect 395439 267921 395505 267924
rect 397122 267982 397617 267984
rect 397122 267926 397556 267982
rect 397612 267926 397617 267982
rect 397122 267924 397617 267926
rect 377007 267834 377406 267836
rect 377007 267778 377012 267834
rect 377068 267778 377406 267834
rect 377007 267776 377406 267778
rect 377967 267836 378033 267839
rect 378735 267836 378801 267839
rect 377967 267834 378801 267836
rect 377967 267778 377972 267834
rect 378028 267778 378740 267834
rect 378796 267778 378801 267834
rect 377967 267776 378801 267778
rect 377007 267773 377073 267776
rect 377967 267773 378033 267776
rect 378735 267773 378801 267776
rect 379311 267836 379377 267839
rect 383439 267836 383505 267839
rect 379311 267834 383505 267836
rect 379311 267778 379316 267834
rect 379372 267778 383444 267834
rect 383500 267778 383505 267834
rect 379311 267776 383505 267778
rect 379311 267773 379377 267776
rect 383439 267773 383505 267776
rect 383674 267774 383680 267838
rect 383744 267836 383750 267838
rect 397122 267836 397182 267924
rect 397551 267921 397617 267924
rect 397698 267982 401745 267984
rect 397698 267926 401684 267982
rect 401740 267926 401745 267982
rect 397698 267924 401745 267926
rect 383744 267776 397182 267836
rect 383744 267774 383750 267776
rect 312512 267628 328062 267688
rect 312512 267626 312518 267628
rect 336442 267626 336448 267690
rect 336512 267688 336518 267690
rect 347194 267688 347200 267690
rect 336512 267628 347200 267688
rect 336512 267626 336518 267628
rect 347194 267626 347200 267628
rect 347264 267626 347270 267690
rect 347578 267626 347584 267690
rect 347648 267688 347654 267690
rect 376770 267688 376830 267773
rect 347648 267628 376830 267688
rect 347648 267626 347654 267628
rect 376954 267626 376960 267690
rect 377024 267688 377030 267690
rect 397698 267688 397758 267924
rect 401679 267921 401745 267924
rect 404751 267984 404817 267987
rect 405370 267984 405376 267986
rect 404751 267982 405376 267984
rect 404751 267926 404756 267982
rect 404812 267926 405376 267982
rect 404751 267924 405376 267926
rect 404751 267921 404817 267924
rect 405370 267922 405376 267924
rect 405440 267922 405446 267986
rect 405615 267984 405681 267987
rect 405754 267984 405760 267986
rect 405615 267982 405760 267984
rect 405615 267926 405620 267982
rect 405676 267926 405760 267982
rect 405615 267924 405760 267926
rect 405615 267921 405681 267924
rect 405754 267922 405760 267924
rect 405824 267922 405830 267986
rect 406330 267922 406336 267986
rect 406400 267984 406406 267986
rect 408591 267984 408657 267987
rect 406400 267982 408657 267984
rect 406400 267926 408596 267982
rect 408652 267926 408657 267982
rect 406400 267924 408657 267926
rect 406400 267922 406406 267924
rect 408591 267921 408657 267924
rect 408783 267984 408849 267987
rect 418959 267984 419025 267987
rect 439119 267984 439185 267987
rect 408783 267982 413118 267984
rect 408783 267926 408788 267982
rect 408844 267926 413118 267982
rect 408783 267924 413118 267926
rect 408783 267921 408849 267924
rect 397839 267836 397905 267839
rect 408783 267836 408849 267839
rect 412911 267836 412977 267839
rect 397839 267834 408702 267836
rect 397839 267778 397844 267834
rect 397900 267778 408702 267834
rect 397839 267776 408702 267778
rect 397839 267773 397905 267776
rect 377024 267628 397758 267688
rect 408642 267688 408702 267776
rect 408783 267834 412977 267836
rect 408783 267778 408788 267834
rect 408844 267778 412916 267834
rect 412972 267778 412977 267834
rect 408783 267776 412977 267778
rect 413058 267836 413118 267924
rect 418959 267982 439185 267984
rect 418959 267926 418964 267982
rect 419020 267926 439124 267982
rect 439180 267926 439185 267982
rect 418959 267924 439185 267926
rect 418959 267921 419025 267924
rect 439119 267921 439185 267924
rect 439311 267984 439377 267987
rect 449199 267984 449265 267987
rect 439311 267982 449265 267984
rect 439311 267926 439316 267982
rect 439372 267926 449204 267982
rect 449260 267926 449265 267982
rect 439311 267924 449265 267926
rect 439311 267921 439377 267924
rect 449199 267921 449265 267924
rect 469455 267984 469521 267987
rect 489519 267984 489585 267987
rect 469455 267982 489585 267984
rect 469455 267926 469460 267982
rect 469516 267926 489524 267982
rect 489580 267926 489585 267982
rect 469455 267924 489585 267926
rect 469455 267921 469521 267924
rect 489519 267921 489585 267924
rect 614223 267836 614289 267839
rect 413058 267834 614289 267836
rect 413058 267778 614228 267834
rect 614284 267778 614289 267834
rect 413058 267776 614289 267778
rect 408783 267773 408849 267776
rect 412911 267773 412977 267776
rect 614223 267773 614289 267776
rect 414927 267688 414993 267691
rect 408642 267686 414993 267688
rect 408642 267630 414932 267686
rect 414988 267630 414993 267686
rect 408642 267628 414993 267630
rect 377024 267626 377030 267628
rect 414927 267625 414993 267628
rect 415119 267688 415185 267691
rect 639087 267688 639153 267691
rect 677442 267690 677502 267880
rect 415119 267686 639153 267688
rect 415119 267630 415124 267686
rect 415180 267630 639092 267686
rect 639148 267630 639153 267686
rect 415119 267628 639153 267630
rect 415119 267625 415185 267628
rect 639087 267625 639153 267628
rect 677434 267626 677440 267690
rect 677504 267626 677510 267690
rect 8158 266560 8584 267360
rect 9384 267359 50926 267360
rect 9384 266561 50127 267359
rect 50925 266561 50931 267359
rect 677058 267098 677118 267362
rect 676858 267034 676864 267098
rect 676928 267034 676934 267098
rect 677050 267034 677056 267098
rect 677120 267034 677126 267098
rect 676866 266770 676926 267034
rect 9384 266560 50926 266561
rect 413679 266208 413745 266211
rect 609423 266208 609489 266211
rect 413679 266206 609489 266208
rect 413679 266150 413684 266206
rect 413740 266150 609428 266206
rect 609484 266150 609489 266206
rect 413679 266148 609489 266150
rect 413679 266145 413745 266148
rect 609423 266145 609489 266148
rect 674607 266060 674673 266063
rect 674754 266060 674814 266252
rect 674607 266058 674814 266060
rect 674607 266002 674612 266058
rect 674668 266002 674814 266058
rect 674607 266000 674814 266002
rect 674607 265997 674673 266000
rect 414927 265912 414993 265915
rect 631791 265912 631857 265915
rect 7814 265112 16354 265912
rect 17154 265911 52718 265912
rect 17154 265113 51919 265911
rect 52717 265113 52723 265911
rect 414927 265910 631857 265912
rect 414927 265854 414932 265910
rect 414988 265854 631796 265910
rect 631852 265854 631857 265910
rect 414927 265852 631857 265854
rect 414927 265849 414993 265852
rect 631791 265849 631857 265852
rect 677250 265471 677310 265734
rect 412911 265468 412977 265471
rect 628431 265468 628497 265471
rect 412911 265466 628497 265468
rect 412911 265410 412916 265466
rect 412972 265410 628436 265466
rect 628492 265410 628497 265466
rect 412911 265408 628497 265410
rect 412911 265405 412977 265408
rect 628431 265405 628497 265408
rect 677199 265466 677310 265471
rect 677199 265410 677204 265466
rect 677260 265410 677310 265466
rect 677199 265408 677310 265410
rect 677199 265405 677265 265408
rect 412815 265320 412881 265323
rect 527343 265320 527409 265323
rect 412815 265318 527409 265320
rect 412815 265262 412820 265318
rect 412876 265262 527348 265318
rect 527404 265262 527409 265318
rect 412815 265260 527409 265262
rect 412815 265257 412881 265260
rect 527343 265257 527409 265260
rect 412719 265172 412785 265175
rect 530895 265172 530961 265175
rect 412719 265170 530961 265172
rect 412719 265114 412724 265170
rect 412780 265114 530900 265170
rect 530956 265114 530961 265170
rect 17154 265112 52718 265113
rect 412719 265112 530961 265114
rect 412719 265109 412785 265112
rect 530895 265109 530961 265112
rect 674946 265027 675006 265142
rect 412623 265024 412689 265027
rect 537999 265024 538065 265027
rect 412623 265022 538065 265024
rect 412623 264966 412628 265022
rect 412684 264966 538004 265022
rect 538060 264966 538065 265022
rect 412623 264964 538065 264966
rect 412623 264961 412689 264964
rect 537999 264961 538065 264964
rect 674895 265022 675006 265027
rect 674895 264966 674900 265022
rect 674956 264966 675006 265022
rect 674895 264964 675006 264966
rect 674895 264961 674961 264964
rect 407089 264945 407182 264949
rect 267565 264922 267635 264927
rect 267565 264896 267570 264922
rect 267564 264862 267570 264896
rect 267630 264896 267635 264922
rect 388974 264913 389044 264918
rect 388974 264896 388979 264913
rect 267630 264862 388979 264896
rect 267564 264853 388979 264862
rect 389039 264853 389044 264913
rect 267564 264848 389044 264853
rect 393009 264899 393079 264904
rect 267564 264836 389024 264848
rect 393009 264839 393014 264899
rect 393074 264896 393079 264899
rect 393074 264839 406994 264896
rect 393009 264836 406994 264839
rect 393009 264834 393079 264836
rect 406934 264728 406994 264836
rect 407089 264875 407098 264945
rect 407168 264875 407182 264945
rect 407701 264935 407771 264939
rect 407665 264934 407771 264935
rect 407089 264811 407182 264875
rect 407290 264814 407296 264878
rect 407360 264876 407366 264878
rect 407665 264876 407706 264934
rect 407360 264874 407706 264876
rect 407766 264874 407771 264934
rect 407360 264869 407771 264874
rect 408065 264938 408188 264946
rect 407360 264816 407725 264869
rect 408065 264868 408109 264938
rect 408179 264868 408188 264938
rect 410528 264941 410598 264946
rect 408065 264860 408188 264868
rect 409991 264921 410061 264926
rect 409991 264861 409996 264921
rect 410056 264876 410061 264921
rect 410528 264881 410533 264941
rect 410593 264929 410598 264941
rect 410593 264881 410622 264929
rect 410362 264876 410368 264878
rect 410056 264861 410368 264876
rect 409991 264856 410368 264861
rect 409995 264816 410368 264856
rect 407360 264814 407366 264816
rect 410362 264814 410368 264816
rect 410432 264814 410438 264878
rect 410528 264876 410622 264881
rect 489519 264876 489585 264879
rect 406934 264668 409854 264728
rect 409794 264284 409854 264668
rect 409978 264666 409984 264730
rect 410048 264728 410054 264730
rect 410562 264728 410622 264876
rect 419010 264816 449214 264876
rect 410048 264668 410622 264728
rect 410048 264666 410054 264668
rect 410746 264666 410752 264730
rect 410816 264728 410822 264730
rect 411514 264728 411520 264730
rect 410816 264668 411520 264728
rect 410816 264666 410822 264668
rect 411514 264666 411520 264668
rect 411584 264666 411590 264730
rect 410554 264518 410560 264582
rect 410624 264580 410630 264582
rect 412047 264580 412113 264583
rect 410624 264578 412113 264580
rect 410624 264522 412052 264578
rect 412108 264522 412113 264578
rect 410624 264520 412113 264522
rect 410624 264518 410630 264520
rect 412047 264517 412113 264520
rect 419010 264284 419070 264816
rect 449154 264728 449214 264816
rect 489519 264874 521214 264876
rect 489519 264818 489524 264874
rect 489580 264818 521214 264874
rect 489519 264816 521214 264818
rect 489519 264813 489585 264816
rect 449391 264728 449457 264731
rect 449154 264726 449457 264728
rect 449154 264670 449396 264726
rect 449452 264670 449457 264726
rect 449154 264668 449457 264670
rect 449391 264665 449457 264668
rect 469359 264728 469425 264731
rect 475791 264728 475857 264731
rect 469359 264726 475857 264728
rect 469359 264670 469364 264726
rect 469420 264670 475796 264726
rect 475852 264670 475857 264726
rect 469359 264668 475857 264670
rect 469359 264665 469425 264668
rect 475791 264665 475857 264668
rect 521154 264432 521214 264816
rect 674415 264654 674481 264657
rect 674415 264652 674784 264654
rect 674415 264596 674420 264652
rect 674476 264596 674784 264652
rect 674415 264594 674784 264596
rect 674415 264591 674481 264594
rect 555855 264580 555921 264583
rect 529986 264578 555921 264580
rect 529986 264522 555860 264578
rect 555916 264522 555921 264578
rect 529986 264520 555921 264522
rect 529986 264432 530046 264520
rect 555855 264517 555921 264520
rect 521154 264372 530046 264432
rect 409794 264224 419070 264284
rect 674170 264074 674176 264138
rect 674240 264136 674246 264138
rect 674240 264076 674784 264136
rect 674240 264074 674246 264076
rect 7202 263216 7374 264016
rect 8174 264015 54502 264016
rect 8174 263217 53703 264015
rect 54501 263217 54507 264015
rect 677634 263251 677694 263514
rect 677583 263246 677694 263251
rect 8174 263216 54502 263217
rect 677583 263190 677588 263246
rect 677644 263190 677694 263246
rect 677583 263188 677694 263190
rect 677583 263185 677649 263188
rect 675138 262807 675198 262996
rect 675138 262802 675249 262807
rect 675138 262746 675188 262802
rect 675244 262746 675249 262802
rect 675138 262744 675249 262746
rect 675183 262741 675249 262744
rect 674319 262508 674385 262511
rect 674319 262506 674784 262508
rect 674319 262450 674324 262506
rect 674380 262450 674784 262506
rect 674319 262448 674784 262450
rect 674319 262445 674385 262448
rect 7296 261322 17562 262122
rect 18362 262121 56068 262122
rect 18362 261323 55269 262121
rect 56067 261323 56073 262121
rect 207183 261324 207249 261327
rect 211842 261324 211902 261812
rect 674754 261771 674814 261886
rect 674703 261766 674814 261771
rect 674703 261710 674708 261766
rect 674764 261710 674814 261766
rect 674703 261708 674814 261710
rect 674703 261705 674769 261708
rect 18362 261322 56068 261323
rect 207183 261322 211902 261324
rect 207183 261266 207188 261322
rect 207244 261266 211902 261322
rect 207183 261264 211902 261266
rect 674127 261324 674193 261327
rect 674754 261324 674814 261368
rect 674127 261322 674814 261324
rect 674127 261266 674132 261322
rect 674188 261266 674814 261322
rect 674127 261264 674814 261266
rect 207183 261261 207249 261264
rect 674127 261261 674193 261264
rect 673978 260818 673984 260882
rect 674048 260880 674054 260882
rect 674048 260820 674784 260880
rect 674048 260818 674054 260820
rect 674754 260143 674814 260258
rect 674754 260138 674865 260143
rect 674754 260082 674804 260138
rect 674860 260082 674865 260138
rect 674754 260080 674865 260082
rect 674799 260077 674865 260080
rect 42447 259696 42513 259699
rect 42447 259694 42558 259696
rect 42447 259638 42452 259694
rect 42508 259638 42558 259694
rect 42447 259633 42558 259638
rect 42498 259518 42558 259633
rect 206844 259544 209180 259720
rect 206844 259536 211458 259544
rect 206844 259496 211282 259536
rect 42831 258956 42897 258959
rect 42528 258954 42897 258956
rect 42528 258898 42836 258954
rect 42892 258898 42897 258954
rect 42528 258896 42897 258898
rect 42831 258893 42897 258896
rect 42447 258660 42513 258663
rect 42447 258658 42558 258660
rect 42447 258602 42452 258658
rect 42508 258602 42558 258658
rect 42447 258597 42558 258602
rect 42498 258334 42558 258597
rect 42306 257624 42366 257890
rect 43215 257624 43281 257627
rect 42306 257622 43281 257624
rect 42306 257566 43220 257622
rect 43276 257566 43281 257622
rect 42306 257564 43281 257566
rect 43215 257561 43281 257564
rect 42447 257476 42513 257479
rect 42447 257474 42558 257476
rect 42447 257418 42452 257474
rect 42508 257418 42558 257474
rect 42447 257413 42558 257418
rect 42498 257298 42558 257413
rect 40378 256970 40384 257034
rect 40448 256970 40454 257034
rect 40386 256736 40446 256970
rect 206844 256926 206998 259496
rect 209004 256926 211282 259496
rect 206844 256878 211282 256926
rect 211434 256878 211458 259536
rect 412810 259516 424188 259554
rect 412810 256884 412836 259516
rect 412992 259382 424188 259516
rect 674946 259551 675006 259740
rect 674946 259546 675057 259551
rect 674946 259490 674996 259546
rect 675052 259490 675057 259546
rect 674946 259488 675057 259490
rect 674991 259485 675057 259488
rect 412992 256980 416548 259382
rect 423896 256980 424188 259382
rect 674031 259252 674097 259255
rect 674031 259250 674784 259252
rect 674031 259194 674036 259250
rect 674092 259194 674784 259250
rect 674031 259192 674784 259194
rect 674031 259189 674097 259192
rect 677058 258367 677118 258630
rect 677058 258362 677169 258367
rect 677058 258306 677108 258362
rect 677164 258306 677169 258362
rect 677058 258304 677169 258306
rect 677103 258301 677169 258304
rect 676866 257775 676926 258112
rect 676866 257770 676977 257775
rect 676866 257714 676916 257770
rect 676972 257714 676977 257770
rect 676866 257712 676977 257714
rect 676911 257709 676977 257712
rect 677058 257331 677118 257594
rect 676911 257328 676977 257331
rect 676866 257326 676977 257328
rect 676866 257270 676916 257326
rect 676972 257270 676977 257326
rect 676866 257265 676977 257270
rect 677058 257326 677169 257331
rect 677058 257270 677108 257326
rect 677164 257270 677169 257326
rect 677058 257268 677169 257270
rect 677103 257265 677169 257268
rect 676866 257002 676926 257265
rect 412992 256884 424188 256980
rect 206844 256796 209180 256878
rect 412810 256870 424188 256884
rect 46191 256736 46257 256739
rect 40386 256734 46257 256736
rect 40386 256706 46196 256734
rect 40416 256678 46196 256706
rect 46252 256678 46257 256734
rect 40416 256676 46257 256678
rect 46191 256673 46257 256676
rect 206446 256362 211188 256376
rect 206446 256326 211020 256362
rect 42159 255996 42225 255999
rect 42306 255998 42366 256262
rect 42298 255996 42304 255998
rect 42159 255994 42304 255996
rect 42159 255938 42164 255994
rect 42220 255938 42304 255994
rect 42159 255936 42304 255938
rect 42159 255933 42225 255936
rect 42298 255934 42304 255936
rect 42368 255934 42374 255998
rect 40578 255406 40638 255670
rect 40570 255342 40576 255406
rect 40640 255342 40646 255406
rect 43023 255108 43089 255111
rect 42528 255106 43089 255108
rect 42528 255050 43028 255106
rect 43084 255050 43089 255106
rect 42528 255048 43089 255050
rect 43023 255045 43089 255048
rect 40386 254222 40446 254560
rect 40378 254158 40384 254222
rect 40448 254158 40454 254222
rect 40770 253778 40830 254042
rect 40762 253714 40768 253778
rect 40832 253714 40838 253778
rect 41154 253334 41214 253450
rect 41146 253270 41152 253334
rect 41216 253270 41222 253334
rect 206446 253276 206478 256326
rect 208996 253276 211020 256326
rect 211164 253276 211188 256362
rect 413090 256348 424314 256438
rect 212034 255407 212094 255880
rect 211983 255402 212094 255407
rect 211983 255346 211988 255402
rect 212044 255346 212094 255402
rect 211983 255344 212094 255346
rect 211983 255341 212049 255344
rect 206446 253250 211188 253276
rect 413090 253274 413114 256348
rect 413240 256270 424314 256348
rect 413240 253412 416506 256270
rect 424074 253412 424314 256270
rect 684932 254958 685646 254996
rect 413240 253274 424314 253412
rect 413090 253256 424314 253274
rect 669318 254778 685834 254958
rect 41922 252595 41982 252932
rect 669318 252610 685012 254778
rect 41871 252590 41982 252595
rect 41871 252534 41876 252590
rect 41932 252534 41982 252590
rect 41871 252532 41982 252534
rect 41871 252529 41937 252532
rect 40962 252150 41022 252414
rect 641196 252276 656316 252608
rect 669318 252276 671666 252610
rect 641196 252222 671666 252276
rect 40954 252086 40960 252150
rect 41024 252086 41030 252150
rect 41346 251706 41406 251822
rect 41338 251642 41344 251706
rect 41408 251642 41414 251706
rect 40194 250967 40254 251304
rect 40143 250962 40254 250967
rect 40143 250906 40148 250962
rect 40204 250906 40254 250962
rect 40143 250904 40254 250906
rect 40143 250901 40209 250904
rect 40194 250523 40254 250786
rect 40194 250518 40305 250523
rect 40194 250462 40244 250518
rect 40300 250462 40305 250518
rect 40194 250460 40305 250462
rect 40239 250457 40305 250460
rect 40002 249931 40062 250194
rect 39951 249926 40062 249931
rect 39951 249870 39956 249926
rect 40012 249870 40062 249926
rect 39951 249868 40062 249870
rect 39951 249865 40017 249868
rect 39810 249339 39870 249676
rect 39810 249334 39921 249339
rect 39810 249278 39860 249334
rect 39916 249278 39921 249334
rect 39810 249276 39921 249278
rect 39855 249273 39921 249276
rect 206991 249336 207057 249339
rect 211842 249336 211902 249896
rect 206991 249334 211902 249336
rect 206991 249278 206996 249334
rect 207052 249278 211902 249334
rect 641196 249864 641918 252222
rect 655400 249928 671666 252222
rect 684932 251802 685012 252610
rect 685600 252610 685834 254778
rect 685600 251802 685772 252610
rect 684932 251722 685772 251802
rect 675898 251642 675904 251706
rect 675968 251704 675974 251706
rect 677583 251704 677649 251707
rect 675968 251702 677649 251704
rect 675968 251646 677588 251702
rect 677644 251646 677649 251702
rect 675968 251644 677649 251646
rect 675968 251642 675974 251644
rect 677583 251641 677649 251644
rect 675706 251494 675712 251558
rect 675776 251556 675782 251558
rect 677199 251556 677265 251559
rect 675776 251554 677265 251556
rect 675776 251498 677204 251554
rect 677260 251498 677265 251554
rect 675776 251496 677265 251498
rect 675776 251494 675782 251496
rect 677199 251493 677265 251496
rect 655400 249864 656316 249928
rect 641196 249286 656316 249864
rect 206991 249276 211902 249278
rect 206991 249273 207057 249276
rect 40002 248895 40062 249158
rect 40002 248890 40113 248895
rect 40002 248834 40052 248890
rect 40108 248834 40113 248890
rect 40002 248832 40113 248834
rect 40047 248829 40113 248832
rect 42114 248303 42174 248566
rect 42063 248298 42174 248303
rect 42063 248242 42068 248298
rect 42124 248242 42174 248298
rect 42063 248240 42174 248242
rect 42063 248237 42129 248240
rect 42498 247708 42558 248048
rect 410746 247794 410752 247858
rect 410816 247856 410822 247858
rect 411514 247856 411520 247858
rect 410816 247796 411520 247856
rect 410816 247794 410822 247796
rect 411514 247794 411520 247796
rect 411584 247794 411590 247858
rect 53295 247708 53361 247711
rect 196815 247708 196881 247711
rect 42498 247648 42750 247708
rect 35202 247267 35262 247530
rect 35151 247262 35262 247267
rect 42690 247264 42750 247648
rect 53295 247706 196881 247708
rect 53295 247650 53300 247706
rect 53356 247650 196820 247706
rect 196876 247650 196881 247706
rect 53295 247648 196881 247650
rect 53295 247645 53361 247648
rect 196815 247645 196881 247648
rect 407482 247646 407488 247710
rect 407552 247708 407558 247710
rect 408442 247708 408448 247710
rect 407552 247648 408448 247708
rect 407552 247646 407558 247648
rect 408442 247646 408448 247648
rect 408512 247646 408518 247710
rect 408634 247646 408640 247710
rect 408704 247708 408710 247710
rect 411130 247708 411136 247710
rect 408704 247648 411136 247708
rect 408704 247646 408710 247648
rect 411130 247646 411136 247648
rect 411200 247646 411206 247710
rect 175503 247560 175569 247563
rect 407290 247560 407296 247562
rect 175503 247558 243006 247560
rect 175503 247502 175508 247558
rect 175564 247502 243006 247558
rect 175503 247500 243006 247502
rect 175503 247497 175569 247500
rect 181263 247412 181329 247415
rect 242946 247412 243006 247500
rect 243138 247500 243966 247560
rect 243138 247412 243198 247500
rect 243906 247412 243966 247500
rect 244098 247500 407296 247560
rect 244098 247412 244158 247500
rect 407290 247498 407296 247500
rect 407360 247498 407366 247562
rect 409786 247498 409792 247562
rect 409856 247560 409862 247562
rect 412143 247560 412209 247563
rect 409856 247558 412209 247560
rect 409856 247502 412148 247558
rect 412204 247502 412209 247558
rect 409856 247500 412209 247502
rect 409856 247498 409862 247500
rect 412143 247497 412209 247500
rect 410362 247412 410368 247414
rect 181263 247410 242814 247412
rect 181263 247354 181268 247410
rect 181324 247354 242814 247410
rect 181263 247352 242814 247354
rect 242946 247352 243198 247412
rect 243330 247352 243774 247412
rect 243906 247352 244158 247412
rect 244290 247352 410368 247412
rect 181263 247349 181329 247352
rect 35151 247206 35156 247262
rect 35212 247206 35262 247262
rect 35151 247204 35262 247206
rect 42498 247204 42750 247264
rect 163983 247264 164049 247267
rect 181455 247264 181521 247267
rect 163983 247262 181521 247264
rect 163983 247206 163988 247262
rect 164044 247206 181460 247262
rect 181516 247206 181521 247262
rect 163983 247204 181521 247206
rect 35151 247201 35217 247204
rect 42498 246823 42558 247204
rect 163983 247201 164049 247204
rect 181455 247201 181521 247204
rect 197199 247264 197265 247267
rect 242754 247264 242814 247352
rect 243330 247264 243390 247352
rect 197199 247262 240510 247264
rect 197199 247206 197204 247262
rect 197260 247206 240510 247262
rect 197199 247204 240510 247206
rect 242754 247204 243390 247264
rect 243714 247264 243774 247352
rect 244290 247264 244350 247352
rect 410362 247350 410368 247352
rect 410432 247350 410438 247414
rect 411322 247350 411328 247414
rect 411392 247412 411398 247414
rect 412431 247412 412497 247415
rect 411392 247410 412497 247412
rect 411392 247354 412436 247410
rect 412492 247354 412497 247410
rect 411392 247352 412497 247354
rect 411392 247350 411398 247352
rect 412431 247349 412497 247352
rect 407098 247264 407104 247266
rect 243714 247204 244350 247264
rect 246210 247204 407104 247264
rect 197199 247201 197265 247204
rect 189999 247116 190065 247119
rect 209871 247116 209937 247119
rect 189999 247114 209937 247116
rect 189999 247058 190004 247114
rect 190060 247058 209876 247114
rect 209932 247058 209937 247114
rect 189999 247056 209937 247058
rect 189999 247053 190065 247056
rect 209871 247053 209937 247056
rect 211599 247116 211665 247119
rect 211599 247114 239934 247116
rect 211599 247058 211604 247114
rect 211660 247058 239934 247114
rect 211599 247056 239934 247058
rect 211599 247053 211665 247056
rect 207226 246906 207232 246970
rect 207296 246968 207302 246970
rect 207296 246908 226686 246968
rect 207296 246906 207302 246908
rect 35151 246820 35217 246823
rect 35151 246818 35262 246820
rect 35151 246762 35156 246818
rect 35212 246762 35262 246818
rect 35151 246757 35262 246762
rect 42447 246818 42558 246823
rect 42447 246762 42452 246818
rect 42508 246762 42558 246818
rect 42447 246760 42558 246762
rect 42447 246757 42513 246760
rect 42874 246758 42880 246822
rect 42944 246820 42950 246822
rect 209967 246820 210033 246823
rect 42944 246818 210033 246820
rect 42944 246762 209972 246818
rect 210028 246762 210033 246818
rect 42944 246760 210033 246762
rect 42944 246758 42950 246760
rect 209967 246757 210033 246760
rect 210255 246820 210321 246823
rect 226383 246820 226449 246823
rect 210255 246818 226449 246820
rect 210255 246762 210260 246818
rect 210316 246762 226388 246818
rect 226444 246762 226449 246818
rect 210255 246760 226449 246762
rect 226626 246820 226686 246908
rect 227202 246908 237774 246968
rect 227202 246820 227262 246908
rect 237714 246823 237774 246908
rect 226626 246760 227262 246820
rect 227343 246820 227409 246823
rect 237039 246820 237105 246823
rect 227343 246818 237105 246820
rect 227343 246762 227348 246818
rect 227404 246762 237044 246818
rect 237100 246762 237105 246818
rect 227343 246760 237105 246762
rect 210255 246757 210321 246760
rect 226383 246757 226449 246760
rect 227343 246757 227409 246760
rect 237039 246757 237105 246760
rect 237711 246818 237777 246823
rect 237711 246762 237716 246818
rect 237772 246762 237777 246818
rect 237711 246757 237777 246762
rect 239874 246820 239934 247056
rect 240450 246823 240510 247204
rect 246210 246968 246270 247204
rect 407098 247202 407104 247204
rect 407168 247202 407174 247266
rect 407290 247202 407296 247266
rect 407360 247264 407366 247266
rect 409978 247264 409984 247266
rect 407360 247204 409984 247264
rect 407360 247202 407366 247204
rect 409978 247202 409984 247204
rect 410048 247202 410054 247266
rect 410170 247202 410176 247266
rect 410240 247264 410246 247266
rect 412047 247264 412113 247267
rect 410240 247262 412113 247264
rect 410240 247206 412052 247262
rect 412108 247206 412113 247262
rect 410240 247204 412113 247206
rect 410240 247202 410246 247204
rect 412047 247201 412113 247204
rect 405754 247116 405760 247118
rect 241746 246908 246270 246968
rect 246402 247056 405760 247116
rect 241746 246823 241806 246908
rect 240015 246820 240081 246823
rect 239874 246818 240081 246820
rect 239874 246762 240020 246818
rect 240076 246762 240081 246818
rect 239874 246760 240081 246762
rect 240450 246818 240561 246823
rect 240450 246762 240500 246818
rect 240556 246762 240561 246818
rect 240450 246760 240561 246762
rect 240015 246757 240081 246760
rect 240495 246757 240561 246760
rect 241743 246818 241809 246823
rect 241743 246762 241748 246818
rect 241804 246762 241809 246818
rect 241743 246757 241809 246762
rect 242511 246820 242577 246823
rect 246402 246820 246462 247056
rect 405754 247054 405760 247056
rect 405824 247054 405830 247118
rect 410554 247116 410560 247118
rect 405954 247056 410560 247116
rect 405954 246968 406014 247056
rect 410554 247054 410560 247056
rect 410624 247054 410630 247118
rect 410746 247054 410752 247118
rect 410816 247116 410822 247118
rect 412239 247116 412305 247119
rect 410816 247114 412305 247116
rect 410816 247058 412244 247114
rect 412300 247058 412305 247114
rect 410816 247056 412305 247058
rect 410816 247054 410822 247056
rect 412239 247053 412305 247056
rect 406714 246968 406720 246970
rect 252546 246908 292014 246968
rect 252546 246823 252606 246908
rect 291954 246823 292014 246908
rect 292290 246908 388590 246968
rect 292290 246823 292350 246908
rect 388530 246823 388590 246908
rect 389634 246908 406014 246968
rect 406098 246908 406720 246968
rect 242511 246818 246462 246820
rect 242511 246762 242516 246818
rect 242572 246762 246462 246818
rect 242511 246760 246462 246762
rect 252495 246818 252606 246823
rect 252495 246762 252500 246818
rect 252556 246762 252606 246818
rect 252495 246760 252606 246762
rect 252687 246820 252753 246823
rect 266703 246820 266769 246823
rect 252687 246818 266769 246820
rect 252687 246762 252692 246818
rect 252748 246762 266708 246818
rect 266764 246762 266769 246818
rect 252687 246760 266769 246762
rect 242511 246757 242577 246760
rect 252495 246757 252561 246760
rect 252687 246757 252753 246760
rect 266703 246757 266769 246760
rect 268623 246820 268689 246823
rect 286095 246820 286161 246823
rect 268623 246818 286161 246820
rect 268623 246762 268628 246818
rect 268684 246762 286100 246818
rect 286156 246762 286161 246818
rect 268623 246760 286161 246762
rect 268623 246757 268689 246760
rect 286095 246757 286161 246760
rect 286287 246820 286353 246823
rect 288879 246820 288945 246823
rect 286287 246818 288945 246820
rect 286287 246762 286292 246818
rect 286348 246762 288884 246818
rect 288940 246762 288945 246818
rect 286287 246760 288945 246762
rect 286287 246757 286353 246760
rect 288879 246757 288945 246760
rect 291951 246818 292017 246823
rect 291951 246762 291956 246818
rect 292012 246762 292017 246818
rect 291951 246757 292017 246762
rect 292239 246818 292350 246823
rect 292239 246762 292244 246818
rect 292300 246762 292350 246818
rect 292239 246760 292350 246762
rect 292623 246820 292689 246823
rect 387375 246820 387441 246823
rect 292623 246818 387441 246820
rect 292623 246762 292628 246818
rect 292684 246762 387380 246818
rect 387436 246762 387441 246818
rect 292623 246760 387441 246762
rect 292239 246757 292305 246760
rect 292623 246757 292689 246760
rect 387375 246757 387441 246760
rect 388527 246818 388593 246823
rect 388527 246762 388532 246818
rect 388588 246762 388593 246818
rect 388527 246757 388593 246762
rect 389487 246820 389553 246823
rect 389634 246820 389694 246908
rect 406098 246823 406158 246908
rect 406714 246906 406720 246908
rect 406784 246906 406790 246970
rect 407290 246968 407296 246970
rect 407058 246908 407296 246968
rect 406462 246834 406614 246844
rect 389487 246818 389694 246820
rect 389487 246762 389492 246818
rect 389548 246762 389694 246818
rect 389487 246760 389694 246762
rect 389775 246820 389841 246823
rect 405903 246820 405969 246823
rect 389775 246818 405969 246820
rect 389775 246762 389780 246818
rect 389836 246762 405908 246818
rect 405964 246762 405969 246818
rect 389775 246760 405969 246762
rect 389487 246757 389553 246760
rect 389775 246757 389841 246760
rect 405903 246757 405969 246760
rect 406095 246818 406161 246823
rect 406095 246762 406100 246818
rect 406156 246762 406161 246818
rect 406095 246757 406161 246762
rect 406462 246758 406520 246834
rect 406598 246758 406614 246834
rect 407058 246823 407118 246908
rect 407290 246906 407296 246908
rect 407360 246906 407366 246970
rect 408826 246968 408832 246970
rect 407682 246908 408832 246968
rect 407682 246823 407742 246908
rect 408826 246906 408832 246908
rect 408896 246906 408902 246970
rect 410938 246968 410944 246970
rect 408978 246908 410944 246968
rect 408978 246823 409038 246908
rect 410938 246906 410944 246908
rect 411008 246906 411014 246970
rect 35202 246420 35262 246757
rect 406462 246746 406614 246758
rect 406767 246820 406833 246823
rect 406906 246820 406912 246822
rect 406767 246818 406912 246820
rect 406767 246762 406772 246818
rect 406828 246762 406912 246818
rect 406767 246760 406912 246762
rect 406767 246757 406833 246760
rect 406906 246758 406912 246760
rect 406976 246758 406982 246822
rect 407055 246818 407121 246823
rect 407055 246762 407060 246818
rect 407116 246762 407121 246818
rect 407055 246757 407121 246762
rect 407247 246820 407313 246823
rect 407482 246820 407488 246822
rect 407247 246818 407488 246820
rect 407247 246762 407252 246818
rect 407308 246762 407488 246818
rect 407247 246760 407488 246762
rect 407247 246757 407313 246760
rect 407482 246758 407488 246760
rect 407552 246758 407558 246822
rect 407631 246818 407742 246823
rect 408111 246822 408177 246823
rect 407631 246762 407636 246818
rect 407692 246762 407742 246818
rect 407631 246760 407742 246762
rect 407631 246757 407697 246760
rect 408058 246758 408064 246822
rect 408128 246820 408177 246822
rect 408128 246818 408220 246820
rect 408172 246762 408220 246818
rect 408128 246760 408220 246762
rect 408128 246758 408177 246760
rect 408442 246758 408448 246822
rect 408512 246820 408518 246822
rect 408591 246820 408657 246823
rect 408783 246822 408849 246823
rect 408783 246820 408832 246822
rect 408512 246818 408657 246820
rect 408512 246762 408596 246818
rect 408652 246762 408657 246818
rect 408512 246760 408657 246762
rect 408740 246818 408832 246820
rect 408740 246762 408788 246818
rect 408740 246760 408832 246762
rect 408512 246758 408518 246760
rect 408111 246757 408177 246758
rect 408591 246757 408657 246760
rect 408783 246758 408832 246760
rect 408896 246758 408902 246822
rect 408975 246818 409041 246823
rect 409167 246822 409233 246823
rect 409167 246820 409216 246822
rect 408975 246762 408980 246818
rect 409036 246762 409041 246818
rect 408783 246757 408849 246758
rect 408975 246757 409041 246762
rect 409124 246818 409216 246820
rect 409124 246762 409172 246818
rect 409124 246760 409216 246762
rect 409167 246758 409216 246760
rect 409280 246758 409286 246822
rect 409359 246820 409425 246823
rect 409594 246820 409600 246822
rect 409359 246818 409600 246820
rect 409359 246762 409364 246818
rect 409420 246762 409600 246818
rect 409359 246760 409600 246762
rect 409167 246757 409233 246758
rect 409359 246757 409425 246760
rect 409594 246758 409600 246760
rect 409664 246758 409670 246822
rect 409839 246820 409905 246823
rect 674554 246820 674560 246822
rect 409839 246818 674560 246820
rect 409839 246762 409844 246818
rect 409900 246762 674560 246818
rect 409839 246760 674560 246762
rect 409839 246757 409905 246760
rect 674554 246758 674560 246760
rect 674624 246758 674630 246822
rect 172719 246672 172785 246675
rect 211599 246672 211665 246675
rect 172719 246670 211665 246672
rect 172719 246614 172724 246670
rect 172780 246614 211604 246670
rect 211660 246614 211665 246670
rect 172719 246612 211665 246614
rect 172719 246609 172785 246612
rect 211599 246609 211665 246612
rect 53583 246524 53649 246527
rect 187695 246524 187761 246527
rect 211023 246524 211089 246527
rect 53583 246522 187761 246524
rect 53583 246466 53588 246522
rect 53644 246466 187700 246522
rect 187756 246466 187761 246522
rect 53583 246464 187761 246466
rect 53583 246461 53649 246464
rect 187695 246461 187761 246464
rect 187842 246522 211089 246524
rect 187842 246466 211028 246522
rect 211084 246466 211089 246522
rect 187842 246464 211089 246466
rect 65103 246376 65169 246379
rect 187842 246376 187902 246464
rect 211023 246461 211089 246464
rect 209775 246376 209841 246379
rect 65103 246374 187902 246376
rect 65103 246318 65108 246374
rect 65164 246318 187902 246374
rect 65103 246316 187902 246318
rect 191490 246374 209841 246376
rect 191490 246318 209780 246374
rect 209836 246318 209841 246374
rect 191490 246316 209841 246318
rect 65103 246313 65169 246316
rect 44559 246228 44625 246231
rect 191490 246228 191550 246316
rect 209775 246313 209841 246316
rect 44559 246226 191550 246228
rect 44559 246170 44564 246226
rect 44620 246170 191550 246226
rect 44559 246168 191550 246170
rect 197583 246228 197649 246231
rect 207226 246228 207232 246230
rect 197583 246226 207232 246228
rect 197583 246170 197588 246226
rect 197644 246170 207232 246226
rect 197583 246168 207232 246170
rect 44559 246165 44625 246168
rect 197583 246165 197649 246168
rect 207226 246166 207232 246168
rect 207296 246166 207302 246230
rect 60495 246080 60561 246083
rect 66255 246080 66321 246083
rect 60495 246078 66321 246080
rect 60495 246022 60500 246078
rect 60556 246022 66260 246078
rect 66316 246022 66321 246078
rect 60495 246020 66321 246022
rect 60495 246017 60561 246020
rect 66255 246017 66321 246020
rect 187023 246080 187089 246083
rect 197199 246080 197265 246083
rect 187023 246078 197265 246080
rect 187023 246022 187028 246078
rect 187084 246022 197204 246078
rect 197260 246022 197265 246078
rect 187023 246020 197265 246022
rect 187023 246017 187089 246020
rect 197199 246017 197265 246020
rect 674554 245870 674560 245934
rect 674624 245932 674630 245934
rect 675183 245932 675249 245935
rect 674624 245930 675249 245932
rect 674624 245874 675188 245930
rect 675244 245874 675249 245930
rect 674624 245872 675249 245874
rect 674624 245870 674630 245872
rect 675183 245869 675249 245872
rect 149583 245784 149649 245787
rect 210831 245784 210897 245787
rect 149583 245782 210897 245784
rect 149583 245726 149588 245782
rect 149644 245726 210836 245782
rect 210892 245726 210897 245782
rect 149583 245724 210897 245726
rect 149583 245721 149649 245724
rect 210831 245721 210897 245724
rect 187695 245636 187761 245639
rect 209967 245636 210033 245639
rect 187695 245634 210033 245636
rect 187695 245578 187700 245634
rect 187756 245578 209972 245634
rect 210028 245578 210033 245634
rect 187695 245576 210033 245578
rect 187695 245573 187761 245576
rect 209967 245573 210033 245576
rect 155343 245488 155409 245491
rect 210543 245488 210609 245491
rect 155343 245486 210609 245488
rect 155343 245430 155348 245486
rect 155404 245430 210548 245486
rect 210604 245430 210609 245486
rect 155343 245428 210609 245430
rect 155343 245425 155409 245428
rect 210543 245425 210609 245428
rect 158319 245192 158385 245195
rect 210255 245192 210321 245195
rect 158319 245190 210321 245192
rect 158319 245134 158324 245190
rect 158380 245134 210260 245190
rect 210316 245134 210321 245190
rect 158319 245132 210321 245134
rect 158319 245129 158385 245132
rect 210255 245129 210321 245132
rect 41530 244982 41536 245046
rect 41600 245044 41606 245046
rect 42874 245044 42880 245046
rect 41600 244984 42880 245044
rect 41600 244982 41606 244984
rect 42874 244982 42880 244984
rect 42944 244982 42950 245046
rect 161103 245044 161169 245047
rect 210063 245044 210129 245047
rect 161103 245042 210129 245044
rect 161103 244986 161108 245042
rect 161164 244986 210068 245042
rect 210124 244986 210129 245042
rect 161103 244984 210129 244986
rect 161103 244981 161169 244984
rect 210063 244981 210129 244984
rect 40143 244896 40209 244899
rect 41722 244896 41728 244898
rect 40143 244894 41728 244896
rect 40143 244838 40148 244894
rect 40204 244838 41728 244894
rect 40143 244836 41728 244838
rect 40143 244833 40209 244836
rect 41722 244834 41728 244836
rect 41792 244834 41798 244898
rect 166863 244896 166929 244899
rect 210063 244896 210129 244899
rect 166863 244894 210129 244896
rect 166863 244838 166868 244894
rect 166924 244838 210068 244894
rect 210124 244838 210129 244894
rect 166863 244836 210129 244838
rect 166863 244833 166929 244836
rect 210063 244833 210129 244836
rect 675375 244750 675441 244751
rect 674362 244686 674368 244750
rect 674432 244748 674438 244750
rect 675322 244748 675328 244750
rect 674432 244688 675328 244748
rect 675392 244746 675441 244750
rect 675436 244690 675441 244746
rect 674432 244686 674438 244688
rect 675322 244686 675328 244688
rect 675392 244686 675441 244690
rect 675375 244685 675441 244686
rect 41914 243798 41920 243862
rect 41984 243860 41990 243862
rect 43119 243860 43185 243863
rect 275586 243860 276030 243897
rect 297090 243860 297534 243897
rect 674362 243860 674368 243862
rect 41984 243858 674368 243860
rect 41984 243802 43124 243858
rect 43180 243837 674368 243858
rect 43180 243802 275646 243837
rect 41984 243800 275646 243802
rect 275970 243800 297150 243837
rect 297474 243800 674368 243837
rect 41984 243798 41990 243800
rect 43119 243797 43185 243800
rect 674362 243798 674368 243800
rect 674432 243798 674438 243862
rect 209967 243712 210033 243715
rect 211023 243714 211089 243715
rect 210298 243712 210304 243714
rect 209967 243710 210304 243712
rect 209967 243654 209972 243710
rect 210028 243654 210304 243710
rect 209967 243652 210304 243654
rect 209967 243649 210033 243652
rect 210298 243650 210304 243652
rect 210368 243650 210374 243714
rect 211023 243710 211072 243714
rect 211136 243712 211142 243714
rect 211503 243712 211569 243715
rect 225999 243712 226065 243715
rect 211023 243654 211028 243710
rect 211023 243650 211072 243654
rect 211136 243652 211180 243712
rect 211503 243710 226065 243712
rect 211503 243654 211508 243710
rect 211564 243654 226004 243710
rect 226060 243654 226065 243710
rect 211503 243652 226065 243654
rect 211136 243650 211142 243652
rect 211023 243649 211089 243650
rect 211503 243649 211569 243652
rect 225999 243649 226065 243652
rect 227439 243712 227505 243715
rect 648015 243712 648081 243715
rect 227439 243710 648081 243712
rect 227439 243654 227444 243710
rect 227500 243654 648020 243710
rect 648076 243654 648081 243710
rect 227439 243652 648081 243654
rect 227439 243649 227505 243652
rect 648015 243649 648081 243652
rect 178383 243564 178449 243567
rect 389295 243564 389361 243567
rect 405562 243564 405568 243566
rect 178383 243562 389118 243564
rect 178383 243506 178388 243562
rect 178444 243506 389118 243562
rect 178383 243504 389118 243506
rect 178383 243501 178449 243504
rect 206607 243416 206673 243419
rect 256047 243416 256113 243419
rect 206607 243414 256113 243416
rect 206607 243358 206612 243414
rect 206668 243358 256052 243414
rect 256108 243358 256113 243414
rect 206607 243356 256113 243358
rect 206607 243353 206673 243356
rect 256047 243353 256113 243356
rect 256239 243416 256305 243419
rect 389058 243416 389118 243504
rect 389295 243562 405568 243564
rect 389295 243506 389300 243562
rect 389356 243506 405568 243562
rect 389295 243504 405568 243506
rect 389295 243501 389361 243504
rect 405562 243502 405568 243504
rect 405632 243502 405638 243566
rect 405711 243564 405777 243567
rect 405946 243564 405952 243566
rect 405711 243562 405952 243564
rect 405711 243506 405716 243562
rect 405772 243506 405952 243562
rect 405711 243504 405952 243506
rect 405711 243501 405777 243504
rect 405946 243502 405952 243504
rect 406016 243502 406022 243566
rect 406191 243564 406257 243567
rect 408250 243564 408256 243566
rect 406191 243562 408256 243564
rect 406191 243506 406196 243562
rect 406252 243506 408256 243562
rect 406191 243504 408256 243506
rect 406191 243501 406257 243504
rect 408250 243502 408256 243504
rect 408320 243502 408326 243566
rect 674170 243502 674176 243566
rect 674240 243564 674246 243566
rect 675471 243564 675537 243567
rect 674240 243562 675537 243564
rect 674240 243506 675476 243562
rect 675532 243506 675537 243562
rect 674240 243504 675537 243506
rect 674240 243502 674246 243504
rect 675471 243501 675537 243504
rect 406330 243416 406336 243418
rect 256239 243414 388926 243416
rect 256239 243358 256244 243414
rect 256300 243358 388926 243414
rect 256239 243356 388926 243358
rect 389058 243356 406336 243416
rect 256239 243353 256305 243356
rect 210639 243268 210705 243271
rect 221199 243268 221265 243271
rect 210639 243266 221265 243268
rect 210639 243210 210644 243266
rect 210700 243210 221204 243266
rect 221260 243210 221265 243266
rect 210639 243208 221265 243210
rect 210639 243205 210705 243208
rect 221199 243205 221265 243208
rect 221391 243268 221457 243271
rect 228207 243268 228273 243271
rect 221391 243266 228273 243268
rect 221391 243210 221396 243266
rect 221452 243210 228212 243266
rect 228268 243210 228273 243266
rect 221391 243208 228273 243210
rect 221391 243205 221457 243208
rect 228207 243205 228273 243208
rect 256239 243268 256305 243271
rect 256527 243268 256593 243271
rect 256239 243266 256593 243268
rect 256239 243210 256244 243266
rect 256300 243210 256532 243266
rect 256588 243210 256593 243266
rect 256239 243208 256593 243210
rect 256239 243205 256305 243208
rect 256527 243205 256593 243208
rect 276399 243268 276465 243271
rect 316527 243268 316593 243271
rect 276399 243266 316593 243268
rect 276399 243210 276404 243266
rect 276460 243210 316532 243266
rect 316588 243210 316593 243266
rect 276399 243208 316593 243210
rect 276399 243205 276465 243208
rect 316527 243205 316593 243208
rect 331119 243268 331185 243271
rect 388866 243268 388926 243356
rect 406330 243354 406336 243356
rect 406400 243354 406406 243418
rect 407674 243268 407680 243270
rect 331119 243266 387198 243268
rect 331119 243210 331124 243266
rect 331180 243210 387198 243266
rect 331119 243208 387198 243210
rect 388866 243208 407680 243268
rect 331119 243205 331185 243208
rect 209775 243120 209841 243123
rect 210682 243120 210688 243122
rect 209775 243118 210688 243120
rect 209775 243062 209780 243118
rect 209836 243062 210688 243118
rect 209775 243060 210688 243062
rect 209775 243057 209841 243060
rect 210682 243058 210688 243060
rect 210752 243058 210758 243122
rect 214959 243120 215025 243123
rect 256335 243120 256401 243123
rect 214959 243118 256401 243120
rect 214959 243062 214964 243118
rect 215020 243062 256340 243118
rect 256396 243062 256401 243118
rect 214959 243060 256401 243062
rect 214959 243057 215025 243060
rect 256335 243057 256401 243060
rect 256719 243120 256785 243123
rect 352239 243120 352305 243123
rect 256719 243118 352305 243120
rect 256719 243062 256724 243118
rect 256780 243062 352244 243118
rect 352300 243062 352305 243118
rect 256719 243060 352305 243062
rect 256719 243057 256785 243060
rect 352239 243057 352305 243060
rect 213231 242972 213297 242975
rect 306447 242972 306513 242975
rect 213231 242970 306513 242972
rect 213231 242914 213236 242970
rect 213292 242914 306452 242970
rect 306508 242914 306513 242970
rect 213231 242912 306513 242914
rect 213231 242909 213297 242912
rect 306447 242909 306513 242912
rect 316719 242972 316785 242975
rect 325071 242972 325137 242975
rect 342063 242972 342129 242975
rect 316719 242970 325137 242972
rect 316719 242914 316724 242970
rect 316780 242914 325076 242970
rect 325132 242914 325137 242970
rect 316719 242912 325137 242914
rect 316719 242909 316785 242912
rect 325071 242909 325137 242912
rect 328578 242970 342129 242972
rect 328578 242914 342068 242970
rect 342124 242914 342129 242970
rect 328578 242912 342129 242914
rect 387138 242972 387198 243208
rect 407674 243206 407680 243208
rect 407744 243206 407750 243270
rect 406138 242972 406144 242974
rect 387138 242912 406144 242972
rect 218895 242824 218961 242827
rect 237711 242824 237777 242827
rect 314991 242824 315057 242827
rect 218895 242822 237630 242824
rect 218895 242766 218900 242822
rect 218956 242766 237630 242822
rect 218895 242764 237630 242766
rect 218895 242761 218961 242764
rect 220815 242676 220881 242679
rect 237423 242676 237489 242679
rect 220815 242674 237489 242676
rect 220815 242618 220820 242674
rect 220876 242618 237428 242674
rect 237484 242618 237489 242674
rect 220815 242616 237489 242618
rect 237570 242676 237630 242764
rect 237711 242822 315057 242824
rect 237711 242766 237716 242822
rect 237772 242766 314996 242822
rect 315052 242766 315057 242822
rect 237711 242764 315057 242766
rect 237711 242761 237777 242764
rect 314991 242761 315057 242764
rect 316719 242824 316785 242827
rect 328578 242824 328638 242912
rect 342063 242909 342129 242912
rect 406138 242910 406144 242912
rect 406208 242910 406214 242974
rect 316719 242822 328638 242824
rect 316719 242766 316724 242822
rect 316780 242766 328638 242822
rect 316719 242764 328638 242766
rect 316719 242761 316785 242764
rect 328762 242762 328768 242826
rect 328832 242824 328838 242826
rect 342927 242824 342993 242827
rect 328832 242822 342993 242824
rect 328832 242766 342932 242822
rect 342988 242766 342993 242822
rect 328832 242764 342993 242766
rect 328832 242762 328838 242764
rect 342927 242761 342993 242764
rect 341199 242676 341265 242679
rect 237570 242674 341265 242676
rect 237570 242618 341204 242674
rect 341260 242618 341265 242674
rect 237570 242616 341265 242618
rect 220815 242613 220881 242616
rect 237423 242613 237489 242616
rect 341199 242613 341265 242616
rect 453615 242676 453681 242679
rect 463695 242676 463761 242679
rect 453615 242674 463761 242676
rect 453615 242618 453620 242674
rect 453676 242618 463700 242674
rect 463756 242618 463761 242674
rect 453615 242616 463761 242618
rect 453615 242613 453681 242616
rect 463695 242613 463761 242616
rect 42159 242528 42225 242531
rect 43503 242528 43569 242531
rect 247503 242528 247569 242531
rect 42159 242526 247569 242528
rect 42159 242470 42164 242526
rect 42220 242470 43508 242526
rect 43564 242470 247508 242526
rect 247564 242470 247569 242526
rect 42159 242468 247569 242470
rect 42159 242465 42225 242468
rect 43503 242465 43569 242468
rect 247503 242465 247569 242468
rect 247695 242528 247761 242531
rect 310479 242528 310545 242531
rect 328143 242528 328209 242531
rect 247695 242526 310398 242528
rect 247695 242470 247700 242526
rect 247756 242470 310398 242526
rect 247695 242468 310398 242470
rect 247695 242465 247761 242468
rect 227727 242380 227793 242383
rect 310191 242380 310257 242383
rect 227727 242378 310257 242380
rect 227727 242322 227732 242378
rect 227788 242322 310196 242378
rect 310252 242322 310257 242378
rect 227727 242320 310257 242322
rect 310338 242380 310398 242468
rect 310479 242526 328209 242528
rect 310479 242470 310484 242526
rect 310540 242470 328148 242526
rect 328204 242470 328209 242526
rect 310479 242468 328209 242470
rect 310479 242465 310545 242468
rect 328143 242465 328209 242468
rect 339759 242528 339825 242531
rect 430479 242528 430545 242531
rect 339759 242526 430545 242528
rect 339759 242470 339764 242526
rect 339820 242470 430484 242526
rect 430540 242470 430545 242526
rect 339759 242468 430545 242470
rect 339759 242465 339825 242468
rect 430479 242465 430545 242468
rect 443439 242528 443505 242531
rect 443631 242528 443697 242531
rect 443439 242526 443697 242528
rect 443439 242470 443444 242526
rect 443500 242470 443636 242526
rect 443692 242470 443697 242526
rect 443439 242468 443697 242470
rect 443439 242465 443505 242468
rect 443631 242465 443697 242468
rect 483759 242528 483825 242531
rect 489519 242528 489585 242531
rect 483759 242526 489585 242528
rect 483759 242470 483764 242526
rect 483820 242470 489524 242526
rect 489580 242470 489585 242526
rect 483759 242468 489585 242470
rect 483759 242465 483825 242468
rect 489519 242465 489585 242468
rect 328378 242380 328384 242382
rect 310338 242320 328384 242380
rect 227727 242317 227793 242320
rect 310191 242317 310257 242320
rect 328378 242318 328384 242320
rect 328448 242318 328454 242382
rect 328527 242380 328593 242383
rect 338991 242380 339057 242383
rect 328527 242378 339057 242380
rect 328527 242322 328532 242378
rect 328588 242322 338996 242378
rect 339052 242322 339057 242378
rect 328527 242320 339057 242322
rect 328527 242317 328593 242320
rect 338991 242317 339057 242320
rect 339567 242380 339633 242383
rect 344271 242380 344337 242383
rect 339567 242378 344337 242380
rect 339567 242322 339572 242378
rect 339628 242322 344276 242378
rect 344332 242322 344337 242378
rect 339567 242320 344337 242322
rect 339567 242317 339633 242320
rect 344271 242317 344337 242320
rect 489711 242380 489777 242383
rect 504015 242380 504081 242383
rect 489711 242378 504081 242380
rect 489711 242322 489716 242378
rect 489772 242322 504020 242378
rect 504076 242322 504081 242378
rect 489711 242320 504081 242322
rect 489711 242317 489777 242320
rect 504015 242317 504081 242320
rect 42063 242084 42129 242087
rect 42447 242084 42513 242087
rect 42063 242082 42513 242084
rect 42063 242026 42068 242082
rect 42124 242026 42452 242082
rect 42508 242026 42513 242082
rect 42063 242024 42513 242026
rect 140802 242084 140862 242276
rect 196815 242232 196881 242235
rect 212026 242232 212032 242234
rect 196815 242230 212032 242232
rect 196815 242174 196820 242230
rect 196876 242174 212032 242230
rect 196815 242172 212032 242174
rect 196815 242169 196881 242172
rect 212026 242170 212032 242172
rect 212096 242170 212102 242234
rect 223695 242232 223761 242235
rect 343407 242232 343473 242235
rect 223695 242230 343473 242232
rect 223695 242174 223700 242230
rect 223756 242174 343412 242230
rect 343468 242174 343473 242230
rect 223695 242172 343473 242174
rect 223695 242169 223761 242172
rect 343407 242169 343473 242172
rect 145402 242084 145408 242086
rect 140802 242024 145408 242084
rect 42063 242021 42129 242024
rect 42447 242021 42513 242024
rect 145402 242022 145408 242024
rect 145472 242022 145478 242086
rect 217167 242084 217233 242087
rect 227343 242084 227409 242087
rect 217167 242082 227409 242084
rect 217167 242026 217172 242082
rect 217228 242026 227348 242082
rect 227404 242026 227409 242082
rect 217167 242024 227409 242026
rect 217167 242021 217233 242024
rect 227343 242021 227409 242024
rect 228207 242084 228273 242087
rect 354639 242084 354705 242087
rect 228207 242082 354705 242084
rect 228207 242026 228212 242082
rect 228268 242026 354644 242082
rect 354700 242026 354705 242082
rect 228207 242024 354705 242026
rect 228207 242021 228273 242024
rect 354639 242021 354705 242024
rect 673978 242022 673984 242086
rect 674048 242084 674054 242086
rect 675375 242084 675441 242087
rect 674048 242082 675441 242084
rect 674048 242026 675380 242082
rect 675436 242026 675441 242082
rect 674048 242024 675441 242026
rect 674048 242022 674054 242024
rect 675375 242021 675441 242024
rect 211119 241936 211185 241939
rect 287727 241936 287793 241939
rect 308943 241936 309009 241939
rect 576207 241936 576273 241939
rect 211119 241934 277950 241936
rect 211119 241878 211124 241934
rect 211180 241878 277950 241934
rect 211119 241876 277950 241878
rect 211119 241873 211185 241876
rect 245391 241788 245457 241791
rect 277743 241788 277809 241791
rect 245391 241786 277809 241788
rect 245391 241730 245396 241786
rect 245452 241730 277748 241786
rect 277804 241730 277809 241786
rect 245391 241728 277809 241730
rect 277890 241788 277950 241876
rect 287727 241934 309009 241936
rect 287727 241878 287732 241934
rect 287788 241878 308948 241934
rect 309004 241878 309009 241934
rect 287727 241876 309009 241878
rect 287727 241873 287793 241876
rect 308943 241873 309009 241876
rect 316098 241934 576273 241936
rect 316098 241878 576212 241934
rect 576268 241878 576273 241934
rect 316098 241876 576273 241878
rect 316098 241788 316158 241876
rect 576207 241873 576273 241876
rect 277890 241728 316158 241788
rect 318255 241788 318321 241791
rect 356751 241788 356817 241791
rect 318255 241786 356817 241788
rect 318255 241730 318260 241786
rect 318316 241730 356756 241786
rect 356812 241730 356817 241786
rect 318255 241728 356817 241730
rect 245391 241725 245457 241728
rect 277743 241725 277809 241728
rect 318255 241725 318321 241728
rect 356751 241725 356817 241728
rect 246735 241640 246801 241643
rect 354447 241640 354513 241643
rect 246735 241638 354513 241640
rect 246735 241582 246740 241638
rect 246796 241582 354452 241638
rect 354508 241582 354513 241638
rect 246735 241580 354513 241582
rect 246735 241577 246801 241580
rect 354447 241577 354513 241580
rect 261231 241492 261297 241495
rect 372879 241492 372945 241495
rect 261231 241490 372945 241492
rect 261231 241434 261236 241490
rect 261292 241434 372884 241490
rect 372940 241434 372945 241490
rect 261231 241432 372945 241434
rect 261231 241429 261297 241432
rect 372879 241429 372945 241432
rect 244527 241344 244593 241347
rect 271503 241344 271569 241347
rect 244527 241342 271569 241344
rect 244527 241286 244532 241342
rect 244588 241286 271508 241342
rect 271564 241286 271569 241342
rect 244527 241284 271569 241286
rect 244527 241281 244593 241284
rect 271503 241281 271569 241284
rect 277743 241344 277809 241347
rect 289647 241344 289713 241347
rect 277743 241342 289713 241344
rect 277743 241286 277748 241342
rect 277804 241286 289652 241342
rect 289708 241286 289713 241342
rect 277743 241284 289713 241286
rect 277743 241281 277809 241284
rect 289647 241281 289713 241284
rect 289839 241344 289905 241347
rect 297807 241344 297873 241347
rect 289839 241342 297873 241344
rect 289839 241286 289844 241342
rect 289900 241286 297812 241342
rect 297868 241286 297873 241342
rect 289839 241284 297873 241286
rect 289839 241281 289905 241284
rect 297807 241281 297873 241284
rect 297999 241344 298065 241347
rect 358959 241344 359025 241347
rect 297999 241342 359025 241344
rect 297999 241286 298004 241342
rect 298060 241286 358964 241342
rect 359020 241286 359025 241342
rect 297999 241284 359025 241286
rect 297999 241281 298065 241284
rect 358959 241281 359025 241284
rect 259599 241196 259665 241199
rect 376815 241196 376881 241199
rect 259599 241194 376881 241196
rect 259599 241138 259604 241194
rect 259660 241138 376820 241194
rect 376876 241138 376881 241194
rect 259599 241136 376881 241138
rect 259599 241133 259665 241136
rect 376815 241133 376881 241136
rect 140802 240604 140862 241092
rect 243183 241048 243249 241051
rect 271311 241048 271377 241051
rect 243183 241046 271377 241048
rect 243183 240990 243188 241046
rect 243244 240990 271316 241046
rect 271372 240990 271377 241046
rect 243183 240988 271377 240990
rect 243183 240985 243249 240988
rect 271311 240985 271377 240988
rect 271503 241048 271569 241051
rect 297999 241048 298065 241051
rect 271503 241046 298065 241048
rect 271503 240990 271508 241046
rect 271564 240990 298004 241046
rect 298060 240990 298065 241046
rect 271503 240988 298065 240990
rect 271503 240985 271569 240988
rect 297999 240985 298065 240988
rect 298191 241048 298257 241051
rect 361647 241048 361713 241051
rect 298191 241046 361713 241048
rect 298191 240990 298196 241046
rect 298252 240990 361652 241046
rect 361708 240990 361713 241046
rect 298191 240988 361713 240990
rect 298191 240985 298257 240988
rect 361647 240985 361713 240988
rect 259023 240900 259089 240903
rect 377871 240900 377937 240903
rect 259023 240898 377937 240900
rect 259023 240842 259028 240898
rect 259084 240842 377876 240898
rect 377932 240842 377937 240898
rect 259023 240840 377937 240842
rect 259023 240837 259089 240840
rect 377871 240837 377937 240840
rect 242703 240752 242769 240755
rect 278031 240752 278097 240755
rect 289839 240752 289905 240755
rect 363087 240752 363153 240755
rect 242703 240750 277950 240752
rect 242703 240694 242708 240750
rect 242764 240694 277950 240750
rect 242703 240692 277950 240694
rect 242703 240689 242769 240692
rect 146127 240604 146193 240607
rect 140802 240602 146193 240604
rect 140802 240546 146132 240602
rect 146188 240546 146193 240602
rect 140802 240544 146193 240546
rect 146127 240541 146193 240544
rect 241743 240604 241809 240607
rect 277890 240604 277950 240692
rect 278031 240750 289905 240752
rect 278031 240694 278036 240750
rect 278092 240694 289844 240750
rect 289900 240694 289905 240750
rect 278031 240692 289905 240694
rect 278031 240689 278097 240692
rect 289839 240689 289905 240692
rect 289986 240750 363153 240752
rect 289986 240694 363092 240750
rect 363148 240694 363153 240750
rect 289986 240692 363153 240694
rect 289986 240604 290046 240692
rect 363087 240689 363153 240692
rect 364815 240604 364881 240607
rect 241743 240602 277758 240604
rect 241743 240546 241748 240602
rect 241804 240546 277758 240602
rect 241743 240544 277758 240546
rect 277890 240544 290046 240604
rect 293442 240602 364881 240604
rect 293442 240546 364820 240602
rect 364876 240546 364881 240602
rect 293442 240544 364881 240546
rect 241743 240541 241809 240544
rect 240975 240456 241041 240459
rect 271119 240456 271185 240459
rect 240975 240454 271185 240456
rect 240975 240398 240980 240454
rect 241036 240398 271124 240454
rect 271180 240398 271185 240454
rect 240975 240396 271185 240398
rect 240975 240393 241041 240396
rect 271119 240393 271185 240396
rect 271311 240456 271377 240459
rect 277551 240456 277617 240459
rect 271311 240454 277617 240456
rect 271311 240398 271316 240454
rect 271372 240398 277556 240454
rect 277612 240398 277617 240454
rect 271311 240396 277617 240398
rect 277698 240456 277758 240544
rect 293442 240456 293502 240544
rect 364815 240541 364881 240544
rect 277698 240396 293502 240456
rect 297999 240456 298065 240459
rect 366543 240456 366609 240459
rect 297999 240454 366609 240456
rect 297999 240398 298004 240454
rect 298060 240398 366548 240454
rect 366604 240398 366609 240454
rect 297999 240396 366609 240398
rect 271311 240393 271377 240396
rect 277551 240393 277617 240396
rect 297999 240393 298065 240396
rect 366543 240393 366609 240396
rect 367599 240456 367665 240459
rect 409743 240456 409809 240459
rect 367599 240454 409809 240456
rect 367599 240398 367604 240454
rect 367660 240398 409748 240454
rect 409804 240398 409809 240454
rect 367599 240396 409809 240398
rect 367599 240393 367665 240396
rect 409743 240393 409809 240396
rect 262959 240308 263025 240311
rect 369807 240308 369873 240311
rect 262959 240306 369873 240308
rect 262959 240250 262964 240306
rect 263020 240250 369812 240306
rect 369868 240250 369873 240306
rect 262959 240248 369873 240250
rect 262959 240245 263025 240248
rect 369807 240245 369873 240248
rect 247695 240160 247761 240163
rect 352815 240160 352881 240163
rect 247695 240158 352881 240160
rect 247695 240102 247700 240158
rect 247756 240102 352820 240158
rect 352876 240102 352881 240158
rect 247695 240100 352881 240102
rect 247695 240097 247761 240100
rect 352815 240097 352881 240100
rect 247983 240012 248049 240015
rect 351279 240012 351345 240015
rect 247983 240010 351345 240012
rect 247983 239954 247988 240010
rect 248044 239954 351284 240010
rect 351340 239954 351345 240010
rect 247983 239952 351345 239954
rect 247983 239949 248049 239952
rect 351279 239949 351345 239952
rect 146607 239864 146673 239867
rect 140832 239862 146673 239864
rect 140832 239806 146612 239862
rect 146668 239806 146673 239862
rect 140832 239804 146673 239806
rect 146607 239801 146673 239804
rect 269295 239864 269361 239867
rect 278223 239864 278289 239867
rect 269295 239862 278289 239864
rect 269295 239806 269300 239862
rect 269356 239806 278228 239862
rect 278284 239806 278289 239862
rect 269295 239804 278289 239806
rect 269295 239801 269361 239804
rect 278223 239801 278289 239804
rect 289647 239864 289713 239867
rect 318255 239864 318321 239867
rect 289647 239862 318321 239864
rect 289647 239806 289652 239862
rect 289708 239806 318260 239862
rect 318316 239806 318321 239862
rect 289647 239804 318321 239806
rect 289647 239801 289713 239804
rect 318255 239801 318321 239804
rect 271119 239716 271185 239719
rect 297999 239716 298065 239719
rect 271119 239714 298065 239716
rect 271119 239658 271124 239714
rect 271180 239658 298004 239714
rect 298060 239658 298065 239714
rect 271119 239656 298065 239658
rect 271119 239653 271185 239656
rect 297999 239653 298065 239656
rect 277935 239568 278001 239571
rect 279759 239568 279825 239571
rect 277935 239566 279825 239568
rect 277935 239510 277940 239566
rect 277996 239510 279764 239566
rect 279820 239510 279825 239566
rect 277935 239508 279825 239510
rect 277935 239505 278001 239508
rect 279759 239505 279825 239508
rect 287631 239568 287697 239571
rect 293775 239568 293841 239571
rect 287631 239566 293841 239568
rect 287631 239510 287636 239566
rect 287692 239510 293780 239566
rect 293836 239510 293841 239566
rect 287631 239508 293841 239510
rect 287631 239505 287697 239508
rect 293775 239505 293841 239508
rect 293391 239420 293457 239423
rect 305295 239420 305361 239423
rect 293391 239418 305361 239420
rect 293391 239362 293396 239418
rect 293452 239362 305300 239418
rect 305356 239362 305361 239418
rect 293391 239360 305361 239362
rect 293391 239357 293457 239360
rect 305295 239357 305361 239360
rect 293967 239272 294033 239275
rect 296271 239272 296337 239275
rect 293967 239270 296337 239272
rect 293967 239214 293972 239270
rect 294028 239214 296276 239270
rect 296332 239214 296337 239270
rect 293967 239212 296337 239214
rect 293967 239209 294033 239212
rect 296271 239209 296337 239212
rect 209391 239124 209457 239127
rect 351375 239124 351441 239127
rect 209391 239122 351441 239124
rect 209391 239066 209396 239122
rect 209452 239066 351380 239122
rect 351436 239066 351441 239122
rect 209391 239064 351441 239066
rect 209391 239061 209457 239064
rect 351375 239061 351441 239064
rect 211311 238976 211377 238979
rect 547503 238976 547569 238979
rect 211311 238974 547569 238976
rect 211311 238918 211316 238974
rect 211372 238918 547508 238974
rect 547564 238918 547569 238974
rect 211311 238916 547569 238918
rect 211311 238913 211377 238916
rect 547503 238913 547569 238916
rect 675183 238976 675249 238979
rect 675514 238976 675520 238978
rect 675183 238974 675520 238976
rect 675183 238918 675188 238974
rect 675244 238918 675520 238974
rect 675183 238916 675520 238918
rect 675183 238913 675249 238916
rect 675514 238914 675520 238916
rect 675584 238914 675590 238978
rect 211215 238828 211281 238831
rect 412623 238828 412689 238831
rect 211215 238826 412689 238828
rect 211215 238770 211220 238826
rect 211276 238770 412628 238826
rect 412684 238770 412689 238826
rect 211215 238768 412689 238770
rect 211215 238765 211281 238768
rect 412623 238765 412689 238768
rect 144111 238680 144177 238683
rect 140832 238678 144177 238680
rect 140832 238622 144116 238678
rect 144172 238622 144177 238678
rect 140832 238620 144177 238622
rect 144111 238617 144177 238620
rect 243567 238680 243633 238683
rect 360687 238680 360753 238683
rect 675759 238682 675825 238683
rect 243567 238678 360753 238680
rect 243567 238622 243572 238678
rect 243628 238622 360692 238678
rect 360748 238622 360753 238678
rect 243567 238620 360753 238622
rect 243567 238617 243633 238620
rect 360687 238617 360753 238620
rect 675706 238618 675712 238682
rect 675776 238680 675825 238682
rect 675776 238678 675868 238680
rect 675820 238622 675868 238678
rect 675776 238620 675868 238622
rect 675776 238618 675825 238620
rect 675759 238617 675825 238618
rect 241359 238532 241425 238535
rect 241786 238532 241792 238534
rect 241359 238530 241792 238532
rect 241359 238474 241364 238530
rect 241420 238474 241792 238530
rect 241359 238472 241792 238474
rect 241359 238469 241425 238472
rect 241786 238470 241792 238472
rect 241856 238470 241862 238534
rect 242319 238532 242385 238535
rect 363855 238532 363921 238535
rect 242319 238530 363921 238532
rect 242319 238474 242324 238530
rect 242380 238474 363860 238530
rect 363916 238474 363921 238530
rect 242319 238472 363921 238474
rect 242319 238469 242385 238472
rect 363855 238469 363921 238472
rect 42298 238322 42304 238386
rect 42368 238384 42374 238386
rect 42543 238384 42609 238387
rect 42368 238382 42609 238384
rect 42368 238326 42548 238382
rect 42604 238326 42609 238382
rect 42368 238324 42609 238326
rect 42368 238322 42374 238324
rect 42543 238321 42609 238324
rect 258639 238384 258705 238387
rect 378831 238384 378897 238387
rect 258639 238382 378897 238384
rect 258639 238326 258644 238382
rect 258700 238326 378836 238382
rect 378892 238326 378897 238382
rect 258639 238324 378897 238326
rect 258639 238321 258705 238324
rect 378831 238321 378897 238324
rect 215823 238236 215889 238239
rect 215823 238234 231870 238236
rect 215823 238178 215828 238234
rect 215884 238178 231870 238234
rect 215823 238176 231870 238178
rect 215823 238173 215889 238176
rect 215247 238088 215313 238091
rect 231810 238088 231870 238176
rect 241786 238174 241792 238238
rect 241856 238236 241862 238238
rect 365775 238236 365841 238239
rect 241856 238234 365841 238236
rect 241856 238178 365780 238234
rect 365836 238178 365841 238234
rect 241856 238176 365841 238178
rect 241856 238174 241862 238176
rect 365775 238173 365841 238176
rect 391407 238088 391473 238091
rect 215247 238086 217086 238088
rect 215247 238030 215252 238086
rect 215308 238030 217086 238086
rect 215247 238028 217086 238030
rect 231810 238086 391473 238088
rect 231810 238030 391412 238086
rect 391468 238030 391473 238086
rect 231810 238028 391473 238030
rect 215247 238025 215313 238028
rect 214863 237940 214929 237943
rect 217026 237940 217086 238028
rect 391407 238025 391473 238028
rect 393135 237940 393201 237943
rect 214863 237938 216894 237940
rect 214863 237882 214868 237938
rect 214924 237882 216894 237938
rect 214863 237880 216894 237882
rect 217026 237938 393201 237940
rect 217026 237882 393140 237938
rect 393196 237882 393201 237938
rect 217026 237880 393201 237882
rect 214863 237877 214929 237880
rect 157743 237792 157809 237795
rect 211450 237792 211456 237794
rect 157743 237790 211456 237792
rect 157743 237734 157748 237790
rect 157804 237734 211456 237790
rect 157743 237732 211456 237734
rect 157743 237729 157809 237732
rect 211450 237730 211456 237732
rect 211520 237792 211526 237794
rect 216687 237792 216753 237795
rect 211520 237790 216753 237792
rect 211520 237734 216692 237790
rect 216748 237734 216753 237790
rect 211520 237732 216753 237734
rect 216834 237792 216894 237880
rect 393135 237877 393201 237880
rect 394671 237792 394737 237795
rect 216834 237790 394737 237792
rect 216834 237734 394676 237790
rect 394732 237734 394737 237790
rect 216834 237732 394737 237734
rect 211520 237730 211526 237732
rect 216687 237729 216753 237732
rect 394671 237729 394737 237732
rect 511119 237792 511185 237795
rect 676474 237792 676480 237794
rect 511119 237790 676480 237792
rect 511119 237734 511124 237790
rect 511180 237734 676480 237790
rect 511119 237732 676480 237734
rect 511119 237729 511185 237732
rect 676474 237730 676480 237732
rect 676544 237730 676550 237794
rect 142479 237644 142545 237647
rect 209583 237644 209649 237647
rect 214767 237644 214833 237647
rect 142479 237642 214833 237644
rect 142479 237586 142484 237642
rect 142540 237586 209588 237642
rect 209644 237586 214772 237642
rect 214828 237586 214833 237642
rect 142479 237584 214833 237586
rect 142479 237581 142545 237584
rect 209583 237581 209649 237584
rect 214767 237581 214833 237584
rect 216207 237644 216273 237647
rect 411951 237644 412017 237647
rect 216207 237642 412017 237644
rect 216207 237586 216212 237642
rect 216268 237586 411956 237642
rect 412012 237586 412017 237642
rect 216207 237584 412017 237586
rect 216207 237581 216273 237584
rect 411951 237581 412017 237584
rect 505359 237644 505425 237647
rect 677050 237644 677056 237646
rect 505359 237642 677056 237644
rect 505359 237586 505364 237642
rect 505420 237586 677056 237642
rect 505359 237584 677056 237586
rect 505359 237581 505425 237584
rect 677050 237582 677056 237584
rect 677120 237582 677126 237646
rect 243951 237496 244017 237499
rect 360015 237496 360081 237499
rect 243951 237494 360081 237496
rect 243951 237438 243956 237494
rect 244012 237438 360020 237494
rect 360076 237438 360081 237494
rect 243951 237436 360081 237438
rect 243951 237433 244017 237436
rect 360015 237433 360081 237436
rect 140802 236904 140862 237392
rect 243087 237348 243153 237351
rect 358479 237348 358545 237351
rect 243087 237346 358545 237348
rect 243087 237290 243092 237346
rect 243148 237290 358484 237346
rect 358540 237290 358545 237346
rect 243087 237288 358545 237290
rect 243087 237285 243153 237288
rect 358479 237285 358545 237288
rect 245295 237200 245361 237203
rect 357807 237200 357873 237203
rect 245295 237198 357873 237200
rect 245295 237142 245300 237198
rect 245356 237142 357812 237198
rect 357868 237142 357873 237198
rect 245295 237140 357873 237142
rect 245295 237137 245361 237140
rect 357807 237137 357873 237140
rect 319887 237052 319953 237055
rect 338127 237052 338193 237055
rect 319887 237050 338193 237052
rect 319887 236994 319892 237050
rect 319948 236994 338132 237050
rect 338188 236994 338193 237050
rect 319887 236992 338193 236994
rect 319887 236989 319953 236992
rect 338127 236989 338193 236992
rect 146319 236904 146385 236907
rect 140802 236902 146385 236904
rect 140802 236846 146324 236902
rect 146380 236846 146385 236902
rect 140802 236844 146385 236846
rect 146319 236841 146385 236844
rect 329775 236904 329841 236907
rect 339759 236904 339825 236907
rect 329775 236902 339825 236904
rect 329775 236846 329780 236902
rect 329836 236846 339764 236902
rect 339820 236846 339825 236902
rect 329775 236844 339825 236846
rect 329775 236841 329841 236844
rect 339759 236841 339825 236844
rect 675759 236904 675825 236907
rect 675898 236904 675904 236906
rect 675759 236902 675904 236904
rect 675759 236846 675764 236902
rect 675820 236846 675904 236902
rect 675759 236844 675904 236846
rect 675759 236841 675825 236844
rect 675898 236842 675904 236844
rect 675968 236842 675974 236906
rect 209679 236756 209745 236759
rect 212175 236756 212241 236759
rect 227439 236756 227505 236759
rect 209679 236754 212094 236756
rect 209679 236698 209684 236754
rect 209740 236698 212094 236754
rect 209679 236696 212094 236698
rect 209679 236693 209745 236696
rect 212034 236460 212094 236696
rect 212175 236754 227505 236756
rect 212175 236698 212180 236754
rect 212236 236698 227444 236754
rect 227500 236698 227505 236754
rect 212175 236696 227505 236698
rect 212175 236693 212241 236696
rect 227439 236693 227505 236696
rect 227631 236756 227697 236759
rect 239098 236756 239104 236758
rect 227631 236754 239104 236756
rect 227631 236698 227636 236754
rect 227692 236698 239104 236754
rect 227631 236696 239104 236698
rect 227631 236693 227697 236696
rect 239098 236694 239104 236696
rect 239168 236694 239174 236758
rect 259119 236756 259185 236759
rect 400335 236756 400401 236759
rect 259119 236754 400401 236756
rect 259119 236698 259124 236754
rect 259180 236698 400340 236754
rect 400396 236698 400401 236754
rect 259119 236696 400401 236698
rect 259119 236693 259185 236696
rect 400335 236693 400401 236696
rect 420399 236756 420465 236759
rect 440655 236756 440721 236759
rect 420399 236754 440721 236756
rect 420399 236698 420404 236754
rect 420460 236698 440660 236754
rect 440716 236698 440721 236754
rect 420399 236696 440721 236698
rect 420399 236693 420465 236696
rect 440655 236693 440721 236696
rect 460719 236756 460785 236759
rect 480975 236756 481041 236759
rect 460719 236754 481041 236756
rect 460719 236698 460724 236754
rect 460780 236698 480980 236754
rect 481036 236698 481041 236754
rect 460719 236696 481041 236698
rect 460719 236693 460785 236696
rect 480975 236693 481041 236696
rect 214767 236608 214833 236611
rect 359247 236608 359313 236611
rect 214767 236606 359313 236608
rect 214767 236550 214772 236606
rect 214828 236550 359252 236606
rect 359308 236550 359313 236606
rect 214767 236548 359313 236550
rect 214767 236545 214833 236548
rect 359247 236545 359313 236548
rect 420591 236460 420657 236463
rect 212034 236458 420657 236460
rect 212034 236402 420596 236458
rect 420652 236402 420657 236458
rect 212034 236400 420657 236402
rect 420591 236397 420657 236400
rect 144015 236312 144081 236315
rect 140802 236310 144081 236312
rect 140802 236254 144020 236310
rect 144076 236254 144081 236310
rect 140802 236252 144081 236254
rect 140802 236210 140862 236252
rect 144015 236249 144081 236252
rect 239098 236250 239104 236314
rect 239168 236312 239174 236314
rect 259119 236312 259185 236315
rect 239168 236310 259185 236312
rect 239168 236254 259124 236310
rect 259180 236254 259185 236310
rect 239168 236252 259185 236254
rect 239168 236250 239174 236252
rect 259119 236249 259185 236252
rect 288975 236312 289041 236315
rect 294063 236312 294129 236315
rect 288975 236310 294129 236312
rect 288975 236254 288980 236310
rect 289036 236254 294068 236310
rect 294124 236254 294129 236310
rect 288975 236252 294129 236254
rect 288975 236249 289041 236252
rect 294063 236249 294129 236252
rect 638415 236312 638481 236315
rect 639279 236312 639345 236315
rect 638415 236310 639345 236312
rect 638415 236254 638420 236310
rect 638476 236254 639284 236310
rect 639340 236254 639345 236310
rect 638415 236252 639345 236254
rect 638415 236249 638481 236252
rect 639279 236249 639345 236252
rect 676474 236250 676480 236314
rect 676544 236312 676550 236314
rect 676858 236312 676864 236314
rect 676544 236252 676864 236312
rect 676544 236250 676550 236252
rect 676858 236250 676864 236252
rect 676928 236250 676934 236314
rect 225807 236164 225873 236167
rect 344751 236164 344817 236167
rect 225807 236162 344817 236164
rect 225807 236106 225812 236162
rect 225868 236106 344756 236162
rect 344812 236106 344817 236162
rect 225807 236104 344817 236106
rect 225807 236101 225873 236104
rect 344751 236101 344817 236104
rect 229551 236016 229617 236019
rect 345999 236016 346065 236019
rect 229551 236014 346065 236016
rect 229551 235958 229556 236014
rect 229612 235958 346004 236014
rect 346060 235958 346065 236014
rect 229551 235956 346065 235958
rect 229551 235953 229617 235956
rect 345999 235953 346065 235956
rect 221295 235868 221361 235871
rect 342543 235868 342609 235871
rect 221295 235866 342609 235868
rect 221295 235810 221300 235866
rect 221356 235810 342548 235866
rect 342604 235810 342609 235866
rect 221295 235808 342609 235810
rect 221295 235805 221361 235808
rect 342543 235805 342609 235808
rect 219759 235720 219825 235723
rect 341583 235720 341649 235723
rect 219759 235718 341649 235720
rect 219759 235662 219764 235718
rect 219820 235662 341588 235718
rect 341644 235662 341649 235718
rect 219759 235660 341649 235662
rect 219759 235657 219825 235660
rect 341583 235657 341649 235660
rect 223023 235572 223089 235575
rect 343311 235572 343377 235575
rect 223023 235570 343377 235572
rect 223023 235514 223028 235570
rect 223084 235514 343316 235570
rect 343372 235514 343377 235570
rect 223023 235512 343377 235514
rect 223023 235509 223089 235512
rect 343311 235509 343377 235512
rect 224463 235424 224529 235427
rect 343791 235424 343857 235427
rect 224463 235422 343857 235424
rect 224463 235366 224468 235422
rect 224524 235366 343796 235422
rect 343852 235366 343857 235422
rect 224463 235364 343857 235366
rect 224463 235361 224529 235364
rect 343791 235361 343857 235364
rect 218223 235276 218289 235279
rect 341103 235276 341169 235279
rect 218223 235274 341169 235276
rect 218223 235218 218228 235274
rect 218284 235218 341108 235274
rect 341164 235218 341169 235274
rect 218223 235216 341169 235218
rect 218223 235213 218289 235216
rect 341103 235213 341169 235216
rect 146511 235128 146577 235131
rect 140832 235126 146577 235128
rect 140832 235070 146516 235126
rect 146572 235070 146577 235126
rect 140832 235068 146577 235070
rect 146511 235065 146577 235068
rect 212367 235128 212433 235131
rect 334959 235128 335025 235131
rect 212367 235126 335025 235128
rect 212367 235070 212372 235126
rect 212428 235070 334964 235126
rect 335020 235070 335025 235126
rect 212367 235068 335025 235070
rect 212367 235065 212433 235068
rect 334959 235065 335025 235068
rect 214191 234980 214257 234983
rect 348207 234980 348273 234983
rect 214191 234978 348273 234980
rect 214191 234922 214196 234978
rect 214252 234922 348212 234978
rect 348268 234922 348273 234978
rect 214191 234920 348273 234922
rect 214191 234917 214257 234920
rect 348207 234917 348273 234920
rect 210159 234832 210225 234835
rect 379407 234832 379473 234835
rect 210159 234830 379473 234832
rect 210159 234774 210164 234830
rect 210220 234774 379412 234830
rect 379468 234774 379473 234830
rect 210159 234772 379473 234774
rect 210159 234769 210225 234772
rect 379407 234769 379473 234772
rect 211642 234622 211648 234686
rect 211712 234684 211718 234686
rect 547119 234684 547185 234687
rect 211712 234682 547185 234684
rect 211712 234626 547124 234682
rect 547180 234626 547185 234682
rect 211712 234624 547185 234626
rect 211712 234622 211718 234624
rect 547119 234621 547185 234624
rect 238959 234536 239025 234539
rect 349167 234536 349233 234539
rect 238959 234534 349233 234536
rect 238959 234478 238964 234534
rect 239020 234478 349172 234534
rect 349228 234478 349233 234534
rect 238959 234476 349233 234478
rect 238959 234473 239025 234476
rect 349167 234473 349233 234476
rect 238671 234388 238737 234391
rect 347727 234388 347793 234391
rect 238671 234386 347793 234388
rect 238671 234330 238676 234386
rect 238732 234330 347732 234386
rect 347788 234330 347793 234386
rect 238671 234328 347793 234330
rect 238671 234325 238737 234328
rect 347727 234325 347793 234328
rect 42063 234092 42129 234095
rect 42298 234092 42304 234094
rect 42063 234090 42304 234092
rect 42063 234034 42068 234090
rect 42124 234034 42304 234090
rect 42063 234032 42304 234034
rect 42063 234029 42129 234032
rect 42298 234030 42304 234032
rect 42368 234030 42374 234094
rect 210298 233882 210304 233946
rect 210368 233944 210374 233946
rect 212559 233944 212625 233947
rect 210368 233942 212625 233944
rect 210368 233886 212564 233942
rect 212620 233886 212625 233942
rect 210368 233884 212625 233886
rect 210368 233882 210374 233884
rect 212559 233881 212625 233884
rect 636922 233882 636928 233946
rect 636992 233944 636998 233946
rect 638031 233944 638097 233947
rect 636992 233942 638097 233944
rect 636992 233886 638036 233942
rect 638092 233886 638097 233942
rect 636992 233884 638097 233886
rect 636992 233882 636998 233884
rect 638031 233881 638097 233884
rect 140802 233648 140862 233840
rect 210061 233811 210131 233816
rect 211298 233811 211368 233816
rect 210061 233751 210066 233811
rect 210126 233751 211303 233811
rect 211363 233751 211368 233811
rect 210061 233746 210131 233751
rect 211298 233746 211368 233751
rect 212026 233734 212032 233798
rect 212096 233796 212102 233798
rect 212271 233796 212337 233799
rect 212986 233796 212992 233798
rect 212096 233794 212992 233796
rect 212096 233738 212276 233794
rect 212332 233738 212992 233794
rect 212096 233736 212992 233738
rect 212096 233734 212102 233736
rect 212271 233733 212337 233736
rect 212986 233734 212992 233736
rect 213056 233734 213062 233798
rect 637690 233734 637696 233798
rect 637760 233796 637766 233798
rect 638799 233796 638865 233799
rect 637760 233794 638865 233796
rect 637760 233738 638804 233794
rect 638860 233738 638865 233794
rect 637760 233736 638865 233738
rect 637760 233734 637766 233736
rect 638799 233733 638865 233736
rect 144015 233648 144081 233651
rect 140802 233646 144081 233648
rect 140802 233590 144020 233646
rect 144076 233590 144081 233646
rect 140802 233588 144081 233590
rect 144015 233585 144081 233588
rect 210682 233586 210688 233650
rect 210752 233648 210758 233650
rect 212079 233648 212145 233651
rect 212559 233650 212625 233651
rect 637167 233650 637233 233651
rect 212559 233648 212608 233650
rect 210752 233646 212430 233648
rect 210752 233590 212084 233646
rect 212140 233590 212430 233646
rect 210752 233588 212430 233590
rect 212516 233646 212608 233648
rect 212516 233590 212564 233646
rect 212516 233588 212608 233590
rect 210752 233586 210758 233588
rect 212079 233585 212145 233588
rect 211066 233438 211072 233502
rect 211136 233500 211142 233502
rect 211695 233500 211761 233503
rect 212218 233500 212224 233502
rect 211136 233498 212224 233500
rect 211136 233442 211700 233498
rect 211756 233442 212224 233498
rect 211136 233440 212224 233442
rect 211136 233438 211142 233440
rect 211695 233437 211761 233440
rect 212218 233438 212224 233440
rect 212288 233438 212294 233502
rect 212370 233500 212430 233588
rect 212559 233586 212608 233588
rect 212672 233586 212678 233650
rect 637114 233648 637120 233650
rect 637076 233588 637120 233648
rect 637184 233646 637233 233650
rect 637228 233590 637233 233646
rect 637114 233586 637120 233588
rect 637184 233586 637233 233590
rect 637498 233586 637504 233650
rect 637568 233648 637574 233650
rect 638895 233648 638961 233651
rect 637568 233646 638961 233648
rect 637568 233590 638900 233646
rect 638956 233590 638961 233646
rect 671682 233636 708937 233637
rect 637568 233588 638961 233590
rect 637568 233586 637574 233588
rect 212559 233585 212625 233586
rect 637167 233585 637233 233586
rect 638895 233585 638961 233588
rect 212794 233500 212800 233502
rect 212370 233440 212800 233500
rect 212794 233438 212800 233440
rect 212864 233438 212870 233502
rect 214287 233498 214353 233503
rect 214287 233442 214292 233498
rect 214348 233442 214353 233498
rect 214287 233437 214353 233442
rect 290895 233500 290961 233503
rect 298191 233500 298257 233503
rect 290895 233498 298257 233500
rect 290895 233442 290900 233498
rect 290956 233442 298196 233498
rect 298252 233442 298257 233498
rect 290895 233440 298257 233442
rect 290895 233437 290961 233440
rect 298191 233437 298257 233440
rect 637306 233438 637312 233502
rect 637376 233500 637382 233502
rect 637455 233500 637521 233503
rect 637376 233498 637521 233500
rect 637376 233442 637460 233498
rect 637516 233442 637521 233498
rect 637376 233440 637521 233442
rect 637376 233438 637382 233440
rect 637455 233437 637521 233440
rect 637882 233438 637888 233502
rect 637952 233500 637958 233502
rect 638223 233500 638289 233503
rect 637952 233498 638289 233500
rect 637952 233442 638228 233498
rect 638284 233442 638289 233498
rect 637952 233440 638289 233442
rect 637952 233438 637958 233440
rect 638223 233437 638289 233440
rect 41146 233290 41152 233354
rect 41216 233352 41222 233354
rect 41775 233352 41841 233355
rect 41216 233350 41841 233352
rect 41216 233294 41780 233350
rect 41836 233294 41841 233350
rect 41216 233292 41841 233294
rect 41216 233290 41222 233292
rect 41775 233289 41841 233292
rect 210682 233290 210688 233354
rect 210752 233352 210758 233354
rect 214290 233352 214350 233437
rect 210752 233292 214350 233352
rect 210752 233290 210758 233292
rect 205071 232760 205137 232763
rect 645807 232760 645873 232763
rect 205071 232758 210558 232760
rect 205071 232702 205076 232758
rect 205132 232702 210558 232758
rect 205071 232700 210558 232702
rect 205071 232697 205137 232700
rect 210498 232656 210558 232700
rect 640386 232758 645873 232760
rect 640386 232702 645812 232758
rect 645868 232702 645873 232758
rect 640386 232700 645873 232702
rect 640386 232656 640446 232700
rect 645807 232697 645873 232700
rect 140802 232168 140862 232656
rect 671677 232544 671683 233636
rect 672775 232544 708937 233636
rect 671682 232543 708937 232544
rect 710031 232543 710037 233637
rect 144111 232168 144177 232171
rect 140802 232166 144177 232168
rect 140802 232110 144116 232166
rect 144172 232110 144177 232166
rect 140802 232108 144177 232110
rect 144111 232105 144177 232108
rect 204687 232168 204753 232171
rect 207951 232168 208017 232171
rect 204687 232166 210528 232168
rect 204687 232110 204692 232166
rect 204748 232110 207956 232166
rect 208012 232110 210528 232166
rect 204687 232108 210528 232110
rect 204687 232105 204753 232108
rect 207951 232105 208017 232108
rect 640386 232020 640446 232138
rect 645711 232020 645777 232023
rect 640386 232018 645777 232020
rect 640386 231962 645716 232018
rect 645772 231962 645777 232018
rect 640386 231960 645777 231962
rect 645711 231957 645777 231960
rect 41530 231662 41536 231726
rect 41600 231724 41606 231726
rect 41775 231724 41841 231727
rect 41600 231722 41841 231724
rect 41600 231666 41780 231722
rect 41836 231666 41841 231722
rect 41600 231664 41841 231666
rect 41600 231662 41606 231664
rect 41775 231661 41841 231664
rect 204783 231576 204849 231579
rect 209295 231576 209361 231579
rect 645231 231576 645297 231579
rect 204783 231574 210528 231576
rect 204783 231518 204788 231574
rect 204844 231518 209300 231574
rect 209356 231518 210528 231574
rect 204783 231516 210528 231518
rect 640416 231574 645297 231576
rect 640416 231518 645236 231574
rect 645292 231518 645297 231574
rect 640416 231516 645297 231518
rect 204783 231513 204849 231516
rect 209295 231513 209361 231516
rect 645231 231513 645297 231516
rect 666066 231435 698422 231436
rect 144015 231428 144081 231431
rect 140832 231426 144081 231428
rect 140832 231370 144020 231426
rect 144076 231370 144081 231426
rect 140832 231368 144081 231370
rect 144015 231365 144081 231368
rect 41967 231134 42033 231135
rect 41914 231070 41920 231134
rect 41984 231132 42033 231134
rect 645135 231132 645201 231135
rect 41984 231130 42076 231132
rect 42028 231074 42076 231130
rect 41984 231072 42076 231074
rect 640386 231130 645201 231132
rect 640386 231074 645140 231130
rect 645196 231074 645201 231130
rect 640386 231072 645201 231074
rect 41984 231070 42033 231072
rect 41967 231069 42033 231070
rect 204879 230984 204945 230987
rect 204879 230982 210528 230984
rect 204879 230926 204884 230982
rect 204940 230926 210528 230982
rect 640386 230954 640446 231072
rect 645135 231069 645201 231072
rect 204879 230924 210528 230926
rect 204879 230921 204945 230924
rect 645327 230688 645393 230691
rect 640194 230686 645393 230688
rect 640194 230630 645332 230686
rect 645388 230630 645393 230686
rect 640194 230628 645393 230630
rect 205455 230540 205521 230543
rect 209487 230540 209553 230543
rect 205455 230538 210528 230540
rect 205455 230482 205460 230538
rect 205516 230482 209492 230538
rect 209548 230482 210528 230538
rect 640194 230510 640254 230628
rect 645327 230625 645393 230628
rect 205455 230480 210528 230482
rect 205455 230477 205521 230480
rect 209487 230477 209553 230480
rect 41775 230394 41841 230395
rect 41722 230392 41728 230394
rect 41684 230332 41728 230392
rect 41792 230390 41841 230394
rect 41836 230334 41841 230390
rect 41722 230330 41728 230332
rect 41792 230330 41841 230334
rect 41775 230329 41841 230330
rect 666061 230253 666067 231435
rect 667249 230253 698422 231435
rect 666066 230252 698422 230253
rect 699606 230252 709750 231436
rect 144207 230244 144273 230247
rect 140832 230242 144273 230244
rect 140832 230186 144212 230242
rect 144268 230186 144273 230242
rect 140832 230184 144273 230186
rect 144207 230181 144273 230184
rect 41338 229738 41344 229802
rect 41408 229800 41414 229802
rect 41775 229800 41841 229803
rect 41408 229798 41841 229800
rect 41408 229742 41780 229798
rect 41836 229742 41841 229798
rect 41408 229740 41841 229742
rect 41408 229738 41414 229740
rect 41775 229737 41841 229740
rect 207087 229800 207153 229803
rect 210498 229800 210558 229918
rect 207087 229798 210558 229800
rect 207087 229742 207092 229798
rect 207148 229742 210558 229798
rect 207087 229740 210558 229742
rect 207087 229737 207153 229740
rect 206031 229356 206097 229359
rect 206031 229354 210528 229356
rect 206031 229298 206036 229354
rect 206092 229298 210528 229354
rect 206031 229296 210528 229298
rect 206031 229293 206097 229296
rect 40762 228998 40768 229062
rect 40832 229060 40838 229062
rect 41775 229060 41841 229063
rect 40832 229058 41841 229060
rect 40832 229002 41780 229058
rect 41836 229002 41841 229058
rect 40832 229000 41841 229002
rect 40832 228998 40838 229000
rect 41775 228997 41841 229000
rect 140802 228468 140862 228956
rect 210159 228912 210225 228915
rect 210159 228910 210528 228912
rect 210159 228854 210164 228910
rect 210220 228854 210528 228910
rect 210159 228852 210528 228854
rect 210159 228849 210225 228852
rect 144111 228468 144177 228471
rect 140802 228466 144177 228468
rect 140802 228410 144116 228466
rect 144172 228410 144177 228466
rect 140802 228408 144177 228410
rect 144111 228405 144177 228408
rect 204591 228320 204657 228323
rect 204591 228318 210528 228320
rect 204591 228262 204596 228318
rect 204652 228262 210528 228318
rect 204591 228260 210528 228262
rect 204591 228257 204657 228260
rect 140802 227876 140862 227914
rect 144015 227876 144081 227879
rect 140802 227874 144081 227876
rect 140802 227818 144020 227874
rect 144076 227818 144081 227874
rect 662173 227873 662179 229055
rect 663361 229000 663367 229055
rect 663361 227873 707214 229000
rect 140802 227816 144081 227818
rect 662472 227816 707214 227873
rect 708398 227816 709618 229000
rect 144015 227813 144081 227816
rect 204495 227728 204561 227731
rect 204495 227726 210528 227728
rect 204495 227670 204500 227726
rect 204556 227670 210528 227726
rect 204495 227668 210528 227670
rect 204495 227665 204561 227668
rect 641087 227314 641093 227365
rect 40570 227222 40576 227286
rect 40640 227284 40646 227286
rect 41775 227284 41841 227287
rect 40640 227282 41841 227284
rect 40640 227226 41780 227282
rect 41836 227226 41841 227282
rect 40640 227224 41841 227226
rect 40640 227222 40646 227224
rect 41775 227221 41841 227224
rect 205647 227284 205713 227287
rect 205647 227282 210528 227284
rect 205647 227226 205652 227282
rect 205708 227226 210528 227282
rect 205647 227224 210528 227226
rect 205647 227221 205713 227224
rect 40954 226630 40960 226694
rect 41024 226692 41030 226694
rect 41775 226692 41841 226695
rect 146799 226692 146865 226695
rect 41024 226690 41841 226692
rect 41024 226634 41780 226690
rect 41836 226634 41841 226690
rect 41024 226632 41841 226634
rect 140832 226690 146865 226692
rect 140832 226634 146804 226690
rect 146860 226634 146865 226690
rect 140832 226632 146865 226634
rect 41024 226630 41030 226632
rect 41775 226629 41841 226632
rect 146799 226629 146865 226632
rect 205167 226692 205233 226695
rect 205167 226690 210528 226692
rect 205167 226634 205172 226690
rect 205228 226634 210528 226690
rect 205167 226632 210528 226634
rect 205167 226629 205233 226632
rect 641018 226130 641093 227314
rect 205359 226100 205425 226103
rect 205359 226098 210528 226100
rect 205359 226042 205364 226098
rect 205420 226042 210528 226098
rect 205359 226040 210528 226042
rect 205359 226037 205425 226040
rect 40378 225890 40384 225954
rect 40448 225952 40454 225954
rect 41775 225952 41841 225955
rect 40448 225950 41841 225952
rect 40448 225894 41780 225950
rect 41836 225894 41841 225950
rect 40448 225892 41841 225894
rect 40448 225890 40454 225892
rect 41775 225889 41841 225892
rect 205551 225656 205617 225659
rect 205551 225654 210528 225656
rect 205551 225598 205556 225654
rect 205612 225598 210528 225654
rect 205551 225596 210528 225598
rect 205551 225593 205617 225596
rect 140802 225064 140862 225466
rect 641087 225131 641093 226130
rect 643327 227314 643333 227365
rect 643327 226130 699854 227314
rect 701038 226130 709224 227314
rect 643327 225131 643333 226130
rect 146799 225064 146865 225067
rect 140802 225062 146865 225064
rect 140802 225006 146804 225062
rect 146860 225006 146865 225062
rect 140802 225004 146865 225006
rect 146799 225001 146865 225004
rect 204975 225064 205041 225067
rect 674703 225064 674769 225067
rect 204975 225062 210528 225064
rect 204975 225006 204980 225062
rect 205036 225006 210528 225062
rect 204975 225004 210528 225006
rect 674703 225062 674814 225064
rect 674703 225006 674708 225062
rect 674764 225006 674814 225062
rect 204975 225001 205041 225004
rect 674703 225001 674814 225006
rect 674754 224886 674814 225001
rect 206799 224472 206865 224475
rect 206799 224470 210528 224472
rect 206799 224414 206804 224470
rect 206860 224414 210528 224470
rect 206799 224412 210528 224414
rect 206799 224409 206865 224412
rect 674415 224324 674481 224327
rect 674415 224322 674784 224324
rect 674415 224266 674420 224322
rect 674476 224266 674784 224322
rect 674415 224264 674784 224266
rect 674415 224261 674481 224264
rect 6672 223084 8730 223884
rect 9530 223883 44490 223884
rect 9530 223085 43691 223883
rect 44489 223085 44495 223883
rect 140802 223732 140862 224220
rect 199695 224028 199761 224031
rect 674703 224028 674769 224031
rect 199695 224026 210528 224028
rect 199695 223970 199700 224026
rect 199756 223970 210528 224026
rect 199695 223968 210528 223970
rect 674703 224026 674814 224028
rect 674703 223970 674708 224026
rect 674764 223970 674814 224026
rect 199695 223965 199761 223968
rect 674703 223965 674814 223970
rect 674754 223776 674814 223965
rect 144399 223732 144465 223735
rect 140802 223730 144465 223732
rect 140802 223674 144404 223730
rect 144460 223674 144465 223730
rect 140802 223672 144465 223674
rect 144399 223669 144465 223672
rect 677434 223522 677440 223586
rect 677504 223522 677510 223586
rect 201711 223436 201777 223439
rect 201711 223434 210528 223436
rect 201711 223378 201716 223434
rect 201772 223378 210528 223434
rect 201711 223376 210528 223378
rect 201711 223373 201777 223376
rect 677442 223258 677502 223522
rect 9530 223084 44490 223085
rect 146799 222992 146865 222995
rect 140832 222990 146865 222992
rect 140832 222934 146804 222990
rect 146860 222934 146865 222990
rect 140832 222932 146865 222934
rect 146799 222929 146865 222932
rect 201615 222844 201681 222847
rect 201615 222842 210528 222844
rect 201615 222786 201620 222842
rect 201676 222786 210528 222842
rect 201615 222784 210528 222786
rect 201615 222781 201681 222784
rect 6714 221940 16292 222740
rect 17092 222739 47736 222740
rect 17092 221941 46937 222739
rect 47735 221941 47741 222739
rect 677050 222486 677056 222550
rect 677120 222486 677126 222550
rect 206991 222400 207057 222403
rect 206991 222398 210528 222400
rect 206991 222342 206996 222398
rect 207052 222342 210528 222398
rect 206991 222340 210528 222342
rect 206991 222337 207057 222340
rect 677058 222148 677118 222486
rect 677442 222402 677502 222666
rect 677434 222338 677440 222402
rect 677504 222338 677510 222402
rect 17092 221940 47736 221941
rect 146703 221808 146769 221811
rect 140832 221806 146769 221808
rect 140832 221750 146708 221806
rect 146764 221750 146769 221806
rect 140832 221748 146769 221750
rect 146703 221745 146769 221748
rect 201807 221808 201873 221811
rect 201807 221806 210528 221808
rect 201807 221750 201812 221806
rect 201868 221750 210528 221806
rect 201807 221748 210528 221750
rect 201807 221745 201873 221748
rect 6730 220730 7364 221530
rect 8164 221529 49518 221530
rect 8164 220731 48719 221529
rect 49517 220731 49523 221529
rect 676866 221366 676926 221630
rect 676858 221302 676864 221366
rect 676928 221364 676934 221366
rect 677242 221364 677248 221366
rect 676928 221304 677248 221364
rect 676928 221302 676934 221304
rect 677242 221302 677248 221304
rect 677312 221302 677318 221366
rect 198831 221216 198897 221219
rect 198831 221214 210528 221216
rect 198831 221158 198836 221214
rect 198892 221158 210528 221214
rect 198831 221156 210528 221158
rect 198831 221153 198897 221156
rect 674946 220923 675006 221038
rect 674946 220918 675057 220923
rect 674946 220862 674996 220918
rect 675052 220862 675057 220918
rect 674946 220860 675057 220862
rect 674991 220857 675057 220860
rect 8164 220730 49518 220731
rect 210159 220698 210225 220701
rect 210159 220696 210528 220698
rect 6688 219456 17702 220256
rect 18502 220255 51402 220256
rect 18502 219457 50603 220255
rect 51401 219457 51407 220255
rect 140802 220180 140862 220668
rect 210159 220640 210164 220696
rect 210220 220640 210528 220696
rect 210159 220638 210528 220640
rect 210159 220635 210225 220638
rect 674170 220488 674176 220552
rect 674240 220550 674246 220552
rect 674240 220490 674784 220550
rect 674240 220488 674246 220490
rect 144399 220180 144465 220183
rect 140802 220178 144465 220180
rect 140802 220122 144404 220178
rect 144460 220122 144465 220178
rect 140802 220120 144465 220122
rect 144399 220117 144465 220120
rect 201711 220180 201777 220183
rect 201711 220178 210528 220180
rect 201711 220122 201716 220178
rect 201772 220122 210528 220178
rect 201711 220120 210528 220122
rect 201711 220117 201777 220120
rect 675522 219739 675582 220002
rect 675471 219734 675582 219739
rect 675471 219678 675476 219734
rect 675532 219678 675582 219734
rect 675471 219676 675582 219678
rect 675471 219673 675537 219676
rect 201615 219588 201681 219591
rect 201615 219586 210528 219588
rect 201615 219530 201620 219586
rect 201676 219530 210528 219586
rect 201615 219528 210528 219530
rect 201615 219525 201681 219528
rect 18502 219456 51402 219457
rect 140802 218996 140862 219482
rect 196047 219440 196113 219443
rect 196047 219438 210558 219440
rect 196047 219382 196052 219438
rect 196108 219382 210558 219438
rect 196047 219380 210558 219382
rect 196047 219377 196113 219380
rect 210498 219040 210558 219380
rect 675138 219295 675198 219410
rect 675087 219290 675198 219295
rect 675087 219234 675092 219290
rect 675148 219234 675198 219290
rect 675087 219232 675198 219234
rect 675087 219229 675153 219232
rect 145594 218996 145600 218998
rect 140802 218936 145600 218996
rect 145594 218934 145600 218936
rect 145664 218934 145670 218998
rect 677058 218703 677118 218892
rect 677058 218698 677169 218703
rect 677058 218642 677108 218698
rect 677164 218642 677169 218698
rect 677058 218640 677169 218642
rect 677103 218637 677169 218640
rect 200655 218552 200721 218555
rect 200655 218550 210528 218552
rect 200655 218494 200660 218550
rect 200716 218494 210528 218550
rect 200655 218492 210528 218494
rect 200655 218489 200721 218492
rect 146799 218256 146865 218259
rect 140832 218254 146865 218256
rect 140832 218198 146804 218254
rect 146860 218198 146865 218254
rect 140832 218196 146865 218198
rect 146799 218193 146865 218196
rect 677250 218111 677310 218374
rect 677199 218106 677310 218111
rect 677199 218050 677204 218106
rect 677260 218050 677310 218106
rect 677199 218048 677310 218050
rect 677199 218045 677265 218048
rect 201711 217960 201777 217963
rect 201711 217958 210528 217960
rect 201711 217902 201716 217958
rect 201772 217902 210528 217958
rect 201711 217900 210528 217902
rect 201711 217897 201777 217900
rect 675330 217667 675390 217782
rect 675279 217662 675390 217667
rect 675279 217606 675284 217662
rect 675340 217606 675390 217662
rect 675279 217604 675390 217606
rect 675279 217601 675345 217604
rect 210159 217442 210225 217445
rect 210159 217440 210528 217442
rect 210159 217384 210164 217440
rect 210220 217384 210528 217440
rect 210159 217382 210528 217384
rect 210159 217379 210225 217382
rect 674946 217075 675006 217264
rect 674895 217070 675006 217075
rect 42447 216480 42513 216483
rect 140802 216480 140862 217034
rect 674895 217014 674900 217070
rect 674956 217014 675006 217070
rect 674895 217012 675006 217014
rect 674895 217009 674961 217012
rect 201615 216924 201681 216927
rect 201615 216922 210528 216924
rect 201615 216866 201620 216922
rect 201676 216866 210528 216922
rect 201615 216864 210528 216866
rect 201615 216861 201681 216864
rect 145786 216480 145792 216482
rect 42447 216478 42558 216480
rect 42447 216422 42452 216478
rect 42508 216422 42558 216478
rect 42447 216417 42558 216422
rect 140802 216420 145792 216480
rect 145786 216418 145792 216420
rect 145856 216418 145862 216482
rect 674511 216480 674577 216483
rect 674754 216480 674814 216746
rect 674511 216478 674814 216480
rect 674511 216422 674516 216478
rect 674572 216422 674814 216478
rect 674511 216420 674814 216422
rect 674511 216417 674577 216420
rect 42498 216302 42558 216417
rect 206703 216332 206769 216335
rect 206703 216330 210528 216332
rect 206703 216274 206708 216330
rect 206764 216274 210528 216330
rect 206703 216272 210528 216274
rect 206703 216269 206769 216272
rect 676866 216039 676926 216154
rect 676866 216034 676977 216039
rect 676866 215978 676916 216034
rect 676972 215978 676977 216034
rect 676866 215976 676977 215978
rect 676911 215973 676977 215976
rect 210159 215814 210225 215817
rect 210159 215812 210528 215814
rect 42831 215740 42897 215743
rect 42528 215738 42897 215740
rect 42528 215682 42836 215738
rect 42892 215682 42897 215738
rect 42528 215680 42897 215682
rect 42831 215677 42897 215680
rect 140802 215296 140862 215784
rect 210159 215756 210164 215812
rect 210220 215756 210528 215812
rect 210159 215754 210528 215756
rect 210159 215751 210225 215754
rect 674511 215444 674577 215447
rect 674754 215444 674814 215562
rect 674511 215442 674814 215444
rect 674511 215386 674516 215442
rect 674572 215386 674814 215442
rect 674511 215384 674814 215386
rect 674511 215381 674577 215384
rect 144207 215296 144273 215299
rect 140802 215294 144273 215296
rect 140802 215238 144212 215294
rect 144268 215238 144273 215294
rect 140802 215236 144273 215238
rect 144207 215233 144273 215236
rect 201711 215296 201777 215299
rect 201711 215294 210528 215296
rect 201711 215238 201716 215294
rect 201772 215238 210528 215294
rect 201711 215236 210528 215238
rect 201711 215233 201777 215236
rect 42831 215222 42897 215225
rect 42528 215220 42897 215222
rect 42528 215164 42836 215220
rect 42892 215164 42897 215220
rect 42528 215162 42897 215164
rect 42831 215159 42897 215162
rect 674754 214855 674814 215118
rect 674754 214850 674865 214855
rect 674754 214794 674804 214850
rect 674860 214794 674865 214850
rect 674754 214792 674865 214794
rect 674799 214789 674865 214792
rect 206415 214704 206481 214707
rect 206415 214702 210528 214704
rect 206415 214646 206420 214702
rect 206476 214646 210528 214702
rect 206415 214644 210528 214646
rect 206415 214641 206481 214644
rect 145978 214556 145984 214558
rect 140832 214496 145984 214556
rect 145978 214494 145984 214496
rect 146048 214494 146054 214558
rect 205935 214556 206001 214559
rect 205935 214554 210558 214556
rect 205935 214498 205940 214554
rect 205996 214498 210558 214554
rect 205935 214496 210558 214498
rect 205935 214493 206001 214496
rect 210498 214156 210558 214496
rect 674754 214411 674814 214526
rect 674703 214406 674814 214411
rect 674703 214350 674708 214406
rect 674764 214350 674814 214406
rect 674703 214348 674814 214350
rect 674703 214345 674769 214348
rect 43215 214112 43281 214115
rect 42528 214110 43281 214112
rect 42528 214054 43220 214110
rect 43276 214054 43281 214110
rect 42528 214052 43281 214054
rect 43215 214049 43281 214052
rect 674607 213816 674673 213819
rect 674754 213816 674814 213934
rect 674607 213814 674814 213816
rect 674607 213758 674612 213814
rect 674668 213758 674814 213814
rect 674607 213756 674814 213758
rect 674607 213753 674673 213756
rect 43407 213668 43473 213671
rect 42498 213666 43473 213668
rect 42498 213610 43412 213666
rect 43468 213610 43473 213666
rect 42498 213608 43473 213610
rect 42498 213490 42558 213608
rect 43407 213605 43473 213608
rect 206319 213668 206385 213671
rect 206319 213666 210528 213668
rect 206319 213610 206324 213666
rect 206380 213610 210528 213666
rect 206319 213608 210528 213610
rect 206319 213605 206385 213608
rect 146799 213372 146865 213375
rect 140832 213370 146865 213372
rect 140832 213314 146804 213370
rect 146860 213314 146865 213370
rect 140832 213312 146865 213314
rect 146799 213309 146865 213312
rect 677058 213227 677118 213490
rect 677007 213222 677118 213227
rect 677007 213166 677012 213222
rect 677068 213166 677118 213222
rect 677007 213164 677118 213166
rect 677007 213161 677073 213164
rect 43311 213076 43377 213079
rect 42528 213074 43377 213076
rect 42528 213018 43316 213074
rect 43372 213018 43377 213074
rect 42528 213016 43377 213018
rect 43311 213013 43377 213016
rect 206319 213076 206385 213079
rect 206319 213074 210528 213076
rect 206319 213018 206324 213074
rect 206380 213018 210528 213074
rect 206319 213016 210528 213018
rect 206319 213013 206385 213016
rect 206127 212780 206193 212783
rect 206127 212778 210558 212780
rect 206127 212722 206132 212778
rect 206188 212722 210558 212778
rect 206127 212720 210558 212722
rect 206127 212717 206193 212720
rect 210498 212528 210558 212720
rect 676866 212635 676926 212898
rect 676815 212630 676926 212635
rect 676815 212574 676820 212630
rect 676876 212574 676926 212630
rect 676815 212572 676926 212574
rect 676815 212569 676881 212572
rect 40578 212190 40638 212454
rect 40570 212126 40576 212190
rect 40640 212126 40646 212190
rect 42498 211747 42558 211862
rect 42447 211742 42558 211747
rect 42447 211686 42452 211742
rect 42508 211686 42558 211742
rect 42447 211684 42558 211686
rect 140802 211744 140862 212232
rect 676815 212188 676881 212191
rect 676815 212186 676926 212188
rect 676815 212130 676820 212186
rect 676876 212130 676926 212186
rect 676815 212125 676926 212130
rect 206607 212040 206673 212043
rect 206607 212038 210528 212040
rect 206607 211982 206612 212038
rect 206668 211982 210528 212038
rect 206607 211980 210528 211982
rect 206607 211977 206673 211980
rect 676866 211862 676926 212125
rect 677058 212043 677118 212306
rect 677007 212038 677118 212043
rect 677007 211982 677012 212038
rect 677068 211982 677118 212038
rect 677007 211980 677118 211982
rect 677007 211977 677073 211980
rect 146799 211744 146865 211747
rect 140802 211742 146865 211744
rect 140802 211686 146804 211742
rect 146860 211686 146865 211742
rect 140802 211684 146865 211686
rect 42447 211681 42513 211684
rect 146799 211681 146865 211684
rect 206895 211448 206961 211451
rect 206895 211446 210528 211448
rect 40386 211154 40446 211418
rect 206895 211390 206900 211446
rect 206956 211390 210528 211446
rect 206895 211388 210528 211390
rect 206895 211385 206961 211388
rect 40378 211090 40384 211154
rect 40448 211090 40454 211154
rect 40962 210562 41022 210826
rect 40954 210498 40960 210562
rect 41024 210498 41030 210562
rect 140802 210560 140862 211048
rect 145359 210560 145425 210563
rect 140802 210558 145425 210560
rect 140802 210502 145364 210558
rect 145420 210502 145425 210558
rect 140802 210500 145425 210502
rect 145359 210497 145425 210500
rect 640194 210412 640254 210826
rect 645615 210412 645681 210415
rect 647919 210412 647985 210415
rect 640194 210410 647985 210412
rect 640194 210354 645620 210410
rect 645676 210354 647924 210410
rect 647980 210354 647985 210410
rect 640194 210352 647985 210354
rect 645615 210349 645681 210352
rect 647919 210349 647985 210352
rect 41538 209970 41598 210234
rect 41530 209906 41536 209970
rect 41600 209906 41606 209970
rect 146703 209820 146769 209823
rect 140832 209818 146769 209820
rect 42114 209527 42174 209790
rect 140832 209762 146708 209818
rect 146764 209762 146769 209818
rect 140832 209760 146769 209762
rect 146703 209757 146769 209760
rect 42063 209522 42174 209527
rect 42063 209466 42068 209522
rect 42124 209466 42174 209522
rect 42063 209464 42174 209466
rect 42063 209461 42129 209464
rect 40770 208934 40830 209198
rect 40762 208870 40768 208934
rect 40832 208870 40838 208934
rect 41154 208342 41214 208606
rect 41146 208278 41152 208342
rect 41216 208278 41222 208342
rect 41346 207898 41406 208162
rect 140802 208044 140862 208602
rect 145455 208044 145521 208047
rect 140802 208042 145521 208044
rect 140802 207986 145460 208042
rect 145516 207986 145521 208042
rect 140802 207984 145521 207986
rect 145455 207981 145521 207984
rect 41338 207834 41344 207898
rect 41408 207834 41414 207898
rect 675706 207686 675712 207750
rect 675776 207748 675782 207750
rect 677103 207748 677169 207751
rect 675776 207746 677169 207748
rect 675776 207690 677108 207746
rect 677164 207690 677169 207746
rect 675776 207688 677169 207690
rect 675776 207686 675782 207688
rect 677103 207685 677169 207688
rect 40002 207307 40062 207570
rect 676666 207538 676672 207602
rect 676736 207600 676742 207602
rect 677199 207600 677265 207603
rect 676736 207598 677265 207600
rect 676736 207542 677204 207598
rect 677260 207542 677265 207598
rect 676736 207540 677265 207542
rect 676736 207538 676742 207540
rect 677199 207537 677265 207540
rect 146799 207452 146865 207455
rect 140832 207450 146865 207452
rect 140832 207394 146804 207450
rect 146860 207394 146865 207450
rect 140832 207392 146865 207394
rect 146799 207389 146865 207392
rect 676474 207390 676480 207454
rect 676544 207452 676550 207454
rect 676911 207452 676977 207455
rect 676544 207450 676977 207452
rect 676544 207394 676916 207450
rect 676972 207394 676977 207450
rect 676544 207392 676977 207394
rect 676544 207390 676550 207392
rect 676911 207389 676977 207392
rect 40002 207302 40113 207307
rect 40002 207246 40052 207302
rect 40108 207246 40113 207302
rect 40002 207244 40113 207246
rect 40047 207241 40113 207244
rect 40194 206715 40254 206978
rect 40143 206710 40254 206715
rect 40143 206654 40148 206710
rect 40204 206654 40254 206710
rect 40143 206652 40254 206654
rect 40143 206649 40209 206652
rect 40002 206123 40062 206534
rect 39951 206118 40062 206123
rect 39951 206062 39956 206118
rect 40012 206062 40062 206118
rect 39951 206060 40062 206062
rect 39951 206057 40017 206060
rect 40194 205679 40254 205942
rect 40194 205674 40305 205679
rect 40194 205618 40244 205674
rect 40300 205618 40305 205674
rect 40194 205616 40305 205618
rect 140802 205676 140862 206154
rect 145551 205676 145617 205679
rect 140802 205674 145617 205676
rect 140802 205618 145556 205674
rect 145612 205618 145617 205674
rect 140802 205616 145617 205618
rect 40239 205613 40305 205616
rect 145551 205613 145617 205616
rect 43023 205380 43089 205383
rect 42528 205378 43089 205380
rect 42528 205322 43028 205378
rect 43084 205322 43089 205378
rect 42528 205320 43089 205322
rect 43023 205317 43089 205320
rect 145743 205084 145809 205087
rect 140832 205082 145809 205084
rect 140832 205026 145748 205082
rect 145804 205026 145809 205082
rect 140832 205024 145809 205026
rect 145743 205021 145809 205024
rect 210159 205084 210225 205087
rect 211066 205084 211072 205086
rect 210159 205082 211072 205084
rect 210159 205026 210164 205082
rect 210220 205026 211072 205082
rect 210159 205024 211072 205026
rect 210159 205021 210225 205024
rect 211066 205022 211072 205024
rect 211136 205022 211142 205086
rect 42498 204495 42558 204832
rect 42447 204490 42558 204495
rect 42447 204434 42452 204490
rect 42508 204434 42558 204490
rect 42447 204432 42558 204434
rect 42447 204429 42513 204432
rect 35202 204051 35262 204314
rect 35151 204046 35262 204051
rect 35151 203990 35156 204046
rect 35212 203990 35262 204046
rect 35151 203988 35262 203990
rect 42447 204048 42513 204051
rect 42447 204046 42558 204048
rect 42447 203990 42452 204046
rect 42508 203990 42558 204046
rect 35151 203985 35217 203988
rect 42447 203985 42558 203990
rect 42498 203722 42558 203985
rect 35151 203604 35217 203607
rect 35151 203602 35262 203604
rect 35151 203546 35156 203602
rect 35212 203546 35262 203602
rect 35151 203541 35262 203546
rect 35202 203204 35262 203541
rect 140802 203308 140862 203796
rect 144975 203308 145041 203311
rect 140802 203306 145041 203308
rect 140802 203250 144980 203306
rect 145036 203250 145041 203306
rect 140802 203248 145041 203250
rect 144975 203245 145041 203248
rect 205743 202716 205809 202719
rect 209199 202716 209265 202719
rect 205743 202714 210528 202716
rect 205743 202658 205748 202714
rect 205804 202658 209204 202714
rect 209260 202658 210528 202714
rect 205743 202656 210528 202658
rect 205743 202653 205809 202656
rect 209199 202653 209265 202656
rect 140802 202124 140862 202612
rect 146799 202124 146865 202127
rect 140802 202122 146865 202124
rect 140802 202066 146804 202122
rect 146860 202066 146865 202122
rect 140802 202064 146865 202066
rect 146799 202061 146865 202064
rect 145647 201384 145713 201387
rect 140832 201382 145713 201384
rect 140832 201326 145652 201382
rect 145708 201326 145713 201382
rect 140832 201324 145713 201326
rect 145647 201321 145713 201324
rect 140802 199608 140862 200142
rect 675375 200054 675441 200055
rect 675322 199990 675328 200054
rect 675392 200052 675441 200054
rect 675392 200050 675484 200052
rect 675436 199994 675484 200050
rect 675392 199992 675484 199994
rect 675392 199990 675441 199992
rect 675375 199989 675441 199990
rect 146799 199608 146865 199611
rect 675471 199610 675537 199611
rect 675471 199608 675520 199610
rect 140802 199606 146865 199608
rect 140802 199550 146804 199606
rect 146860 199550 146865 199606
rect 140802 199548 146865 199550
rect 675428 199606 675520 199608
rect 675428 199550 675476 199606
rect 675428 199548 675520 199550
rect 146799 199545 146865 199548
rect 675471 199546 675520 199548
rect 675584 199546 675590 199610
rect 675471 199545 675537 199546
rect 145071 199016 145137 199019
rect 140832 199014 145137 199016
rect 140832 198958 145076 199014
rect 145132 198958 145137 199014
rect 140832 198956 145137 198958
rect 145071 198953 145137 198956
rect 675759 198426 675825 198427
rect 675706 198362 675712 198426
rect 675776 198424 675825 198426
rect 675776 198422 675868 198424
rect 675820 198366 675868 198422
rect 675776 198364 675868 198366
rect 675776 198362 675825 198364
rect 675759 198361 675825 198362
rect 146799 197832 146865 197835
rect 41116 197827 41186 197832
rect 140832 197830 146865 197832
rect 41116 197767 41121 197827
rect 41181 197767 41188 197827
rect 140832 197774 146804 197830
rect 146860 197774 146865 197830
rect 140832 197772 146865 197774
rect 146799 197769 146865 197772
rect 41116 197762 41188 197767
rect 41128 197684 41188 197762
rect 42106 197684 42112 197686
rect 41128 197624 42112 197684
rect 42106 197622 42112 197624
rect 42176 197622 42182 197686
rect 144591 196648 144657 196651
rect 140832 196646 144657 196648
rect 140832 196590 144596 196646
rect 144652 196590 144657 196646
rect 140832 196588 144657 196590
rect 144591 196585 144657 196588
rect 140802 194872 140862 195360
rect 675759 195316 675825 195319
rect 676474 195316 676480 195318
rect 675759 195314 676480 195316
rect 675759 195258 675764 195314
rect 675820 195258 676480 195314
rect 675759 195256 676480 195258
rect 675759 195253 675825 195256
rect 676474 195254 676480 195256
rect 676544 195254 676550 195318
rect 210874 194958 210880 195022
rect 210944 194958 210950 195022
rect 211066 194958 211072 195022
rect 211136 194958 211142 195022
rect 144399 194872 144465 194875
rect 140802 194870 144465 194872
rect 140802 194814 144404 194870
rect 144460 194814 144465 194870
rect 140802 194812 144465 194814
rect 144399 194809 144465 194812
rect 210882 194578 210942 194958
rect 210874 194514 210880 194578
rect 210944 194514 210950 194578
rect 140802 193688 140862 194176
rect 211074 194134 211134 194958
rect 211066 194070 211072 194134
rect 211136 194070 211142 194134
rect 145839 193688 145905 193691
rect 140802 193686 145905 193688
rect 140802 193630 145844 193686
rect 145900 193630 145905 193686
rect 140802 193628 145905 193630
rect 145839 193625 145905 193628
rect 674170 193478 674176 193542
rect 674240 193540 674246 193542
rect 675375 193540 675441 193543
rect 674240 193538 675441 193540
rect 674240 193482 675380 193538
rect 675436 193482 675441 193538
rect 674240 193480 675441 193482
rect 674240 193478 674246 193480
rect 675375 193477 675441 193480
rect 675087 193096 675153 193099
rect 675322 193096 675328 193098
rect 675087 193094 675328 193096
rect 675087 193038 675092 193094
rect 675148 193038 675328 193094
rect 675087 193036 675328 193038
rect 675087 193033 675153 193036
rect 675322 193034 675328 193036
rect 675392 193034 675398 193098
rect 146703 192948 146769 192951
rect 140832 192946 146769 192948
rect 140832 192890 146708 192946
rect 146764 192890 146769 192946
rect 140832 192888 146769 192890
rect 146703 192885 146769 192888
rect 146799 191764 146865 191767
rect 140832 191762 146865 191764
rect 140832 191706 146804 191762
rect 146860 191706 146865 191762
rect 140832 191704 146865 191706
rect 146799 191701 146865 191704
rect 675759 191616 675825 191619
rect 676666 191616 676672 191618
rect 675759 191614 676672 191616
rect 675759 191558 675764 191614
rect 675820 191558 676672 191614
rect 675759 191556 676672 191558
rect 675759 191553 675825 191556
rect 676666 191554 676672 191556
rect 676736 191554 676742 191618
rect 42159 191026 42225 191027
rect 42106 191024 42112 191026
rect 42068 190964 42112 191024
rect 42176 191022 42225 191026
rect 42220 190966 42225 191022
rect 42106 190962 42112 190964
rect 42176 190962 42225 190966
rect 42159 190961 42225 190962
rect 41530 190074 41536 190138
rect 41600 190136 41606 190138
rect 41775 190136 41841 190139
rect 41600 190134 41841 190136
rect 41600 190078 41780 190134
rect 41836 190078 41841 190134
rect 41600 190076 41841 190078
rect 140802 190136 140862 190476
rect 145935 190136 146001 190139
rect 140802 190134 146001 190136
rect 140802 190078 145940 190134
rect 145996 190078 146001 190134
rect 140802 190076 146001 190078
rect 41600 190074 41606 190076
rect 41775 190073 41841 190076
rect 145935 190073 146001 190076
rect 210106 190074 210112 190138
rect 210176 190136 210182 190138
rect 211066 190136 211072 190138
rect 210176 190076 211072 190136
rect 210176 190074 210182 190076
rect 211066 190074 211072 190076
rect 211136 190074 211142 190138
rect 671682 189502 708777 189503
rect 146031 189396 146097 189399
rect 140832 189394 146097 189396
rect 140832 189338 146036 189394
rect 146092 189338 146097 189394
rect 140832 189336 146097 189338
rect 146031 189333 146097 189336
rect 41775 189102 41841 189103
rect 41722 189100 41728 189102
rect 41684 189040 41728 189100
rect 41792 189098 41841 189102
rect 41836 189042 41841 189098
rect 41722 189038 41728 189040
rect 41792 189038 41841 189042
rect 41775 189037 41841 189038
rect 671677 188410 671683 189502
rect 672775 188410 708777 189502
rect 671682 188409 708777 188410
rect 709871 188409 711275 189503
rect 41967 188362 42033 188363
rect 41914 188298 41920 188362
rect 41984 188360 42033 188362
rect 42927 188360 42993 188363
rect 41984 188358 42993 188360
rect 42028 188302 42932 188358
rect 42988 188302 42993 188358
rect 41984 188300 42993 188302
rect 41984 188298 42033 188300
rect 41967 188297 42033 188298
rect 42927 188297 42993 188300
rect 146799 188212 146865 188215
rect 140832 188210 146865 188212
rect 140832 188154 146804 188210
rect 146860 188154 146865 188210
rect 140832 188152 146865 188154
rect 146799 188149 146865 188152
rect 666066 187433 698514 187434
rect 41338 187114 41344 187178
rect 41408 187176 41414 187178
rect 41775 187176 41841 187179
rect 41408 187174 41841 187176
rect 41408 187118 41780 187174
rect 41836 187118 41841 187174
rect 41408 187116 41841 187118
rect 41408 187114 41414 187116
rect 41775 187113 41841 187116
rect 41146 186374 41152 186438
rect 41216 186436 41222 186438
rect 41775 186436 41841 186439
rect 41216 186434 41841 186436
rect 41216 186378 41780 186434
rect 41836 186378 41841 186434
rect 41216 186376 41841 186378
rect 140802 186436 140862 186924
rect 146415 186436 146481 186439
rect 140802 186434 146481 186436
rect 140802 186378 146420 186434
rect 146476 186378 146481 186434
rect 140802 186376 146481 186378
rect 41216 186374 41222 186376
rect 41775 186373 41841 186376
rect 146415 186373 146481 186376
rect 666061 186251 666067 187433
rect 667249 186251 698514 187433
rect 666066 186250 698514 186251
rect 699698 186250 710266 187434
rect 40954 185782 40960 185846
rect 41024 185844 41030 185846
rect 41775 185844 41841 185847
rect 41024 185842 41841 185844
rect 41024 185786 41780 185842
rect 41836 185786 41841 185842
rect 41024 185784 41841 185786
rect 41024 185782 41030 185784
rect 41775 185781 41841 185784
rect 140802 185252 140862 185740
rect 146223 185252 146289 185255
rect 140802 185250 146289 185252
rect 140802 185194 146228 185250
rect 146284 185194 146289 185250
rect 140802 185192 146289 185194
rect 146223 185189 146289 185192
rect 146799 184512 146865 184515
rect 140832 184510 146865 184512
rect 140832 184454 146804 184510
rect 146860 184454 146865 184510
rect 140832 184452 146865 184454
rect 146799 184449 146865 184452
rect 40570 184154 40576 184218
rect 40640 184216 40646 184218
rect 41775 184216 41841 184219
rect 40640 184214 41841 184216
rect 40640 184158 41780 184214
rect 41836 184158 41841 184214
rect 40640 184156 41841 184158
rect 40640 184154 40646 184156
rect 41775 184153 41841 184156
rect 645415 183647 645421 185881
rect 647655 185084 647661 185881
rect 647655 183900 700656 185084
rect 701840 183900 710016 185084
rect 647655 183647 647661 183900
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 144495 183328 144561 183331
rect 140832 183326 144561 183328
rect 140832 183270 144500 183326
rect 144556 183270 144561 183326
rect 140832 183268 144561 183270
rect 144495 183265 144561 183268
rect 40378 182822 40384 182886
rect 40448 182884 40454 182886
rect 41775 182884 41841 182887
rect 40448 182882 41841 182884
rect 40448 182826 41780 182882
rect 41836 182826 41841 182882
rect 40448 182824 41841 182826
rect 40448 182822 40454 182824
rect 41775 182821 41841 182824
rect 140802 181848 140862 182188
rect 144015 181848 144081 181851
rect 140802 181846 144081 181848
rect 140802 181790 144020 181846
rect 144076 181790 144081 181846
rect 140802 181788 144081 181790
rect 144015 181785 144081 181788
rect 140802 180516 140862 180994
rect 641087 180957 641093 183191
rect 643327 182394 643333 183191
rect 643327 181210 706104 182394
rect 707288 181210 710404 182394
rect 643327 180957 643333 181210
rect 146607 180516 146673 180519
rect 140802 180514 146673 180516
rect 140802 180458 146612 180514
rect 146668 180458 146673 180514
rect 140802 180456 146673 180458
rect 146607 180453 146673 180456
rect 145263 179776 145329 179779
rect 140832 179774 145329 179776
rect 140832 179718 145268 179774
rect 145324 179718 145329 179774
rect 140832 179716 145329 179718
rect 145263 179713 145329 179716
rect 674607 179628 674673 179631
rect 674754 179628 674814 179894
rect 674607 179626 674814 179628
rect 674607 179570 674612 179626
rect 674668 179570 674814 179626
rect 674607 179568 674814 179570
rect 674607 179565 674673 179568
rect 674415 179332 674481 179335
rect 674415 179330 674784 179332
rect 674415 179274 674420 179330
rect 674476 179274 674784 179330
rect 674415 179272 674784 179274
rect 674415 179269 674481 179272
rect 674415 178814 674481 178817
rect 674415 178812 674784 178814
rect 674415 178756 674420 178812
rect 674476 178756 674784 178812
rect 674415 178754 674784 178756
rect 674415 178751 674481 178754
rect 146799 178592 146865 178595
rect 140832 178590 146865 178592
rect 140832 178534 146804 178590
rect 146860 178534 146865 178590
rect 140832 178532 146865 178534
rect 146799 178529 146865 178532
rect 677434 178382 677440 178446
rect 677504 178382 677510 178446
rect 677442 178266 677502 178382
rect 677442 177410 677502 177674
rect 677050 177346 677056 177410
rect 677120 177346 677126 177410
rect 677434 177346 677440 177410
rect 677504 177346 677510 177410
rect 140802 176816 140862 177304
rect 677058 177156 677118 177346
rect 144111 176816 144177 176819
rect 140802 176814 144177 176816
rect 140802 176758 144116 176814
rect 144172 176758 144177 176814
rect 140802 176756 144177 176758
rect 144111 176753 144177 176756
rect 677250 176374 677310 176638
rect 677242 176310 677248 176374
rect 677312 176310 677318 176374
rect 146799 176076 146865 176079
rect 140832 176074 146865 176076
rect 140832 176018 146804 176074
rect 146860 176018 146865 176074
rect 140832 176016 146865 176018
rect 146799 176013 146865 176016
rect 675138 175931 675198 176046
rect 675087 175926 675198 175931
rect 675087 175870 675092 175926
rect 675148 175870 675198 175926
rect 675087 175868 675198 175870
rect 675087 175865 675153 175868
rect 209914 175718 209920 175782
rect 209984 175780 209990 175782
rect 211066 175780 211072 175782
rect 209984 175720 211072 175780
rect 209984 175718 209990 175720
rect 211066 175718 211072 175720
rect 211136 175718 211142 175782
rect 676866 175191 676926 175528
rect 676866 175186 676977 175191
rect 676866 175130 676916 175186
rect 676972 175130 676977 175186
rect 676866 175128 676977 175130
rect 676911 175125 676977 175128
rect 140802 174448 140862 174982
rect 675522 174747 675582 175010
rect 675471 174742 675582 174747
rect 675471 174686 675476 174742
rect 675532 174686 675582 174742
rect 675471 174684 675582 174686
rect 675471 174681 675537 174684
rect 144975 174448 145041 174451
rect 140802 174446 145041 174448
rect 140802 174390 144980 174446
rect 145036 174390 145041 174446
rect 140802 174388 145041 174390
rect 144975 174385 145041 174388
rect 210682 174386 210688 174450
rect 210752 174448 210758 174450
rect 211066 174448 211072 174450
rect 210752 174388 211072 174448
rect 210752 174386 210758 174388
rect 211066 174386 211072 174388
rect 211136 174386 211142 174450
rect 675138 174303 675198 174418
rect 675138 174298 675249 174303
rect 675138 174242 675188 174298
rect 675244 174242 675249 174298
rect 675138 174240 675249 174242
rect 675183 174237 675249 174240
rect 210298 173942 210304 174006
rect 210368 174004 210374 174006
rect 210874 174004 210880 174006
rect 210368 173944 210880 174004
rect 210368 173942 210374 173944
rect 210874 173942 210880 173944
rect 210944 173942 210950 174006
rect 674031 173856 674097 173859
rect 674031 173854 674784 173856
rect 674031 173798 674036 173854
rect 674092 173798 674784 173854
rect 674031 173796 674784 173798
rect 674031 173793 674097 173796
rect 140802 173412 140862 173752
rect 144783 173412 144849 173415
rect 140802 173410 144849 173412
rect 140802 173354 144788 173410
rect 144844 173354 144849 173410
rect 140802 173352 144849 173354
rect 144783 173349 144849 173352
rect 676866 173119 676926 173382
rect 676815 173114 676926 173119
rect 676815 173058 676820 173114
rect 676876 173058 676926 173114
rect 676815 173056 676926 173058
rect 676815 173053 676881 173056
rect 675330 172675 675390 172790
rect 675279 172670 675390 172675
rect 675279 172614 675284 172670
rect 675340 172614 675390 172670
rect 675279 172612 675390 172614
rect 675279 172609 675345 172612
rect 140802 172080 140862 172562
rect 674946 172083 675006 172198
rect 145263 172080 145329 172083
rect 140802 172078 145329 172080
rect 140802 172022 145268 172078
rect 145324 172022 145329 172078
rect 140802 172020 145329 172022
rect 674946 172078 675057 172083
rect 674946 172022 674996 172078
rect 675052 172022 675057 172078
rect 674946 172020 675057 172022
rect 145263 172017 145329 172020
rect 674991 172017 675057 172020
rect 674946 171491 675006 171754
rect 674895 171486 675006 171491
rect 674895 171430 674900 171486
rect 674956 171430 675006 171486
rect 674895 171428 675006 171430
rect 674895 171425 674961 171428
rect 146799 171340 146865 171343
rect 140832 171338 146865 171340
rect 140832 171282 146804 171338
rect 146860 171282 146865 171338
rect 140832 171280 146865 171282
rect 146799 171277 146865 171280
rect 209914 171278 209920 171342
rect 209984 171340 209990 171342
rect 211066 171340 211072 171342
rect 209984 171280 211072 171340
rect 209984 171278 209990 171280
rect 211066 171278 211072 171280
rect 211136 171278 211142 171342
rect 673978 171130 673984 171194
rect 674048 171192 674054 171194
rect 674048 171132 674784 171192
rect 674048 171130 674054 171132
rect 210106 170538 210112 170602
rect 210176 170600 210182 170602
rect 211066 170600 211072 170602
rect 210176 170540 211072 170600
rect 210176 170538 210182 170540
rect 211066 170538 211072 170540
rect 211136 170538 211142 170602
rect 673935 170600 674001 170603
rect 673935 170598 674784 170600
rect 673935 170542 673940 170598
rect 673996 170542 674784 170598
rect 673935 170540 674784 170542
rect 673935 170537 674001 170540
rect 146703 170156 146769 170159
rect 140832 170154 146769 170156
rect 140832 170098 146708 170154
rect 146764 170098 146769 170154
rect 140832 170096 146769 170098
rect 146703 170093 146769 170096
rect 674415 170156 674481 170159
rect 674415 170154 674784 170156
rect 674415 170098 674420 170154
rect 674476 170098 674784 170154
rect 674415 170096 674784 170098
rect 674415 170093 674481 170096
rect 674223 169564 674289 169567
rect 674223 169562 674784 169564
rect 674223 169506 674228 169562
rect 674284 169506 674784 169562
rect 674223 169504 674784 169506
rect 674223 169501 674289 169504
rect 674127 168972 674193 168975
rect 674127 168970 674784 168972
rect 674127 168914 674132 168970
rect 674188 168914 674784 168970
rect 674127 168912 674784 168914
rect 674127 168909 674193 168912
rect 140802 168380 140862 168868
rect 144783 168380 144849 168383
rect 140802 168378 144849 168380
rect 140802 168322 144788 168378
rect 144844 168322 144849 168378
rect 140802 168320 144849 168322
rect 144783 168317 144849 168320
rect 674754 168235 674814 168498
rect 674703 168230 674814 168235
rect 674703 168174 674708 168230
rect 674764 168174 674814 168230
rect 674703 168172 674814 168174
rect 674703 168169 674769 168172
rect 146799 167640 146865 167643
rect 140832 167638 146865 167640
rect 140832 167582 146804 167638
rect 146860 167582 146865 167638
rect 140832 167580 146865 167582
rect 146799 167577 146865 167580
rect 674607 167640 674673 167643
rect 674754 167640 674814 167906
rect 674607 167638 674814 167640
rect 674607 167582 674612 167638
rect 674668 167582 674814 167638
rect 674607 167580 674814 167582
rect 674607 167577 674673 167580
rect 674754 167199 674814 167314
rect 674703 167194 674814 167199
rect 674703 167138 674708 167194
rect 674764 167138 674814 167194
rect 674703 167136 674814 167138
rect 674703 167133 674769 167136
rect 647919 167048 647985 167051
rect 640194 167046 647985 167048
rect 640194 166990 647924 167046
rect 647980 166990 647985 167046
rect 640194 166988 647985 166990
rect 640194 166870 640254 166988
rect 647919 166985 647985 166988
rect 144783 166604 144849 166607
rect 140832 166602 144849 166604
rect 140832 166546 144788 166602
rect 144844 166546 144849 166602
rect 140832 166544 144849 166546
rect 144783 166541 144849 166544
rect 646287 166308 646353 166311
rect 640416 166306 646353 166308
rect 640416 166250 646292 166306
rect 646348 166250 646353 166306
rect 640416 166248 646353 166250
rect 646287 166245 646353 166248
rect 646863 166012 646929 166015
rect 640386 166010 646929 166012
rect 640386 165954 646868 166010
rect 646924 165954 646929 166010
rect 640386 165952 646929 165954
rect 640386 165686 640446 165952
rect 646863 165949 646929 165952
rect 140802 164828 140862 165316
rect 145167 164828 145233 164831
rect 140802 164826 145233 164828
rect 140802 164770 145172 164826
rect 145228 164770 145233 164826
rect 140802 164768 145233 164770
rect 145167 164765 145233 164768
rect 210159 164236 210225 164239
rect 211066 164236 211072 164238
rect 210159 164234 211072 164236
rect 210159 164178 210164 164234
rect 210220 164178 211072 164234
rect 210159 164176 211072 164178
rect 210159 164173 210225 164176
rect 211066 164174 211072 164176
rect 211136 164174 211142 164238
rect 140802 163644 140862 164130
rect 144207 163644 144273 163647
rect 140802 163642 144273 163644
rect 140802 163586 144212 163642
rect 144268 163586 144273 163642
rect 140802 163584 144273 163586
rect 144207 163581 144273 163584
rect 144879 162904 144945 162907
rect 140832 162902 144945 162904
rect 140832 162846 144884 162902
rect 144940 162846 144945 162902
rect 140832 162844 144945 162846
rect 144879 162841 144945 162844
rect 140802 161424 140862 161682
rect 675706 161510 675712 161574
rect 675776 161572 675782 161574
rect 676911 161572 676977 161575
rect 675776 161570 676977 161572
rect 675776 161514 676916 161570
rect 676972 161514 676977 161570
rect 675776 161512 676977 161514
rect 675776 161510 675782 161512
rect 676911 161509 676977 161512
rect 144975 161424 145041 161427
rect 140802 161422 145041 161424
rect 140802 161366 144980 161422
rect 145036 161366 145041 161422
rect 140802 161364 145041 161366
rect 144975 161361 145041 161364
rect 676666 161362 676672 161426
rect 676736 161424 676742 161426
rect 676815 161424 676881 161427
rect 676736 161422 676881 161424
rect 676736 161366 676820 161422
rect 676876 161366 676881 161422
rect 676736 161364 676881 161366
rect 676736 161362 676742 161364
rect 676815 161361 676881 161364
rect 140802 159944 140862 160432
rect 144015 159944 144081 159947
rect 140802 159942 144081 159944
rect 140802 159886 144020 159942
rect 144076 159886 144081 159942
rect 140802 159884 144081 159886
rect 144015 159881 144081 159884
rect 144879 159352 144945 159355
rect 140832 159350 144945 159352
rect 140832 159294 144884 159350
rect 144940 159294 144945 159350
rect 140832 159292 144945 159294
rect 144879 159289 144945 159292
rect 144111 158168 144177 158171
rect 140832 158166 144177 158168
rect 140832 158110 144116 158166
rect 144172 158110 144177 158166
rect 140832 158108 144177 158110
rect 144111 158105 144177 158108
rect 140802 156392 140862 156880
rect 144879 156392 144945 156395
rect 140802 156390 144945 156392
rect 140802 156334 144884 156390
rect 144940 156334 144945 156390
rect 140802 156332 144945 156334
rect 144879 156329 144945 156332
rect 140802 155652 140862 155696
rect 144303 155652 144369 155655
rect 140802 155650 144369 155652
rect 140802 155594 144308 155650
rect 144364 155594 144369 155650
rect 140802 155592 144369 155594
rect 144303 155589 144369 155592
rect 675279 155210 675345 155211
rect 675279 155208 675328 155210
rect 675236 155206 675328 155208
rect 675236 155150 675284 155206
rect 675236 155148 675328 155150
rect 675279 155146 675328 155148
rect 675392 155146 675398 155210
rect 675279 155145 675345 155146
rect 144783 154468 144849 154471
rect 675471 154470 675537 154471
rect 675471 154468 675520 154470
rect 140832 154466 144849 154468
rect 140832 154410 144788 154466
rect 144844 154410 144849 154466
rect 140832 154408 144849 154410
rect 675428 154466 675520 154468
rect 675428 154410 675476 154466
rect 675428 154408 675520 154410
rect 144783 154405 144849 154408
rect 675471 154406 675520 154408
rect 675584 154406 675590 154470
rect 675471 154405 675537 154406
rect 140802 152988 140862 153250
rect 144879 152988 144945 152991
rect 140802 152986 144945 152988
rect 140802 152930 144884 152986
rect 144940 152930 144945 152986
rect 140802 152928 144945 152930
rect 144879 152925 144945 152928
rect 140802 151656 140862 152144
rect 210106 151890 210112 151954
rect 210176 151952 210182 151954
rect 210874 151952 210880 151954
rect 210176 151892 210880 151952
rect 210176 151890 210182 151892
rect 210874 151890 210880 151892
rect 210944 151890 210950 151954
rect 144495 151656 144561 151659
rect 140802 151654 144561 151656
rect 140802 151598 144500 151654
rect 144556 151598 144561 151654
rect 140802 151596 144561 151598
rect 144495 151593 144561 151596
rect 144879 150916 144945 150919
rect 140832 150914 144945 150916
rect 140832 150858 144884 150914
rect 144940 150858 144945 150914
rect 140832 150856 144945 150858
rect 144879 150853 144945 150856
rect 673978 150262 673984 150326
rect 674048 150324 674054 150326
rect 675471 150324 675537 150327
rect 674048 150322 675537 150324
rect 674048 150266 675476 150322
rect 675532 150266 675537 150322
rect 674048 150264 675537 150266
rect 674048 150262 674054 150264
rect 675471 150261 675537 150264
rect 144783 149732 144849 149735
rect 140832 149730 144849 149732
rect 140832 149674 144788 149730
rect 144844 149674 144849 149730
rect 140832 149672 144849 149674
rect 144783 149669 144849 149672
rect 675759 148550 675825 148551
rect 675706 148486 675712 148550
rect 675776 148548 675825 148550
rect 675776 148546 675868 148548
rect 675820 148490 675868 148546
rect 675776 148488 675868 148490
rect 675776 148486 675825 148488
rect 675759 148485 675825 148486
rect 140802 147956 140862 148444
rect 144879 147956 144945 147959
rect 140802 147954 144945 147956
rect 140802 147898 144884 147954
rect 144940 147898 144945 147954
rect 140802 147896 144945 147898
rect 144879 147893 144945 147896
rect 140802 146920 140862 147260
rect 144687 146920 144753 146923
rect 140802 146918 144753 146920
rect 140802 146862 144692 146918
rect 144748 146862 144753 146918
rect 140802 146860 144753 146862
rect 144687 146857 144753 146860
rect 675759 146624 675825 146627
rect 676666 146624 676672 146626
rect 675759 146622 676672 146624
rect 675759 146566 675764 146622
rect 675820 146566 676672 146622
rect 675759 146564 676672 146566
rect 675759 146561 675825 146564
rect 676666 146562 676672 146564
rect 676736 146562 676742 146626
rect 144495 146032 144561 146035
rect 140832 146030 144561 146032
rect 140832 145974 144500 146030
rect 144556 145974 144561 146030
rect 140832 145972 144561 145974
rect 144495 145969 144561 145972
rect 140802 144404 140862 144790
rect 144826 144786 144832 144850
rect 144896 144848 144902 144850
rect 146319 144848 146385 144851
rect 144896 144846 146385 144848
rect 144896 144790 146324 144846
rect 146380 144790 146385 144846
rect 144896 144788 146385 144790
rect 144896 144786 144902 144788
rect 146319 144785 146385 144788
rect 144303 144404 144369 144407
rect 140802 144402 144369 144404
rect 140802 144346 144308 144402
rect 144364 144346 144369 144402
rect 140802 144344 144369 144346
rect 144303 144341 144369 144344
rect 671682 143722 708743 143723
rect 140802 143220 140862 143708
rect 144495 143220 144561 143223
rect 140802 143218 144561 143220
rect 140802 143162 144500 143218
rect 144556 143162 144561 143218
rect 140802 143160 144561 143162
rect 144495 143157 144561 143160
rect 671677 142630 671683 143722
rect 672775 142630 708743 143722
rect 671682 142629 708743 142630
rect 709837 142629 709843 143723
rect 144303 142480 144369 142483
rect 140832 142478 144369 142480
rect 140832 142422 144308 142478
rect 144364 142422 144369 142478
rect 140832 142420 144369 142422
rect 144303 142417 144369 142420
rect 666066 141405 698402 141406
rect 144303 141296 144369 141299
rect 140832 141294 144369 141296
rect 140832 141238 144308 141294
rect 144364 141238 144369 141294
rect 140832 141236 144369 141238
rect 144303 141233 144369 141236
rect 645327 141148 645393 141151
rect 645186 141146 645393 141148
rect 645186 141090 645332 141146
rect 645388 141090 645393 141146
rect 645186 141088 645393 141090
rect 645186 140852 645246 141088
rect 645327 141085 645393 141088
rect 645327 140852 645393 140855
rect 645186 140850 645393 140852
rect 645186 140794 645332 140850
rect 645388 140794 645393 140850
rect 645186 140792 645393 140794
rect 645327 140789 645393 140792
rect 666061 140223 666067 141405
rect 667249 140223 698402 141405
rect 666066 140222 698402 140223
rect 699586 140222 703644 141406
rect 140802 139520 140862 140008
rect 144303 139520 144369 139523
rect 140802 139518 144369 139520
rect 140802 139462 144308 139518
rect 144364 139462 144369 139518
rect 140802 139460 144369 139462
rect 144303 139457 144369 139460
rect 140802 138336 140862 138824
rect 645415 138676 645421 139451
rect 146319 138336 146385 138339
rect 140802 138334 146385 138336
rect 140802 138278 146324 138334
rect 146380 138278 146385 138334
rect 140802 138276 146385 138278
rect 146319 138273 146385 138276
rect 144303 137596 144369 137599
rect 140832 137594 144369 137596
rect 140832 137538 144308 137594
rect 144364 137538 144369 137594
rect 140832 137536 144369 137538
rect 144303 137533 144369 137536
rect 210298 137238 210304 137302
rect 210368 137300 210374 137302
rect 211066 137300 211072 137302
rect 210368 137240 211072 137300
rect 210368 137238 210374 137240
rect 211066 137238 211072 137240
rect 211136 137238 211142 137302
rect 140802 136116 140862 136522
rect 146895 136116 146961 136119
rect 140802 136114 146961 136116
rect 140802 136058 146900 136114
rect 146956 136058 146961 136114
rect 140802 136056 146961 136058
rect 146895 136053 146961 136056
rect 641087 135469 641093 137703
rect 643327 136690 643333 137703
rect 645306 137492 645421 138676
rect 645415 137217 645421 137492
rect 647655 138676 647661 139451
rect 647655 137492 700550 138676
rect 701734 137492 701740 138676
rect 647655 137217 647661 137492
rect 643327 135506 706922 136690
rect 708106 135506 710558 136690
rect 643327 135469 643333 135506
rect 140802 134784 140862 135272
rect 144303 134784 144369 134787
rect 140802 134782 144369 134784
rect 140802 134726 144308 134782
rect 144364 134726 144369 134782
rect 140802 134724 144369 134726
rect 144303 134721 144369 134724
rect 676866 134343 676926 134680
rect 676866 134338 676977 134343
rect 676866 134282 676916 134338
rect 676972 134282 676977 134338
rect 676866 134280 676977 134282
rect 676911 134277 676977 134280
rect 144495 134044 144561 134047
rect 140832 134042 144561 134044
rect 140832 133986 144500 134042
rect 144556 133986 144561 134042
rect 140832 133984 144561 133986
rect 144495 133981 144561 133984
rect 676866 133899 676926 134162
rect 676815 133894 676926 133899
rect 676815 133838 676820 133894
rect 676876 133838 676926 133894
rect 676815 133836 676926 133838
rect 676815 133833 676881 133836
rect 674415 133600 674481 133603
rect 674415 133598 674784 133600
rect 674415 133542 674420 133598
rect 674476 133542 674784 133598
rect 674415 133540 674784 133542
rect 674415 133537 674481 133540
rect 677434 133390 677440 133454
rect 677504 133390 677510 133454
rect 677442 132978 677502 133390
rect 144303 132860 144369 132863
rect 140832 132858 144369 132860
rect 140832 132802 144308 132858
rect 144364 132802 144369 132858
rect 140832 132800 144369 132802
rect 144303 132797 144369 132800
rect 674415 132564 674481 132567
rect 674415 132562 674784 132564
rect 674415 132506 674420 132562
rect 674476 132506 674784 132562
rect 674415 132504 674784 132506
rect 674415 132501 674481 132504
rect 677050 132206 677056 132270
rect 677120 132206 677126 132270
rect 677058 131942 677118 132206
rect 677242 131762 677248 131826
rect 677312 131762 677318 131826
rect 140802 131084 140862 131572
rect 677250 131350 677310 131762
rect 144495 131084 144561 131087
rect 140802 131082 144561 131084
rect 140802 131026 144500 131082
rect 144556 131026 144561 131082
rect 140802 131024 144561 131026
rect 144495 131021 144561 131024
rect 674511 130640 674577 130643
rect 674754 130640 674814 130906
rect 674511 130638 674814 130640
rect 674511 130582 674516 130638
rect 674572 130582 674814 130638
rect 674511 130580 674814 130582
rect 674511 130577 674577 130580
rect 140802 130048 140862 130388
rect 677058 130051 677118 130314
rect 144303 130048 144369 130051
rect 140802 130046 144369 130048
rect 140802 129990 144308 130046
rect 144364 129990 144369 130046
rect 140802 129988 144369 129990
rect 677058 130046 677169 130051
rect 677058 129990 677108 130046
rect 677164 129990 677169 130046
rect 677058 129988 677169 129990
rect 144303 129985 144369 129988
rect 677103 129985 677169 129988
rect 675138 129607 675198 129722
rect 675138 129602 675249 129607
rect 675138 129546 675188 129602
rect 675244 129546 675249 129602
rect 675138 129544 675249 129546
rect 675183 129541 675249 129544
rect 144303 129308 144369 129311
rect 140832 129306 144369 129308
rect 140832 129250 144308 129306
rect 144364 129250 144369 129306
rect 140832 129248 144369 129250
rect 144303 129245 144369 129248
rect 674319 129308 674385 129311
rect 674319 129306 674784 129308
rect 674319 129250 674324 129306
rect 674380 129250 674784 129306
rect 674319 129248 674784 129250
rect 674319 129245 674385 129248
rect 673978 128654 673984 128718
rect 674048 128716 674054 128718
rect 674048 128656 674784 128716
rect 674048 128654 674054 128656
rect 140802 127680 140862 128090
rect 677058 127831 677118 128094
rect 677007 127826 677118 127831
rect 677007 127770 677012 127826
rect 677068 127770 677118 127826
rect 677007 127768 677118 127770
rect 677007 127765 677073 127768
rect 146511 127680 146577 127683
rect 140802 127678 146577 127680
rect 140802 127622 146516 127678
rect 146572 127622 146577 127678
rect 140802 127620 146577 127622
rect 146511 127617 146577 127620
rect 675138 127387 675198 127650
rect 675087 127382 675198 127387
rect 675087 127326 675092 127382
rect 675148 127326 675198 127382
rect 675087 127324 675198 127326
rect 675087 127321 675153 127324
rect 674223 127088 674289 127091
rect 674223 127086 674784 127088
rect 674223 127030 674228 127086
rect 674284 127030 674784 127086
rect 674223 127028 674784 127030
rect 674223 127025 674289 127028
rect 146991 126940 147057 126943
rect 140832 126938 147057 126940
rect 140832 126882 146996 126938
rect 147052 126882 147057 126938
rect 140832 126880 147057 126882
rect 146991 126877 147057 126880
rect 144303 126792 144369 126795
rect 144826 126792 144832 126794
rect 144303 126790 144832 126792
rect 144303 126734 144308 126790
rect 144364 126734 144832 126790
rect 144303 126732 144832 126734
rect 144303 126729 144369 126732
rect 144826 126730 144832 126732
rect 144896 126730 144902 126794
rect 674607 126348 674673 126351
rect 674754 126348 674814 126466
rect 674607 126346 674814 126348
rect 674607 126290 674612 126346
rect 674668 126290 674814 126346
rect 674607 126288 674814 126290
rect 674607 126285 674673 126288
rect 674170 125990 674176 126054
rect 674240 126052 674246 126054
rect 674240 125992 674784 126052
rect 674240 125990 674246 125992
rect 39855 125312 39921 125315
rect 39810 125310 39921 125312
rect 39810 125254 39860 125310
rect 39916 125254 39921 125310
rect 39810 125249 39921 125254
rect 39810 125058 39870 125249
rect 140802 125164 140862 125642
rect 673935 125460 674001 125463
rect 673935 125458 674784 125460
rect 673935 125402 673940 125458
rect 673996 125402 674784 125458
rect 673935 125400 674784 125402
rect 673935 125397 674001 125400
rect 144399 125164 144465 125167
rect 140802 125162 144465 125164
rect 140802 125106 144404 125162
rect 144460 125106 144465 125162
rect 140802 125104 144465 125106
rect 144399 125101 144465 125104
rect 210159 125164 210225 125167
rect 210490 125164 210496 125166
rect 210159 125162 210496 125164
rect 210159 125106 210164 125162
rect 210220 125106 210496 125162
rect 210159 125104 210496 125106
rect 210159 125101 210225 125104
rect 210490 125102 210496 125104
rect 210560 125102 210566 125166
rect 39593 124850 39999 125058
rect 44554 124850 51364 124890
rect 39593 120616 51364 124850
rect 674754 124723 674814 124838
rect 674754 124718 674865 124723
rect 674754 124662 674804 124718
rect 674860 124662 674865 124718
rect 674754 124660 674865 124662
rect 674799 124657 674865 124660
rect 144303 124572 144369 124575
rect 144634 124572 144640 124574
rect 144303 124570 144640 124572
rect 144303 124514 144308 124570
rect 144364 124514 144640 124570
rect 144303 124512 144640 124514
rect 144303 124509 144369 124512
rect 144634 124510 144640 124512
rect 144704 124510 144710 124574
rect 144303 124424 144369 124427
rect 140832 124422 144369 124424
rect 140832 124366 144308 124422
rect 144364 124366 144369 124422
rect 140832 124364 144369 124366
rect 144303 124361 144369 124364
rect 674946 124131 675006 124320
rect 674895 124126 675006 124131
rect 674895 124070 674900 124126
rect 674956 124070 675006 124126
rect 674895 124068 675006 124070
rect 674895 124065 674961 124068
rect 674415 123832 674481 123835
rect 674415 123830 674784 123832
rect 674415 123774 674420 123830
rect 674476 123774 674784 123830
rect 674415 123772 674784 123774
rect 674415 123769 674481 123772
rect 140802 122648 140862 123136
rect 210298 123030 210304 123094
rect 210368 123092 210374 123094
rect 211066 123092 211072 123094
rect 210368 123032 211072 123092
rect 210368 123030 210374 123032
rect 211066 123030 211072 123032
rect 211136 123030 211142 123094
rect 676866 122947 676926 123210
rect 676815 122942 676926 122947
rect 676815 122886 676820 122942
rect 676876 122886 676926 122942
rect 676815 122884 676926 122886
rect 676815 122881 676881 122884
rect 144399 122648 144465 122651
rect 140802 122646 144465 122648
rect 140802 122590 144404 122646
rect 144460 122590 144465 122646
rect 140802 122588 144465 122590
rect 144399 122585 144465 122588
rect 676866 122355 676926 122692
rect 676866 122350 676977 122355
rect 676866 122294 676916 122350
rect 676972 122294 676977 122350
rect 676866 122292 676977 122294
rect 676911 122289 676977 122292
rect 140802 121612 140862 121952
rect 674754 121911 674814 122174
rect 674703 121906 674814 121911
rect 674703 121850 674708 121906
rect 674764 121850 674814 121906
rect 674703 121848 674814 121850
rect 674703 121845 674769 121848
rect 210298 121698 210304 121762
rect 210368 121698 210374 121762
rect 144303 121612 144369 121615
rect 140802 121610 144369 121612
rect 140802 121554 144308 121610
rect 144364 121554 144369 121610
rect 140802 121552 144369 121554
rect 144303 121549 144369 121552
rect 210159 121318 210225 121319
rect 210306 121318 210366 121698
rect 640386 121464 640446 121730
rect 645903 121464 645969 121467
rect 640386 121462 645969 121464
rect 640386 121406 645908 121462
rect 645964 121406 645969 121462
rect 640386 121404 645969 121406
rect 645903 121401 645969 121404
rect 210106 121316 210112 121318
rect 210068 121256 210112 121316
rect 210176 121314 210225 121318
rect 210220 121258 210225 121314
rect 210106 121254 210112 121256
rect 210176 121254 210225 121258
rect 210298 121254 210304 121318
rect 210368 121254 210374 121318
rect 210159 121253 210225 121254
rect 645807 121168 645873 121171
rect 640416 121166 645873 121168
rect 640416 121110 645812 121166
rect 645868 121110 645873 121166
rect 640416 121108 645873 121110
rect 645807 121105 645873 121108
rect 144591 120872 144657 120875
rect 645999 120872 646065 120875
rect 140832 120870 144657 120872
rect 140832 120814 144596 120870
rect 144652 120814 144657 120870
rect 140832 120812 144657 120814
rect 144591 120809 144657 120812
rect 640386 120870 646065 120872
rect 640386 120814 646004 120870
rect 646060 120814 646065 120870
rect 640386 120812 646065 120814
rect 39593 120592 48196 120616
rect 39593 120278 39999 120592
rect 44554 115126 48196 120592
rect 51046 115126 51364 120616
rect 640386 120546 640446 120812
rect 645999 120809 646065 120812
rect 647631 120428 647697 120431
rect 640386 120426 647697 120428
rect 640386 120370 647636 120426
rect 647692 120370 647697 120426
rect 640386 120368 647697 120370
rect 640386 120028 640446 120368
rect 647631 120365 647697 120368
rect 140802 119096 140862 119630
rect 144399 119096 144465 119099
rect 140802 119094 144465 119096
rect 140802 119038 144404 119094
rect 144460 119038 144465 119094
rect 140802 119036 144465 119038
rect 144399 119033 144465 119036
rect 140610 118208 140670 118400
rect 144303 118208 144369 118211
rect 140610 118206 144369 118208
rect 140610 118150 144308 118206
rect 144364 118150 144369 118206
rect 140610 118148 144369 118150
rect 144303 118145 144369 118148
rect 210298 117998 210304 118062
rect 210368 118060 210374 118062
rect 211066 118060 211072 118062
rect 210368 118000 211072 118060
rect 210368 117998 210374 118000
rect 211066 117998 211072 118000
rect 211136 117998 211142 118062
rect 676474 117998 676480 118062
rect 676544 118060 676550 118062
rect 677007 118060 677073 118063
rect 676544 118058 677073 118060
rect 676544 118002 677012 118058
rect 677068 118002 677073 118058
rect 676544 118000 677073 118002
rect 676544 117998 676550 118000
rect 677007 117997 677073 118000
rect 675898 117850 675904 117914
rect 675968 117912 675974 117914
rect 677103 117912 677169 117915
rect 675968 117910 677169 117912
rect 675968 117854 677108 117910
rect 677164 117854 677169 117910
rect 675968 117852 677169 117854
rect 675968 117850 675974 117852
rect 677103 117849 677169 117852
rect 140802 116728 140862 117210
rect 144303 116728 144369 116731
rect 140802 116726 144369 116728
rect 140802 116670 144308 116726
rect 144364 116670 144369 116726
rect 140802 116668 144369 116670
rect 144303 116665 144369 116668
rect 144303 115988 144369 115991
rect 140832 115986 144369 115988
rect 140832 115930 144308 115986
rect 144364 115930 144369 115986
rect 140832 115928 144369 115930
rect 144303 115925 144369 115928
rect 44554 114966 51364 115126
rect 39802 110902 51364 114966
rect 140802 114212 140862 114762
rect 144399 114212 144465 114215
rect 140802 114210 144465 114212
rect 140802 114154 144404 114210
rect 144460 114154 144465 114210
rect 140802 114152 144465 114154
rect 144399 114149 144465 114152
rect 140802 113176 140862 113664
rect 144303 113326 144369 113327
rect 144250 113324 144256 113326
rect 144212 113264 144256 113324
rect 144320 113322 144369 113326
rect 144364 113266 144369 113322
rect 144250 113262 144256 113264
rect 144320 113262 144369 113266
rect 144303 113261 144369 113262
rect 144303 113176 144369 113179
rect 140802 113174 144369 113176
rect 140802 113118 144308 113174
rect 144364 113118 144369 113174
rect 140802 113116 144369 113118
rect 144303 113113 144369 113116
rect 144303 112436 144369 112439
rect 140832 112434 144369 112436
rect 140832 112378 144308 112434
rect 144364 112378 144369 112434
rect 140832 112376 144369 112378
rect 144303 112373 144369 112376
rect 144399 111252 144465 111255
rect 140832 111250 144465 111252
rect 140832 111194 144404 111250
rect 144460 111194 144465 111250
rect 140832 111192 144465 111194
rect 144399 111189 144465 111192
rect 44554 110824 51364 110902
rect 675375 110070 675441 110071
rect 675322 110068 675328 110070
rect 675284 110008 675328 110068
rect 675392 110066 675441 110070
rect 675436 110010 675441 110066
rect 675322 110006 675328 110008
rect 675392 110006 675441 110010
rect 675375 110005 675441 110006
rect 140802 109772 140862 109964
rect 144303 109772 144369 109775
rect 140802 109770 144369 109772
rect 140802 109714 144308 109770
rect 144364 109714 144369 109770
rect 140802 109712 144369 109714
rect 144303 109709 144369 109712
rect 675471 109330 675537 109331
rect 675471 109326 675520 109330
rect 675584 109328 675590 109330
rect 675471 109270 675476 109326
rect 675471 109266 675520 109270
rect 675584 109268 675628 109328
rect 675584 109266 675590 109268
rect 675471 109265 675537 109266
rect 140802 108292 140862 108778
rect 144591 108292 144657 108295
rect 140802 108290 144657 108292
rect 140802 108234 144596 108290
rect 144652 108234 144657 108290
rect 140802 108232 144657 108234
rect 144591 108229 144657 108232
rect 673978 108082 673984 108146
rect 674048 108144 674054 108146
rect 675375 108144 675441 108147
rect 674048 108142 675441 108144
rect 674048 108086 675380 108142
rect 675436 108086 675441 108142
rect 674048 108084 675441 108086
rect 674048 108082 674054 108084
rect 675375 108081 675441 108084
rect 144303 107552 144369 107555
rect 140832 107550 144369 107552
rect 140832 107494 144308 107550
rect 144364 107494 144369 107550
rect 140832 107492 144369 107494
rect 144303 107489 144369 107492
rect 144250 106750 144256 106814
rect 144320 106812 144326 106814
rect 144399 106812 144465 106815
rect 144320 106810 144465 106812
rect 144320 106754 144404 106810
rect 144460 106754 144465 106810
rect 144320 106752 144465 106754
rect 144320 106750 144326 106752
rect 144399 106749 144465 106752
rect 144634 106602 144640 106666
rect 144704 106664 144710 106666
rect 145071 106664 145137 106667
rect 144704 106662 145137 106664
rect 144704 106606 145076 106662
rect 145132 106606 145137 106662
rect 144704 106604 145137 106606
rect 144704 106602 144710 106604
rect 145071 106601 145137 106604
rect 146511 106516 146577 106519
rect 140832 106514 146577 106516
rect 140832 106458 146516 106514
rect 146572 106458 146577 106514
rect 140832 106456 146577 106458
rect 146511 106453 146577 106456
rect 209722 106454 209728 106518
rect 209792 106516 209798 106518
rect 210490 106516 210496 106518
rect 209792 106456 210496 106516
rect 209792 106454 209798 106456
rect 210490 106454 210496 106456
rect 210560 106454 210566 106518
rect 668175 106516 668241 106519
rect 665346 106514 668241 106516
rect 665346 106458 668180 106514
rect 668236 106458 668241 106514
rect 665346 106456 668241 106458
rect 665346 106082 665406 106456
rect 668175 106453 668241 106456
rect 140802 104740 140862 105228
rect 665346 105187 665406 105361
rect 665295 105182 665406 105187
rect 665295 105126 665300 105182
rect 665356 105126 665406 105182
rect 665295 105124 665406 105126
rect 665295 105121 665361 105124
rect 674170 105122 674176 105186
rect 674240 105184 674246 105186
rect 675375 105184 675441 105187
rect 674240 105182 675441 105184
rect 674240 105126 675380 105182
rect 675436 105126 675441 105182
rect 674240 105124 675441 105126
rect 674240 105122 674246 105124
rect 675375 105121 675441 105124
rect 146319 104740 146385 104743
rect 140802 104738 146385 104740
rect 140802 104682 146324 104738
rect 146380 104682 146385 104738
rect 140802 104680 146385 104682
rect 146319 104677 146385 104680
rect 665154 104595 665214 104996
rect 665154 104590 665265 104595
rect 665154 104534 665204 104590
rect 665260 104534 665265 104590
rect 665154 104532 665265 104534
rect 665199 104529 665265 104532
rect 645423 104296 645489 104299
rect 640416 104294 645489 104296
rect 640416 104238 645428 104294
rect 645484 104238 645489 104294
rect 640416 104236 645489 104238
rect 645423 104233 645489 104236
rect 141039 104148 141105 104151
rect 146511 104148 146577 104151
rect 141039 104146 146577 104148
rect 141039 104090 141044 104146
rect 141100 104090 146516 104146
rect 146572 104090 146577 104146
rect 141039 104088 146577 104090
rect 141039 104085 141105 104088
rect 146511 104085 146577 104088
rect 140610 103852 140670 103970
rect 141039 103852 141105 103855
rect 140610 103850 141105 103852
rect 140610 103794 141044 103850
rect 141100 103794 141105 103850
rect 140610 103792 141105 103794
rect 141039 103789 141105 103792
rect 675759 103260 675825 103263
rect 675898 103260 675904 103262
rect 675759 103258 675904 103260
rect 675759 103202 675764 103258
rect 675820 103202 675904 103258
rect 675759 103200 675904 103202
rect 675759 103197 675825 103200
rect 675898 103198 675904 103200
rect 675968 103198 675974 103262
rect 146319 102816 146385 102819
rect 140832 102814 146385 102816
rect 140832 102758 146324 102814
rect 146380 102758 146385 102814
rect 140832 102756 146385 102758
rect 146319 102753 146385 102756
rect 204591 102076 204657 102079
rect 204591 102074 210528 102076
rect 204591 102018 204596 102074
rect 204652 102018 210528 102074
rect 204591 102016 210528 102018
rect 204591 102013 204657 102016
rect 146511 101632 146577 101635
rect 140832 101630 146577 101632
rect 140832 101574 146516 101630
rect 146572 101574 146577 101630
rect 140832 101572 146577 101574
rect 146511 101569 146577 101572
rect 204687 101632 204753 101635
rect 204687 101630 210528 101632
rect 204687 101574 204692 101630
rect 204748 101574 210528 101630
rect 204687 101572 210528 101574
rect 204687 101569 204753 101572
rect 675759 101484 675825 101487
rect 676474 101484 676480 101486
rect 675759 101482 676480 101484
rect 675759 101426 675764 101482
rect 675820 101426 676480 101482
rect 675759 101424 676480 101426
rect 675759 101421 675825 101424
rect 676474 101422 676480 101424
rect 676544 101422 676550 101486
rect 204495 101040 204561 101043
rect 204495 101038 210528 101040
rect 204495 100982 204500 101038
rect 204556 100982 210528 101038
rect 204495 100980 210528 100982
rect 204495 100977 204561 100980
rect 198351 100448 198417 100451
rect 198351 100446 210528 100448
rect 198351 100390 198356 100446
rect 198412 100390 210528 100446
rect 198351 100388 210528 100390
rect 198351 100385 198417 100388
rect 140802 99856 140862 100344
rect 210159 99930 210225 99933
rect 210159 99928 210528 99930
rect 210159 99872 210164 99928
rect 210220 99872 210528 99928
rect 210159 99870 210528 99872
rect 210159 99867 210225 99870
rect 146127 99856 146193 99859
rect 140802 99854 146193 99856
rect 140802 99798 146132 99854
rect 146188 99798 146193 99854
rect 140802 99796 146193 99798
rect 146127 99793 146193 99796
rect 201711 99412 201777 99415
rect 201711 99410 210528 99412
rect 201711 99354 201716 99410
rect 201772 99354 210528 99410
rect 201711 99352 210528 99354
rect 201711 99349 201777 99352
rect 146319 99116 146385 99119
rect 140832 99114 146385 99116
rect 140832 99058 146324 99114
rect 146380 99058 146385 99114
rect 140832 99056 146385 99058
rect 146319 99053 146385 99056
rect 204591 98820 204657 98823
rect 204591 98818 210528 98820
rect 204591 98762 204596 98818
rect 204652 98762 210528 98818
rect 204591 98760 210528 98762
rect 204591 98757 204657 98760
rect 194703 98672 194769 98675
rect 194703 98670 210558 98672
rect 194703 98614 194708 98670
rect 194764 98614 210558 98670
rect 194703 98612 210558 98614
rect 194703 98609 194769 98612
rect 210498 98272 210558 98612
rect 146511 98080 146577 98083
rect 140832 98078 146577 98080
rect 140832 98022 146516 98078
rect 146572 98022 146577 98078
rect 140832 98020 146577 98022
rect 146511 98017 146577 98020
rect 207183 97932 207249 97935
rect 208047 97932 208113 97935
rect 207183 97930 208113 97932
rect 207183 97874 207188 97930
rect 207244 97874 208052 97930
rect 208108 97874 208113 97930
rect 207183 97872 208113 97874
rect 207183 97869 207249 97872
rect 208047 97869 208113 97872
rect 200559 97784 200625 97787
rect 200559 97782 210528 97784
rect 200559 97726 200564 97782
rect 200620 97726 210528 97782
rect 200559 97724 210528 97726
rect 200559 97721 200625 97724
rect 201039 97192 201105 97195
rect 201039 97190 210528 97192
rect 201039 97134 201044 97190
rect 201100 97134 210528 97190
rect 201039 97132 210528 97134
rect 201039 97129 201105 97132
rect 140802 96304 140862 96792
rect 210159 96674 210225 96677
rect 210159 96672 210528 96674
rect 210159 96616 210164 96672
rect 210220 96616 210528 96672
rect 210159 96614 210528 96616
rect 210159 96611 210225 96614
rect 146319 96304 146385 96307
rect 140802 96302 146385 96304
rect 140802 96246 146324 96302
rect 146380 96246 146385 96302
rect 140802 96244 146385 96246
rect 146319 96241 146385 96244
rect 200751 96156 200817 96159
rect 200751 96154 210528 96156
rect 200751 96098 200756 96154
rect 200812 96098 210528 96154
rect 200751 96096 210528 96098
rect 200751 96093 200817 96096
rect 146511 95564 146577 95567
rect 140832 95562 146577 95564
rect 140832 95506 146516 95562
rect 146572 95506 146577 95562
rect 140832 95504 146577 95506
rect 146511 95501 146577 95504
rect 201711 95564 201777 95567
rect 201711 95562 210528 95564
rect 201711 95506 201716 95562
rect 201772 95506 210528 95562
rect 201711 95504 210528 95506
rect 201711 95501 201777 95504
rect 210159 95046 210225 95049
rect 210159 95044 210528 95046
rect 210159 94988 210164 95044
rect 210220 94988 210528 95044
rect 210159 94986 210528 94988
rect 210159 94983 210225 94986
rect 201711 94528 201777 94531
rect 201711 94526 210528 94528
rect 201711 94470 201716 94526
rect 201772 94470 210528 94526
rect 201711 94468 210528 94470
rect 201711 94465 201777 94468
rect 146319 94380 146385 94383
rect 140832 94378 146385 94380
rect 140832 94322 146324 94378
rect 146380 94322 146385 94378
rect 140832 94320 146385 94322
rect 146319 94317 146385 94320
rect 203055 93936 203121 93939
rect 203055 93934 210528 93936
rect 203055 93878 203060 93934
rect 203116 93878 210528 93934
rect 203055 93876 210528 93878
rect 203055 93873 203121 93876
rect 195471 93788 195537 93791
rect 195471 93786 210558 93788
rect 195471 93730 195476 93786
rect 195532 93730 210558 93786
rect 195471 93728 210558 93730
rect 195471 93725 195537 93728
rect 210498 93388 210558 93728
rect 140802 92752 140862 93092
rect 201615 92900 201681 92903
rect 201615 92898 210528 92900
rect 201615 92842 201620 92898
rect 201676 92842 210528 92898
rect 201615 92840 210528 92842
rect 201615 92837 201681 92840
rect 146511 92752 146577 92755
rect 140802 92750 146577 92752
rect 140802 92694 146516 92750
rect 146572 92694 146577 92750
rect 140802 92692 146577 92694
rect 146511 92689 146577 92692
rect 194799 92308 194865 92311
rect 194799 92306 210528 92308
rect 194799 92250 194804 92306
rect 194860 92250 210528 92306
rect 194799 92248 210528 92250
rect 194799 92245 194865 92248
rect 140802 91420 140862 91908
rect 210159 91790 210225 91793
rect 210159 91788 210528 91790
rect 210159 91732 210164 91788
rect 210220 91732 210528 91788
rect 210159 91730 210528 91732
rect 210159 91727 210225 91730
rect 146319 91420 146385 91423
rect 140802 91418 146385 91420
rect 140802 91362 146324 91418
rect 146380 91362 146385 91418
rect 140802 91360 146385 91362
rect 146319 91357 146385 91360
rect 200175 91272 200241 91275
rect 200175 91270 210528 91272
rect 200175 91214 200180 91270
rect 200236 91214 210528 91270
rect 200175 91212 210528 91214
rect 200175 91209 200241 91212
rect 210106 90914 210112 90978
rect 210176 90976 210182 90978
rect 210490 90976 210496 90978
rect 210176 90916 210496 90976
rect 210176 90914 210182 90916
rect 210490 90914 210496 90916
rect 210560 90914 210566 90978
rect 146511 90828 146577 90831
rect 140832 90826 146577 90828
rect 140832 90770 146516 90826
rect 146572 90770 146577 90826
rect 140832 90768 146577 90770
rect 146511 90765 146577 90768
rect 197295 90680 197361 90683
rect 197295 90678 210528 90680
rect 197295 90622 197300 90678
rect 197356 90622 210528 90678
rect 197295 90620 210528 90622
rect 197295 90617 197361 90620
rect 210106 90322 210112 90386
rect 210176 90384 210182 90386
rect 211066 90384 211072 90386
rect 210176 90324 211072 90384
rect 210176 90322 210182 90324
rect 211066 90322 211072 90324
rect 211136 90322 211142 90386
rect 194415 90088 194481 90091
rect 194415 90086 210528 90088
rect 194415 90030 194420 90086
rect 194476 90030 210528 90086
rect 194415 90028 210528 90030
rect 194415 90025 194481 90028
rect 146127 89644 146193 89647
rect 140832 89642 146193 89644
rect 140832 89586 146132 89642
rect 146188 89586 146193 89642
rect 140832 89584 146193 89586
rect 146127 89581 146193 89584
rect 201711 89644 201777 89647
rect 201711 89642 210528 89644
rect 201711 89586 201716 89642
rect 201772 89586 210528 89642
rect 201711 89584 210528 89586
rect 201711 89581 201777 89584
rect 210682 89286 210688 89350
rect 210752 89348 210758 89350
rect 211066 89348 211072 89350
rect 210752 89288 211072 89348
rect 210752 89286 210758 89288
rect 211066 89286 211072 89288
rect 211136 89286 211142 89350
rect 201711 89052 201777 89055
rect 647535 89052 647601 89055
rect 201711 89050 210528 89052
rect 201711 88994 201716 89050
rect 201772 88994 210528 89050
rect 201711 88992 210528 88994
rect 640416 89050 647601 89052
rect 640416 88994 647540 89050
rect 647596 88994 647601 89050
rect 640416 88992 647601 88994
rect 201711 88989 201777 88992
rect 647535 88989 647601 88992
rect 201327 88460 201393 88463
rect 201327 88458 210528 88460
rect 201327 88402 201332 88458
rect 201388 88402 210528 88458
rect 201327 88400 210528 88402
rect 201327 88397 201393 88400
rect 140802 87868 140862 88356
rect 640194 88164 640254 88430
rect 645807 88164 645873 88167
rect 640194 88162 645873 88164
rect 640194 88106 645812 88162
rect 645868 88106 645873 88162
rect 640194 88104 645873 88106
rect 645807 88101 645873 88104
rect 201615 88016 201681 88019
rect 201615 88014 210528 88016
rect 201615 87958 201620 88014
rect 201676 87958 210528 88014
rect 201615 87956 210528 87958
rect 201615 87953 201681 87956
rect 144207 87868 144273 87871
rect 140802 87866 144273 87868
rect 140802 87810 144212 87866
rect 144268 87810 144273 87866
rect 140802 87808 144273 87810
rect 144207 87805 144273 87808
rect 210298 87658 210304 87722
rect 210368 87720 210374 87722
rect 211066 87720 211072 87722
rect 210368 87660 211072 87720
rect 210368 87658 210374 87660
rect 211066 87658 211072 87660
rect 211136 87658 211142 87722
rect 640386 87720 640446 87986
rect 645423 87720 645489 87723
rect 640386 87718 645489 87720
rect 640386 87662 645428 87718
rect 645484 87662 645489 87718
rect 640386 87660 645489 87662
rect 645423 87657 645489 87660
rect 201807 87424 201873 87427
rect 647631 87424 647697 87427
rect 201807 87422 210528 87424
rect 201807 87366 201812 87422
rect 201868 87366 210528 87422
rect 201807 87364 210528 87366
rect 640416 87422 647697 87424
rect 640416 87366 647636 87422
rect 647692 87366 647697 87422
rect 640416 87364 647697 87366
rect 201807 87361 201873 87364
rect 647631 87361 647697 87364
rect 210682 87214 210688 87278
rect 210752 87276 210758 87278
rect 211066 87276 211072 87278
rect 210752 87216 211072 87276
rect 210752 87214 210758 87216
rect 211066 87214 211072 87216
rect 211136 87214 211142 87278
rect 144111 87128 144177 87131
rect 140832 87126 144177 87128
rect 140832 87070 144116 87126
rect 144172 87070 144177 87126
rect 140832 87068 144177 87070
rect 144111 87065 144177 87068
rect 650895 86980 650961 86983
rect 650895 86978 656736 86980
rect 650895 86922 650900 86978
rect 650956 86922 656736 86978
rect 650895 86920 656736 86922
rect 650895 86917 650961 86920
rect 197871 86832 197937 86835
rect 197871 86830 210528 86832
rect 197871 86774 197876 86830
rect 197932 86774 210528 86830
rect 197871 86772 210528 86774
rect 197871 86769 197937 86772
rect 640194 86684 640254 86802
rect 645807 86684 645873 86687
rect 640194 86682 645873 86684
rect 640194 86626 645812 86682
rect 645868 86626 645873 86682
rect 640194 86624 645873 86626
rect 645807 86621 645873 86624
rect 201615 86388 201681 86391
rect 201615 86386 210528 86388
rect 201615 86330 201620 86386
rect 201676 86330 210528 86386
rect 201615 86328 210528 86330
rect 201615 86325 201681 86328
rect 640386 86240 640446 86358
rect 647823 86240 647889 86243
rect 640386 86238 647889 86240
rect 640386 86182 647828 86238
rect 647884 86182 647889 86238
rect 640386 86180 647889 86182
rect 647823 86177 647889 86180
rect 651183 86240 651249 86243
rect 651183 86238 656736 86240
rect 651183 86182 651188 86238
rect 651244 86182 656736 86238
rect 651183 86180 656736 86182
rect 651183 86177 651249 86180
rect 146511 85944 146577 85947
rect 140832 85942 146577 85944
rect 140832 85886 146516 85942
rect 146572 85886 146577 85942
rect 140832 85884 146577 85886
rect 146511 85881 146577 85884
rect 197775 85796 197841 85799
rect 647247 85796 647313 85799
rect 197775 85794 210528 85796
rect 197775 85738 197780 85794
rect 197836 85738 210528 85794
rect 197775 85736 210528 85738
rect 640416 85794 647313 85796
rect 640416 85738 647252 85794
rect 647308 85738 647313 85794
rect 640416 85736 647313 85738
rect 197775 85733 197841 85736
rect 647247 85733 647313 85736
rect 663426 85651 663486 86210
rect 663426 85646 663537 85651
rect 663426 85590 663476 85646
rect 663532 85590 663537 85646
rect 663426 85588 663537 85590
rect 663471 85585 663537 85588
rect 647727 85500 647793 85503
rect 640386 85498 647793 85500
rect 640386 85442 647732 85498
rect 647788 85442 647793 85498
rect 640386 85440 647793 85442
rect 201711 85204 201777 85207
rect 201711 85202 210528 85204
rect 201711 85146 201716 85202
rect 201772 85146 210528 85202
rect 640386 85174 640446 85440
rect 647727 85437 647793 85440
rect 650991 85352 651057 85355
rect 650991 85350 656736 85352
rect 650991 85294 650996 85350
rect 651052 85294 656736 85350
rect 650991 85292 656736 85294
rect 650991 85289 651057 85292
rect 663279 85204 663345 85207
rect 663234 85202 663345 85204
rect 201711 85144 210528 85146
rect 663234 85146 663284 85202
rect 663340 85146 663345 85202
rect 201711 85141 201777 85144
rect 663234 85141 663345 85146
rect 645423 85056 645489 85059
rect 640194 85054 645489 85056
rect 640194 84998 645428 85054
rect 645484 84998 645489 85054
rect 640194 84996 645489 84998
rect 198735 84760 198801 84763
rect 198735 84758 210528 84760
rect 198735 84702 198740 84758
rect 198796 84702 210528 84758
rect 640194 84730 640254 84996
rect 645423 84993 645489 84996
rect 198735 84700 210528 84702
rect 198735 84697 198801 84700
rect 140802 84168 140862 84656
rect 663234 84582 663294 85141
rect 663426 84763 663486 85322
rect 663375 84758 663486 84763
rect 663375 84702 663380 84758
rect 663436 84702 663486 84758
rect 663375 84700 663486 84702
rect 663375 84697 663441 84700
rect 650991 84316 651057 84319
rect 650991 84314 656736 84316
rect 650991 84258 650996 84314
rect 651052 84258 656736 84314
rect 650991 84256 656736 84258
rect 650991 84253 651057 84256
rect 145071 84168 145137 84171
rect 140802 84166 145137 84168
rect 140802 84110 145076 84166
rect 145132 84110 145137 84166
rect 140802 84108 145137 84110
rect 145071 84105 145137 84108
rect 201807 84168 201873 84171
rect 645807 84168 645873 84171
rect 201807 84166 210528 84168
rect 201807 84110 201812 84166
rect 201868 84110 210528 84166
rect 201807 84108 210528 84110
rect 640416 84166 645873 84168
rect 640416 84110 645812 84166
rect 645868 84110 645873 84166
rect 640416 84108 645873 84110
rect 201807 84105 201873 84108
rect 645807 84105 645873 84108
rect 650607 83872 650673 83875
rect 640386 83870 650673 83872
rect 640386 83814 650612 83870
rect 650668 83814 650673 83870
rect 640386 83812 650673 83814
rect 140802 83576 140862 83618
rect 146127 83576 146193 83579
rect 140802 83574 146193 83576
rect 140802 83518 146132 83574
rect 146188 83518 146193 83574
rect 140802 83516 146193 83518
rect 146127 83513 146193 83516
rect 196047 83576 196113 83579
rect 196047 83574 210528 83576
rect 196047 83518 196052 83574
rect 196108 83518 210528 83574
rect 640386 83546 640446 83812
rect 650607 83809 650673 83812
rect 196047 83516 210528 83518
rect 196047 83513 196113 83516
rect 651087 83428 651153 83431
rect 651087 83426 656736 83428
rect 651087 83370 651092 83426
rect 651148 83370 656736 83426
rect 651087 83368 656736 83370
rect 651087 83365 651153 83368
rect 645423 83280 645489 83283
rect 640194 83278 645489 83280
rect 640194 83222 645428 83278
rect 645484 83222 645489 83278
rect 640194 83220 645489 83222
rect 201711 83132 201777 83135
rect 201711 83130 210528 83132
rect 201711 83074 201716 83130
rect 201772 83074 210528 83130
rect 640194 83102 640254 83220
rect 645423 83217 645489 83220
rect 201711 83072 210528 83074
rect 201711 83069 201777 83072
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 210106 82626 210112 82690
rect 210176 82688 210182 82690
rect 210874 82688 210880 82690
rect 210176 82628 210880 82688
rect 210176 82626 210182 82628
rect 210874 82626 210880 82628
rect 210944 82626 210950 82690
rect 650895 82688 650961 82691
rect 650895 82686 656736 82688
rect 650895 82630 650900 82686
rect 650956 82630 656736 82686
rect 650895 82628 656736 82630
rect 650895 82625 650961 82628
rect 201615 82540 201681 82543
rect 645423 82540 645489 82543
rect 201615 82538 210528 82540
rect 201615 82482 201620 82538
rect 201676 82482 210528 82538
rect 201615 82480 210528 82482
rect 640416 82538 645489 82540
rect 640416 82482 645428 82538
rect 645484 82482 645489 82538
rect 640416 82480 645489 82482
rect 201615 82477 201681 82480
rect 645423 82477 645489 82480
rect 146511 82392 146577 82395
rect 140832 82390 146577 82392
rect 42252 82360 45378 82362
rect 40792 82346 45378 82360
rect 38346 82236 45378 82346
rect 140832 82334 146516 82390
rect 146572 82334 146577 82390
rect 140832 82332 146577 82334
rect 146511 82329 146577 82332
rect 647439 82244 647505 82247
rect 38346 78432 40974 82236
rect 40792 72776 40974 78432
rect 38544 69066 40974 72776
rect 45006 69066 45378 82236
rect 640386 82242 647505 82244
rect 640386 82186 647444 82242
rect 647500 82186 647505 82242
rect 640386 82184 647505 82186
rect 201711 81948 201777 81951
rect 201711 81946 210528 81948
rect 201711 81890 201716 81946
rect 201772 81890 210528 81946
rect 640386 81918 640446 82184
rect 647439 82181 647505 82184
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 201711 81888 210528 81890
rect 201711 81885 201777 81888
rect 201807 81504 201873 81507
rect 201807 81502 210528 81504
rect 201807 81446 201812 81502
rect 201868 81446 210528 81502
rect 201807 81444 210528 81446
rect 201807 81441 201873 81444
rect 640386 81356 640446 81474
rect 645423 81356 645489 81359
rect 640386 81354 645489 81356
rect 640386 81298 645428 81354
rect 645484 81298 645489 81354
rect 640386 81296 645489 81298
rect 645423 81293 645489 81296
rect 662895 81208 662961 81211
rect 663042 81208 663102 81770
rect 662895 81206 663102 81208
rect 140802 80764 140862 81170
rect 662895 81150 662900 81206
rect 662956 81150 663102 81206
rect 662895 81148 663102 81150
rect 662895 81145 662961 81148
rect 201519 80912 201585 80915
rect 646191 80912 646257 80915
rect 201519 80910 210528 80912
rect 201519 80854 201524 80910
rect 201580 80854 210528 80910
rect 201519 80852 210528 80854
rect 640416 80910 646257 80912
rect 640416 80854 646196 80910
rect 646252 80854 646257 80910
rect 640416 80852 646257 80854
rect 201519 80849 201585 80852
rect 646191 80849 646257 80852
rect 144591 80764 144657 80767
rect 140802 80762 144657 80764
rect 140802 80706 144596 80762
rect 144652 80706 144657 80762
rect 140802 80704 144657 80706
rect 144591 80701 144657 80704
rect 203151 80320 203217 80323
rect 203151 80318 210528 80320
rect 203151 80262 203156 80318
rect 203212 80262 210528 80318
rect 203151 80260 210528 80262
rect 203151 80257 203217 80260
rect 200271 80172 200337 80175
rect 640194 80172 640254 80290
rect 645999 80172 646065 80175
rect 200271 80170 210558 80172
rect 200271 80114 200276 80170
rect 200332 80114 210558 80170
rect 200271 80112 210558 80114
rect 640194 80170 646065 80172
rect 640194 80114 646004 80170
rect 646060 80114 646065 80170
rect 640194 80112 646065 80114
rect 200271 80109 200337 80112
rect 140802 79432 140862 79920
rect 210498 79772 210558 80112
rect 645999 80109 646065 80112
rect 645423 80024 645489 80027
rect 640386 80022 645489 80024
rect 640386 79966 645428 80022
rect 645484 79966 645489 80022
rect 640386 79964 645489 79966
rect 640386 79772 640446 79964
rect 645423 79961 645489 79964
rect 146319 79432 146385 79435
rect 140802 79430 146385 79432
rect 140802 79374 146324 79430
rect 146380 79374 146385 79430
rect 140802 79372 146385 79374
rect 146319 79369 146385 79372
rect 197391 79284 197457 79287
rect 645807 79284 645873 79287
rect 197391 79282 210528 79284
rect 197391 79226 197396 79282
rect 197452 79226 210528 79282
rect 197391 79224 210528 79226
rect 640416 79282 645873 79284
rect 640416 79226 645812 79282
rect 645868 79226 645873 79282
rect 640416 79224 645873 79226
rect 197391 79221 197457 79224
rect 645807 79221 645873 79224
rect 146511 78692 146577 78695
rect 140832 78690 146577 78692
rect 140832 78634 146516 78690
rect 146572 78634 146577 78690
rect 140832 78632 146577 78634
rect 146511 78629 146577 78632
rect 194511 78692 194577 78695
rect 645423 78692 645489 78695
rect 194511 78690 210528 78692
rect 194511 78634 194516 78690
rect 194572 78634 210528 78690
rect 194511 78632 210528 78634
rect 640416 78690 645489 78692
rect 640416 78634 645428 78690
rect 645484 78634 645489 78690
rect 640416 78632 645489 78634
rect 194511 78629 194577 78632
rect 645423 78629 645489 78632
rect 645903 78544 645969 78547
rect 640386 78542 645969 78544
rect 640386 78486 645908 78542
rect 645964 78486 645969 78542
rect 640386 78484 645969 78486
rect 210159 78174 210225 78177
rect 210159 78172 210528 78174
rect 210159 78116 210164 78172
rect 210220 78116 210528 78172
rect 640386 78144 640446 78484
rect 645903 78481 645969 78484
rect 210159 78114 210528 78116
rect 210159 78111 210225 78114
rect 201711 77656 201777 77659
rect 645423 77656 645489 77659
rect 201711 77654 210528 77656
rect 201711 77598 201716 77654
rect 201772 77598 210528 77654
rect 201711 77596 210528 77598
rect 640416 77654 645489 77656
rect 640416 77598 645428 77654
rect 645484 77598 645489 77654
rect 640416 77596 645489 77598
rect 201711 77593 201777 77596
rect 645423 77593 645489 77596
rect 144399 77508 144465 77511
rect 140832 77506 144465 77508
rect 140832 77450 144404 77506
rect 144460 77450 144465 77506
rect 140832 77448 144465 77450
rect 144399 77445 144465 77448
rect 201711 77064 201777 77067
rect 645423 77064 645489 77067
rect 201711 77062 210528 77064
rect 201711 77006 201716 77062
rect 201772 77006 210528 77062
rect 201711 77004 210528 77006
rect 640416 77062 645489 77064
rect 640416 77006 645428 77062
rect 645484 77006 645489 77062
rect 640416 77004 645489 77006
rect 201711 77001 201777 77004
rect 645423 77001 645489 77004
rect 645423 76768 645489 76771
rect 640386 76766 645489 76768
rect 640386 76710 645428 76766
rect 645484 76710 645489 76766
rect 640386 76708 645489 76710
rect 210159 76546 210225 76549
rect 210159 76544 210528 76546
rect 210159 76488 210164 76544
rect 210220 76488 210528 76544
rect 640386 76516 640446 76708
rect 645423 76705 645489 76708
rect 210159 76486 210528 76488
rect 210159 76483 210225 76486
rect 140802 75732 140862 76220
rect 200271 76028 200337 76031
rect 645807 76028 645873 76031
rect 200271 76026 210528 76028
rect 200271 75970 200276 76026
rect 200332 75970 210528 76026
rect 200271 75968 210528 75970
rect 640416 76026 645873 76028
rect 640416 75970 645812 76026
rect 645868 75970 645873 76026
rect 640416 75968 645873 75970
rect 200271 75965 200337 75968
rect 645807 75965 645873 75968
rect 146319 75732 146385 75735
rect 140802 75730 146385 75732
rect 140802 75674 146324 75730
rect 146380 75674 146385 75730
rect 140802 75672 146385 75674
rect 146319 75669 146385 75672
rect 201615 75436 201681 75439
rect 645423 75436 645489 75439
rect 201615 75434 210528 75436
rect 201615 75378 201620 75434
rect 201676 75378 210528 75434
rect 201615 75376 210528 75378
rect 640416 75434 645489 75436
rect 640416 75378 645428 75434
rect 645484 75378 645489 75434
rect 640416 75376 645489 75378
rect 201615 75373 201681 75376
rect 645423 75373 645489 75376
rect 196911 75288 196977 75291
rect 645903 75288 645969 75291
rect 196911 75286 210558 75288
rect 196911 75230 196916 75286
rect 196972 75230 210558 75286
rect 196911 75228 210558 75230
rect 196911 75225 196977 75228
rect 140802 75140 140862 75184
rect 144015 75140 144081 75143
rect 140802 75138 144081 75140
rect 140802 75082 144020 75138
rect 144076 75082 144081 75138
rect 140802 75080 144081 75082
rect 144015 75077 144081 75080
rect 210498 74888 210558 75228
rect 640386 75286 645969 75288
rect 640386 75230 645908 75286
rect 645964 75230 645969 75286
rect 640386 75228 645969 75230
rect 640386 74888 640446 75228
rect 645903 75225 645969 75228
rect 201711 74400 201777 74403
rect 645423 74400 645489 74403
rect 201711 74398 210528 74400
rect 201711 74342 201716 74398
rect 201772 74342 210528 74398
rect 201711 74340 210528 74342
rect 640416 74398 645489 74400
rect 640416 74342 645428 74398
rect 645484 74342 645489 74398
rect 640416 74340 645489 74342
rect 201711 74337 201777 74340
rect 645423 74337 645489 74340
rect 146703 73956 146769 73959
rect 140832 73954 146769 73956
rect 140832 73898 146708 73954
rect 146764 73898 146769 73954
rect 140832 73896 146769 73898
rect 146703 73893 146769 73896
rect 201615 73808 201681 73811
rect 645807 73808 645873 73811
rect 201615 73806 210528 73808
rect 201615 73750 201620 73806
rect 201676 73750 210528 73806
rect 201615 73748 210528 73750
rect 640416 73806 645873 73808
rect 640416 73750 645812 73806
rect 645868 73750 645873 73806
rect 640416 73748 645873 73750
rect 201615 73745 201681 73748
rect 645807 73745 645873 73748
rect 210159 73290 210225 73293
rect 210159 73288 210528 73290
rect 210159 73232 210164 73288
rect 210220 73232 210528 73288
rect 210159 73230 210528 73232
rect 210159 73227 210225 73230
rect 210106 72858 210112 72922
rect 210176 72920 210182 72922
rect 211066 72920 211072 72922
rect 210176 72860 211072 72920
rect 210176 72858 210182 72860
rect 211066 72858 211072 72860
rect 211136 72858 211142 72922
rect 640386 72920 640446 73260
rect 645423 72920 645489 72923
rect 640386 72918 645489 72920
rect 640386 72862 645428 72918
rect 645484 72862 645489 72918
rect 640386 72860 645489 72862
rect 645423 72857 645489 72860
rect 144399 72772 144465 72775
rect 140832 72770 144465 72772
rect 140832 72714 144404 72770
rect 144460 72714 144465 72770
rect 140832 72712 144465 72714
rect 144399 72709 144465 72712
rect 201807 72772 201873 72775
rect 646383 72772 646449 72775
rect 201807 72770 210528 72772
rect 201807 72714 201812 72770
rect 201868 72714 210528 72770
rect 201807 72712 210528 72714
rect 640416 72770 646449 72772
rect 640416 72714 646388 72770
rect 646444 72714 646449 72770
rect 640416 72712 646449 72714
rect 201807 72709 201873 72712
rect 646383 72709 646449 72712
rect 201519 72180 201585 72183
rect 646671 72180 646737 72183
rect 201519 72178 210528 72180
rect 201519 72122 201524 72178
rect 201580 72122 210528 72178
rect 201519 72120 210528 72122
rect 640416 72178 646737 72180
rect 640416 72122 646676 72178
rect 646732 72122 646737 72178
rect 640416 72120 646737 72122
rect 201519 72117 201585 72120
rect 646671 72117 646737 72120
rect 209967 71662 210033 71665
rect 209967 71660 210528 71662
rect 209967 71604 209972 71660
rect 210028 71604 210528 71660
rect 209967 71602 210528 71604
rect 209967 71599 210033 71602
rect 140802 70996 140862 71484
rect 201711 71144 201777 71147
rect 201711 71142 210528 71144
rect 201711 71086 201716 71142
rect 201772 71086 210528 71142
rect 201711 71084 210528 71086
rect 201711 71081 201777 71084
rect 146703 70996 146769 70999
rect 140802 70994 146769 70996
rect 140802 70938 146708 70994
rect 146764 70938 146769 70994
rect 140802 70936 146769 70938
rect 146703 70933 146769 70936
rect 201615 70552 201681 70555
rect 201615 70550 210528 70552
rect 201615 70494 201620 70550
rect 201676 70494 210528 70550
rect 201615 70492 210528 70494
rect 201615 70489 201681 70492
rect 140802 69812 140862 70290
rect 200367 69960 200433 69963
rect 200367 69958 210528 69960
rect 200367 69902 200372 69958
rect 200428 69902 210528 69958
rect 200367 69900 210528 69902
rect 200367 69897 200433 69900
rect 144015 69812 144081 69815
rect 140802 69810 144081 69812
rect 140802 69754 144020 69810
rect 144076 69754 144081 69810
rect 140802 69752 144081 69754
rect 144015 69749 144081 69752
rect 201807 69516 201873 69519
rect 201807 69514 210528 69516
rect 201807 69458 201812 69514
rect 201868 69458 210528 69514
rect 201807 69456 210528 69458
rect 201807 69453 201873 69456
rect 145839 69072 145905 69075
rect 38544 68996 45378 69066
rect 140832 69070 145905 69072
rect 140832 69014 145844 69070
rect 145900 69014 145905 69070
rect 140832 69012 145905 69014
rect 145839 69009 145905 69012
rect 40792 68974 45378 68996
rect 40792 68966 45220 68974
rect 195471 68924 195537 68927
rect 195471 68922 210528 68924
rect 195471 68866 195476 68922
rect 195532 68866 210528 68922
rect 195471 68864 210528 68866
rect 195471 68861 195537 68864
rect 196239 68332 196305 68335
rect 196239 68330 210528 68332
rect 196239 68274 196244 68330
rect 196300 68274 210528 68330
rect 196239 68272 210528 68274
rect 196239 68269 196305 68272
rect 140802 67444 140862 67932
rect 201711 67888 201777 67891
rect 201711 67886 210528 67888
rect 201711 67830 201716 67886
rect 201772 67830 210528 67886
rect 201711 67828 210528 67830
rect 201711 67825 201777 67828
rect 146703 67444 146769 67447
rect 140802 67442 146769 67444
rect 140802 67386 146708 67442
rect 146764 67386 146769 67442
rect 140802 67384 146769 67386
rect 146703 67381 146769 67384
rect 201615 67296 201681 67299
rect 201615 67294 210528 67296
rect 201615 67238 201620 67294
rect 201676 67238 210528 67294
rect 201615 67236 210528 67238
rect 201615 67233 201681 67236
rect 140802 66408 140862 66748
rect 201807 66704 201873 66707
rect 201807 66702 210528 66704
rect 201807 66646 201812 66702
rect 201868 66646 210528 66702
rect 201807 66644 210528 66646
rect 201807 66641 201873 66644
rect 146799 66408 146865 66411
rect 140802 66406 146865 66408
rect 140802 66350 146804 66406
rect 146860 66350 146865 66406
rect 140802 66348 146865 66350
rect 146799 66345 146865 66348
rect 193647 66260 193713 66263
rect 193647 66258 210528 66260
rect 193647 66202 193652 66258
rect 193708 66202 210528 66258
rect 193647 66200 210528 66202
rect 193647 66197 193713 66200
rect 198543 65668 198609 65671
rect 198543 65666 210528 65668
rect 198543 65610 198548 65666
rect 198604 65610 210528 65666
rect 198543 65608 210528 65610
rect 198543 65605 198609 65608
rect 146703 65520 146769 65523
rect 140832 65518 146769 65520
rect 140832 65462 146708 65518
rect 146764 65462 146769 65518
rect 140832 65460 146769 65462
rect 146703 65457 146769 65460
rect 201711 65076 201777 65079
rect 201711 65074 210528 65076
rect 201711 65018 201716 65074
rect 201772 65018 210528 65074
rect 201711 65016 210528 65018
rect 201711 65013 201777 65016
rect 146799 64780 146865 64783
rect 140802 64778 146865 64780
rect 140802 64722 146804 64778
rect 146860 64722 146865 64778
rect 140802 64720 146865 64722
rect 140802 64334 140862 64720
rect 146799 64717 146865 64720
rect 201711 64632 201777 64635
rect 201711 64630 210528 64632
rect 201711 64574 201716 64630
rect 201772 64574 210528 64630
rect 201711 64572 210528 64574
rect 201711 64569 201777 64572
rect 201807 64040 201873 64043
rect 201807 64038 210528 64040
rect 201807 63982 201812 64038
rect 201868 63982 210528 64038
rect 201807 63980 210528 63982
rect 201807 63977 201873 63980
rect 195471 63448 195537 63451
rect 195471 63446 210528 63448
rect 195471 63390 195476 63446
rect 195532 63390 210528 63446
rect 195471 63388 210528 63390
rect 195471 63385 195537 63388
rect 140802 62560 140862 63048
rect 201711 63004 201777 63007
rect 201711 63002 210528 63004
rect 201711 62946 201716 63002
rect 201772 62946 210528 63002
rect 201711 62944 210528 62946
rect 201711 62941 201777 62944
rect 209487 62856 209553 62859
rect 209914 62856 209920 62858
rect 209487 62854 209920 62856
rect 209487 62798 209492 62854
rect 209548 62798 209920 62854
rect 209487 62796 209920 62798
rect 209487 62793 209553 62796
rect 209914 62794 209920 62796
rect 209984 62794 209990 62858
rect 146799 62560 146865 62563
rect 140802 62558 146865 62560
rect 140802 62502 146804 62558
rect 146860 62502 146865 62558
rect 140802 62500 146865 62502
rect 146799 62497 146865 62500
rect 210159 62560 210225 62563
rect 210298 62560 210304 62562
rect 210159 62558 210304 62560
rect 210159 62502 210164 62558
rect 210220 62502 210304 62558
rect 210159 62500 210304 62502
rect 210159 62497 210225 62500
rect 210298 62498 210304 62500
rect 210368 62498 210374 62562
rect 146895 62412 146961 62415
rect 140802 62410 146961 62412
rect 140802 62354 146900 62410
rect 146956 62354 146961 62410
rect 140802 62352 146961 62354
rect 140802 61864 140862 62352
rect 146895 62349 146961 62352
rect 201615 62412 201681 62415
rect 201615 62410 210528 62412
rect 201615 62354 201620 62410
rect 201676 62354 210528 62410
rect 201615 62352 210528 62354
rect 201615 62349 201681 62352
rect 201519 61820 201585 61823
rect 201519 61818 210528 61820
rect 201519 61762 201524 61818
rect 201580 61762 210528 61818
rect 201519 61760 210528 61762
rect 201519 61757 201585 61760
rect 201807 61376 201873 61379
rect 201807 61374 210528 61376
rect 201807 61318 201812 61374
rect 201868 61318 210528 61374
rect 201807 61316 210528 61318
rect 201807 61313 201873 61316
rect 146895 60784 146961 60787
rect 140832 60782 146961 60784
rect 140832 60726 146900 60782
rect 146956 60726 146961 60782
rect 140832 60724 146961 60726
rect 146895 60721 146961 60724
rect 195471 60784 195537 60787
rect 195471 60782 210528 60784
rect 195471 60726 195476 60782
rect 195532 60726 210528 60782
rect 195471 60724 210528 60726
rect 195471 60721 195537 60724
rect 201711 60192 201777 60195
rect 201711 60190 210528 60192
rect 201711 60134 201716 60190
rect 201772 60134 210528 60190
rect 201711 60132 210528 60134
rect 201711 60129 201777 60132
rect 209967 59674 210033 59677
rect 209967 59672 210528 59674
rect 209967 59616 209972 59672
rect 210028 59616 210528 59672
rect 209967 59614 210528 59616
rect 209967 59611 210033 59614
rect 146799 59600 146865 59603
rect 140832 59598 146865 59600
rect 140832 59542 146804 59598
rect 146860 59542 146865 59598
rect 140832 59540 146865 59542
rect 146799 59537 146865 59540
rect 198351 59156 198417 59159
rect 198351 59154 210528 59156
rect 198351 59098 198356 59154
rect 198412 59098 210528 59154
rect 198351 59096 210528 59098
rect 198351 59093 198417 59096
rect 146799 58712 146865 58715
rect 140802 58710 146865 58712
rect 140802 58654 146804 58710
rect 146860 58654 146865 58710
rect 140802 58652 146865 58654
rect 140802 58322 140862 58652
rect 146799 58649 146865 58652
rect 211074 58270 211134 58534
rect 211066 58206 211072 58270
rect 211136 58206 211142 58270
rect 210255 58046 210321 58049
rect 210255 58044 210528 58046
rect 210255 57988 210260 58044
rect 210316 57988 210528 58044
rect 210255 57986 210528 57988
rect 210255 57983 210321 57986
rect 206991 57528 207057 57531
rect 206991 57526 210528 57528
rect 206991 57470 206996 57526
rect 207052 57470 210528 57526
rect 206991 57468 210528 57470
rect 206991 57465 207057 57468
rect 146799 57084 146865 57087
rect 140832 57082 146865 57084
rect 140832 57026 146804 57082
rect 146860 57026 146865 57082
rect 140832 57024 146865 57026
rect 146799 57021 146865 57024
rect 210255 56936 210321 56939
rect 210255 56934 210528 56936
rect 210255 56878 210260 56934
rect 210316 56878 210528 56934
rect 210255 56876 210528 56878
rect 210255 56873 210321 56876
rect 144015 56492 144081 56495
rect 140802 56490 144081 56492
rect 140802 56434 144020 56490
rect 144076 56434 144081 56490
rect 140802 56432 144081 56434
rect 140802 55874 140862 56432
rect 144015 56429 144081 56432
rect 209967 56418 210033 56421
rect 209967 56416 210528 56418
rect 209967 56360 209972 56416
rect 210028 56360 210528 56416
rect 209967 56358 210528 56360
rect 209967 56355 210033 56358
rect 206895 55900 206961 55903
rect 206895 55898 210528 55900
rect 206895 55842 206900 55898
rect 206956 55842 210528 55898
rect 206895 55840 210528 55842
rect 206895 55837 206961 55840
rect 210159 55308 210225 55311
rect 210159 55306 210528 55308
rect 210159 55250 210164 55306
rect 210220 55250 210528 55306
rect 210159 55248 210528 55250
rect 210159 55245 210225 55248
rect 144783 54716 144849 54719
rect 140832 54714 144849 54716
rect 140832 54658 144788 54714
rect 144844 54658 144849 54714
rect 140832 54656 144849 54658
rect 144783 54653 144849 54656
rect 210690 54275 210750 54760
rect 210298 54210 210304 54274
rect 210368 54272 210374 54274
rect 210447 54272 210513 54275
rect 210368 54270 210513 54272
rect 210368 54214 210452 54270
rect 210508 54214 210513 54270
rect 210368 54212 210513 54214
rect 210368 54210 210374 54212
rect 210447 54209 210513 54212
rect 210639 54270 210750 54275
rect 210639 54214 210644 54270
rect 210700 54214 210750 54270
rect 210639 54212 210750 54214
rect 210639 54209 210705 54212
rect 211642 54210 211648 54274
rect 211712 54272 211718 54274
rect 214767 54272 214833 54275
rect 211712 54270 214833 54272
rect 211712 54214 214772 54270
rect 214828 54214 214833 54270
rect 211712 54212 214833 54214
rect 211712 54210 211718 54212
rect 214767 54209 214833 54212
rect 144495 54124 144561 54127
rect 140802 54122 144561 54124
rect 140802 54066 144500 54122
rect 144556 54066 144561 54122
rect 140802 54064 144561 54066
rect 140802 53576 140862 54064
rect 144495 54061 144561 54064
rect 209914 54062 209920 54126
rect 209984 54124 209990 54126
rect 210255 54124 210321 54127
rect 209984 54122 210321 54124
rect 209984 54066 210260 54122
rect 210316 54066 210321 54122
rect 209984 54064 210321 54066
rect 209984 54062 209990 54064
rect 210255 54061 210321 54064
rect 212794 54062 212800 54126
rect 212864 54124 212870 54126
rect 216975 54124 217041 54127
rect 212864 54122 217041 54124
rect 212864 54066 216980 54122
rect 217036 54066 217041 54122
rect 212864 54064 217041 54066
rect 212864 54062 212870 54064
rect 216975 54061 217041 54064
rect 211066 53914 211072 53978
rect 211136 53976 211142 53978
rect 216975 53976 217041 53979
rect 211136 53974 217041 53976
rect 211136 53918 216980 53974
rect 217036 53918 217041 53974
rect 211136 53916 217041 53918
rect 211136 53914 211142 53916
rect 216975 53913 217041 53916
rect 209722 53766 209728 53830
rect 209792 53828 209798 53830
rect 209792 53768 221166 53828
rect 209792 53766 209798 53768
rect 212218 53618 212224 53682
rect 212288 53680 212294 53682
rect 212288 53620 216030 53680
rect 212288 53618 212294 53620
rect 215970 53535 216030 53620
rect 221106 53535 221166 53768
rect 213039 53534 213105 53535
rect 212986 53532 212992 53534
rect 212948 53472 212992 53532
rect 213056 53530 213105 53534
rect 213100 53474 213105 53530
rect 212986 53470 212992 53472
rect 213056 53470 213105 53474
rect 213039 53469 213105 53470
rect 214959 53532 215025 53535
rect 215775 53532 215841 53535
rect 214959 53530 215841 53532
rect 214959 53474 214964 53530
rect 215020 53474 215780 53530
rect 215836 53474 215841 53530
rect 214959 53472 215841 53474
rect 214959 53469 215025 53472
rect 215775 53469 215841 53472
rect 215967 53530 216033 53535
rect 215967 53474 215972 53530
rect 216028 53474 216033 53530
rect 215967 53469 216033 53474
rect 221103 53530 221169 53535
rect 221103 53474 221108 53530
rect 221164 53474 221169 53530
rect 221103 53469 221169 53474
rect 212410 53322 212416 53386
rect 212480 53384 212486 53386
rect 216687 53384 216753 53387
rect 212480 53382 216753 53384
rect 212480 53326 216692 53382
rect 216748 53326 216753 53382
rect 212480 53324 216753 53326
rect 212480 53322 212486 53324
rect 216687 53321 216753 53324
rect 211450 53174 211456 53238
rect 211520 53236 211526 53238
rect 217839 53236 217905 53239
rect 211520 53234 217905 53236
rect 211520 53178 217844 53234
rect 217900 53178 217905 53234
rect 211520 53176 217905 53178
rect 211520 53174 211526 53176
rect 217839 53173 217905 53176
rect 223311 52348 223377 52351
rect 637306 52348 637312 52350
rect 223311 52346 637312 52348
rect 223311 52290 223316 52346
rect 223372 52290 637312 52346
rect 223311 52288 637312 52290
rect 223311 52285 223377 52288
rect 637306 52286 637312 52288
rect 637376 52286 637382 52350
rect 221871 52200 221937 52203
rect 637882 52200 637888 52202
rect 221871 52198 637888 52200
rect 221871 52142 221876 52198
rect 221932 52142 637888 52198
rect 221871 52140 637888 52142
rect 221871 52137 221937 52140
rect 637882 52138 637888 52140
rect 637952 52138 637958 52202
rect 211887 52052 211953 52055
rect 637498 52052 637504 52054
rect 211887 52050 637504 52052
rect 211887 51994 211892 52050
rect 211948 51994 637504 52050
rect 211887 51992 637504 51994
rect 211887 51989 211953 51992
rect 637498 51990 637504 51992
rect 637568 51990 637574 52054
rect 212655 51904 212721 51907
rect 637690 51904 637696 51906
rect 212655 51902 637696 51904
rect 212655 51846 212660 51902
rect 212716 51846 637696 51902
rect 212655 51844 637696 51846
rect 212655 51841 212721 51844
rect 637690 51842 637696 51844
rect 637760 51842 637766 51906
rect 223695 51756 223761 51759
rect 637114 51756 637120 51758
rect 223695 51754 637120 51756
rect 223695 51698 223700 51754
rect 223756 51698 637120 51754
rect 223695 51696 637120 51698
rect 223695 51693 223761 51696
rect 637114 51694 637120 51696
rect 637184 51694 637190 51758
rect 222639 51608 222705 51611
rect 636922 51608 636928 51610
rect 222639 51606 636928 51608
rect 222639 51550 222644 51606
rect 222700 51550 636928 51606
rect 222639 51548 636928 51550
rect 222639 51545 222705 51548
rect 636922 51546 636928 51548
rect 636992 51546 636998 51610
rect 145402 51398 145408 51462
rect 145472 51460 145478 51462
rect 243759 51460 243825 51463
rect 145472 51458 243825 51460
rect 145472 51402 243764 51458
rect 243820 51402 243825 51458
rect 145472 51400 243825 51402
rect 145472 51398 145478 51400
rect 243759 51397 243825 51400
rect 145786 51250 145792 51314
rect 145856 51312 145862 51314
rect 237519 51312 237585 51315
rect 145856 51310 237585 51312
rect 145856 51254 237524 51310
rect 237580 51254 237585 51310
rect 145856 51252 237585 51254
rect 145856 51250 145862 51252
rect 237519 51249 237585 51252
rect 145594 51102 145600 51166
rect 145664 51164 145670 51166
rect 237615 51164 237681 51167
rect 145664 51162 237681 51164
rect 145664 51106 237620 51162
rect 237676 51106 237681 51162
rect 145664 51104 237681 51106
rect 145664 51102 145670 51104
rect 237615 51101 237681 51104
rect 145978 50954 145984 51018
rect 146048 51016 146054 51018
rect 236751 51016 236817 51019
rect 146048 51014 236817 51016
rect 146048 50958 236756 51014
rect 236812 50958 236817 51014
rect 146048 50956 236817 50958
rect 146048 50954 146054 50956
rect 236751 50953 236817 50956
rect 467439 49092 467505 49095
rect 471034 49092 471040 49094
rect 467439 49090 471040 49092
rect 467439 49034 467444 49090
rect 467500 49034 471040 49090
rect 467439 49032 471040 49034
rect 467439 49029 467505 49032
rect 471034 49030 471040 49032
rect 471104 49030 471110 49094
rect 168399 48796 168465 48799
rect 242991 48796 243057 48799
rect 168399 48794 243057 48796
rect 168399 48738 168404 48794
rect 168460 48738 242996 48794
rect 243052 48738 243057 48794
rect 168399 48736 243057 48738
rect 168399 48733 168465 48736
rect 242991 48733 243057 48736
rect 171279 48648 171345 48651
rect 242415 48648 242481 48651
rect 171279 48646 242481 48648
rect 171279 48590 171284 48646
rect 171340 48590 242420 48646
rect 242476 48590 242481 48646
rect 171279 48588 242481 48590
rect 171279 48585 171345 48588
rect 242415 48585 242481 48588
rect 174159 48500 174225 48503
rect 243375 48500 243441 48503
rect 174159 48498 243441 48500
rect 174159 48442 174164 48498
rect 174220 48442 243380 48498
rect 243436 48442 243441 48498
rect 174159 48440 243441 48442
rect 174159 48437 174225 48440
rect 243375 48437 243441 48440
rect 202959 48352 203025 48355
rect 241935 48352 242001 48355
rect 202959 48350 242001 48352
rect 202959 48294 202964 48350
rect 203020 48294 241940 48350
rect 241996 48294 242001 48350
rect 202959 48292 242001 48294
rect 202959 48289 203025 48292
rect 241935 48289 242001 48292
rect 165519 48204 165585 48207
rect 242031 48204 242097 48207
rect 165519 48202 242097 48204
rect 165519 48146 165524 48202
rect 165580 48146 242036 48202
rect 242092 48146 242097 48202
rect 165519 48144 242097 48146
rect 165519 48141 165585 48144
rect 242031 48141 242097 48144
rect 213231 45244 213297 45247
rect 411087 45244 411153 45247
rect 213231 45242 411153 45244
rect 213231 45186 213236 45242
rect 213292 45186 411092 45242
rect 411148 45186 411153 45242
rect 213231 45184 411153 45186
rect 213231 45181 213297 45184
rect 411087 45181 411153 45184
rect 214671 45096 214737 45099
rect 521338 45096 521344 45098
rect 214671 45094 521344 45096
rect 214671 45038 214676 45094
rect 214732 45038 521344 45094
rect 214671 45036 521344 45038
rect 214671 45033 214737 45036
rect 521338 45034 521344 45036
rect 521408 45034 521414 45098
rect 215439 44948 215505 44951
rect 527098 44948 527104 44950
rect 215439 44946 527104 44948
rect 215439 44890 215444 44946
rect 215500 44890 527104 44946
rect 215439 44888 527104 44890
rect 215439 44885 215505 44888
rect 527098 44886 527104 44888
rect 527168 44886 527174 44950
rect 212847 44800 212913 44803
rect 416559 44800 416625 44803
rect 212847 44798 416625 44800
rect 212847 44742 212852 44798
rect 212908 44742 416564 44798
rect 416620 44742 416625 44798
rect 212847 44740 416625 44742
rect 212847 44737 212913 44740
rect 416559 44737 416625 44740
rect 521338 43258 521344 43322
rect 521408 43320 521414 43322
rect 521583 43320 521649 43323
rect 521408 43318 521649 43320
rect 521408 43262 521588 43318
rect 521644 43262 521649 43318
rect 521408 43260 521649 43262
rect 521408 43258 521414 43260
rect 521583 43257 521649 43260
rect 527098 43258 527104 43322
rect 527168 43320 527174 43322
rect 529263 43320 529329 43323
rect 527168 43318 529329 43320
rect 527168 43262 529268 43318
rect 529324 43262 529329 43318
rect 527168 43260 529329 43262
rect 527168 43258 527174 43260
rect 529263 43257 529329 43260
rect 297231 43172 297297 43175
rect 302415 43172 302481 43175
rect 297231 43170 302481 43172
rect 297231 43114 297236 43170
rect 297292 43114 302420 43170
rect 302476 43114 302481 43170
rect 297231 43112 302481 43114
rect 297231 43109 297297 43112
rect 302415 43109 302481 43112
rect 351375 43172 351441 43175
rect 357135 43172 357201 43175
rect 351375 43170 357201 43172
rect 351375 43114 351380 43170
rect 351436 43114 357140 43170
rect 357196 43114 357201 43170
rect 351375 43112 357201 43114
rect 351375 43109 351441 43112
rect 357135 43109 357201 43112
rect 455727 43172 455793 43175
rect 463983 43172 464049 43175
rect 455727 43170 464049 43172
rect 455727 43114 455732 43170
rect 455788 43114 463988 43170
rect 464044 43114 464049 43170
rect 455727 43112 464049 43114
rect 455727 43109 455793 43112
rect 463983 43109 464049 43112
rect 567226 42740 622300 42800
rect 282351 42136 282417 42139
rect 306735 42136 306801 42139
rect 282351 42134 306801 42136
rect 282351 42078 282356 42134
rect 282412 42078 306740 42134
rect 306796 42078 306801 42134
rect 282351 42076 306801 42078
rect 282351 42073 282417 42076
rect 306735 42073 306801 42076
rect 362799 42136 362865 42139
rect 364623 42136 364689 42139
rect 471087 42138 471153 42139
rect 362799 42134 364689 42136
rect 362799 42078 362804 42134
rect 362860 42078 364628 42134
rect 364684 42078 364689 42134
rect 362799 42076 364689 42078
rect 362799 42073 362865 42076
rect 364623 42073 364689 42076
rect 471034 42074 471040 42138
rect 471104 42136 471153 42138
rect 471104 42134 471196 42136
rect 471148 42078 471196 42134
rect 471104 42076 471196 42078
rect 471104 42074 471153 42076
rect 471087 42073 471153 42074
rect 187599 41840 187665 41843
rect 189946 41840 189952 41842
rect 187599 41838 189952 41840
rect 187599 41782 187604 41838
rect 187660 41782 189952 41838
rect 187599 41780 189952 41782
rect 187599 41777 187665 41780
rect 189946 41778 189952 41780
rect 190016 41778 190022 41842
rect 194319 41840 194385 41843
rect 211599 41840 211665 41843
rect 194319 41838 334174 41840
rect 194319 41782 194324 41838
rect 194380 41782 334174 41838
rect 194319 41780 334174 41782
rect 194319 41777 194385 41780
rect 211599 41777 211665 41780
rect 241536 41696 245458 41698
rect 241536 41648 255708 41696
rect 189946 40594 189952 40658
rect 190016 40656 190022 40658
rect 211023 40656 211089 40659
rect 190016 40654 211089 40656
rect 190016 40598 211028 40654
rect 211084 40598 211089 40654
rect 190016 40596 211089 40598
rect 190016 40594 190022 40596
rect 211023 40593 211089 40596
rect 142095 40212 142161 40215
rect 141718 40210 142161 40212
rect 141718 40154 142100 40210
rect 142156 40154 142161 40210
rect 241536 40190 245742 41648
rect 141718 40152 142161 40154
rect 141718 39959 141778 40152
rect 142095 40149 142161 40152
rect 241556 40136 245742 40190
rect 251484 40136 255708 41648
rect 334114 41308 334174 41780
rect 333882 41248 334174 41308
rect 374319 41248 374385 41251
rect 333882 40952 333942 41248
rect 334114 41246 334174 41248
rect 354306 41246 374385 41248
rect 354306 41190 374324 41246
rect 374380 41190 374385 41246
rect 354306 41188 374385 41190
rect 334094 40952 334190 40976
rect 333880 40950 334190 40952
rect 333880 40894 334100 40950
rect 334156 40894 334190 40950
rect 333880 40892 334190 40894
rect 334094 40880 334190 40892
rect 344175 40952 344241 40955
rect 354306 40952 354366 41188
rect 374319 41185 374385 41188
rect 344175 40950 354366 40952
rect 344175 40894 344180 40950
rect 344236 40894 354366 40950
rect 344175 40892 354366 40894
rect 344175 40889 344241 40892
rect 374319 40804 374385 40807
rect 374319 40802 388734 40804
rect 374319 40746 374324 40802
rect 374380 40746 388734 40802
rect 374319 40744 388734 40746
rect 374319 40741 374385 40744
rect 388674 40508 388734 40744
rect 397506 40744 409086 40804
rect 397506 40508 397566 40744
rect 409026 40656 409086 40744
rect 469498 40742 469504 40806
rect 469568 40804 469574 40806
rect 469568 40744 489726 40804
rect 469568 40742 469574 40744
rect 443439 40656 443505 40659
rect 409026 40654 443505 40656
rect 409026 40598 443444 40654
rect 443500 40598 443505 40654
rect 409026 40596 443505 40598
rect 443439 40593 443505 40596
rect 453519 40656 453585 40659
rect 469306 40656 469312 40658
rect 453519 40654 469312 40656
rect 453519 40598 453524 40654
rect 453580 40598 469312 40654
rect 453519 40596 469312 40598
rect 453519 40593 453585 40596
rect 469306 40594 469312 40596
rect 469376 40594 469382 40658
rect 489666 40656 489726 40744
rect 529794 40744 538494 40804
rect 529794 40656 529854 40744
rect 489666 40596 509694 40656
rect 388674 40448 397566 40508
rect 509634 40508 509694 40596
rect 509826 40596 529854 40656
rect 509826 40508 509886 40596
rect 509634 40448 509886 40508
rect 538434 40508 538494 40744
rect 567226 40508 567286 42740
rect 569358 42478 583544 42550
rect 569358 42122 573642 42478
rect 538434 40448 567298 40508
rect 567226 40444 567286 40448
rect 443439 40360 443505 40363
rect 453519 40360 453585 40363
rect 443439 40358 453585 40360
rect 443439 40302 443444 40358
rect 443500 40302 453524 40358
rect 453580 40302 453585 40358
rect 443439 40300 453585 40302
rect 443439 40297 443505 40300
rect 453519 40297 453585 40300
rect 569350 40312 573642 42122
rect 579070 40312 583544 42478
rect 622240 40508 622300 42740
rect 623439 40508 623505 40511
rect 622232 40506 623505 40508
rect 622232 40450 623444 40506
rect 623500 40450 623505 40506
rect 622232 40448 623505 40450
rect 623439 40445 623505 40448
rect 241556 40090 255708 40136
rect 241556 39480 245706 40090
rect 251548 39430 255708 40090
rect 569350 40254 583544 40312
rect 569350 39694 573656 40254
rect 579222 39664 583540 40254
<< via3 >>
rect 121358 1022108 121958 1022708
rect 60258 999438 62730 1000238
rect 60276 996948 62750 997622
rect 122816 1021442 123416 1022042
rect 124006 1030258 124606 1030858
rect 121359 996961 121957 997559
rect 122817 997035 123415 997633
rect 125334 1031010 125934 1031610
rect 173268 1022188 173868 1022788
rect 124007 997007 124605 997605
rect 125335 997065 125933 997663
rect 174520 1021450 175120 1022050
rect 173269 997025 173867 997623
rect 174521 996931 175119 997529
rect 176204 1020668 176804 1021268
rect 177460 1020102 178060 1020702
rect 176205 996839 176803 997437
rect 223906 1022192 224506 1022792
rect 177461 996835 178059 997433
rect 225484 1021496 226084 1022096
rect 223907 996797 224505 997395
rect 227324 1020798 227924 1021398
rect 228774 1020014 229374 1020614
rect 274880 1022126 275480 1022726
rect 225485 996707 226083 997305
rect 227325 996883 227923 997481
rect 228775 996981 229373 997579
rect 276374 1021510 276974 1022110
rect 277780 1020716 278380 1021316
rect 278922 1020056 279522 1020656
rect 327774 1022084 328374 1022684
rect 274881 996865 275479 997463
rect 276375 996953 276973 997551
rect 277781 996997 278379 997595
rect 278923 996997 279521 997595
rect 329332 1021334 329932 1021934
rect 298157 997528 298227 997533
rect 298157 997468 298162 997528
rect 298162 997468 298222 997528
rect 298222 997468 298227 997528
rect 298157 997463 298227 997468
rect 327775 996991 328373 997589
rect 330888 1020762 331488 1021362
rect 332436 1020100 333036 1020700
rect 377196 1022158 377796 1022758
rect 378530 1021496 379130 1022096
rect 380080 1020654 380680 1021254
rect 329333 996843 329931 997441
rect 330889 996947 331487 997545
rect 332437 997005 333035 997603
rect 377197 997007 377795 997605
rect 378531 997021 379129 997619
rect 381548 1020080 382148 1020680
rect 410146 1022032 410746 1022632
rect 380081 996997 380679 997595
rect 381549 997011 382147 997609
rect 412148 1021102 412748 1021702
rect 410147 996827 410745 997425
rect 414358 1020556 414958 1021156
rect 415922 1019966 416522 1020566
rect 491650 1021972 492250 1022572
rect 412149 996815 412747 997413
rect 414359 996933 414957 997531
rect 415923 996949 416521 997547
rect 493070 1021282 493670 1021882
rect 494582 1020566 495182 1021166
rect 496096 1019950 496696 1020550
rect 568178 1022164 568778 1022764
rect 491651 996783 492249 997381
rect 493071 996783 493669 997381
rect 494583 996925 495181 997523
rect 496097 996973 496695 997571
rect 570328 1021442 570928 1022042
rect 571834 1020844 572434 1021444
rect 573446 1019996 574046 1020596
rect 568179 996853 568777 997451
rect 570329 996945 570927 997543
rect 571835 996987 572433 997585
rect 573447 996929 574045 997527
rect 298159 996740 298229 996745
rect 298159 996680 298164 996740
rect 298164 996680 298224 996740
rect 298224 996680 298229 996740
rect 298159 996675 298229 996680
rect 476608 996082 476672 996146
rect 580256 996004 585666 997072
rect 476608 995786 476672 995850
rect 30806 984370 31614 988352
rect 41196 984584 42102 988042
rect 42112 968762 42176 968766
rect 42112 968706 42124 968762
rect 42124 968706 42176 968762
rect 42112 968702 42176 968706
rect 675712 967370 675776 967434
rect 41344 967074 41408 967138
rect 676096 965594 676160 965658
rect 42304 965002 42368 965066
rect 674368 965002 674432 965066
rect 675136 964914 675200 964918
rect 675136 964858 675188 964914
rect 675188 964858 675200 964914
rect 675136 964854 675200 964858
rect 40960 963966 41024 964030
rect 41152 963226 41216 963290
rect 674944 962782 675008 962846
rect 40768 962634 40832 962698
rect 674560 962486 674624 962550
rect 676288 962190 676352 962254
rect 40384 962042 40448 962106
rect 42688 961894 42752 961958
rect 674752 961450 674816 961514
rect 675712 961066 675776 961070
rect 675712 961010 675724 961066
rect 675724 961010 675776 961066
rect 675712 961006 675776 961010
rect 42688 960414 42752 960478
rect 675904 960118 675968 960182
rect 41536 959674 41600 959738
rect 41728 959142 41792 959146
rect 41728 959086 41780 959142
rect 41780 959086 41792 959142
rect 41728 959082 41792 959086
rect 675328 959082 675392 959146
rect 40576 958490 40640 958554
rect 41920 957810 41984 957814
rect 41920 957754 41932 957810
rect 41932 957754 41984 957810
rect 41920 957750 41984 957754
rect 675520 957662 675584 957666
rect 675520 957606 675532 957662
rect 675532 957606 675584 957662
rect 675520 957602 675584 957606
rect 673984 955974 674048 956038
rect 42496 955826 42560 955890
rect 677056 953458 677120 953522
rect 676864 953310 676928 953374
rect 8752 952032 9552 952832
rect 50127 952033 50925 952831
rect 16320 950306 17120 951106
rect 51919 950307 52717 951105
rect 671683 949780 672775 950872
rect 699411 949779 700505 950873
rect 7286 948482 8086 949282
rect 53703 948483 54501 949281
rect 666067 948219 667249 949401
rect 709356 948218 710540 949402
rect 17618 946946 18418 947746
rect 55269 946947 56067 947745
rect 662179 946233 663361 947415
rect 700802 946232 701986 947416
rect 42304 945614 42368 945678
rect 42880 945614 42944 945678
rect 659369 944309 660551 945491
rect 708038 944308 709222 945492
rect 40192 941322 40256 941386
rect 42496 941322 42560 941386
rect 41344 940878 41408 940942
rect 41920 939694 41984 939758
rect 40384 939102 40448 939166
rect 42112 938658 42176 938722
rect 40576 937622 40640 937686
rect 674368 937474 674432 937538
rect 41728 937030 41792 937094
rect 675136 936586 675200 936650
rect 42880 936142 42944 936206
rect 674944 935994 675008 936058
rect 41152 935846 41216 935910
rect 675328 935550 675392 935614
rect 41536 935402 41600 935466
rect 40768 934810 40832 934874
rect 676096 934514 676160 934578
rect 40960 934366 41024 934430
rect 674560 933922 674624 933986
rect 676288 933330 676352 933394
rect 673984 932590 674048 932654
rect 675520 932294 675584 932358
rect 674752 931702 674816 931766
rect 677056 931258 677120 931322
rect 676864 930666 676928 930730
rect 43192 916604 44420 922378
rect 671794 912320 674916 917844
rect 674752 876942 674816 877006
rect 673984 876498 674048 876562
rect 675712 875906 675776 875970
rect 674560 875758 674624 875822
rect 675904 875610 675968 875674
rect 674176 874130 674240 874194
rect 674944 873390 675008 873454
rect 674368 872798 674432 872862
rect 675136 869838 675200 869902
rect 675328 864718 675392 864722
rect 675328 864662 675380 864718
rect 675380 864662 675392 864718
rect 675328 864658 675392 864662
rect 44902 828278 45730 841394
rect 8804 825720 9604 826520
rect 50127 825721 50925 826519
rect 16354 824258 17154 825058
rect 51919 824259 52717 825057
rect 7284 822700 8084 823500
rect 53703 822701 54501 823499
rect 17446 821426 18246 822226
rect 55269 821427 56067 822225
rect 668858 819526 670730 832382
rect 40384 815966 40448 816030
rect 40576 813894 40640 813958
rect 40768 811674 40832 811738
rect 40960 802054 41024 802118
rect 41920 800426 41984 800490
rect 42304 800278 42368 800342
rect 42496 799686 42560 799750
rect 42112 797614 42176 797678
rect 42496 797526 42560 797530
rect 42496 797470 42508 797526
rect 42508 797470 42560 797526
rect 42496 797466 42560 797470
rect 42304 797022 42368 797086
rect 41920 792582 41984 792646
rect 40768 791842 40832 791906
rect 40576 791694 40640 791758
rect 42112 791310 42176 791314
rect 42112 791254 42124 791310
rect 42124 791254 42176 791310
rect 42112 791250 42176 791254
rect 41728 791102 41792 791166
rect 42688 791102 42752 791166
rect 675904 787994 675968 788058
rect 675520 787166 675584 787170
rect 675520 787110 675532 787166
rect 675532 787110 675584 787166
rect 675520 787106 675584 787110
rect 676096 786662 676160 786726
rect 676288 784886 676352 784950
rect 675712 784206 675776 784210
rect 675712 784150 675724 784206
rect 675724 784150 675776 784206
rect 675712 784146 675776 784150
rect 8578 782976 9378 783776
rect 50127 782977 50925 783775
rect 16310 781848 17110 782648
rect 51919 781849 52717 782647
rect 676672 781926 676736 781990
rect 7234 780440 8034 781240
rect 53703 780441 54501 781239
rect 676480 780594 676544 780658
rect 17582 778984 18382 779784
rect 55269 778985 56067 779783
rect 677056 777486 677120 777550
rect 677056 776894 677120 776958
rect 677056 776154 677120 776218
rect 676864 774822 676928 774886
rect 40960 773342 41024 773406
rect 677632 773046 677696 773110
rect 40384 772750 40448 772814
rect 40576 772306 40640 772370
rect 671683 770828 672775 771920
rect 699229 770827 700323 771921
rect 666067 769345 667249 770527
rect 709390 769344 710574 770528
rect 41344 768606 41408 768670
rect 662179 767447 663361 768629
rect 700828 767446 702012 768630
rect 659369 765777 660551 766959
rect 707978 765776 709162 766960
rect 42304 765202 42368 765266
rect 677056 760318 677120 760382
rect 40768 760170 40832 760234
rect 42496 760170 42560 760234
rect 677824 759934 677888 759938
rect 677824 759878 677876 759934
rect 677876 759878 677888 759934
rect 677824 759874 677888 759878
rect 674560 759282 674624 759346
rect 43072 759134 43136 759198
rect 675328 758838 675392 758902
rect 674752 758246 674816 758310
rect 41536 757418 41600 757422
rect 41536 757362 41588 757418
rect 41588 757362 41600 757418
rect 41536 757358 41600 757362
rect 674176 757358 674240 757422
rect 675136 757210 675200 757274
rect 41920 757122 41984 757126
rect 41920 757066 41932 757122
rect 41932 757066 41984 757122
rect 41920 757062 41984 757066
rect 42688 757062 42752 757126
rect 676864 756618 676928 756682
rect 676864 756086 676928 756090
rect 676864 756030 676916 756086
rect 676916 756030 676928 756086
rect 676864 756026 676928 756030
rect 673984 755730 674048 755794
rect 674944 755582 675008 755646
rect 42496 754842 42560 754906
rect 674368 754694 674432 754758
rect 677440 754398 677504 754462
rect 677632 753954 677696 754018
rect 677248 753362 677312 753426
rect 677632 753422 677696 753426
rect 677632 753366 677644 753422
rect 677644 753366 677696 753422
rect 677632 753362 677696 753366
rect 677824 752770 677888 752834
rect 42880 751882 42944 751946
rect 41536 751734 41600 751798
rect 42688 751646 42752 751650
rect 42688 751590 42740 751646
rect 42740 751590 42752 751646
rect 42688 751586 42752 751590
rect 41920 751054 41984 751058
rect 41920 750998 41932 751054
rect 41932 750998 41984 751054
rect 41920 750994 41984 750998
rect 42304 750550 42368 750614
rect 43072 750314 43136 750318
rect 43072 750258 43084 750314
rect 43084 750258 43136 750314
rect 43072 750254 43136 750258
rect 42880 749722 42944 749726
rect 42880 749666 42892 749722
rect 42892 749666 42944 749722
rect 42880 749662 42944 749666
rect 41920 748686 41984 748690
rect 41920 748630 41972 748686
rect 41972 748630 41984 748686
rect 41920 748626 41984 748630
rect 41536 747146 41600 747210
rect 40768 746850 40832 746914
rect 41344 746110 41408 746174
rect 676864 744482 676928 744546
rect 677248 744482 677312 744546
rect 676864 744334 676928 744398
rect 677632 744334 677696 744398
rect 674176 743150 674240 743214
rect 673984 742410 674048 742474
rect 674368 741670 674432 741734
rect 8760 739788 9560 740588
rect 50127 739789 50925 740587
rect 676672 740338 676736 740402
rect 675136 740042 675200 740106
rect 16424 738434 17224 739234
rect 51919 738435 52717 739233
rect 674944 739154 675008 739218
rect 674752 738562 674816 738626
rect 7422 737032 8222 737832
rect 53703 737033 54501 737831
rect 17528 735350 18328 736150
rect 55269 735351 56067 736149
rect 675328 734478 675392 734482
rect 675328 734422 675380 734478
rect 675380 734422 675392 734478
rect 675328 734418 675392 734422
rect 40576 729534 40640 729598
rect 41152 729090 41216 729154
rect 677248 728054 677312 728118
rect 41344 727462 41408 727526
rect 671683 726632 672775 727724
rect 699315 726631 700409 727725
rect 676672 725982 676736 726046
rect 677440 725834 677504 725898
rect 40960 725242 41024 725306
rect 42880 725020 42944 725084
rect 666067 724223 667249 725405
rect 709350 724222 710534 725406
rect 662179 722189 663361 723371
rect 700686 722188 701870 723372
rect 41728 721986 41792 722050
rect 659369 720099 660551 721281
rect 708076 720098 709260 721282
rect 41920 715770 41984 715834
rect 43270 715770 43334 715834
rect 41536 715622 41600 715686
rect 42496 715622 42560 715686
rect 676864 715474 676928 715538
rect 677440 714882 677504 714946
rect 677632 714882 677696 714946
rect 43072 714290 43136 714354
rect 676096 714290 676160 714354
rect 677056 714290 677120 714354
rect 40768 714202 40832 714206
rect 40768 714146 40780 714202
rect 40780 714146 40832 714202
rect 40768 714142 40832 714146
rect 41728 714142 41792 714206
rect 41920 713906 41984 713910
rect 41920 713850 41932 713906
rect 41932 713850 41984 713906
rect 41920 713846 41984 713850
rect 42112 713906 42176 713910
rect 42112 713850 42164 713906
rect 42164 713850 42176 713906
rect 42112 713846 42176 713850
rect 675904 713254 675968 713318
rect 676288 712662 676352 712726
rect 676480 712218 676544 712282
rect 41920 711626 41984 711690
rect 42304 711626 42368 711690
rect 677248 711626 677312 711690
rect 41728 711182 41792 711246
rect 41728 711034 41792 711098
rect 42496 711034 42560 711098
rect 675520 711034 675584 711098
rect 42304 710886 42368 710950
rect 675712 710590 675776 710654
rect 42112 709910 42176 709914
rect 42112 709854 42164 709910
rect 42164 709854 42176 709910
rect 42112 709850 42176 709854
rect 41536 707334 41600 707398
rect 40768 707186 40832 707250
rect 42688 706890 42752 706954
rect 43268 706890 43332 706954
rect 42880 706446 42944 706510
rect 41344 705114 41408 705178
rect 42496 704522 42560 704586
rect 41728 704138 41792 704142
rect 41728 704082 41780 704138
rect 41780 704082 41792 704138
rect 41728 704078 41792 704082
rect 40960 703338 41024 703402
rect 43072 700526 43136 700590
rect 675520 697922 675584 697926
rect 675520 697866 675532 697922
rect 675532 697866 675584 697922
rect 675520 697862 675584 697866
rect 676672 697270 676736 697334
rect 8706 696342 9506 697142
rect 50127 696343 50925 697141
rect 675328 696974 675392 697038
rect 676288 696974 676352 697038
rect 675328 696886 675392 696890
rect 675328 696830 675380 696886
rect 675380 696830 675392 696886
rect 675328 696826 675392 696830
rect 16332 695068 17132 695868
rect 51919 695069 52717 695867
rect 675712 694814 675776 694818
rect 675712 694758 675724 694814
rect 675724 694758 675776 694814
rect 675712 694754 675776 694758
rect 7212 693954 8012 694754
rect 53703 693955 54501 694753
rect 674560 694310 674624 694374
rect 17798 692284 18598 693084
rect 55269 692285 56067 693083
rect 676480 691942 676544 692006
rect 675904 689130 675968 689194
rect 676096 688242 676160 688306
rect 40576 686910 40640 686974
rect 42112 686466 42176 686530
rect 40384 685874 40448 685938
rect 41152 685874 41216 685938
rect 40576 684246 40640 684310
rect 43072 683062 43136 683126
rect 40768 682026 40832 682090
rect 671683 681224 672775 682316
rect 699121 681223 700215 682317
rect 666067 679621 667249 680803
rect 709418 679620 710602 680804
rect 41536 678178 41600 678242
rect 662179 677785 663361 678967
rect 700498 677784 701682 678968
rect 659369 676061 660551 677243
rect 708330 676060 709514 677244
rect 41728 675574 41792 675578
rect 41728 675518 41740 675574
rect 41740 675518 41792 675574
rect 41728 675514 41792 675518
rect 41344 670926 41408 670990
rect 42304 670926 42368 670990
rect 42496 670630 42560 670694
rect 43072 670690 43136 670694
rect 43072 670634 43084 670690
rect 43084 670634 43136 670690
rect 43072 670630 43136 670634
rect 41920 670482 41984 670546
rect 677248 670186 677312 670250
rect 677440 670186 677504 670250
rect 677056 669594 677120 669658
rect 674368 668854 674432 668918
rect 674176 667744 674240 667808
rect 675136 667522 675200 667586
rect 673984 665598 674048 665662
rect 41536 665302 41600 665366
rect 674944 665302 675008 665366
rect 674752 664858 674816 664922
rect 42304 664710 42368 664774
rect 41344 663970 41408 664034
rect 676288 663674 676352 663738
rect 42496 662786 42560 662850
rect 40768 662342 40832 662406
rect 41728 662194 41792 662258
rect 42688 662194 42752 662258
rect 41920 661070 41984 661074
rect 41920 661014 41932 661070
rect 41932 661014 41984 661070
rect 41920 661010 41984 661014
rect 40576 660862 40640 660926
rect 8566 653016 9366 653816
rect 50127 653017 50925 653815
rect 676480 653610 676544 653674
rect 16290 651820 17090 652620
rect 51919 651821 52717 652619
rect 674752 652574 674816 652638
rect 674176 652130 674240 652194
rect 7184 650716 7984 651516
rect 53703 650717 54501 651515
rect 675136 651390 675200 651454
rect 17672 649150 18472 649950
rect 55269 649151 56067 649949
rect 673984 649762 674048 649826
rect 674752 649762 674816 649826
rect 674752 649614 674816 649678
rect 674368 648874 674432 648938
rect 42112 647098 42176 647162
rect 40384 646950 40448 647014
rect 676288 645322 676352 645386
rect 40960 641030 41024 641094
rect 673984 640290 674048 640354
rect 40576 638810 40640 638874
rect 676480 638514 676544 638578
rect 671683 635880 672775 636972
rect 699309 635879 700403 636973
rect 666067 634303 667249 635485
rect 709374 634302 710558 635486
rect 662179 632443 663361 633625
rect 700650 632442 701834 633626
rect 673792 630818 673856 630882
rect 674944 630818 675008 630882
rect 674368 630670 674432 630734
rect 675136 630670 675200 630734
rect 659369 628833 660551 630015
rect 708128 628832 709312 630016
rect 41536 627770 41600 627774
rect 41536 627714 41548 627770
rect 41548 627714 41600 627770
rect 41536 627710 41600 627714
rect 42112 627622 42176 627626
rect 42112 627566 42124 627622
rect 42124 627566 42176 627622
rect 42112 627562 42176 627566
rect 42304 627414 42368 627478
rect 42496 626970 42560 627034
rect 677248 626378 677312 626442
rect 677440 625157 677504 625221
rect 677056 624602 677120 624666
rect 42496 624514 42560 624518
rect 42496 624458 42508 624514
rect 42508 624458 42560 624514
rect 42496 624454 42560 624458
rect 675328 624158 675392 624222
rect 675520 623122 675584 623186
rect 675712 622530 675776 622594
rect 42304 622086 42368 622150
rect 42112 621494 42176 621558
rect 676672 620902 676736 620966
rect 674944 620814 675008 620818
rect 674944 620758 674996 620814
rect 674996 620758 675008 620814
rect 674944 620754 675008 620758
rect 674560 620310 674624 620374
rect 674560 619866 674624 619930
rect 676096 619866 676160 619930
rect 41536 619570 41600 619634
rect 675904 618682 675968 618746
rect 41728 618238 41792 618302
rect 42304 618238 42368 618302
rect 41920 617706 41984 617710
rect 41920 617650 41972 617706
rect 41972 617650 41984 617706
rect 41920 617646 41984 617650
rect 42496 617646 42560 617710
rect 40960 617202 41024 617266
rect 40576 616462 40640 616526
rect 674752 613798 674816 613862
rect 676096 613798 676160 613862
rect 673984 613650 674048 613714
rect 675520 613650 675584 613714
rect 8736 609926 9536 610726
rect 50127 609927 50925 610725
rect 16282 608646 17082 609446
rect 51919 608647 52717 609445
rect 7318 607092 8118 607892
rect 53703 607093 54501 607891
rect 673984 607730 674048 607794
rect 675136 607138 675200 607202
rect 675328 606546 675392 606610
rect 675904 606546 675968 606610
rect 675328 606398 675392 606462
rect 17654 605356 18454 606156
rect 55269 605357 56067 606155
rect 42304 605066 42368 605130
rect 42496 605066 42560 605130
rect 42304 604918 42368 604982
rect 42496 604918 42560 604982
rect 674368 604770 674432 604834
rect 675520 600478 675584 600542
rect 676672 600478 676736 600542
rect 42880 599220 42944 599284
rect 40384 597814 40448 597878
rect 40576 595594 40640 595658
rect 676096 595446 676160 595510
rect 676096 595298 676160 595362
rect 674752 594706 674816 594770
rect 675904 594706 675968 594770
rect 675904 593374 675968 593438
rect 42112 592930 42176 592994
rect 42496 591894 42560 591958
rect 671683 591550 672775 592642
rect 699395 591549 700489 592643
rect 30592 590710 30656 590774
rect 674944 590858 675008 590922
rect 676672 590858 676736 590922
rect 674560 590562 674624 590626
rect 675712 590414 675776 590478
rect 30592 590266 30656 590330
rect 674560 590266 674624 590330
rect 675136 590266 675200 590330
rect 675520 590326 675584 590330
rect 675520 590270 675532 590326
rect 675532 590270 675584 590326
rect 675520 590266 675584 590270
rect 674752 590118 674816 590182
rect 675136 589970 675200 590034
rect 676480 589970 676544 590034
rect 676480 589822 676544 589886
rect 676864 589822 676928 589886
rect 41920 588934 41984 588998
rect 42688 588934 42752 588998
rect 666067 587955 667249 589137
rect 709314 587954 710498 589138
rect 662179 586173 663361 587355
rect 700810 586172 701994 587356
rect 42304 584198 42368 584262
rect 659369 583903 660551 585085
rect 708068 583902 709252 585086
rect 42304 581238 42368 581302
rect 41728 579166 41792 579230
rect 41920 579166 41984 579230
rect 677248 579462 677312 579526
rect 41536 579018 41600 579082
rect 42112 579018 42176 579082
rect 42304 579018 42368 579082
rect 677056 579018 677120 579082
rect 41920 578870 41984 578934
rect 42688 578870 42752 578934
rect 676672 578870 676736 578934
rect 676480 578426 676544 578490
rect 674944 577834 675008 577898
rect 675520 577242 675584 577306
rect 42880 577006 42944 577010
rect 42880 576950 42932 577006
rect 42932 576950 42944 577006
rect 42880 576946 42944 576950
rect 676288 576798 676352 576862
rect 675136 576206 675200 576270
rect 41920 575970 41984 575974
rect 41920 575914 41972 575970
rect 41972 575914 41984 575970
rect 41920 575910 41984 575914
rect 674176 575318 674240 575382
rect 674752 575170 674816 575234
rect 42112 574638 42176 574642
rect 42112 574582 42124 574638
rect 42124 574582 42176 574638
rect 42112 574578 42176 574582
rect 41728 574490 41792 574494
rect 41728 574434 41780 574490
rect 41780 574434 41792 574490
rect 41728 574430 41792 574434
rect 40384 573838 40448 573902
rect 40576 573098 40640 573162
rect 8620 566846 9420 567646
rect 50127 566847 50925 567645
rect 16256 565744 17056 566544
rect 51919 565745 52717 566543
rect 7348 564474 8148 565274
rect 53703 564475 54501 565273
rect 17620 563022 18420 563822
rect 55269 563023 56067 563821
rect 674944 562442 675008 562506
rect 674176 561998 674240 562062
rect 41920 561554 41984 561618
rect 42496 561554 42560 561618
rect 675136 561406 675200 561470
rect 40192 560518 40256 560582
rect 674752 558890 674816 558954
rect 40192 556818 40256 556882
rect 40384 554598 40448 554662
rect 676864 554450 676928 554514
rect 40576 552378 40640 552442
rect 671683 546058 672775 547150
rect 699205 546057 700299 547151
rect 666067 544313 667249 545495
rect 709418 544312 710602 545496
rect 662179 542719 663361 543901
rect 700596 542718 701780 543902
rect 42880 541634 42944 541638
rect 42880 541578 42932 541634
rect 42932 541578 42944 541634
rect 42880 541574 42944 541578
rect 42688 541278 42752 541342
rect 42304 541130 42368 541194
rect 41920 541042 41984 541046
rect 41920 540986 41932 541042
rect 41932 540986 41984 541042
rect 41920 540982 41984 540986
rect 659369 540699 660551 541881
rect 707930 540698 709114 541882
rect 41920 536838 41984 536902
rect 42880 535654 42944 535718
rect 677248 535062 677312 535126
rect 677056 534470 677120 534534
rect 42688 534322 42752 534386
rect 675328 533878 675392 533942
rect 676096 533434 676160 533498
rect 42304 533346 42368 533350
rect 42304 533290 42356 533346
rect 42356 533290 42368 533346
rect 42304 533286 42368 533290
rect 42496 532694 42560 532758
rect 673984 532546 674048 532610
rect 674368 531954 674432 532018
rect 41920 531806 41984 531870
rect 675712 531806 675776 531870
rect 41728 531718 41792 531722
rect 41728 531662 41780 531718
rect 41780 531662 41792 531718
rect 41728 531658 41792 531662
rect 40576 531214 40640 531278
rect 675904 531214 675968 531278
rect 40384 530622 40448 530686
rect 674560 530622 674624 530686
rect 669372 518422 670344 518424
rect 669368 514106 670344 518422
rect 669372 508462 670344 514106
rect 669372 504232 670350 508462
rect 671683 501996 672775 503088
rect 699153 501995 700247 503089
rect 666067 500091 667249 501273
rect 709152 500090 710336 501274
rect 662179 498231 663361 499413
rect 700596 498230 701780 499414
rect 45974 483786 46716 497304
rect 659369 496317 660551 497499
rect 708036 496316 709220 497500
rect 677824 490958 677888 491022
rect 677632 490514 677696 490578
rect 675136 489922 675200 489986
rect 677440 489922 677504 489986
rect 674944 488886 675008 488950
rect 674176 486370 674240 486434
rect 674752 486074 674816 486138
rect 676864 483410 676928 483474
rect 665144 460522 668046 473848
rect 47166 441662 49188 454744
rect 8774 439190 9574 439990
rect 50127 439191 50925 439989
rect 16250 437824 17050 438624
rect 51919 437825 52717 438623
rect 7356 436296 8156 437096
rect 53703 436297 54501 437095
rect 17690 434948 18490 435748
rect 55269 434949 56067 435747
rect 40384 429242 40448 429306
rect 40576 428650 40640 428714
rect 40960 428058 41024 428122
rect 40768 427022 40832 427086
rect 41344 426430 41408 426494
rect 41536 425986 41600 426050
rect 41152 424802 41216 424866
rect 42112 424358 42176 424422
rect 42304 423914 42368 423978
rect 671683 413856 672775 414948
rect 699209 413855 700303 414949
rect 666067 411817 667249 412999
rect 709366 411816 710550 413000
rect 662179 410033 663361 411215
rect 700720 410032 701904 411216
rect 659369 408249 660551 409431
rect 708100 408248 709284 409432
rect 41536 406006 41600 406070
rect 41920 405178 41984 405182
rect 41920 405122 41932 405178
rect 41932 405122 41984 405178
rect 41920 405118 41984 405122
rect 41728 404438 41792 404442
rect 41728 404382 41780 404438
rect 41780 404382 41792 404438
rect 41728 404378 41792 404382
rect 677824 403934 677888 403998
rect 42304 403046 42368 403110
rect 677632 402750 677696 402814
rect 42112 402662 42176 402666
rect 42112 402606 42164 402662
rect 42164 402606 42176 402662
rect 42112 402602 42176 402606
rect 677440 402158 677504 402222
rect 41344 401862 41408 401926
rect 674560 400530 674624 400594
rect 40960 400086 41024 400150
rect 41152 399494 41216 399558
rect 674368 399198 674432 399262
rect 40768 398754 40832 398818
rect 674176 398754 674240 398818
rect 8624 396038 9424 396838
rect 50127 396039 50925 396837
rect 16362 394606 17162 395406
rect 51919 394607 52717 395405
rect 7322 393086 8122 393886
rect 53703 393087 54501 393885
rect 17528 391566 18328 392366
rect 55269 391567 56067 392365
rect 40384 386026 40448 386090
rect 40576 386026 40640 386090
rect 40960 384842 41024 384906
rect 40768 383806 40832 383870
rect 41344 383214 41408 383278
rect 41536 382770 41600 382834
rect 41152 381586 41216 381650
rect 674368 378774 674432 378838
rect 42112 375074 42176 375138
rect 675328 374482 675392 374546
rect 677056 374334 677120 374398
rect 675520 374038 675584 374102
rect 674560 373890 674624 373954
rect 677056 373002 677120 373066
rect 42304 372854 42368 372918
rect 674176 371966 674240 372030
rect 671683 368888 672775 369980
rect 699307 368887 700401 369981
rect 666067 366733 667249 367915
rect 709268 366732 710452 367916
rect 662179 364879 663361 366061
rect 700568 364878 701752 366062
rect 659369 363129 660551 364311
rect 707888 363128 709072 364312
rect 41536 362790 41600 362854
rect 41920 360866 41984 360930
rect 42496 360866 42560 360930
rect 41728 360570 41792 360634
rect 42688 360570 42752 360634
rect 42304 359830 42368 359894
rect 42112 359446 42176 359450
rect 42112 359390 42124 359446
rect 42124 359390 42176 359446
rect 42112 359386 42176 359390
rect 41344 358646 41408 358710
rect 676864 357610 676928 357674
rect 677056 357610 677120 357674
rect 40960 356870 41024 356934
rect 41152 356426 41216 356490
rect 677440 356426 677504 356490
rect 673984 355686 674048 355750
rect 40768 355538 40832 355602
rect 8636 352300 9436 353100
rect 50127 352301 50925 353099
rect 16348 351238 17148 352038
rect 51919 351239 52717 352037
rect 7236 350088 8036 350888
rect 53703 350089 54501 350887
rect 17548 348586 18348 349386
rect 55269 348587 56067 349385
rect 676480 345474 676544 345538
rect 676672 345326 676736 345390
rect 40384 342958 40448 343022
rect 40576 342810 40640 342874
rect 40768 341774 40832 341838
rect 40960 340590 41024 340654
rect 41344 340146 41408 340210
rect 41536 339554 41600 339618
rect 42496 338962 42560 339026
rect 42880 338962 42944 339026
rect 41152 338518 41216 338582
rect 43072 338222 43136 338286
rect 675328 335026 675392 335030
rect 675328 334970 675340 335026
rect 675340 334970 675392 335026
rect 675328 334966 675392 334970
rect 675520 333842 675584 333846
rect 675520 333786 675532 333842
rect 675532 333786 675584 333842
rect 675520 333782 675584 333786
rect 32020 330486 32604 331648
rect 44906 330504 45450 331636
rect 676480 330526 676544 330590
rect 42304 329786 42368 329850
rect 675328 329490 675392 329554
rect 673984 328306 674048 328370
rect 676672 326826 676736 326890
rect 42496 326530 42560 326594
rect 671683 323144 672775 324236
rect 699295 323143 700389 324237
rect 41920 322534 41984 322598
rect 42880 322534 42944 322598
rect 666067 321423 667249 322605
rect 709502 321422 710686 322606
rect 42496 320966 42560 320970
rect 42496 320910 42508 320966
rect 42508 320910 42560 320966
rect 42496 320906 42560 320910
rect 41536 319722 41600 319786
rect 662179 319289 663361 320471
rect 700628 319288 701812 320472
rect 41920 318746 41984 318750
rect 41920 318690 41972 318746
rect 41972 318690 41984 318746
rect 41920 318686 41984 318690
rect 41920 317858 41984 317862
rect 41920 317802 41972 317858
rect 41972 317802 41984 317858
rect 41920 317798 41984 317802
rect 42112 317058 42176 317122
rect 43072 317058 43136 317122
rect 659369 317003 660551 318185
rect 707920 317002 709104 318186
rect 42304 316614 42368 316678
rect 42112 316082 42176 316086
rect 42112 316026 42124 316082
rect 42124 316026 42176 316082
rect 42112 316022 42176 316026
rect 41344 315430 41408 315494
rect 40768 313654 40832 313718
rect 676864 313654 676928 313718
rect 41152 313210 41216 313274
rect 677248 312470 677312 312534
rect 40960 312322 41024 312386
rect 677056 312026 677120 312090
rect 677440 312026 677504 312090
rect 676864 311434 676928 311498
rect 673984 310694 674048 310758
rect 8738 309136 9538 309936
rect 50127 309137 50925 309935
rect 16328 307998 17128 308798
rect 51919 307999 52717 308797
rect 7378 306336 8178 307136
rect 53703 306337 54501 307135
rect 17732 304848 18532 305648
rect 55269 304849 56067 305647
rect 40384 299742 40448 299806
rect 40576 299594 40640 299658
rect 42304 299594 42368 299658
rect 675904 299446 675968 299510
rect 676672 299298 676736 299362
rect 40768 298558 40832 298622
rect 40960 297374 41024 297438
rect 41344 296930 41408 296994
rect 41536 296486 41600 296550
rect 41152 295302 41216 295366
rect 42112 294858 42176 294922
rect 42688 293378 42752 293442
rect 675328 290034 675392 290038
rect 675328 289978 675340 290034
rect 675340 289978 675392 290034
rect 675328 289974 675392 289978
rect 675520 289590 675584 289594
rect 675520 289534 675532 289590
rect 675532 289534 675584 289590
rect 675520 289530 675584 289534
rect 36346 286660 36976 287744
rect 46158 286664 46718 287742
rect 41920 285534 41984 285598
rect 42496 285534 42560 285598
rect 41728 285090 41792 285154
rect 674560 284942 674624 285006
rect 674368 284794 674432 284858
rect 675904 284794 675968 284858
rect 673984 283610 674048 283674
rect 676672 281834 676736 281898
rect 671683 278476 672775 279568
rect 699329 278475 700423 279569
rect 42688 277986 42752 278050
rect 666067 276817 667249 277999
rect 709390 276816 710574 278000
rect 41536 276506 41600 276570
rect 674560 276358 674624 276422
rect 41920 275530 41984 275534
rect 41920 275474 41972 275530
rect 41972 275474 41984 275530
rect 41920 275470 41984 275474
rect 42496 274730 42560 274794
rect 662179 274045 663361 275227
rect 700624 274044 701808 275228
rect 41728 273606 41792 273610
rect 41728 273550 41780 273606
rect 41780 273550 41792 273606
rect 41728 273546 41792 273550
rect 374464 273546 374528 273610
rect 409408 273398 409472 273462
rect 384064 273250 384128 273314
rect 409792 273250 409856 273314
rect 42112 273014 42176 273018
rect 42112 272958 42124 273014
rect 42124 272958 42176 273014
rect 42112 272954 42176 272958
rect 374464 272954 374528 273018
rect 408256 272954 408320 273018
rect 135232 272510 135296 272574
rect 410560 272806 410624 272870
rect 409600 272658 409664 272722
rect 41344 272214 41408 272278
rect 378304 272066 378368 272130
rect 407872 271770 407936 271834
rect 406144 271622 406208 271686
rect 407488 271474 407552 271538
rect 410176 272214 410240 272278
rect 410944 271918 411008 271982
rect 659369 271927 660551 273109
rect 707924 271926 709108 273110
rect 411136 271622 411200 271686
rect 411328 271474 411392 271538
rect 377920 271178 377984 271242
rect 406528 271178 406592 271242
rect 409216 271178 409280 271242
rect 406720 271030 406784 271094
rect 348544 270882 348608 270946
rect 391744 270882 391808 270946
rect 406912 270882 406976 270946
rect 135232 270734 135296 270798
rect 407680 270734 407744 270798
rect 40768 270586 40832 270650
rect 41920 270586 41984 270650
rect 42880 270586 42944 270650
rect 369472 270646 369536 270650
rect 369472 270590 369484 270646
rect 369484 270590 369536 270646
rect 369472 270586 369536 270590
rect 369856 270646 369920 270650
rect 369856 270590 369868 270646
rect 369868 270590 369920 270646
rect 369856 270586 369920 270590
rect 41152 269994 41216 270058
rect 40960 269106 41024 269170
rect 290752 269106 290816 269170
rect 316672 269106 316736 269170
rect 347200 269166 347264 269170
rect 347200 269110 347252 269166
rect 347252 269110 347264 269166
rect 347200 269106 347264 269110
rect 347584 269166 347648 269170
rect 347584 269110 347596 269166
rect 347596 269110 347648 269166
rect 347584 269106 347648 269110
rect 677248 268662 677312 268726
rect 290752 268366 290816 268430
rect 348352 268366 348416 268430
rect 377536 268366 377600 268430
rect 405952 268366 406016 268430
rect 292288 268070 292352 268134
rect 312448 268070 312512 268134
rect 316672 268070 316736 268134
rect 336448 268130 336512 268134
rect 336448 268074 336460 268130
rect 336460 268074 336512 268130
rect 336448 268070 336512 268074
rect 267904 267774 267968 267838
rect 307840 267774 307904 267838
rect 308416 267774 308480 267838
rect 312448 267626 312512 267690
rect 376576 267774 376640 267838
rect 383680 267774 383744 267838
rect 336448 267626 336512 267690
rect 347200 267626 347264 267690
rect 347584 267626 347648 267690
rect 376960 267626 377024 267690
rect 405376 267922 405440 267986
rect 405760 267922 405824 267986
rect 406336 267922 406400 267986
rect 677440 267626 677504 267690
rect 8584 266560 9384 267360
rect 50127 266561 50925 267359
rect 676864 267034 676928 267098
rect 677056 267034 677120 267098
rect 16354 265112 17154 265912
rect 51919 265113 52717 265911
rect 407098 264940 407168 264945
rect 407098 264880 407103 264940
rect 407103 264880 407163 264940
rect 407163 264880 407168 264940
rect 407098 264875 407168 264880
rect 407296 264814 407360 264878
rect 408109 264933 408179 264938
rect 408109 264873 408114 264933
rect 408114 264873 408174 264933
rect 408174 264873 408179 264933
rect 408109 264868 408179 264873
rect 410368 264814 410432 264878
rect 409984 264666 410048 264730
rect 410752 264666 410816 264730
rect 411520 264666 411584 264730
rect 410560 264518 410624 264582
rect 674176 264074 674240 264138
rect 7374 263216 8174 264016
rect 53703 263217 54501 264015
rect 17562 261322 18362 262122
rect 55269 261323 56067 262121
rect 673984 260818 674048 260882
rect 40384 256970 40448 257034
rect 206998 256926 209004 259496
rect 211282 256878 211434 259536
rect 412836 256884 412992 259516
rect 416548 256980 423896 259382
rect 42304 255934 42368 255998
rect 40576 255342 40640 255406
rect 40384 254158 40448 254222
rect 40768 253714 40832 253778
rect 41152 253270 41216 253334
rect 206478 253276 208996 256326
rect 211020 253276 211164 256362
rect 413114 253274 413240 256348
rect 416506 253412 424074 256270
rect 40960 252086 41024 252150
rect 41344 251642 41408 251706
rect 641918 249864 655400 252222
rect 685012 251802 685600 254778
rect 675904 251642 675968 251706
rect 675712 251494 675776 251558
rect 410752 247794 410816 247858
rect 411520 247794 411584 247858
rect 407488 247646 407552 247710
rect 408448 247646 408512 247710
rect 408640 247646 408704 247710
rect 411136 247646 411200 247710
rect 407296 247498 407360 247562
rect 409792 247498 409856 247562
rect 410368 247350 410432 247414
rect 411328 247350 411392 247414
rect 207232 246906 207296 246970
rect 42880 246758 42944 246822
rect 407104 247202 407168 247266
rect 407296 247202 407360 247266
rect 409984 247202 410048 247266
rect 410176 247202 410240 247266
rect 405760 247054 405824 247118
rect 410560 247054 410624 247118
rect 410752 247054 410816 247118
rect 406720 246906 406784 246970
rect 406520 246758 406598 246834
rect 407296 246906 407360 246970
rect 408832 246906 408896 246970
rect 410944 246906 411008 246970
rect 406912 246758 406976 246822
rect 407488 246758 407552 246822
rect 408064 246818 408128 246822
rect 408064 246762 408116 246818
rect 408116 246762 408128 246818
rect 408064 246758 408128 246762
rect 408448 246758 408512 246822
rect 408832 246818 408896 246822
rect 408832 246762 408844 246818
rect 408844 246762 408896 246818
rect 408832 246758 408896 246762
rect 409216 246818 409280 246822
rect 409216 246762 409228 246818
rect 409228 246762 409280 246818
rect 409216 246758 409280 246762
rect 409600 246758 409664 246822
rect 674560 246758 674624 246822
rect 207232 246166 207296 246230
rect 674560 245870 674624 245934
rect 41536 244982 41600 245046
rect 42880 244982 42944 245046
rect 41728 244834 41792 244898
rect 674368 244686 674432 244750
rect 675328 244746 675392 244750
rect 675328 244690 675380 244746
rect 675380 244690 675392 244746
rect 675328 244686 675392 244690
rect 41920 243798 41984 243862
rect 674368 243798 674432 243862
rect 210304 243650 210368 243714
rect 211072 243710 211136 243714
rect 211072 243654 211084 243710
rect 211084 243654 211136 243710
rect 211072 243650 211136 243654
rect 405568 243502 405632 243566
rect 405952 243502 406016 243566
rect 408256 243502 408320 243566
rect 674176 243502 674240 243566
rect 406336 243354 406400 243418
rect 210688 243058 210752 243122
rect 407680 243206 407744 243270
rect 406144 242910 406208 242974
rect 328768 242762 328832 242826
rect 328384 242318 328448 242382
rect 212032 242170 212096 242234
rect 145408 242022 145472 242086
rect 673984 242022 674048 242086
rect 675520 238914 675584 238978
rect 675712 238678 675776 238682
rect 675712 238622 675764 238678
rect 675764 238622 675776 238678
rect 675712 238618 675776 238622
rect 241792 238470 241856 238534
rect 42304 238322 42368 238386
rect 241792 238174 241856 238238
rect 211456 237730 211520 237794
rect 676480 237730 676544 237794
rect 677056 237582 677120 237646
rect 675904 236842 675968 236906
rect 239104 236694 239168 236758
rect 239104 236250 239168 236314
rect 676480 236250 676544 236314
rect 676864 236250 676928 236314
rect 211648 234622 211712 234686
rect 42304 234030 42368 234094
rect 210304 233882 210368 233946
rect 636928 233882 636992 233946
rect 212032 233734 212096 233798
rect 212992 233734 213056 233798
rect 637696 233734 637760 233798
rect 210688 233586 210752 233650
rect 212608 233646 212672 233650
rect 212608 233590 212620 233646
rect 212620 233590 212672 233646
rect 211072 233438 211136 233502
rect 212224 233438 212288 233502
rect 212608 233586 212672 233590
rect 637120 233646 637184 233650
rect 637120 233590 637172 233646
rect 637172 233590 637184 233646
rect 637120 233586 637184 233590
rect 637504 233586 637568 233650
rect 212800 233438 212864 233502
rect 637312 233438 637376 233502
rect 637888 233438 637952 233502
rect 41152 233290 41216 233354
rect 210688 233290 210752 233354
rect 671683 232544 672775 233636
rect 708937 232543 710031 233637
rect 41536 231662 41600 231726
rect 41920 231130 41984 231134
rect 41920 231074 41972 231130
rect 41972 231074 41984 231130
rect 41920 231070 41984 231074
rect 41728 230390 41792 230394
rect 41728 230334 41780 230390
rect 41780 230334 41792 230390
rect 41728 230330 41792 230334
rect 666067 230253 667249 231435
rect 698422 230252 699606 231436
rect 41344 229738 41408 229802
rect 40768 228998 40832 229062
rect 662179 227873 663361 229055
rect 707214 227816 708398 229000
rect 40576 227222 40640 227286
rect 40960 226630 41024 226694
rect 40384 225890 40448 225954
rect 641093 225131 643327 227365
rect 699854 226130 701038 227314
rect 8730 223084 9530 223884
rect 43691 223085 44489 223883
rect 677440 223522 677504 223586
rect 16292 221940 17092 222740
rect 46937 221941 47735 222739
rect 677056 222486 677120 222550
rect 677440 222338 677504 222402
rect 7364 220730 8164 221530
rect 48719 220731 49517 221529
rect 676864 221302 676928 221366
rect 677248 221302 677312 221366
rect 17702 219456 18502 220256
rect 50603 219457 51401 220255
rect 674176 220488 674240 220552
rect 145600 218934 145664 218998
rect 145792 216418 145856 216482
rect 145984 214494 146048 214558
rect 40576 212126 40640 212190
rect 40384 211090 40448 211154
rect 40960 210498 41024 210562
rect 41536 209906 41600 209970
rect 40768 208870 40832 208934
rect 41152 208278 41216 208342
rect 41344 207834 41408 207898
rect 675712 207686 675776 207750
rect 676672 207538 676736 207602
rect 676480 207390 676544 207454
rect 211072 205022 211136 205086
rect 675328 200050 675392 200054
rect 675328 199994 675380 200050
rect 675380 199994 675392 200050
rect 675328 199990 675392 199994
rect 675520 199606 675584 199610
rect 675520 199550 675532 199606
rect 675532 199550 675584 199606
rect 675520 199546 675584 199550
rect 675712 198422 675776 198426
rect 675712 198366 675764 198422
rect 675764 198366 675776 198422
rect 675712 198362 675776 198366
rect 42112 197622 42176 197686
rect 676480 195254 676544 195318
rect 210880 194958 210944 195022
rect 211072 194958 211136 195022
rect 210880 194514 210944 194578
rect 211072 194070 211136 194134
rect 674176 193478 674240 193542
rect 675328 193034 675392 193098
rect 676672 191554 676736 191618
rect 42112 191022 42176 191026
rect 42112 190966 42164 191022
rect 42164 190966 42176 191022
rect 42112 190962 42176 190966
rect 41536 190074 41600 190138
rect 210112 190074 210176 190138
rect 211072 190074 211136 190138
rect 41728 189098 41792 189102
rect 41728 189042 41780 189098
rect 41780 189042 41792 189098
rect 41728 189038 41792 189042
rect 671683 188410 672775 189502
rect 708777 188409 709871 189503
rect 41920 188358 41984 188362
rect 41920 188302 41972 188358
rect 41972 188302 41984 188358
rect 41920 188298 41984 188302
rect 41344 187114 41408 187178
rect 41152 186374 41216 186438
rect 666067 186251 667249 187433
rect 698514 186250 699698 187434
rect 40960 185782 41024 185846
rect 40576 184154 40640 184218
rect 645421 183647 647655 185881
rect 700656 183900 701840 185084
rect 40768 183562 40832 183626
rect 40384 182822 40448 182886
rect 641093 180957 643327 183191
rect 706104 181210 707288 182394
rect 677440 178382 677504 178446
rect 677056 177346 677120 177410
rect 677440 177346 677504 177410
rect 677248 176310 677312 176374
rect 209920 175718 209984 175782
rect 211072 175718 211136 175782
rect 210688 174386 210752 174450
rect 211072 174386 211136 174450
rect 210304 173942 210368 174006
rect 210880 173942 210944 174006
rect 209920 171278 209984 171342
rect 211072 171278 211136 171342
rect 673984 171130 674048 171194
rect 210112 170538 210176 170602
rect 211072 170538 211136 170602
rect 211072 164174 211136 164238
rect 675712 161510 675776 161574
rect 676672 161362 676736 161426
rect 675328 155206 675392 155210
rect 675328 155150 675340 155206
rect 675340 155150 675392 155206
rect 675328 155146 675392 155150
rect 675520 154466 675584 154470
rect 675520 154410 675532 154466
rect 675532 154410 675584 154466
rect 675520 154406 675584 154410
rect 210112 151890 210176 151954
rect 210880 151890 210944 151954
rect 673984 150262 674048 150326
rect 675712 148546 675776 148550
rect 675712 148490 675764 148546
rect 675764 148490 675776 148546
rect 675712 148486 675776 148490
rect 676672 146562 676736 146626
rect 144832 144786 144896 144850
rect 671683 142630 672775 143722
rect 708743 142629 709837 143723
rect 666067 140223 667249 141405
rect 698402 140222 699586 141406
rect 210304 137238 210368 137302
rect 211072 137238 211136 137302
rect 641093 135469 643327 137703
rect 645421 137217 647655 139451
rect 700550 137492 701734 138676
rect 706922 135506 708106 136690
rect 677440 133390 677504 133454
rect 677056 132206 677120 132270
rect 677248 131762 677312 131826
rect 673984 128654 674048 128718
rect 144832 126730 144896 126794
rect 674176 125990 674240 126054
rect 210496 125102 210560 125166
rect 144640 124510 144704 124574
rect 210304 123030 210368 123094
rect 211072 123030 211136 123094
rect 210304 121698 210368 121762
rect 210112 121314 210176 121318
rect 210112 121258 210164 121314
rect 210164 121258 210176 121314
rect 210112 121254 210176 121258
rect 210304 121254 210368 121318
rect 48196 115126 51046 120616
rect 210304 117998 210368 118062
rect 211072 117998 211136 118062
rect 676480 117998 676544 118062
rect 675904 117850 675968 117914
rect 144256 113322 144320 113326
rect 144256 113266 144308 113322
rect 144308 113266 144320 113322
rect 144256 113262 144320 113266
rect 675328 110066 675392 110070
rect 675328 110010 675380 110066
rect 675380 110010 675392 110066
rect 675328 110006 675392 110010
rect 675520 109326 675584 109330
rect 675520 109270 675532 109326
rect 675532 109270 675584 109326
rect 675520 109266 675584 109270
rect 673984 108082 674048 108146
rect 144256 106750 144320 106814
rect 144640 106602 144704 106666
rect 209728 106454 209792 106518
rect 210496 106454 210560 106518
rect 674176 105122 674240 105186
rect 675904 103198 675968 103262
rect 676480 101422 676544 101486
rect 210112 90914 210176 90978
rect 210496 90914 210560 90978
rect 210112 90322 210176 90386
rect 211072 90322 211136 90386
rect 210688 89286 210752 89350
rect 211072 89286 211136 89350
rect 210304 87658 210368 87722
rect 211072 87658 211136 87722
rect 210688 87214 210752 87278
rect 211072 87214 211136 87278
rect 210112 82626 210176 82690
rect 210880 82626 210944 82690
rect 40974 69066 45006 82236
rect 210112 72858 210176 72922
rect 211072 72858 211136 72922
rect 209920 62794 209984 62858
rect 210304 62498 210368 62562
rect 211072 58206 211136 58270
rect 210304 54210 210368 54274
rect 211648 54210 211712 54274
rect 209920 54062 209984 54126
rect 212800 54062 212864 54126
rect 211072 53914 211136 53978
rect 209728 53766 209792 53830
rect 212224 53618 212288 53682
rect 212992 53530 213056 53534
rect 212992 53474 213044 53530
rect 213044 53474 213056 53530
rect 212992 53470 213056 53474
rect 212416 53322 212480 53386
rect 211456 53174 211520 53238
rect 637312 52286 637376 52350
rect 637888 52138 637952 52202
rect 637504 51990 637568 52054
rect 637696 51842 637760 51906
rect 637120 51694 637184 51758
rect 636928 51546 636992 51610
rect 145408 51398 145472 51462
rect 145792 51250 145856 51314
rect 145600 51102 145664 51166
rect 145984 50954 146048 51018
rect 471040 49030 471104 49094
rect 521344 45034 521408 45098
rect 527104 44886 527168 44950
rect 521344 43258 521408 43322
rect 527104 43258 527168 43322
rect 471040 42134 471104 42138
rect 471040 42078 471092 42134
rect 471092 42078 471104 42134
rect 471040 42074 471104 42078
rect 189952 41778 190016 41842
rect 189952 40594 190016 40658
rect 245742 40136 251484 41648
rect 469504 40742 469568 40806
rect 469312 40594 469376 40658
rect 573642 40312 579070 42478
<< metal4 >>
rect 125333 1031610 125935 1031611
rect 125333 1031433 125334 1031610
rect 109840 1031113 125334 1031433
rect 125333 1031010 125334 1031113
rect 125934 1031010 125935 1031610
rect 125333 1031009 125935 1031010
rect 124005 1030858 124607 1030859
rect 124005 1030773 124006 1030858
rect 109282 1030453 124006 1030773
rect 124005 1030258 124006 1030453
rect 124606 1030773 124607 1030858
rect 124606 1030453 124620 1030773
rect 124606 1030258 124607 1030453
rect 124005 1030257 124607 1030258
rect 223905 1022792 224507 1022793
rect 173267 1022788 173869 1022789
rect 121357 1022708 121959 1022709
rect 121357 1022489 121358 1022708
rect 108124 1022169 121358 1022489
rect 121357 1022108 121358 1022169
rect 121958 1022489 121959 1022708
rect 173267 1022489 173268 1022788
rect 121958 1022169 122024 1022489
rect 159562 1022188 173268 1022489
rect 173868 1022188 173869 1022788
rect 223905 1022489 223906 1022792
rect 159562 1022187 173869 1022188
rect 211082 1022192 223906 1022489
rect 224506 1022489 224507 1022792
rect 568177 1022764 568779 1022765
rect 377195 1022758 377797 1022759
rect 274879 1022726 275481 1022727
rect 274879 1022489 274880 1022726
rect 224506 1022192 224648 1022489
rect 159562 1022169 173832 1022187
rect 211082 1022169 224648 1022192
rect 262308 1022169 274880 1022489
rect 121958 1022108 121959 1022169
rect 274879 1022126 274880 1022169
rect 275480 1022126 275481 1022726
rect 327773 1022684 328375 1022685
rect 327773 1022489 327774 1022684
rect 313756 1022169 327774 1022489
rect 274879 1022125 275481 1022126
rect 121357 1022107 121959 1022108
rect 276373 1022110 276975 1022111
rect 225483 1022096 226085 1022097
rect 174519 1022050 175121 1022051
rect 122815 1022042 123417 1022043
rect 122815 1021829 122816 1022042
rect 108618 1021509 122816 1021829
rect 122815 1021442 122816 1021509
rect 123416 1021829 123417 1022042
rect 174519 1021829 174520 1022050
rect 123416 1021509 123418 1021829
rect 160040 1021509 174520 1021829
rect 123416 1021442 123417 1021509
rect 174519 1021450 174520 1021509
rect 175120 1021450 175121 1022050
rect 225483 1021829 225484 1022096
rect 211604 1021509 225484 1021829
rect 225483 1021496 225484 1021509
rect 226084 1021829 226085 1022096
rect 276373 1021829 276374 1022110
rect 226084 1021509 226130 1021829
rect 262704 1021510 276374 1021829
rect 276974 1021510 276975 1022110
rect 327773 1022084 327774 1022169
rect 328374 1022084 328375 1022684
rect 377195 1022489 377196 1022758
rect 364336 1022169 377196 1022489
rect 377195 1022158 377196 1022169
rect 377796 1022489 377797 1022758
rect 410145 1022632 410747 1022633
rect 410145 1022489 410146 1022632
rect 377796 1022169 377844 1022489
rect 409988 1022169 410146 1022489
rect 377796 1022158 377797 1022169
rect 377195 1022157 377797 1022158
rect 327773 1022083 328375 1022084
rect 378529 1022096 379131 1022097
rect 329331 1021934 329933 1021935
rect 329331 1021829 329332 1021934
rect 262704 1021509 276975 1021510
rect 314504 1021509 329332 1021829
rect 226084 1021496 226085 1021509
rect 225483 1021495 226085 1021496
rect 174519 1021449 175121 1021450
rect 122815 1021441 123417 1021442
rect 227323 1021398 227925 1021399
rect 176203 1021268 176805 1021269
rect 176203 1021169 176204 1021268
rect 160344 1020849 176204 1021169
rect 176203 1020668 176204 1020849
rect 176804 1021169 176805 1021268
rect 227323 1021169 227324 1021398
rect 176804 1020849 176830 1021169
rect 211126 1020849 227324 1021169
rect 176804 1020668 176805 1020849
rect 227323 1020798 227324 1020849
rect 227924 1021169 227925 1021398
rect 329331 1021334 329332 1021509
rect 329932 1021334 329933 1021934
rect 378529 1021829 378530 1022096
rect 364602 1021509 378530 1021829
rect 378529 1021496 378530 1021509
rect 379130 1021496 379131 1022096
rect 410145 1022032 410146 1022169
rect 410746 1022489 410747 1022632
rect 491649 1022572 492251 1022573
rect 491649 1022489 491650 1022572
rect 410746 1022169 423200 1022489
rect 491646 1022169 491650 1022489
rect 410746 1022032 410747 1022169
rect 410145 1022031 410747 1022032
rect 491649 1021972 491650 1022169
rect 492250 1022489 492251 1022572
rect 568177 1022489 568178 1022764
rect 492250 1022169 500480 1022489
rect 560340 1022169 568178 1022489
rect 492250 1021972 492251 1022169
rect 568177 1022164 568178 1022169
rect 568778 1022489 568779 1022764
rect 568778 1022169 568814 1022489
rect 568778 1022164 568779 1022169
rect 568177 1022163 568779 1022164
rect 491649 1021971 492251 1021972
rect 570327 1022042 570929 1022043
rect 493069 1021882 493671 1021883
rect 412096 1021702 422760 1021829
rect 412096 1021509 412148 1021702
rect 378529 1021495 379131 1021496
rect 329331 1021333 329933 1021334
rect 330887 1021362 331489 1021363
rect 277779 1021316 278381 1021317
rect 277779 1021169 277780 1021316
rect 227924 1020849 227960 1021169
rect 263012 1020849 277780 1021169
rect 227924 1020798 227925 1020849
rect 227323 1020797 227925 1020798
rect 277779 1020716 277780 1020849
rect 278380 1021169 278381 1021316
rect 330887 1021169 330888 1021362
rect 278380 1020849 278396 1021169
rect 315254 1020849 330888 1021169
rect 278380 1020716 278381 1020849
rect 330887 1020762 330888 1020849
rect 331488 1020762 331489 1021362
rect 380079 1021254 380681 1021255
rect 380079 1021169 380080 1021254
rect 364646 1020849 380080 1021169
rect 330887 1020761 331489 1020762
rect 277779 1020715 278381 1020716
rect 176203 1020667 176805 1020668
rect 177459 1020702 178061 1020703
rect 177459 1020509 177460 1020702
rect 160648 1020189 177460 1020509
rect 177459 1020102 177460 1020189
rect 178060 1020102 178061 1020702
rect 332435 1020700 333037 1020701
rect 278921 1020656 279523 1020657
rect 228773 1020614 229375 1020615
rect 228773 1020509 228774 1020614
rect 212128 1020189 228774 1020509
rect 177459 1020101 178061 1020102
rect 228773 1020014 228774 1020189
rect 229374 1020509 229375 1020614
rect 278921 1020509 278922 1020656
rect 229374 1020189 229442 1020509
rect 263012 1020189 278922 1020509
rect 229374 1020014 229375 1020189
rect 278921 1020056 278922 1020189
rect 279522 1020056 279523 1020656
rect 332435 1020509 332436 1020700
rect 314946 1020189 332436 1020509
rect 332435 1020100 332436 1020189
rect 333036 1020100 333037 1020700
rect 380079 1020654 380080 1020849
rect 380680 1020654 380681 1021254
rect 412147 1021102 412148 1021509
rect 412748 1021509 422760 1021702
rect 412748 1021102 412749 1021509
rect 493069 1021282 493070 1021882
rect 493670 1021829 493671 1021882
rect 570327 1021829 570328 1022042
rect 493670 1021509 500084 1021829
rect 560964 1021509 570328 1021829
rect 493670 1021282 493671 1021509
rect 570327 1021442 570328 1021509
rect 570928 1021829 570929 1022042
rect 570928 1021509 570934 1021829
rect 570928 1021442 570929 1021509
rect 570327 1021441 570929 1021442
rect 571833 1021444 572435 1021445
rect 493069 1021281 493671 1021282
rect 571833 1021169 571834 1021444
rect 412147 1021101 412749 1021102
rect 414312 1021156 423450 1021169
rect 414312 1020849 414358 1021156
rect 380079 1020653 380681 1020654
rect 381547 1020680 382149 1020681
rect 381547 1020509 381548 1020680
rect 364912 1020189 381548 1020509
rect 332435 1020099 333037 1020100
rect 381547 1020080 381548 1020189
rect 382148 1020509 382149 1020680
rect 414357 1020556 414358 1020849
rect 414958 1020849 423450 1021156
rect 494534 1021166 499320 1021169
rect 494534 1020849 494582 1021166
rect 414958 1020556 414959 1020849
rect 414357 1020555 414959 1020556
rect 415921 1020566 416523 1020567
rect 382148 1020189 382268 1020509
rect 382148 1020080 382149 1020189
rect 381547 1020079 382149 1020080
rect 278921 1020055 279523 1020056
rect 228773 1020013 229375 1020014
rect 415921 1019966 415922 1020566
rect 416522 1020509 416523 1020566
rect 494581 1020566 494582 1020849
rect 495182 1020849 499320 1021166
rect 561438 1020849 571834 1021169
rect 495182 1020566 495183 1020849
rect 571833 1020844 571834 1020849
rect 572434 1021169 572435 1021444
rect 572434 1020849 572580 1021169
rect 572434 1020844 572435 1020849
rect 571833 1020843 572435 1020844
rect 494581 1020565 495183 1020566
rect 573445 1020596 574047 1020597
rect 496095 1020550 496697 1020551
rect 416522 1020189 422174 1020509
rect 416522 1019966 416523 1020189
rect 415921 1019965 416523 1019966
rect 496095 1019950 496096 1020550
rect 496696 1020509 496697 1020550
rect 573445 1020509 573446 1020596
rect 496696 1020189 499862 1020509
rect 560738 1020189 573446 1020509
rect 496696 1019950 496697 1020189
rect 573445 1019996 573446 1020189
rect 574046 1019996 574047 1020596
rect 573445 1019995 574047 1019996
rect 496095 1019949 496697 1019950
rect 60222 1000238 62794 1000290
rect 60222 999438 60258 1000238
rect 62730 999438 62794 1000238
rect 60222 999380 62794 999438
rect 125334 997663 125934 997664
rect 60236 997622 62784 997650
rect 54692 997038 56068 997236
rect 54692 996198 54718 997038
rect 60236 996948 60276 997622
rect 62750 996948 62784 997622
rect 122816 997633 123416 997634
rect 60236 996908 62784 996948
rect 121358 997559 121958 997560
rect 121358 996961 121359 997559
rect 121957 996961 121958 997559
rect 53092 995752 54534 995978
rect 53092 994938 53140 995752
rect 54504 994938 54534 995752
rect 51584 994554 52914 994654
rect 51584 993544 51620 994554
rect 52878 993544 52914 994554
rect 49632 993104 51436 993248
rect 49632 992148 49664 993104
rect 51396 992148 51436 993104
rect 44866 990200 45466 990402
rect 30764 988352 31690 988390
rect 30764 984370 30806 988352
rect 31614 984370 31690 988352
rect 41094 988148 42430 988188
rect 41094 984514 41134 988148
rect 42390 984514 42430 988148
rect 41094 984474 42430 984514
rect 43272 985556 44476 985638
rect 43272 985550 44494 985556
rect 30764 984328 31690 984370
rect 43272 983126 43290 985550
rect 44470 985138 44494 985550
rect 44470 983126 44492 985138
rect 43272 983088 44492 983126
rect 42111 968766 42177 968767
rect 42111 968702 42112 968766
rect 42176 968702 42177 968766
rect 42111 968701 42177 968702
rect 41343 967138 41409 967139
rect 41343 967074 41344 967138
rect 41408 967074 41409 967138
rect 41343 967073 41409 967074
rect 40959 964030 41025 964031
rect 40959 963966 40960 964030
rect 41024 963966 41025 964030
rect 40959 963965 41025 963966
rect 40767 962698 40833 962699
rect 40767 962634 40768 962698
rect 40832 962634 40833 962698
rect 40767 962633 40833 962634
rect 40383 962106 40449 962107
rect 40383 962042 40384 962106
rect 40448 962042 40449 962106
rect 40383 962041 40449 962042
rect 8927 952833 9247 952998
rect 8751 952832 9553 952833
rect 8751 952032 8752 952832
rect 9552 952032 9553 952832
rect 8751 952031 9553 952032
rect 7607 949283 7927 949324
rect 7285 949282 8087 949283
rect 7285 948482 7286 949282
rect 8086 948482 8087 949282
rect 7285 948481 8087 948482
rect 7607 944198 7927 948481
rect 8927 942590 9247 952031
rect 16551 951107 16871 951150
rect 16319 951106 17121 951107
rect 16319 950306 16320 951106
rect 17120 950306 17121 951106
rect 16319 950305 17121 950306
rect 16551 943166 16871 950305
rect 17871 947747 18191 947762
rect 17617 947746 18419 947747
rect 17617 946946 17618 947746
rect 18418 946946 18419 947746
rect 17617 946945 18419 946946
rect 17871 944632 18191 946945
rect 40191 941386 40257 941387
rect 40191 941322 40192 941386
rect 40256 941322 40257 941386
rect 40191 941321 40257 941322
rect 40194 938757 40254 941321
rect 40386 939167 40446 962041
rect 40575 958554 40641 958555
rect 40575 958490 40576 958554
rect 40640 958490 40641 958554
rect 40575 958489 40641 958490
rect 40383 939166 40449 939167
rect 40383 939102 40384 939166
rect 40448 939102 40449 939166
rect 40383 939101 40449 939102
rect 40194 938697 40446 938757
rect 8927 826521 9247 826642
rect 8803 826520 9605 826521
rect 8803 825720 8804 826520
rect 9604 825720 9605 826520
rect 8803 825719 9605 825720
rect 7607 823501 7927 823628
rect 7283 823500 8085 823501
rect 7283 822700 7284 823500
rect 8084 822700 8085 823500
rect 7283 822699 8085 822700
rect 7607 818178 7927 822699
rect 8927 816920 9247 825719
rect 16551 825059 16871 825146
rect 16353 825058 17155 825059
rect 16353 824258 16354 825058
rect 17154 824258 17155 825058
rect 16353 824257 17155 824258
rect 16551 817490 16871 824257
rect 17871 822227 18191 822322
rect 17445 822226 18247 822227
rect 17445 821426 17446 822226
rect 18246 821426 18247 822226
rect 17445 821425 18247 821426
rect 17871 818772 18191 821425
rect 40386 816031 40446 938697
rect 40578 937687 40638 958489
rect 40575 937686 40641 937687
rect 40575 937622 40576 937686
rect 40640 937622 40641 937686
rect 40575 937621 40641 937622
rect 40770 934875 40830 962633
rect 40767 934874 40833 934875
rect 40767 934810 40768 934874
rect 40832 934810 40833 934874
rect 40767 934809 40833 934810
rect 40962 934431 41022 963965
rect 41151 963290 41217 963291
rect 41151 963226 41152 963290
rect 41216 963226 41217 963290
rect 41151 963225 41217 963226
rect 41154 935911 41214 963225
rect 41346 940943 41406 967073
rect 41535 959738 41601 959739
rect 41535 959674 41536 959738
rect 41600 959674 41601 959738
rect 41535 959673 41601 959674
rect 41343 940942 41409 940943
rect 41343 940878 41344 940942
rect 41408 940878 41409 940942
rect 41343 940877 41409 940878
rect 41151 935910 41217 935911
rect 41151 935846 41152 935910
rect 41216 935846 41217 935910
rect 41151 935845 41217 935846
rect 41538 935467 41598 959673
rect 41727 959146 41793 959147
rect 41727 959082 41728 959146
rect 41792 959082 41793 959146
rect 41727 959081 41793 959082
rect 41730 937095 41790 959081
rect 41919 957814 41985 957815
rect 41919 957750 41920 957814
rect 41984 957750 41985 957814
rect 41919 957749 41985 957750
rect 41922 939759 41982 957749
rect 41919 939758 41985 939759
rect 41919 939694 41920 939758
rect 41984 939694 41985 939758
rect 41919 939693 41985 939694
rect 42114 938723 42174 968701
rect 42303 965066 42369 965067
rect 42303 965002 42304 965066
rect 42368 965002 42369 965066
rect 42303 965001 42369 965002
rect 42306 945679 42366 965001
rect 42687 961958 42753 961959
rect 42687 961894 42688 961958
rect 42752 961894 42753 961958
rect 42687 961893 42753 961894
rect 42690 960479 42750 961893
rect 42687 960478 42753 960479
rect 42687 960414 42688 960478
rect 42752 960414 42753 960478
rect 42687 960413 42753 960414
rect 42495 955890 42561 955891
rect 42495 955826 42496 955890
rect 42560 955826 42561 955890
rect 42495 955825 42561 955826
rect 42303 945678 42369 945679
rect 42303 945614 42304 945678
rect 42368 945614 42369 945678
rect 42303 945613 42369 945614
rect 42498 941387 42558 955825
rect 42495 941386 42561 941387
rect 42495 941322 42496 941386
rect 42560 941322 42561 941386
rect 42495 941321 42561 941322
rect 42111 938722 42177 938723
rect 42111 938658 42112 938722
rect 42176 938658 42177 938722
rect 42111 938657 42177 938658
rect 41727 937094 41793 937095
rect 41727 937030 41728 937094
rect 41792 937030 41793 937094
rect 41727 937029 41793 937030
rect 41535 935466 41601 935467
rect 41535 935402 41536 935466
rect 41600 935402 41601 935466
rect 41535 935401 41601 935402
rect 40959 934430 41025 934431
rect 40959 934366 40960 934430
rect 41024 934366 41025 934430
rect 40959 934365 41025 934366
rect 40383 816030 40449 816031
rect 40383 815966 40384 816030
rect 40448 815966 40449 816030
rect 40383 815965 40449 815966
rect 8927 783777 9247 783970
rect 8577 783776 9379 783777
rect 8577 782976 8578 783776
rect 9378 782976 9379 783776
rect 8577 782975 9379 782976
rect 7233 781240 8035 781241
rect 7233 780440 7234 781240
rect 8034 780440 8035 781240
rect 7233 780439 8035 780440
rect 7607 774692 7927 780439
rect 8927 773772 9247 782975
rect 16551 782649 16871 782720
rect 16309 782648 17111 782649
rect 16309 781848 16310 782648
rect 17110 781848 17111 782648
rect 16309 781847 17111 781848
rect 16551 774268 16871 781847
rect 17871 779785 18191 779820
rect 17581 779784 18383 779785
rect 17581 778984 17582 779784
rect 18382 778984 18383 779784
rect 17581 778983 18383 778984
rect 17871 775800 18191 778983
rect 40386 773589 40446 815965
rect 40575 813958 40641 813959
rect 40575 813894 40576 813958
rect 40640 813894 40641 813958
rect 40575 813893 40641 813894
rect 40578 791759 40638 813893
rect 40767 811738 40833 811739
rect 40767 811674 40768 811738
rect 40832 811674 40833 811738
rect 40767 811673 40833 811674
rect 40770 791907 40830 811673
rect 40959 802118 41025 802119
rect 40959 802054 40960 802118
rect 41024 802054 41025 802118
rect 40959 802053 41025 802054
rect 40767 791906 40833 791907
rect 40767 791842 40768 791906
rect 40832 791842 40833 791906
rect 40767 791841 40833 791842
rect 40575 791758 40641 791759
rect 40575 791694 40576 791758
rect 40640 791694 40641 791758
rect 40575 791693 40641 791694
rect 40386 773529 40638 773589
rect 40383 772814 40449 772815
rect 40383 772750 40384 772814
rect 40448 772750 40449 772814
rect 40383 772749 40449 772750
rect 8927 740589 9247 740660
rect 8759 740588 9561 740589
rect 8759 739788 8760 740588
rect 9560 739788 9561 740588
rect 8759 739787 9561 739788
rect 7607 737833 7927 737840
rect 7421 737832 8223 737833
rect 7421 737032 7422 737832
rect 8222 737032 8223 737832
rect 7421 737031 8223 737032
rect 7607 731808 7927 737031
rect 8927 730350 9247 739787
rect 16551 739235 16871 739322
rect 16423 739234 17225 739235
rect 16423 738434 16424 739234
rect 17224 738434 17225 739234
rect 16423 738433 17225 738434
rect 16551 731102 16871 738433
rect 17871 736151 18191 736172
rect 17527 736150 18329 736151
rect 17527 735350 17528 736150
rect 18328 735350 18329 736150
rect 17527 735349 18329 735350
rect 17871 731972 18191 735349
rect 40386 729633 40446 772749
rect 40578 772371 40638 773529
rect 40962 773407 41022 802053
rect 41919 800490 41985 800491
rect 41919 800426 41920 800490
rect 41984 800426 41985 800490
rect 41919 800425 41985 800426
rect 41922 792647 41982 800425
rect 42303 800342 42369 800343
rect 42303 800278 42304 800342
rect 42368 800278 42369 800342
rect 42303 800277 42369 800278
rect 42111 797678 42177 797679
rect 42111 797614 42112 797678
rect 42176 797614 42177 797678
rect 42111 797613 42177 797614
rect 41919 792646 41985 792647
rect 41919 792582 41920 792646
rect 41984 792582 41985 792646
rect 41919 792581 41985 792582
rect 42114 791315 42174 797613
rect 42306 797087 42366 800277
rect 42495 799750 42561 799751
rect 42495 799686 42496 799750
rect 42560 799686 42561 799750
rect 42495 799685 42561 799686
rect 42498 797531 42558 799685
rect 42495 797530 42561 797531
rect 42495 797466 42496 797530
rect 42560 797466 42561 797530
rect 42495 797465 42561 797466
rect 42303 797086 42369 797087
rect 42303 797022 42304 797086
rect 42368 797022 42369 797086
rect 42303 797021 42369 797022
rect 42111 791314 42177 791315
rect 42111 791250 42112 791314
rect 42176 791250 42177 791314
rect 42111 791249 42177 791250
rect 41727 791166 41793 791167
rect 41727 791102 41728 791166
rect 41792 791102 41793 791166
rect 41727 791101 41793 791102
rect 40959 773406 41025 773407
rect 40959 773342 40960 773406
rect 41024 773342 41025 773406
rect 40959 773341 41025 773342
rect 40575 772370 40641 772371
rect 40575 772306 40576 772370
rect 40640 772306 40641 772370
rect 40575 772305 40641 772306
rect 40578 730299 40638 772305
rect 41343 768670 41409 768671
rect 41343 768606 41344 768670
rect 41408 768606 41409 768670
rect 41343 768605 41409 768606
rect 40767 760234 40833 760235
rect 40767 760170 40768 760234
rect 40832 760170 40833 760234
rect 40767 760169 40833 760170
rect 40770 746915 40830 760169
rect 40767 746914 40833 746915
rect 40767 746850 40768 746914
rect 40832 746850 40833 746914
rect 40767 746849 40833 746850
rect 41346 746175 41406 768605
rect 41535 757422 41601 757423
rect 41535 757358 41536 757422
rect 41600 757358 41601 757422
rect 41535 757357 41601 757358
rect 41538 751799 41598 757357
rect 41535 751798 41601 751799
rect 41535 751734 41536 751798
rect 41600 751734 41601 751798
rect 41535 751733 41601 751734
rect 41730 747615 41790 791101
rect 41919 757126 41985 757127
rect 41919 757062 41920 757126
rect 41984 757062 41985 757126
rect 41919 757061 41985 757062
rect 41922 751059 41982 757061
rect 41919 751058 41985 751059
rect 41919 750994 41920 751058
rect 41984 750994 41985 751058
rect 41919 750993 41985 750994
rect 42114 750612 42174 791249
rect 42690 791167 42750 960413
rect 42879 945678 42945 945679
rect 42879 945614 42880 945678
rect 42944 945614 42945 945678
rect 42879 945613 42945 945614
rect 42882 936207 42942 945613
rect 42879 936206 42945 936207
rect 42879 936142 42880 936206
rect 42944 936142 42945 936206
rect 42879 936141 42945 936142
rect 43272 922410 44476 983088
rect 43126 922378 44496 922410
rect 43126 916604 43192 922378
rect 44420 916604 44496 922378
rect 43126 916538 44496 916604
rect 42687 791166 42753 791167
rect 42687 791102 42688 791166
rect 42752 791102 42753 791166
rect 42687 791101 42753 791102
rect 42303 765266 42369 765267
rect 42303 765202 42304 765266
rect 42368 765202 42369 765266
rect 42303 765201 42369 765202
rect 42306 750615 42366 765201
rect 42495 760234 42561 760235
rect 42495 760170 42496 760234
rect 42560 760170 42561 760234
rect 42495 760169 42561 760170
rect 42498 754907 42558 760169
rect 43071 759198 43137 759199
rect 43071 759134 43072 759198
rect 43136 759134 43137 759198
rect 43071 759133 43137 759134
rect 42687 757126 42753 757127
rect 42687 757062 42688 757126
rect 42752 757062 42753 757126
rect 42687 757061 42753 757062
rect 42495 754906 42561 754907
rect 42495 754842 42496 754906
rect 42560 754842 42561 754906
rect 42495 754841 42561 754842
rect 42690 751651 42750 757061
rect 42879 751946 42945 751947
rect 42879 751882 42880 751946
rect 42944 751882 42945 751946
rect 42879 751881 42945 751882
rect 42687 751650 42753 751651
rect 42687 751586 42688 751650
rect 42752 751586 42753 751650
rect 42687 751585 42753 751586
rect 41922 750552 42174 750612
rect 42303 750614 42369 750615
rect 41922 748691 41982 750552
rect 42303 750550 42304 750614
rect 42368 750550 42369 750614
rect 42303 750549 42369 750550
rect 42882 749727 42942 751881
rect 43074 750319 43134 759133
rect 43071 750318 43137 750319
rect 43071 750254 43072 750318
rect 43136 750254 43137 750318
rect 43071 750253 43137 750254
rect 42879 749726 42945 749727
rect 42879 749662 42880 749726
rect 42944 749662 42945 749726
rect 42879 749661 42945 749662
rect 41919 748690 41985 748691
rect 41919 748626 41920 748690
rect 41984 748626 41985 748690
rect 41919 748625 41985 748626
rect 41538 747555 41790 747615
rect 41538 747211 41598 747555
rect 41535 747210 41601 747211
rect 41535 747146 41536 747210
rect 41600 747146 41601 747210
rect 41535 747145 41601 747146
rect 41343 746174 41409 746175
rect 41343 746110 41344 746174
rect 41408 746110 41409 746174
rect 41343 746109 41409 746110
rect 40578 730239 41214 730299
rect 40386 729599 40638 729633
rect 40386 729598 40641 729599
rect 40386 729573 40576 729598
rect 40575 729534 40576 729573
rect 40640 729534 40641 729598
rect 40575 729533 40641 729534
rect 8927 697143 9247 697246
rect 8705 697142 9507 697143
rect 8705 696342 8706 697142
rect 9506 696342 9507 697142
rect 8705 696341 9507 696342
rect 7607 694755 7927 694864
rect 7211 694754 8013 694755
rect 7211 693954 7212 694754
rect 8012 693954 8013 694754
rect 7211 693953 8013 693954
rect 7607 688640 7927 693953
rect 8927 687332 9247 696341
rect 16551 695869 16871 695906
rect 16331 695868 17133 695869
rect 16331 695068 16332 695868
rect 17132 695068 17133 695868
rect 16331 695067 17133 695068
rect 16551 687896 16871 695067
rect 17871 693085 18191 693170
rect 17797 693084 18599 693085
rect 17797 692284 17798 693084
rect 18598 692284 18599 693084
rect 17797 692283 18599 692284
rect 17871 688886 18191 692283
rect 40578 686975 40638 729533
rect 41154 729155 41214 730239
rect 41151 729154 41217 729155
rect 41151 729090 41152 729154
rect 41216 729090 41217 729154
rect 41151 729089 41217 729090
rect 40959 725306 41025 725307
rect 40959 725242 40960 725306
rect 41024 725242 41025 725306
rect 40959 725241 41025 725242
rect 40767 714206 40833 714207
rect 40767 714142 40768 714206
rect 40832 714142 40833 714206
rect 40767 714141 40833 714142
rect 40770 707251 40830 714141
rect 40767 707250 40833 707251
rect 40767 707186 40768 707250
rect 40832 707186 40833 707250
rect 40767 707185 40833 707186
rect 40962 703403 41022 725241
rect 40959 703402 41025 703403
rect 40959 703338 40960 703402
rect 41024 703338 41025 703402
rect 40959 703337 41025 703338
rect 40575 686974 40641 686975
rect 40575 686910 40576 686974
rect 40640 686910 40641 686974
rect 40575 686909 40641 686910
rect 41154 685939 41214 729089
rect 41343 727526 41409 727527
rect 41343 727462 41344 727526
rect 41408 727462 41409 727526
rect 41343 727461 41409 727462
rect 41346 705179 41406 727461
rect 41538 715687 41598 747145
rect 41727 722050 41793 722051
rect 41727 721986 41728 722050
rect 41792 721986 41793 722050
rect 41727 721985 41793 721986
rect 41535 715686 41601 715687
rect 41535 715622 41536 715686
rect 41600 715622 41601 715686
rect 41535 715621 41601 715622
rect 41730 714981 41790 721985
rect 41922 715835 41982 748625
rect 42879 725084 42945 725085
rect 42879 725020 42880 725084
rect 42944 725020 42945 725084
rect 42879 725019 42945 725020
rect 41919 715834 41985 715835
rect 41919 715770 41920 715834
rect 41984 715770 41985 715834
rect 41919 715769 41985 715770
rect 42495 715686 42561 715687
rect 42495 715622 42496 715686
rect 42560 715622 42561 715686
rect 42495 715621 42561 715622
rect 41538 714921 41790 714981
rect 41538 707399 41598 714921
rect 41727 714206 41793 714207
rect 41727 714142 41728 714206
rect 41792 714142 41793 714206
rect 41727 714141 41793 714142
rect 41730 711247 41790 714141
rect 41919 713910 41985 713911
rect 41919 713846 41920 713910
rect 41984 713846 41985 713910
rect 41919 713845 41985 713846
rect 42111 713910 42177 713911
rect 42111 713846 42112 713910
rect 42176 713846 42177 713910
rect 42111 713845 42177 713846
rect 41922 711691 41982 713845
rect 41919 711690 41985 711691
rect 41919 711626 41920 711690
rect 41984 711626 41985 711690
rect 41919 711625 41985 711626
rect 41727 711246 41793 711247
rect 41727 711182 41728 711246
rect 41792 711182 41793 711246
rect 41727 711181 41793 711182
rect 41727 711098 41793 711099
rect 41727 711034 41728 711098
rect 41792 711034 41793 711098
rect 41727 711033 41793 711034
rect 41535 707398 41601 707399
rect 41535 707334 41536 707398
rect 41600 707334 41601 707398
rect 41535 707333 41601 707334
rect 41343 705178 41409 705179
rect 41343 705114 41344 705178
rect 41408 705114 41409 705178
rect 41343 705113 41409 705114
rect 41730 704143 41790 711033
rect 42114 709915 42174 713845
rect 42303 711690 42369 711691
rect 42303 711626 42304 711690
rect 42368 711626 42369 711690
rect 42303 711625 42369 711626
rect 42306 710951 42366 711625
rect 42498 711099 42558 715621
rect 42495 711098 42561 711099
rect 42495 711034 42496 711098
rect 42560 711034 42561 711098
rect 42495 711033 42561 711034
rect 42303 710950 42369 710951
rect 42303 710886 42304 710950
rect 42368 710886 42369 710950
rect 42303 710885 42369 710886
rect 42111 709914 42177 709915
rect 42111 709850 42112 709914
rect 42176 709850 42177 709914
rect 42111 709849 42177 709850
rect 42687 706954 42753 706955
rect 42687 706890 42688 706954
rect 42752 706890 42753 706954
rect 42687 706889 42753 706890
rect 42690 705657 42750 706889
rect 42882 706511 42942 725019
rect 43272 716550 44476 916538
rect 44866 841528 45466 989600
rect 46142 989156 46742 989724
rect 44818 841394 45864 841528
rect 44818 828278 44902 841394
rect 45730 828278 45864 841394
rect 44818 828210 45864 828278
rect 43272 716056 44488 716550
rect 43244 715834 43342 715848
rect 43244 715770 43270 715834
rect 43334 715770 43342 715834
rect 43244 715748 43342 715770
rect 43071 714354 43137 714355
rect 43071 714290 43072 714354
rect 43136 714290 43137 714354
rect 43071 714289 43137 714290
rect 42879 706510 42945 706511
rect 42879 706446 42880 706510
rect 42944 706446 42945 706510
rect 42879 706445 42945 706446
rect 42498 705597 42750 705657
rect 42498 704587 42558 705597
rect 42495 704586 42561 704587
rect 42495 704522 42496 704586
rect 42560 704522 42561 704586
rect 42495 704521 42561 704522
rect 41727 704142 41793 704143
rect 41727 704078 41728 704142
rect 41792 704078 41793 704142
rect 41727 704077 41793 704078
rect 40383 685938 40449 685939
rect 40383 685874 40384 685938
rect 40448 685874 40449 685938
rect 40383 685873 40449 685874
rect 41151 685938 41217 685939
rect 41151 685874 41152 685938
rect 41216 685874 41217 685938
rect 41151 685873 41217 685874
rect 8927 653817 9247 653936
rect 8565 653816 9367 653817
rect 8565 653016 8566 653816
rect 9366 653016 9367 653816
rect 8565 653015 9367 653016
rect 7607 651517 7927 651584
rect 7183 651516 7985 651517
rect 7183 650716 7184 651516
rect 7984 650716 7985 651516
rect 7183 650715 7985 650716
rect 7607 645224 7927 650715
rect 8927 643864 9247 653015
rect 16551 652621 16871 652644
rect 16289 652620 17091 652621
rect 16289 651820 16290 652620
rect 17090 651820 17091 652620
rect 16289 651819 17091 651820
rect 16551 644510 16871 651819
rect 17871 649951 18191 649970
rect 17671 649950 18473 649951
rect 17671 649150 17672 649950
rect 18472 649150 18473 649950
rect 17671 649149 18473 649150
rect 17871 646124 18191 649149
rect 40386 647015 40446 685873
rect 40575 684310 40641 684311
rect 40575 684246 40576 684310
rect 40640 684246 40641 684310
rect 40575 684245 40641 684246
rect 40578 660927 40638 684245
rect 40767 682090 40833 682091
rect 40767 682026 40768 682090
rect 40832 682026 40833 682090
rect 40767 682025 40833 682026
rect 40770 662407 40830 682025
rect 41535 678242 41601 678243
rect 41535 678178 41536 678242
rect 41600 678178 41601 678242
rect 41535 678177 41601 678178
rect 41343 670990 41409 670991
rect 41343 670926 41344 670990
rect 41408 670926 41409 670990
rect 41343 670925 41409 670926
rect 41346 664035 41406 670925
rect 41538 665367 41598 678177
rect 41730 675579 41790 704077
rect 42111 686530 42177 686531
rect 42111 686466 42112 686530
rect 42176 686466 42177 686530
rect 42111 686465 42177 686466
rect 41727 675578 41793 675579
rect 41727 675514 41728 675578
rect 41792 675514 41793 675578
rect 41727 675513 41793 675514
rect 41919 670546 41985 670547
rect 41919 670482 41920 670546
rect 41984 670482 41985 670546
rect 41919 670481 41985 670482
rect 41535 665366 41601 665367
rect 41535 665302 41536 665366
rect 41600 665302 41601 665366
rect 41535 665301 41601 665302
rect 41343 664034 41409 664035
rect 41343 663970 41344 664034
rect 41408 663970 41409 664034
rect 41343 663969 41409 663970
rect 40767 662406 40833 662407
rect 40767 662342 40768 662406
rect 40832 662342 40833 662406
rect 40767 662341 40833 662342
rect 41727 662258 41793 662259
rect 41727 662194 41728 662258
rect 41792 662194 41793 662258
rect 41727 662193 41793 662194
rect 40575 660926 40641 660927
rect 40575 660862 40576 660926
rect 40640 660862 40641 660926
rect 40575 660861 40641 660862
rect 40383 647014 40449 647015
rect 40383 646950 40384 647014
rect 40448 646950 40449 647014
rect 40383 646949 40449 646950
rect 40959 641094 41025 641095
rect 40959 641030 40960 641094
rect 41024 641030 41025 641094
rect 40959 641029 41025 641030
rect 40575 638874 40641 638875
rect 40575 638810 40576 638874
rect 40640 638810 40641 638874
rect 40575 638809 40641 638810
rect 40578 616527 40638 638809
rect 40962 617267 41022 641029
rect 41535 627774 41601 627775
rect 41535 627710 41536 627774
rect 41600 627710 41601 627774
rect 41535 627709 41601 627710
rect 41538 619635 41598 627709
rect 41535 619634 41601 619635
rect 41535 619570 41536 619634
rect 41600 619570 41601 619634
rect 41535 619569 41601 619570
rect 41730 618303 41790 662193
rect 41922 661075 41982 670481
rect 41919 661074 41985 661075
rect 41919 661010 41920 661074
rect 41984 661010 41985 661074
rect 41919 661009 41985 661010
rect 41727 618302 41793 618303
rect 41727 618238 41728 618302
rect 41792 618238 41793 618302
rect 41727 618237 41793 618238
rect 41922 617711 41982 661009
rect 42114 647163 42174 686465
rect 42303 670990 42369 670991
rect 42303 670926 42304 670990
rect 42368 670926 42369 670990
rect 42498 670988 42558 704521
rect 43074 700591 43134 714289
rect 43270 706955 43334 715748
rect 43267 706954 43334 706955
rect 43267 706890 43268 706954
rect 43332 706890 43334 706954
rect 43267 706889 43333 706890
rect 43422 706690 44488 716056
rect 43272 706576 44488 706690
rect 43071 700590 43137 700591
rect 43071 700526 43072 700590
rect 43136 700526 43137 700590
rect 43071 700525 43137 700526
rect 43071 683126 43137 683127
rect 43071 683062 43072 683126
rect 43136 683062 43137 683126
rect 43071 683061 43137 683062
rect 42498 670928 42750 670988
rect 42303 670925 42369 670926
rect 42306 664775 42366 670925
rect 42495 670694 42561 670695
rect 42495 670630 42496 670694
rect 42560 670630 42561 670694
rect 42495 670629 42561 670630
rect 42303 664774 42369 664775
rect 42303 664710 42304 664774
rect 42368 664710 42369 664774
rect 42303 664709 42369 664710
rect 42498 662851 42558 670629
rect 42495 662850 42561 662851
rect 42495 662786 42496 662850
rect 42560 662786 42561 662850
rect 42495 662785 42561 662786
rect 42690 662259 42750 670928
rect 43074 670695 43134 683061
rect 43071 670694 43137 670695
rect 43071 670630 43072 670694
rect 43136 670630 43137 670694
rect 43071 670629 43137 670630
rect 42687 662258 42753 662259
rect 42687 662194 42688 662258
rect 42752 662194 42753 662258
rect 42687 662193 42753 662194
rect 42111 647162 42177 647163
rect 42111 647098 42112 647162
rect 42176 647098 42177 647162
rect 42111 647097 42177 647098
rect 42111 627626 42177 627627
rect 42111 627562 42112 627626
rect 42176 627562 42177 627626
rect 42111 627561 42177 627562
rect 42114 621559 42174 627561
rect 42303 627478 42369 627479
rect 42303 627414 42304 627478
rect 42368 627414 42369 627478
rect 42303 627413 42369 627414
rect 42306 622151 42366 627413
rect 42495 627034 42561 627035
rect 42495 626970 42496 627034
rect 42560 626970 42561 627034
rect 42495 626969 42561 626970
rect 42498 624519 42558 626969
rect 42495 624518 42561 624519
rect 42495 624454 42496 624518
rect 42560 624454 42561 624518
rect 42495 624453 42561 624454
rect 42303 622150 42369 622151
rect 42303 622086 42304 622150
rect 42368 622086 42369 622150
rect 42303 622085 42369 622086
rect 42111 621558 42177 621559
rect 42111 621494 42112 621558
rect 42176 621494 42177 621558
rect 42111 621493 42177 621494
rect 42303 618302 42369 618303
rect 42303 618238 42304 618302
rect 42368 618238 42369 618302
rect 42303 618237 42369 618238
rect 41919 617710 41985 617711
rect 41919 617646 41920 617710
rect 41984 617646 41985 617710
rect 41919 617645 41985 617646
rect 40959 617266 41025 617267
rect 40959 617202 40960 617266
rect 41024 617202 41025 617266
rect 40959 617201 41025 617202
rect 40575 616526 40641 616527
rect 40575 616462 40576 616526
rect 40640 616462 40641 616526
rect 40575 616461 40641 616462
rect 8927 610727 9247 610828
rect 8735 610726 9537 610727
rect 8735 609926 8736 610726
rect 9536 609926 9537 610726
rect 8735 609925 9537 609926
rect 7607 607893 7927 607948
rect 7317 607892 8119 607893
rect 7317 607092 7318 607892
rect 8118 607092 8119 607892
rect 7317 607091 8119 607092
rect 7607 601498 7927 607091
rect 8927 600812 9247 609925
rect 16551 609447 16871 609502
rect 16281 609446 17083 609447
rect 16281 608646 16282 609446
rect 17082 608646 17083 609446
rect 16281 608645 17083 608646
rect 16551 601224 16871 608645
rect 17871 606157 18191 606164
rect 17653 606156 18455 606157
rect 17653 605356 17654 606156
rect 18454 605356 18455 606156
rect 17653 605355 18455 605356
rect 17871 602368 18191 605355
rect 42306 605131 42366 618237
rect 42495 617710 42561 617711
rect 42495 617646 42496 617710
rect 42560 617646 42561 617710
rect 42495 617645 42561 617646
rect 42498 605131 42558 617645
rect 42303 605130 42369 605131
rect 42303 605066 42304 605130
rect 42368 605066 42369 605130
rect 42303 605065 42369 605066
rect 42495 605130 42561 605131
rect 42495 605066 42496 605130
rect 42560 605066 42561 605130
rect 42495 605065 42561 605066
rect 42303 604982 42369 604983
rect 42303 604918 42304 604982
rect 42368 604918 42369 604982
rect 42303 604917 42369 604918
rect 42495 604982 42561 604983
rect 42495 604918 42496 604982
rect 42560 604918 42561 604982
rect 42495 604917 42561 604918
rect 40383 597878 40449 597879
rect 40383 597814 40384 597878
rect 40448 597814 40449 597878
rect 40383 597813 40449 597814
rect 30591 590774 30657 590775
rect 30591 590710 30592 590774
rect 30656 590710 30657 590774
rect 30591 590709 30657 590710
rect 30594 590331 30654 590709
rect 30591 590330 30657 590331
rect 30591 590266 30592 590330
rect 30656 590266 30657 590330
rect 30591 590265 30657 590266
rect 40386 573903 40446 597813
rect 40575 595658 40641 595659
rect 40575 595594 40576 595658
rect 40640 595594 40641 595658
rect 40575 595593 40641 595594
rect 40383 573902 40449 573903
rect 40383 573838 40384 573902
rect 40448 573838 40449 573902
rect 40383 573837 40449 573838
rect 40578 573163 40638 595593
rect 42306 593769 42366 604917
rect 42498 601761 42558 604917
rect 42498 601701 42750 601761
rect 41538 593709 42366 593769
rect 41538 579083 41598 593709
rect 42111 592994 42177 592995
rect 42111 592930 42112 592994
rect 42176 592930 42177 592994
rect 42111 592929 42177 592930
rect 41919 588998 41985 588999
rect 41919 588934 41920 588998
rect 41984 588934 41985 588998
rect 41919 588933 41985 588934
rect 41922 579231 41982 588933
rect 42114 580449 42174 592929
rect 42495 591958 42561 591959
rect 42495 591894 42496 591958
rect 42560 591894 42561 591958
rect 42495 591893 42561 591894
rect 42303 584262 42369 584263
rect 42303 584198 42304 584262
rect 42368 584198 42369 584262
rect 42303 584197 42369 584198
rect 42306 581303 42366 584197
rect 42498 582447 42558 591893
rect 42690 588999 42750 601701
rect 42879 599284 42945 599285
rect 42879 599220 42880 599284
rect 42944 599220 42945 599284
rect 42879 599219 42945 599220
rect 42687 588998 42753 588999
rect 42687 588934 42688 588998
rect 42752 588934 42753 588998
rect 42687 588933 42753 588934
rect 42498 582387 42750 582447
rect 42303 581302 42369 581303
rect 42303 581238 42304 581302
rect 42368 581238 42369 581302
rect 42303 581237 42369 581238
rect 42114 580389 42366 580449
rect 41727 579230 41793 579231
rect 41727 579166 41728 579230
rect 41792 579166 41793 579230
rect 41727 579165 41793 579166
rect 41919 579230 41985 579231
rect 41919 579166 41920 579230
rect 41984 579166 41985 579230
rect 41919 579165 41985 579166
rect 41535 579082 41601 579083
rect 41535 579018 41536 579082
rect 41600 579018 41601 579082
rect 41535 579017 41601 579018
rect 41730 574495 41790 579165
rect 42306 579083 42366 580389
rect 42111 579082 42177 579083
rect 42111 579018 42112 579082
rect 42176 579018 42177 579082
rect 42111 579017 42177 579018
rect 42303 579082 42369 579083
rect 42303 579018 42304 579082
rect 42368 579018 42369 579082
rect 42303 579017 42369 579018
rect 41919 578934 41985 578935
rect 41919 578870 41920 578934
rect 41984 578870 41985 578934
rect 41919 578869 41985 578870
rect 41922 575975 41982 578869
rect 41919 575974 41985 575975
rect 41919 575910 41920 575974
rect 41984 575910 41985 575974
rect 41919 575909 41985 575910
rect 41727 574494 41793 574495
rect 41727 574430 41728 574494
rect 41792 574430 41793 574494
rect 41727 574429 41793 574430
rect 40575 573162 40641 573163
rect 40575 573098 40576 573162
rect 40640 573098 40641 573162
rect 40575 573097 40641 573098
rect 8619 567646 9421 567647
rect 8619 566846 8620 567646
rect 9420 566846 9421 567646
rect 8619 566845 9421 566846
rect 7607 565275 7927 565356
rect 7347 565274 8149 565275
rect 7347 564474 7348 565274
rect 8148 564474 8149 565274
rect 7347 564473 8149 564474
rect 7607 558900 7927 564473
rect 8927 557720 9247 566845
rect 16551 566545 16871 566584
rect 16255 566544 17057 566545
rect 16255 565744 16256 566544
rect 17056 565744 17057 566544
rect 16255 565743 17057 565744
rect 16551 558310 16871 565743
rect 17871 563823 18191 563856
rect 17619 563822 18421 563823
rect 17619 563022 17620 563822
rect 18420 563022 18421 563822
rect 17619 563021 18421 563022
rect 17871 559356 18191 563021
rect 40191 560582 40257 560583
rect 40191 560518 40192 560582
rect 40256 560518 40257 560582
rect 40191 560517 40257 560518
rect 40194 556883 40254 560517
rect 40191 556882 40257 556883
rect 40191 556818 40192 556882
rect 40256 556818 40257 556882
rect 40191 556817 40257 556818
rect 40383 554662 40449 554663
rect 40383 554598 40384 554662
rect 40448 554598 40449 554662
rect 40383 554597 40449 554598
rect 40386 530687 40446 554597
rect 40575 552442 40641 552443
rect 40575 552378 40576 552442
rect 40640 552378 40641 552442
rect 40575 552377 40641 552378
rect 40578 531279 40638 552377
rect 41730 531723 41790 574429
rect 41922 561619 41982 575909
rect 42114 574643 42174 579017
rect 42690 578935 42750 582387
rect 42687 578934 42753 578935
rect 42687 578870 42688 578934
rect 42752 578870 42753 578934
rect 42687 578869 42753 578870
rect 42882 577011 42942 599219
rect 42879 577010 42945 577011
rect 42879 576946 42880 577010
rect 42944 576946 42945 577010
rect 42879 576945 42945 576946
rect 42111 574642 42177 574643
rect 42111 574578 42112 574642
rect 42176 574578 42177 574642
rect 42111 574577 42177 574578
rect 41919 561618 41985 561619
rect 41919 561554 41920 561618
rect 41984 561554 41985 561618
rect 41919 561553 41985 561554
rect 42495 561618 42561 561619
rect 42495 561554 42496 561618
rect 42560 561554 42561 561618
rect 42495 561553 42561 561554
rect 42303 541194 42369 541195
rect 42303 541130 42304 541194
rect 42368 541130 42369 541194
rect 42303 541129 42369 541130
rect 41919 541046 41985 541047
rect 41919 540982 41920 541046
rect 41984 540982 41985 541046
rect 41919 540981 41985 540982
rect 41922 536903 41982 540981
rect 41919 536902 41985 536903
rect 41919 536838 41920 536902
rect 41984 536838 41985 536902
rect 41919 536837 41985 536838
rect 42306 533351 42366 541129
rect 42303 533350 42369 533351
rect 42303 533286 42304 533350
rect 42368 533286 42369 533350
rect 42303 533285 42369 533286
rect 42498 532759 42558 561553
rect 42879 541638 42945 541639
rect 42879 541574 42880 541638
rect 42944 541574 42945 541638
rect 42879 541573 42945 541574
rect 42687 541342 42753 541343
rect 42687 541278 42688 541342
rect 42752 541278 42753 541342
rect 42687 541277 42753 541278
rect 42690 534387 42750 541277
rect 42882 535719 42942 541573
rect 42879 535718 42945 535719
rect 42879 535654 42880 535718
rect 42944 535654 42945 535718
rect 42879 535653 42945 535654
rect 42687 534386 42753 534387
rect 42687 534322 42688 534386
rect 42752 534322 42753 534386
rect 42687 534321 42753 534322
rect 42495 532758 42561 532759
rect 42495 532694 42496 532758
rect 42560 532694 42561 532758
rect 42495 532693 42561 532694
rect 41919 531870 41985 531871
rect 41919 531806 41920 531870
rect 41984 531806 41985 531870
rect 41919 531805 41985 531806
rect 41727 531722 41793 531723
rect 41727 531658 41728 531722
rect 41792 531658 41793 531722
rect 41727 531657 41793 531658
rect 40575 531278 40641 531279
rect 40575 531214 40576 531278
rect 40640 531214 40641 531278
rect 40575 531213 40641 531214
rect 40383 530686 40449 530687
rect 40383 530622 40384 530686
rect 40448 530622 40449 530686
rect 40383 530621 40449 530622
rect 8927 439991 9247 440020
rect 8773 439990 9575 439991
rect 8773 439190 8774 439990
rect 9574 439190 9575 439990
rect 8773 439189 9575 439190
rect 7355 437096 8157 437097
rect 7355 436296 7356 437096
rect 8156 436296 8157 437096
rect 7355 436295 8157 436296
rect 7607 431392 7927 436295
rect 8927 430264 9247 439189
rect 16249 438624 17051 438625
rect 16249 437824 16250 438624
rect 17050 437824 17051 438624
rect 16249 437823 17051 437824
rect 16551 430672 16871 437823
rect 17689 435748 18491 435749
rect 17689 434948 17690 435748
rect 18490 434948 18491 435748
rect 17689 434947 18491 434948
rect 17871 432046 18191 434947
rect 40383 429306 40449 429307
rect 40383 429242 40384 429306
rect 40448 429242 40449 429306
rect 40383 429241 40449 429242
rect 8623 396838 9425 396839
rect 8623 396038 8624 396838
rect 9424 396038 9425 396838
rect 8623 396037 9425 396038
rect 7607 393887 7927 394018
rect 7321 393886 8123 393887
rect 7321 393086 7322 393886
rect 8122 393086 8123 393886
rect 7321 393085 8123 393086
rect 7607 387776 7927 393085
rect 8927 386924 9247 396037
rect 16361 395406 17163 395407
rect 16361 394606 16362 395406
rect 17162 394606 17163 395406
rect 16361 394605 17163 394606
rect 16551 387508 16871 394605
rect 17871 392367 18191 392380
rect 17527 392366 18329 392367
rect 17527 391566 17528 392366
rect 18328 391566 18329 392366
rect 17527 391565 18329 391566
rect 17871 388952 18191 391565
rect 40386 386091 40446 429241
rect 40575 428714 40641 428715
rect 40575 428650 40576 428714
rect 40640 428650 40641 428714
rect 40575 428649 40641 428650
rect 40578 386091 40638 428649
rect 40959 428122 41025 428123
rect 40959 428058 40960 428122
rect 41024 428058 41025 428122
rect 40959 428057 41025 428058
rect 40767 427086 40833 427087
rect 40767 427022 40768 427086
rect 40832 427022 40833 427086
rect 40767 427021 40833 427022
rect 40770 398819 40830 427021
rect 40962 400151 41022 428057
rect 41343 426494 41409 426495
rect 41343 426430 41344 426494
rect 41408 426430 41409 426494
rect 41343 426429 41409 426430
rect 41151 424866 41217 424867
rect 41151 424802 41152 424866
rect 41216 424802 41217 424866
rect 41151 424801 41217 424802
rect 40959 400150 41025 400151
rect 40959 400086 40960 400150
rect 41024 400086 41025 400150
rect 40959 400085 41025 400086
rect 41154 399559 41214 424801
rect 41346 401927 41406 426429
rect 41535 426050 41601 426051
rect 41535 425986 41536 426050
rect 41600 425986 41601 426050
rect 41535 425985 41601 425986
rect 41538 406071 41598 425985
rect 41535 406070 41601 406071
rect 41535 406006 41536 406070
rect 41600 406006 41601 406070
rect 41535 406005 41601 406006
rect 41730 404443 41790 531657
rect 41922 405183 41982 531805
rect 42111 424422 42177 424423
rect 42111 424358 42112 424422
rect 42176 424358 42177 424422
rect 42111 424357 42177 424358
rect 41919 405182 41985 405183
rect 41919 405118 41920 405182
rect 41984 405118 41985 405182
rect 41919 405117 41985 405118
rect 41727 404442 41793 404443
rect 41727 404378 41728 404442
rect 41792 404378 41793 404442
rect 41727 404377 41793 404378
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40767 398818 40833 398819
rect 40767 398754 40768 398818
rect 40832 398754 40833 398818
rect 40767 398753 40833 398754
rect 40383 386090 40449 386091
rect 40383 386026 40384 386090
rect 40448 386026 40449 386090
rect 40383 386025 40449 386026
rect 40575 386090 40641 386091
rect 40575 386026 40576 386090
rect 40640 386026 40641 386090
rect 40575 386025 40641 386026
rect 8927 353101 9247 353182
rect 8635 353100 9437 353101
rect 8635 352300 8636 353100
rect 9436 352300 9437 353100
rect 8635 352299 9437 352300
rect 7607 350889 7927 350982
rect 7235 350888 8037 350889
rect 7235 350088 7236 350888
rect 8036 350088 8037 350888
rect 7235 350087 8037 350088
rect 7607 344818 7927 350087
rect 8927 343816 9247 352299
rect 16347 352038 17149 352039
rect 16347 351238 16348 352038
rect 17148 351238 17149 352038
rect 16347 351237 17149 351238
rect 16551 344484 16871 351237
rect 17871 349387 18191 349404
rect 17547 349386 18349 349387
rect 17547 348586 17548 349386
rect 18348 348586 18349 349386
rect 17547 348585 18349 348586
rect 17871 345484 18191 348585
rect 40386 343023 40446 386025
rect 40383 343022 40449 343023
rect 40383 342958 40384 343022
rect 40448 342958 40449 343022
rect 40383 342957 40449 342958
rect 31982 331648 32638 331686
rect 31982 330486 32020 331648
rect 32604 330486 32638 331648
rect 31982 330460 32638 330486
rect 8927 309937 9247 309952
rect 8737 309936 9539 309937
rect 8737 309136 8738 309936
rect 9538 309136 9539 309936
rect 8737 309135 9539 309136
rect 7607 307137 7927 307234
rect 7377 307136 8179 307137
rect 7377 306336 7378 307136
rect 8178 306336 8179 307136
rect 7377 306335 8179 306336
rect 7607 301518 7927 306335
rect 8927 300664 9247 309135
rect 16551 308799 16871 308812
rect 16327 308798 17129 308799
rect 16327 307998 16328 308798
rect 17128 307998 17129 308798
rect 16327 307997 17129 307998
rect 16551 300772 16871 307997
rect 17871 305649 18191 305698
rect 17731 305648 18533 305649
rect 17731 304848 17732 305648
rect 18532 304848 18533 305648
rect 17731 304847 18533 304848
rect 17871 302308 18191 304847
rect 40386 299807 40446 342957
rect 40578 342875 40638 386025
rect 40959 384906 41025 384907
rect 40959 384842 40960 384906
rect 41024 384842 41025 384906
rect 40959 384841 41025 384842
rect 40767 383870 40833 383871
rect 40767 383806 40768 383870
rect 40832 383806 40833 383870
rect 40767 383805 40833 383806
rect 40770 355603 40830 383805
rect 40962 356935 41022 384841
rect 41343 383278 41409 383279
rect 41343 383214 41344 383278
rect 41408 383214 41409 383278
rect 41343 383213 41409 383214
rect 41151 381650 41217 381651
rect 41151 381586 41152 381650
rect 41216 381586 41217 381650
rect 41151 381585 41217 381586
rect 40959 356934 41025 356935
rect 40959 356870 40960 356934
rect 41024 356870 41025 356934
rect 40959 356869 41025 356870
rect 41154 356491 41214 381585
rect 41346 358711 41406 383213
rect 41535 382834 41601 382835
rect 41535 382770 41536 382834
rect 41600 382770 41601 382834
rect 41535 382769 41601 382770
rect 41538 362855 41598 382769
rect 41535 362854 41601 362855
rect 41535 362790 41536 362854
rect 41600 362790 41601 362854
rect 41535 362789 41601 362790
rect 41730 360635 41790 404377
rect 41922 360931 41982 405117
rect 42114 402667 42174 424357
rect 42303 423978 42369 423979
rect 42303 423914 42304 423978
rect 42368 423914 42369 423978
rect 42303 423913 42369 423914
rect 42306 403111 42366 423913
rect 42303 403110 42369 403111
rect 42303 403046 42304 403110
rect 42368 403046 42369 403110
rect 42303 403045 42369 403046
rect 42111 402666 42177 402667
rect 42111 402602 42112 402666
rect 42176 402602 42177 402666
rect 42111 402601 42177 402602
rect 42111 375138 42177 375139
rect 42111 375074 42112 375138
rect 42176 375074 42177 375138
rect 42111 375073 42177 375074
rect 41919 360930 41985 360931
rect 41919 360866 41920 360930
rect 41984 360866 41985 360930
rect 41919 360865 41985 360866
rect 41727 360634 41793 360635
rect 41727 360570 41728 360634
rect 41792 360570 41793 360634
rect 41727 360569 41793 360570
rect 42114 359451 42174 375073
rect 42303 372918 42369 372919
rect 42303 372854 42304 372918
rect 42368 372854 42369 372918
rect 42303 372853 42369 372854
rect 42306 359895 42366 372853
rect 42495 360930 42561 360931
rect 42495 360866 42496 360930
rect 42560 360866 42561 360930
rect 42495 360865 42561 360866
rect 42303 359894 42369 359895
rect 42303 359830 42304 359894
rect 42368 359830 42369 359894
rect 42303 359829 42369 359830
rect 42111 359450 42177 359451
rect 42111 359386 42112 359450
rect 42176 359386 42177 359450
rect 42111 359385 42177 359386
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40767 355602 40833 355603
rect 40767 355538 40768 355602
rect 40832 355538 40833 355602
rect 40767 355537 40833 355538
rect 40575 342874 40641 342875
rect 40575 342810 40576 342874
rect 40640 342810 40641 342874
rect 40575 342809 40641 342810
rect 40383 299806 40449 299807
rect 40383 299742 40384 299806
rect 40448 299742 40449 299806
rect 40383 299741 40449 299742
rect 36324 287744 37012 287818
rect 36324 286660 36346 287744
rect 36976 286660 37012 287744
rect 36324 286598 37012 286660
rect 8927 267361 9247 267494
rect 8583 267360 9385 267361
rect 8583 266560 8584 267360
rect 9384 266560 9385 267360
rect 8583 266559 9385 266560
rect 7607 264017 7927 264128
rect 7373 264016 8175 264017
rect 7373 263216 7374 264016
rect 8174 263216 8175 264016
rect 7373 263215 8175 263216
rect 7607 258584 7927 263215
rect 8927 257116 9247 266559
rect 16353 265912 17155 265913
rect 16353 265112 16354 265912
rect 17154 265112 17155 265912
rect 16353 265111 17155 265112
rect 16551 257460 16871 265111
rect 17561 262122 18363 262123
rect 17561 261322 17562 262122
rect 18362 261322 18363 262122
rect 17561 261321 18363 261322
rect 17871 258324 18191 261321
rect 40386 257035 40446 299741
rect 40578 299659 40638 342809
rect 40767 341838 40833 341839
rect 40767 341774 40768 341838
rect 40832 341774 40833 341838
rect 40767 341773 40833 341774
rect 40770 313719 40830 341773
rect 40959 340654 41025 340655
rect 40959 340590 40960 340654
rect 41024 340590 41025 340654
rect 40959 340589 41025 340590
rect 40767 313718 40833 313719
rect 40767 313654 40768 313718
rect 40832 313654 40833 313718
rect 40767 313653 40833 313654
rect 40962 312387 41022 340589
rect 41343 340210 41409 340211
rect 41343 340146 41344 340210
rect 41408 340146 41409 340210
rect 41343 340145 41409 340146
rect 41151 338582 41217 338583
rect 41151 338518 41152 338582
rect 41216 338518 41217 338582
rect 41151 338517 41217 338518
rect 41154 313275 41214 338517
rect 41346 315495 41406 340145
rect 41535 339618 41601 339619
rect 41535 339554 41536 339618
rect 41600 339554 41601 339618
rect 41535 339553 41601 339554
rect 41538 319787 41598 339553
rect 42498 339027 42558 360865
rect 42687 360634 42753 360635
rect 42687 360570 42688 360634
rect 42752 360570 42753 360634
rect 42687 360569 42753 360570
rect 42495 339026 42561 339027
rect 42495 338962 42496 339026
rect 42560 338962 42561 339026
rect 42495 338961 42561 338962
rect 42690 338691 42750 360569
rect 42879 339026 42945 339027
rect 42879 338962 42880 339026
rect 42944 338962 42945 339026
rect 42879 338961 42945 338962
rect 42114 338631 42750 338691
rect 41919 322598 41985 322599
rect 41919 322534 41920 322598
rect 41984 322534 41985 322598
rect 41919 322533 41985 322534
rect 41535 319786 41601 319787
rect 41535 319722 41536 319786
rect 41600 319722 41601 319786
rect 41535 319721 41601 319722
rect 41922 318751 41982 322533
rect 41919 318750 41985 318751
rect 41919 318711 41920 318750
rect 41730 318686 41920 318711
rect 41984 318686 41985 318750
rect 41730 318685 41985 318686
rect 41730 318651 41982 318685
rect 41343 315494 41409 315495
rect 41343 315430 41344 315494
rect 41408 315430 41409 315494
rect 41343 315429 41409 315430
rect 41151 313274 41217 313275
rect 41151 313210 41152 313274
rect 41216 313210 41217 313274
rect 41151 313209 41217 313210
rect 40959 312386 41025 312387
rect 40959 312322 40960 312386
rect 41024 312322 41025 312386
rect 40959 312321 41025 312322
rect 40575 299658 40641 299659
rect 40575 299594 40576 299658
rect 40640 299594 40641 299658
rect 40575 299593 40641 299594
rect 40767 298622 40833 298623
rect 40767 298558 40768 298622
rect 40832 298558 40833 298622
rect 40767 298557 40833 298558
rect 40770 270651 40830 298557
rect 40959 297438 41025 297439
rect 40959 297374 40960 297438
rect 41024 297374 41025 297438
rect 40959 297373 41025 297374
rect 40767 270650 40833 270651
rect 40767 270586 40768 270650
rect 40832 270586 40833 270650
rect 40767 270585 40833 270586
rect 40962 269171 41022 297373
rect 41343 296994 41409 296995
rect 41343 296930 41344 296994
rect 41408 296930 41409 296994
rect 41343 296929 41409 296930
rect 41151 295366 41217 295367
rect 41151 295302 41152 295366
rect 41216 295302 41217 295366
rect 41151 295301 41217 295302
rect 41154 270059 41214 295301
rect 41346 272279 41406 296929
rect 41535 296550 41601 296551
rect 41535 296486 41536 296550
rect 41600 296486 41601 296550
rect 41535 296485 41601 296486
rect 41538 276571 41598 296485
rect 41730 285411 41790 318651
rect 42114 318045 42174 338631
rect 42303 329850 42369 329851
rect 42303 329786 42304 329850
rect 42368 329786 42369 329850
rect 42303 329785 42369 329786
rect 41922 317985 42174 318045
rect 41922 317863 41982 317985
rect 41919 317862 41985 317863
rect 41919 317798 41920 317862
rect 41984 317798 41985 317862
rect 41919 317797 41985 317798
rect 41922 285599 41982 317797
rect 42111 317122 42177 317123
rect 42111 317058 42112 317122
rect 42176 317058 42177 317122
rect 42111 317057 42177 317058
rect 42114 316087 42174 317057
rect 42306 316679 42366 329785
rect 42495 326594 42561 326595
rect 42495 326530 42496 326594
rect 42560 326530 42561 326594
rect 42495 326529 42561 326530
rect 42498 320971 42558 326529
rect 42882 322599 42942 338961
rect 43071 338286 43137 338287
rect 43071 338222 43072 338286
rect 43136 338222 43137 338286
rect 43071 338221 43137 338222
rect 42879 322598 42945 322599
rect 42879 322534 42880 322598
rect 42944 322534 42945 322598
rect 42879 322533 42945 322534
rect 42495 320970 42561 320971
rect 42495 320906 42496 320970
rect 42560 320906 42561 320970
rect 42495 320905 42561 320906
rect 43074 317123 43134 338221
rect 43071 317122 43137 317123
rect 43071 317058 43072 317122
rect 43136 317058 43137 317122
rect 43071 317057 43137 317058
rect 42303 316678 42369 316679
rect 42303 316614 42304 316678
rect 42368 316614 42369 316678
rect 42303 316613 42369 316614
rect 42111 316086 42177 316087
rect 42111 316022 42112 316086
rect 42176 316022 42177 316086
rect 42111 316021 42177 316022
rect 42303 299658 42369 299659
rect 42303 299594 42304 299658
rect 42368 299594 42369 299658
rect 42303 299593 42369 299594
rect 42111 294922 42177 294923
rect 42111 294858 42112 294922
rect 42176 294858 42177 294922
rect 42111 294857 42177 294858
rect 41919 285598 41985 285599
rect 41919 285534 41920 285598
rect 41984 285534 41985 285598
rect 41919 285533 41985 285534
rect 41730 285351 41982 285411
rect 41727 285154 41793 285155
rect 41727 285090 41728 285154
rect 41792 285090 41793 285154
rect 41727 285089 41793 285090
rect 41535 276570 41601 276571
rect 41535 276506 41536 276570
rect 41600 276506 41601 276570
rect 41535 276505 41601 276506
rect 41730 273611 41790 285089
rect 41922 275535 41982 285351
rect 41919 275534 41985 275535
rect 41919 275470 41920 275534
rect 41984 275470 41985 275534
rect 41919 275469 41985 275470
rect 41727 273610 41793 273611
rect 41727 273546 41728 273610
rect 41792 273546 41793 273610
rect 41727 273545 41793 273546
rect 41343 272278 41409 272279
rect 41343 272214 41344 272278
rect 41408 272214 41409 272278
rect 41343 272213 41409 272214
rect 41922 270651 41982 275469
rect 42114 273019 42174 294857
rect 42111 273018 42177 273019
rect 42111 272954 42112 273018
rect 42176 272954 42177 273018
rect 42111 272953 42177 272954
rect 41919 270650 41985 270651
rect 41919 270586 41920 270650
rect 41984 270586 41985 270650
rect 41919 270585 41985 270586
rect 41151 270058 41217 270059
rect 41151 269994 41152 270058
rect 41216 269994 41217 270058
rect 41151 269993 41217 269994
rect 40959 269170 41025 269171
rect 40959 269106 40960 269170
rect 41024 269106 41025 269170
rect 40959 269105 41025 269106
rect 40383 257034 40449 257035
rect 40383 256970 40384 257034
rect 40448 256970 40449 257034
rect 40383 256969 40449 256970
rect 42306 255999 42366 299593
rect 42687 293442 42753 293443
rect 42687 293378 42688 293442
rect 42752 293378 42753 293442
rect 42687 293377 42753 293378
rect 42495 285598 42561 285599
rect 42495 285534 42496 285598
rect 42560 285534 42561 285598
rect 42495 285533 42561 285534
rect 42498 274795 42558 285533
rect 42690 278051 42750 293377
rect 42687 278050 42753 278051
rect 42687 277986 42688 278050
rect 42752 277986 42753 278050
rect 42687 277985 42753 277986
rect 43272 277114 44476 706576
rect 43272 275482 43906 277114
rect 44432 275482 44476 277114
rect 42495 274794 42561 274795
rect 42495 274730 42496 274794
rect 42560 274730 42561 274794
rect 42495 274729 42561 274730
rect 42879 270650 42945 270651
rect 42879 270586 42880 270650
rect 42944 270586 42945 270650
rect 42879 270585 42945 270586
rect 42303 255998 42369 255999
rect 42303 255934 42304 255998
rect 42368 255934 42369 255998
rect 42303 255933 42369 255934
rect 40575 255406 40641 255407
rect 40575 255342 40576 255406
rect 40640 255342 40641 255406
rect 40575 255341 40641 255342
rect 40383 254222 40449 254223
rect 40383 254158 40384 254222
rect 40448 254158 40449 254222
rect 40383 254157 40449 254158
rect 40386 225955 40446 254157
rect 40578 227287 40638 255341
rect 40767 253778 40833 253779
rect 40767 253714 40768 253778
rect 40832 253714 40833 253778
rect 40767 253713 40833 253714
rect 40770 229063 40830 253713
rect 41151 253334 41217 253335
rect 41151 253270 41152 253334
rect 41216 253270 41217 253334
rect 41151 253269 41217 253270
rect 40959 252150 41025 252151
rect 40959 252086 40960 252150
rect 41024 252086 41025 252150
rect 40959 252085 41025 252086
rect 40767 229062 40833 229063
rect 40767 228998 40768 229062
rect 40832 228998 40833 229062
rect 40767 228997 40833 228998
rect 40575 227286 40641 227287
rect 40575 227222 40576 227286
rect 40640 227222 40641 227286
rect 40575 227221 40641 227222
rect 40962 226695 41022 252085
rect 41154 233355 41214 253269
rect 41343 251706 41409 251707
rect 41343 251642 41344 251706
rect 41408 251642 41409 251706
rect 41343 251641 41409 251642
rect 41151 233354 41217 233355
rect 41151 233290 41152 233354
rect 41216 233290 41217 233354
rect 41151 233289 41217 233290
rect 41346 229803 41406 251641
rect 42882 246823 42942 270585
rect 43272 266848 44476 275482
rect 44866 331636 45466 828210
rect 46142 497400 46742 988556
rect 47232 986974 49272 987022
rect 47232 985814 47268 986974
rect 49228 985814 49272 986974
rect 47232 985786 49272 985814
rect 45902 497304 46764 497400
rect 45902 483786 45974 497304
rect 46716 483786 46764 497304
rect 45902 483666 46764 483786
rect 44866 330504 44906 331636
rect 45450 330504 45466 331636
rect 44866 267378 45466 330504
rect 46142 287742 46742 483666
rect 47244 454802 49272 985786
rect 47140 454744 49272 454802
rect 47140 441662 47166 454744
rect 49188 441662 49272 454744
rect 47140 441590 49272 441662
rect 46142 286664 46158 287742
rect 46718 286664 46742 287742
rect 46142 268394 46742 286664
rect 47244 275590 49272 441590
rect 47196 275552 49272 275590
rect 47196 269828 47242 275552
rect 49208 269828 49272 275552
rect 47196 269792 49272 269828
rect 47244 269762 49272 269792
rect 49632 952831 51436 992148
rect 49632 952033 50127 952831
rect 50925 952033 51436 952831
rect 49632 826519 51436 952033
rect 49632 825721 50127 826519
rect 50925 825721 51436 826519
rect 49632 783775 51436 825721
rect 49632 782977 50127 783775
rect 50925 782977 51436 783775
rect 49632 740587 51436 782977
rect 49632 739789 50127 740587
rect 50925 739789 51436 740587
rect 49632 697141 51436 739789
rect 49632 696343 50127 697141
rect 50925 696343 51436 697141
rect 49632 653815 51436 696343
rect 49632 653017 50127 653815
rect 50925 653017 51436 653815
rect 49632 610725 51436 653017
rect 49632 609927 50127 610725
rect 50925 609927 51436 610725
rect 49632 567645 51436 609927
rect 49632 566847 50127 567645
rect 50925 566847 51436 567645
rect 49632 439989 51436 566847
rect 49632 439191 50127 439989
rect 50925 439191 51436 439989
rect 49632 396837 51436 439191
rect 49632 396039 50127 396837
rect 50925 396039 51436 396837
rect 49632 353099 51436 396039
rect 49632 352301 50127 353099
rect 50925 352301 51436 353099
rect 49632 309935 51436 352301
rect 49632 309137 50127 309935
rect 50925 309137 51436 309935
rect 44866 266996 44912 267378
rect 45430 266996 45466 267378
rect 44866 266886 45466 266996
rect 49632 267359 51436 309137
rect 43272 266248 43870 266848
rect 44470 266248 44476 266848
rect 43272 266084 44476 266248
rect 49632 266561 50127 267359
rect 50925 266561 51436 267359
rect 49632 265760 51436 266561
rect 51584 951105 52914 993544
rect 51584 950307 51919 951105
rect 52717 950307 52914 951105
rect 51584 825057 52914 950307
rect 51584 824259 51919 825057
rect 52717 824259 52914 825057
rect 51584 782647 52914 824259
rect 51584 781849 51919 782647
rect 52717 781849 52914 782647
rect 51584 739233 52914 781849
rect 51584 738435 51919 739233
rect 52717 738435 52914 739233
rect 51584 695867 52914 738435
rect 51584 695069 51919 695867
rect 52717 695069 52914 695867
rect 51584 652619 52914 695069
rect 51584 651821 51919 652619
rect 52717 651821 52914 652619
rect 51584 609445 52914 651821
rect 51584 608647 51919 609445
rect 52717 608647 52914 609445
rect 51584 566543 52914 608647
rect 51584 565745 51919 566543
rect 52717 565745 52914 566543
rect 51584 438623 52914 565745
rect 51584 437825 51919 438623
rect 52717 437825 52914 438623
rect 51584 395405 52914 437825
rect 51584 394607 51919 395405
rect 52717 394607 52914 395405
rect 51584 352037 52914 394607
rect 51584 351239 51919 352037
rect 52717 351239 52914 352037
rect 51584 308797 52914 351239
rect 51584 307999 51919 308797
rect 52717 307999 52914 308797
rect 51584 265911 52914 307999
rect 48980 265720 51440 265760
rect 48980 265646 49020 265720
rect 43258 262254 49020 265646
rect 51400 262254 51440 265720
rect 43258 262214 51440 262254
rect 51584 265113 51919 265911
rect 52717 265113 52914 265911
rect 43258 262212 51436 262214
rect 42879 246822 42945 246823
rect 42879 246758 42880 246822
rect 42944 246758 42945 246822
rect 42879 246757 42945 246758
rect 42882 245047 42942 246757
rect 41535 245046 41601 245047
rect 41535 244982 41536 245046
rect 41600 244982 41601 245046
rect 41535 244981 41601 244982
rect 42879 245046 42945 245047
rect 42879 244982 42880 245046
rect 42944 244982 42945 245046
rect 42879 244981 42945 244982
rect 41538 231727 41598 244981
rect 41727 244898 41793 244899
rect 41727 244834 41728 244898
rect 41792 244834 41793 244898
rect 41727 244833 41793 244834
rect 41535 231726 41601 231727
rect 41535 231662 41536 231726
rect 41600 231662 41601 231726
rect 41535 231661 41601 231662
rect 41538 230133 41598 231661
rect 41730 230395 41790 244833
rect 41919 243862 41985 243863
rect 41919 243798 41920 243862
rect 41984 243798 41985 243862
rect 41919 243797 41985 243798
rect 41922 231135 41982 243797
rect 43258 241906 45132 262212
rect 49632 262190 51436 262212
rect 51584 261564 52914 265113
rect 45498 259733 52914 261564
rect 53092 949281 54534 994938
rect 53092 948483 53703 949281
rect 54501 948483 54534 949281
rect 53092 823499 54534 948483
rect 53092 822701 53703 823499
rect 54501 822701 54534 823499
rect 53092 781239 54534 822701
rect 53092 780441 53703 781239
rect 54501 780441 54534 781239
rect 53092 737831 54534 780441
rect 53092 737033 53703 737831
rect 54501 737033 54534 737831
rect 53092 694753 54534 737033
rect 53092 693955 53703 694753
rect 54501 693955 54534 694753
rect 53092 651515 54534 693955
rect 53092 650717 53703 651515
rect 54501 650717 54534 651515
rect 53092 607891 54534 650717
rect 53092 607093 53703 607891
rect 54501 607093 54534 607891
rect 53092 565273 54534 607093
rect 53092 564475 53703 565273
rect 54501 564475 54534 565273
rect 53092 437095 54534 564475
rect 53092 436297 53703 437095
rect 54501 436297 54534 437095
rect 53092 393885 54534 436297
rect 53092 393087 53703 393885
rect 54501 393087 54534 393885
rect 53092 350887 54534 393087
rect 53092 350089 53703 350887
rect 54501 350089 54534 350887
rect 53092 307135 54534 350089
rect 53092 306337 53703 307135
rect 54501 306337 54534 307135
rect 53092 264015 54534 306337
rect 53092 263217 53703 264015
rect 54501 263217 54534 264015
rect 45498 259724 52908 259733
rect 45504 259702 52718 259724
rect 45504 248530 47748 259702
rect 53092 259488 54534 263217
rect 48222 259448 54534 259488
rect 48222 256860 48262 259448
rect 54378 259316 54534 259448
rect 54692 947745 56068 996198
rect 61432 984246 62032 996908
rect 121358 992918 121958 996961
rect 122816 997035 122817 997633
rect 123415 997035 123416 997633
rect 122816 994298 123416 997035
rect 124006 997605 124606 997606
rect 124006 997007 124007 997605
rect 124605 997007 124606 997605
rect 124006 995470 124606 997007
rect 125334 997065 125335 997663
rect 125933 997065 125934 997663
rect 125334 996724 125934 997065
rect 125334 996172 125358 996724
rect 125910 996172 125934 996724
rect 125334 996148 125934 996172
rect 173268 997623 173868 997624
rect 173268 997025 173269 997623
rect 173867 997025 173868 997623
rect 378530 997619 379130 997620
rect 377196 997605 377796 997606
rect 332436 997603 333036 997604
rect 277780 997595 278380 997596
rect 228774 997579 229374 997580
rect 124006 994918 124030 995470
rect 124582 994918 124606 995470
rect 124006 994894 124606 994918
rect 122816 993746 122840 994298
rect 123392 993746 123416 994298
rect 122816 993722 123416 993746
rect 121358 992366 121382 992918
rect 121934 992366 121958 992918
rect 121358 992342 121958 992366
rect 173268 992918 173868 997025
rect 174520 997529 175120 997530
rect 174520 996931 174521 997529
rect 175119 996931 175120 997529
rect 227324 997481 227924 997482
rect 174520 994298 175120 996931
rect 176204 997437 176804 997438
rect 176204 996839 176205 997437
rect 176803 996839 176804 997437
rect 176204 995470 176804 996839
rect 177460 997433 178060 997434
rect 177460 996835 177461 997433
rect 178059 996835 178060 997433
rect 177460 996724 178060 996835
rect 177460 996172 177484 996724
rect 178036 996172 178060 996724
rect 177460 996148 178060 996172
rect 223906 997395 224506 997396
rect 223906 996797 223907 997395
rect 224505 996797 224506 997395
rect 176204 994918 176228 995470
rect 176780 994918 176804 995470
rect 176204 994894 176804 994918
rect 174520 993746 174544 994298
rect 175096 993746 175120 994298
rect 174520 993722 175120 993746
rect 173268 992366 173292 992918
rect 173844 992366 173868 992918
rect 173268 992342 173868 992366
rect 223906 992918 224506 996797
rect 225484 997305 226084 997306
rect 225484 996707 225485 997305
rect 226083 996707 226084 997305
rect 225484 994298 226084 996707
rect 227324 996883 227325 997481
rect 227923 996883 227924 997481
rect 227324 995470 227924 996883
rect 228774 996981 228775 997579
rect 229373 996981 229374 997579
rect 276374 997551 276974 997552
rect 228774 996724 229374 996981
rect 228774 996172 228798 996724
rect 229350 996172 229374 996724
rect 228774 996148 229374 996172
rect 274880 997463 275480 997464
rect 274880 996865 274881 997463
rect 275479 996865 275480 997463
rect 227324 994918 227348 995470
rect 227900 994918 227924 995470
rect 227324 994894 227924 994918
rect 225484 993746 225508 994298
rect 226060 993746 226084 994298
rect 225484 993722 226084 993746
rect 223906 992366 223930 992918
rect 224482 992366 224506 992918
rect 223906 992342 224506 992366
rect 274880 992918 275480 996865
rect 276374 996953 276375 997551
rect 276973 996953 276974 997551
rect 276374 994298 276974 996953
rect 277780 996997 277781 997595
rect 278379 996997 278380 997595
rect 277780 995470 278380 996997
rect 278922 997595 279522 997596
rect 278922 996997 278923 997595
rect 279521 996997 279522 997595
rect 327774 997589 328374 997590
rect 298156 997533 298228 997534
rect 298156 997463 298157 997533
rect 298227 997463 298228 997533
rect 298156 997462 298228 997463
rect 278922 996724 279522 996997
rect 298162 996746 298222 997462
rect 327774 996991 327775 997589
rect 328373 996991 328374 997589
rect 330888 997545 331488 997546
rect 278922 996172 278946 996724
rect 279498 996172 279522 996724
rect 298158 996745 298230 996746
rect 298158 996675 298159 996745
rect 298229 996675 298230 996745
rect 298158 996674 298230 996675
rect 298162 996636 298222 996674
rect 278922 996148 279522 996172
rect 277780 994918 277804 995470
rect 278356 994918 278380 995470
rect 277780 994894 278380 994918
rect 276374 993746 276398 994298
rect 276950 993746 276974 994298
rect 276374 993722 276974 993746
rect 274880 992366 274904 992918
rect 275456 992366 275480 992918
rect 274880 992342 275480 992366
rect 327774 992918 328374 996991
rect 329332 997441 329932 997442
rect 329332 996843 329333 997441
rect 329931 996843 329932 997441
rect 329332 994298 329932 996843
rect 330888 996947 330889 997545
rect 331487 996947 331488 997545
rect 330888 995470 331488 996947
rect 332436 997005 332437 997603
rect 333035 997005 333036 997603
rect 332436 996724 333036 997005
rect 332436 996172 332460 996724
rect 333012 996172 333036 996724
rect 332436 996148 333036 996172
rect 377196 997007 377197 997605
rect 377795 997007 377796 997605
rect 330888 994918 330912 995470
rect 331464 994918 331488 995470
rect 330888 994894 331488 994918
rect 329332 993746 329356 994298
rect 329908 993746 329932 994298
rect 329332 993722 329932 993746
rect 327774 992366 327798 992918
rect 328350 992366 328374 992918
rect 327774 992342 328374 992366
rect 377196 992918 377796 997007
rect 378530 997021 378531 997619
rect 379129 997021 379130 997619
rect 381548 997609 382148 997610
rect 378530 994298 379130 997021
rect 380080 997595 380680 997596
rect 380080 996997 380081 997595
rect 380679 996997 380680 997595
rect 380080 995470 380680 996997
rect 381548 997011 381549 997609
rect 382147 997011 382148 997609
rect 571834 997585 572434 997586
rect 496096 997571 496696 997572
rect 415922 997547 416522 997548
rect 414358 997531 414958 997532
rect 381548 996724 382148 997011
rect 381548 996172 381572 996724
rect 382124 996172 382148 996724
rect 381548 996148 382148 996172
rect 410146 997425 410746 997426
rect 410146 996827 410147 997425
rect 410745 996827 410746 997425
rect 380080 994918 380104 995470
rect 380656 994918 380680 995470
rect 380080 994894 380680 994918
rect 378530 993746 378554 994298
rect 379106 993746 379130 994298
rect 378530 993722 379130 993746
rect 377196 992366 377220 992918
rect 377772 992366 377796 992918
rect 377196 992342 377796 992366
rect 410146 992918 410746 996827
rect 412148 997413 412748 997414
rect 412148 996815 412149 997413
rect 412747 996815 412748 997413
rect 412148 994298 412748 996815
rect 414358 996933 414359 997531
rect 414957 996933 414958 997531
rect 414358 995470 414958 996933
rect 415922 996949 415923 997547
rect 416521 996949 416522 997547
rect 494582 997523 495182 997524
rect 415922 996724 416522 996949
rect 415922 996172 415946 996724
rect 416498 996172 416522 996724
rect 415922 996148 416522 996172
rect 491650 997381 492250 997382
rect 491650 996783 491651 997381
rect 492249 996783 492250 997381
rect 476607 996146 476673 996147
rect 476607 996082 476608 996146
rect 476672 996082 476673 996146
rect 476607 996081 476673 996082
rect 476610 995851 476670 996081
rect 476607 995850 476673 995851
rect 476607 995786 476608 995850
rect 476672 995786 476673 995850
rect 476607 995785 476673 995786
rect 414358 994918 414382 995470
rect 414934 994918 414958 995470
rect 414358 994894 414958 994918
rect 412148 993746 412172 994298
rect 412724 993746 412748 994298
rect 412148 993722 412748 993746
rect 410146 992366 410170 992918
rect 410722 992366 410746 992918
rect 410146 992342 410746 992366
rect 491650 992918 492250 996783
rect 493070 997381 493670 997382
rect 493070 996783 493071 997381
rect 493669 996783 493670 997381
rect 493070 994298 493670 996783
rect 494582 996925 494583 997523
rect 495181 996925 495182 997523
rect 494582 995470 495182 996925
rect 496096 996973 496097 997571
rect 496695 996973 496696 997571
rect 570328 997543 570928 997544
rect 496096 996724 496696 996973
rect 496096 996172 496120 996724
rect 496672 996172 496696 996724
rect 496096 996148 496696 996172
rect 568178 997451 568778 997452
rect 568178 996853 568179 997451
rect 568777 996853 568778 997451
rect 494582 994918 494606 995470
rect 495158 994918 495182 995470
rect 494582 994894 495182 994918
rect 493070 993746 493094 994298
rect 493646 993746 493670 994298
rect 493070 993722 493670 993746
rect 491650 992366 491674 992918
rect 492226 992366 492250 992918
rect 491650 992342 492250 992366
rect 568178 992918 568778 996853
rect 570328 996945 570329 997543
rect 570927 996945 570928 997543
rect 570328 994298 570928 996945
rect 571834 996987 571835 997585
rect 572433 996987 572434 997585
rect 571834 995470 572434 996987
rect 573446 997527 574046 997528
rect 573446 996929 573447 997527
rect 574045 996929 574046 997527
rect 573446 996724 574046 996929
rect 573446 996172 573470 996724
rect 574022 996172 574046 996724
rect 573446 996148 574046 996172
rect 580184 997096 585702 997132
rect 580184 995988 580186 997096
rect 585676 995988 585702 997096
rect 665024 996748 668306 996837
rect 580184 995918 585702 995988
rect 651552 996686 656548 996746
rect 651552 996024 651576 996686
rect 656490 996024 656548 996686
rect 651552 996022 655360 996024
rect 655902 996022 656548 996024
rect 651552 995984 656548 996022
rect 571834 994918 571858 995470
rect 572410 994918 572434 995470
rect 651568 995030 652168 995122
rect 571834 994894 572434 994918
rect 650536 995000 653634 995030
rect 650536 994470 650578 995000
rect 653584 994470 653634 995000
rect 650536 994440 653634 994470
rect 570328 993746 570352 994298
rect 570904 993746 570928 994298
rect 650628 994094 651228 994098
rect 650256 994084 651292 994094
rect 570328 993722 570928 993746
rect 648658 994070 651292 994084
rect 648658 993536 648716 994070
rect 648658 993472 651292 993536
rect 568178 992366 568202 992918
rect 568754 992366 568778 992918
rect 568178 992342 568778 992366
rect 650628 982236 651228 993472
rect 651568 982290 652168 994440
rect 655328 985376 655928 995984
rect 665024 994456 665102 996748
rect 668240 994456 668306 996748
rect 658682 993126 660572 993138
rect 658682 993070 660610 993126
rect 658682 992298 659386 993070
rect 660564 992298 660610 993070
rect 658682 992280 660610 992298
rect 661102 992954 664196 993397
rect 54692 946947 55269 947745
rect 56067 946947 56068 947745
rect 54692 822225 56068 946947
rect 54692 821427 55269 822225
rect 56067 821427 56068 822225
rect 54692 779783 56068 821427
rect 54692 778985 55269 779783
rect 56067 778985 56068 779783
rect 54692 736149 56068 778985
rect 54692 735351 55269 736149
rect 56067 735351 56068 736149
rect 54692 693083 56068 735351
rect 54692 692285 55269 693083
rect 56067 692285 56068 693083
rect 54692 649949 56068 692285
rect 54692 649151 55269 649949
rect 56067 649151 56068 649949
rect 54692 606155 56068 649151
rect 54692 605357 55269 606155
rect 56067 605357 56068 606155
rect 54692 563821 56068 605357
rect 54692 563023 55269 563821
rect 56067 563023 56068 563821
rect 54692 435747 56068 563023
rect 54692 434949 55269 435747
rect 56067 434949 56068 435747
rect 54692 392365 56068 434949
rect 54692 391567 55269 392365
rect 56067 391567 56068 392365
rect 54692 349385 56068 391567
rect 54692 348587 55269 349385
rect 56067 348587 56068 349385
rect 54692 305647 56068 348587
rect 54692 304849 55269 305647
rect 56067 304849 56068 305647
rect 54692 262121 56068 304849
rect 658682 945491 660572 992280
rect 658682 944309 659369 945491
rect 660551 944309 660572 945491
rect 658682 766959 660572 944309
rect 658682 765777 659369 766959
rect 660551 765777 660572 766959
rect 658682 721281 660572 765777
rect 658682 720099 659369 721281
rect 660551 720099 660572 721281
rect 658682 677243 660572 720099
rect 658682 676061 659369 677243
rect 660551 676061 660572 677243
rect 658682 630015 660572 676061
rect 658682 628833 659369 630015
rect 660551 628833 660572 630015
rect 658682 585085 660572 628833
rect 658682 583903 659369 585085
rect 660551 583903 660572 585085
rect 658682 541881 660572 583903
rect 658682 540699 659369 541881
rect 660551 540699 660572 541881
rect 658682 497499 660572 540699
rect 658682 496317 659369 497499
rect 660551 496317 660572 497499
rect 658682 409431 660572 496317
rect 658682 408249 659369 409431
rect 660551 408249 660572 409431
rect 658682 364311 660572 408249
rect 658682 363129 659369 364311
rect 660551 363129 660572 364311
rect 658682 318185 660572 363129
rect 658682 317003 659369 318185
rect 660551 317003 660572 318185
rect 56732 267352 57332 272482
rect 57672 268876 58272 273540
rect 60492 270646 61092 277178
rect 59062 270606 61094 270646
rect 59062 270210 59102 270606
rect 61054 270210 61094 270606
rect 59062 270170 61094 270210
rect 57648 268836 59514 268876
rect 57648 267890 57688 268836
rect 59474 267890 59514 268836
rect 57648 267850 59514 267890
rect 56332 267312 58946 267352
rect 56332 267052 56474 267312
rect 58874 267052 58946 267312
rect 56332 267028 58946 267052
rect 56732 266994 57332 267028
rect 61432 266700 62032 277168
rect 374463 273610 374529 273611
rect 374463 273546 374464 273610
rect 374528 273546 374529 273610
rect 374463 273545 374529 273546
rect 374466 273019 374526 273545
rect 409407 273462 409473 273463
rect 409407 273398 409408 273462
rect 409472 273398 409473 273462
rect 409407 273397 409473 273398
rect 384063 273314 384129 273315
rect 384063 273250 384064 273314
rect 384128 273250 384129 273314
rect 384063 273249 384129 273250
rect 374463 273018 374529 273019
rect 374463 272954 374464 273018
rect 374528 272954 374529 273018
rect 374463 272953 374529 272954
rect 135231 272574 135297 272575
rect 135231 272510 135232 272574
rect 135296 272510 135297 272574
rect 135231 272509 135297 272510
rect 135234 270799 135294 272509
rect 378303 272130 378369 272131
rect 378303 272066 378304 272130
rect 378368 272066 378369 272130
rect 378303 272065 378369 272066
rect 378306 271425 378366 272065
rect 377922 271365 378366 271425
rect 377922 271243 377982 271365
rect 377919 271242 377985 271243
rect 377919 271178 377920 271242
rect 377984 271178 377985 271242
rect 377919 271177 377985 271178
rect 348543 270946 348609 270947
rect 348543 270882 348544 270946
rect 348608 270882 348609 270946
rect 348543 270881 348609 270882
rect 135231 270798 135297 270799
rect 135231 270734 135232 270798
rect 135296 270734 135297 270798
rect 135231 270733 135297 270734
rect 208870 270248 210654 270428
rect 60436 266660 62802 266700
rect 60436 266096 60476 266660
rect 62762 266096 62802 266660
rect 60436 266056 62802 266096
rect 54692 261323 55269 262121
rect 56067 262000 56068 262121
rect 181802 265614 193604 269723
rect 56067 261323 56082 262000
rect 54692 260586 56082 261323
rect 181802 261204 181826 265614
rect 193584 261204 193604 265614
rect 54378 257056 54550 259316
rect 54378 256860 54418 257056
rect 48222 256820 54418 256860
rect 45496 248490 47796 248530
rect 45496 247160 45536 248490
rect 45480 247120 45536 247160
rect 45480 244696 45520 247120
rect 45480 244656 45536 244696
rect 45496 244520 45536 244656
rect 47756 244520 47796 248490
rect 45496 244480 47796 244520
rect 45504 241982 47748 244480
rect 45504 241906 47850 241982
rect 42490 239682 45168 241906
rect 42490 239410 45170 239682
rect 42490 239408 43732 239410
rect 42490 239398 43722 239408
rect 42490 239366 43714 239398
rect 44458 239366 45170 239410
rect 42303 238386 42369 238387
rect 42303 238322 42304 238386
rect 42368 238322 42369 238386
rect 42303 238321 42369 238322
rect 42306 234095 42366 238321
rect 42490 237972 42530 239366
rect 45096 237972 45170 239366
rect 42490 237844 45170 237972
rect 42303 234094 42369 234095
rect 42303 234030 42304 234094
rect 42368 234030 42369 234094
rect 42303 234029 42369 234030
rect 41919 231134 41985 231135
rect 41919 231070 41920 231134
rect 41984 231070 41985 231134
rect 41919 231069 41985 231070
rect 41727 230394 41793 230395
rect 41727 230330 41728 230394
rect 41792 230330 41793 230394
rect 41727 230329 41793 230330
rect 41538 230073 41790 230133
rect 41343 229802 41409 229803
rect 41343 229738 41344 229802
rect 41408 229738 41409 229802
rect 41343 229737 41409 229738
rect 40959 226694 41025 226695
rect 40959 226630 40960 226694
rect 41024 226630 41025 226694
rect 40959 226629 41025 226630
rect 40383 225954 40449 225955
rect 40383 225890 40384 225954
rect 40448 225890 40449 225954
rect 40383 225889 40449 225890
rect 8927 223885 9247 223996
rect 8729 223884 9531 223885
rect 8729 223084 8730 223884
rect 9530 223084 9531 223884
rect 8729 223083 9531 223084
rect 7607 221531 7927 221604
rect 7363 221530 8165 221531
rect 7363 220730 7364 221530
rect 8164 220730 8165 221530
rect 7363 220729 8165 220730
rect 7607 214832 7927 220729
rect 8927 213678 9247 223083
rect 16551 222741 16871 222928
rect 16291 222740 17093 222741
rect 16291 221940 16292 222740
rect 17092 221940 17093 222740
rect 16291 221939 17093 221940
rect 16551 214276 16871 221939
rect 17871 220257 18191 220322
rect 17701 220256 18503 220257
rect 17701 219456 17702 220256
rect 18502 219456 18503 220256
rect 17701 219455 18503 219456
rect 17871 215430 18191 219455
rect 40575 212190 40641 212191
rect 40575 212126 40576 212190
rect 40640 212126 40641 212190
rect 40575 212125 40641 212126
rect 40383 211154 40449 211155
rect 40383 211090 40384 211154
rect 40448 211090 40449 211154
rect 40383 211089 40449 211090
rect 40386 182887 40446 211089
rect 40578 184219 40638 212125
rect 40959 210562 41025 210563
rect 40959 210498 40960 210562
rect 41024 210498 41025 210562
rect 40959 210497 41025 210498
rect 40767 208934 40833 208935
rect 40767 208870 40768 208934
rect 40832 208870 40833 208934
rect 40767 208869 40833 208870
rect 40575 184218 40641 184219
rect 40575 184154 40576 184218
rect 40640 184154 40641 184218
rect 40575 184153 40641 184154
rect 40770 183627 40830 208869
rect 40962 185847 41022 210497
rect 41535 209970 41601 209971
rect 41535 209906 41536 209970
rect 41600 209906 41601 209970
rect 41535 209905 41601 209906
rect 41151 208342 41217 208343
rect 41151 208278 41152 208342
rect 41216 208278 41217 208342
rect 41151 208277 41217 208278
rect 41154 186439 41214 208277
rect 41343 207898 41409 207899
rect 41343 207834 41344 207898
rect 41408 207834 41409 207898
rect 41343 207833 41409 207834
rect 41346 187179 41406 207833
rect 41538 190139 41598 209905
rect 41535 190138 41601 190139
rect 41535 190074 41536 190138
rect 41600 190074 41601 190138
rect 41535 190073 41601 190074
rect 41730 189103 41790 230073
rect 41727 189102 41793 189103
rect 41727 189038 41728 189102
rect 41792 189038 41793 189102
rect 41727 189037 41793 189038
rect 41922 188363 41982 231069
rect 42490 229356 45168 237844
rect 45562 234028 47850 241906
rect 45548 233890 47850 234028
rect 45548 232804 45600 233890
rect 47800 232804 47850 233890
rect 45548 232682 47850 232804
rect 42462 229100 45168 229356
rect 42458 229084 45168 229100
rect 42458 229082 43698 229084
rect 42458 229072 43688 229082
rect 42458 229040 43680 229072
rect 44424 229040 45168 229084
rect 42458 227646 42496 229040
rect 45062 227646 45168 229040
rect 42458 227562 45168 227646
rect 42462 227518 45168 227562
rect 42490 223883 45168 227518
rect 45562 224106 47850 232682
rect 42490 223085 43691 223883
rect 44489 223085 45168 223883
rect 42490 219030 45168 223085
rect 45536 223968 47850 224106
rect 45536 222882 45588 223968
rect 47788 222882 47850 223968
rect 45536 222760 47850 222882
rect 42484 218774 45168 219030
rect 42480 218758 45168 218774
rect 42480 218756 43720 218758
rect 42480 218746 43710 218756
rect 42480 218714 43702 218746
rect 44446 218714 45168 218758
rect 42480 217320 42518 218714
rect 45084 217320 45168 218714
rect 42480 217236 45168 217320
rect 42484 217192 45168 217236
rect 42490 209350 45168 217192
rect 45562 222739 47850 222760
rect 45562 221941 46937 222739
rect 47735 221941 47850 222739
rect 45562 214028 47850 221941
rect 48226 221529 50152 256820
rect 54692 256322 56068 260586
rect 50528 256282 56090 256322
rect 50528 253286 50568 256282
rect 56050 253286 56090 256282
rect 50528 253246 56090 253286
rect 48226 220731 48719 221529
rect 49517 220731 50152 221529
rect 48226 220042 50152 220731
rect 50570 220255 52270 253246
rect 145407 242086 145473 242087
rect 145407 242022 145408 242086
rect 145472 242022 145473 242086
rect 145407 242021 145473 242022
rect 50570 219457 50603 220255
rect 51401 219457 52270 220255
rect 50570 219272 52270 219457
rect 45562 213990 47858 214028
rect 45562 212904 45614 213990
rect 47814 212904 47858 213990
rect 45562 212842 47858 212904
rect 42490 209078 45182 209350
rect 42490 209076 43744 209078
rect 42490 209066 43734 209076
rect 42490 209034 43726 209066
rect 44470 209034 45182 209078
rect 42490 207640 42542 209034
rect 45108 207640 45182 209034
rect 42490 207512 45182 207640
rect 42490 199410 45168 207512
rect 42486 199154 45168 199410
rect 42482 199138 45168 199154
rect 42482 199136 43722 199138
rect 42482 199126 43712 199136
rect 42482 199094 43704 199126
rect 44448 199094 45168 199138
rect 42482 197700 42520 199094
rect 45086 197700 45168 199094
rect 42111 197686 42177 197687
rect 42111 197622 42112 197686
rect 42176 197622 42177 197686
rect 42111 197621 42177 197622
rect 42114 191027 42174 197621
rect 42482 197616 45168 197700
rect 42486 197572 45168 197616
rect 42111 191026 42177 191027
rect 42111 190962 42112 191026
rect 42176 190962 42177 191026
rect 42111 190961 42177 190962
rect 42490 189066 45168 197572
rect 42486 189050 45168 189066
rect 42486 189048 43726 189050
rect 42486 189038 43716 189048
rect 42486 189006 43708 189038
rect 44452 189006 45168 189050
rect 41919 188362 41985 188363
rect 41919 188298 41920 188362
rect 41984 188298 41985 188362
rect 41919 188297 41985 188298
rect 42486 187612 42524 189006
rect 45090 187612 45168 189006
rect 42486 187528 45168 187612
rect 41343 187178 41409 187179
rect 41343 187114 41344 187178
rect 41408 187114 41409 187178
rect 41343 187113 41409 187114
rect 41151 186438 41217 186439
rect 41151 186374 41152 186438
rect 41216 186374 41217 186438
rect 41151 186373 41217 186374
rect 40959 185846 41025 185847
rect 40959 185782 40960 185846
rect 41024 185782 41025 185846
rect 40959 185781 41025 185782
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40383 182886 40449 182887
rect 40383 182822 40384 182886
rect 40448 182822 40449 182886
rect 40383 182821 40449 182822
rect 42490 179118 45168 187528
rect 45562 203700 47850 212842
rect 45562 203662 47858 203700
rect 45562 202576 45614 203662
rect 47814 202576 47858 203662
rect 45562 202514 47858 202576
rect 45562 193916 47850 202514
rect 45562 193878 47858 193916
rect 45562 192792 45614 193878
rect 47814 192792 47858 193878
rect 45562 192730 47858 192792
rect 45562 184130 47850 192730
rect 45562 184092 47858 184130
rect 45562 183006 45614 184092
rect 47814 183006 47858 184092
rect 45562 182944 47858 183006
rect 42490 179102 45174 179118
rect 42490 179100 43738 179102
rect 42490 179090 43728 179100
rect 42490 179058 43720 179090
rect 44464 179058 45174 179102
rect 42490 177664 42536 179058
rect 45102 177664 45174 179058
rect 42490 177580 45174 177664
rect 42490 169192 45168 177580
rect 42486 169176 45168 169192
rect 42486 169174 43726 169176
rect 42486 169132 43716 169174
rect 44452 169132 45168 169176
rect 42486 167738 42524 169132
rect 45090 167738 45168 169132
rect 42486 167654 45168 167738
rect 42490 159104 45168 167654
rect 42474 159088 45168 159104
rect 42474 159044 43714 159088
rect 44440 159044 45168 159088
rect 42474 157650 42512 159044
rect 45078 157650 45168 159044
rect 42474 157566 45168 157650
rect 42490 149120 45168 157566
rect 42464 149060 45168 149120
rect 42464 147666 42502 149060
rect 45068 147666 45168 149060
rect 42464 147582 45168 147666
rect 42490 139298 45168 147582
rect 42474 139238 45168 139298
rect 42474 137844 42512 139238
rect 45078 137844 45168 139238
rect 42474 137760 45168 137844
rect 42490 129430 45168 137760
rect 42464 129370 45168 129430
rect 42464 127976 42502 129370
rect 45068 127976 45168 129370
rect 42464 127892 45168 127976
rect 42490 119330 45168 127892
rect 42490 117936 42528 119330
rect 45094 117936 45168 119330
rect 42490 109324 45168 117936
rect 45562 173802 47850 182944
rect 45562 173764 47858 173802
rect 45562 172678 45614 173764
rect 47814 172678 47858 173764
rect 45562 172616 47858 172678
rect 45562 164018 47850 172616
rect 45562 163980 47858 164018
rect 45562 162894 45614 163980
rect 47814 162894 47858 163980
rect 45562 162832 47858 162894
rect 45562 154234 47850 162832
rect 45562 154196 47858 154234
rect 45562 153110 45614 154196
rect 47814 153110 47858 154196
rect 45562 153048 47858 153110
rect 45562 143906 47850 153048
rect 144831 144850 144897 144851
rect 144831 144786 144832 144850
rect 144896 144786 144897 144850
rect 144831 144785 144897 144786
rect 45562 143868 47858 143906
rect 45562 142782 45614 143868
rect 47814 142782 47858 143868
rect 45562 142720 47858 142782
rect 45562 134120 47850 142720
rect 45562 134082 47858 134120
rect 45562 132996 45614 134082
rect 47814 132996 47858 134082
rect 45562 132934 47858 132996
rect 45562 123792 47850 132934
rect 144834 126795 144894 144785
rect 144831 126794 144897 126795
rect 144831 126730 144832 126794
rect 144896 126730 144897 126794
rect 144831 126729 144897 126730
rect 144639 124574 144705 124575
rect 144639 124510 144640 124574
rect 144704 124510 144705 124574
rect 144639 124509 144705 124510
rect 45562 123754 47858 123792
rect 45562 122668 45614 123754
rect 47814 122668 47858 123754
rect 45562 122606 47858 122668
rect 45562 114212 47850 122606
rect 48038 120616 51232 120774
rect 48038 115126 48196 120616
rect 51046 115126 51232 120616
rect 48038 114888 51232 115126
rect 45562 114174 47926 114212
rect 45562 113122 45682 114174
rect 45638 113088 45682 113122
rect 47882 113734 47926 114174
rect 47882 113088 47942 113734
rect 45638 113026 47942 113088
rect 42430 109068 45168 109324
rect 42426 109052 45168 109068
rect 42426 109050 43666 109052
rect 42426 109040 43656 109050
rect 42426 109008 43648 109040
rect 44392 109008 45168 109052
rect 42426 107614 42464 109008
rect 45030 107614 45168 109008
rect 42426 107530 45168 107614
rect 42430 107486 45168 107530
rect 42490 99238 45168 107486
rect 45654 103884 47942 113026
rect 45638 103846 47942 103884
rect 45638 102760 45682 103846
rect 47882 102760 47942 103846
rect 45638 102698 47942 102760
rect 42454 98982 45168 99238
rect 42450 98966 45168 98982
rect 42450 98964 43690 98966
rect 42450 98954 43680 98964
rect 42450 98922 43672 98954
rect 44416 98922 45168 98966
rect 42450 97528 42488 98922
rect 45054 97528 45168 98922
rect 42450 97444 45168 97528
rect 42454 97400 45168 97444
rect 42490 89412 45168 97400
rect 45654 93906 47942 102698
rect 45626 93868 47942 93906
rect 45626 92782 45670 93868
rect 47870 92782 47942 93868
rect 45626 92720 47942 92782
rect 42478 89156 45168 89412
rect 42474 89142 45168 89156
rect 42474 89140 43720 89142
rect 42474 89138 43714 89140
rect 42474 89128 43704 89138
rect 42474 89096 43696 89128
rect 44446 89096 45168 89142
rect 42474 87702 42512 89096
rect 45078 87702 45168 89096
rect 42474 87618 45168 87702
rect 42478 87574 45168 87618
rect 42490 83634 45168 87574
rect 42372 83084 45168 83634
rect 45654 83916 47942 92720
rect 40836 82236 45208 83084
rect 40836 79346 40974 82236
rect 40820 79288 40974 79346
rect 45006 79288 45208 82236
rect 40820 77556 40888 79288
rect 45134 77556 45208 79288
rect 40820 77498 40974 77556
rect 40836 69384 40974 77498
rect 45006 69384 45208 77556
rect 45654 82830 45698 83916
rect 47898 82830 47942 83916
rect 45654 73970 47942 82830
rect 45628 73834 47942 73970
rect 45628 72892 45668 73834
rect 47790 72892 47942 73834
rect 45628 72808 47942 72892
rect 40836 67906 40900 69384
rect 45180 67906 45208 69384
rect 40836 59148 45208 67906
rect 40728 59078 45208 59148
rect 40728 57596 40844 59078
rect 45106 57596 45208 59078
rect 40728 57480 45208 57596
rect 40836 45628 45208 57480
rect 45654 64006 47942 72808
rect 45654 63064 45694 64006
rect 47816 63064 47942 64006
rect 45654 49658 47942 63064
rect 48564 55910 50852 114888
rect 144255 113326 144321 113327
rect 144255 113262 144256 113326
rect 144320 113262 144321 113326
rect 144255 113261 144321 113262
rect 144258 106815 144318 113261
rect 144255 106814 144321 106815
rect 144255 106750 144256 106814
rect 144320 106750 144321 106814
rect 144255 106749 144321 106750
rect 144642 106667 144702 124509
rect 144639 106666 144705 106667
rect 144639 106602 144640 106666
rect 144704 106602 144705 106666
rect 144639 106601 144705 106602
rect 50830 52944 50852 55910
rect 144462 51598 144938 51680
rect 144462 50716 144490 51598
rect 144898 50716 144938 51598
rect 145410 51463 145470 242021
rect 145599 218998 145665 218999
rect 145599 218934 145600 218998
rect 145664 218934 145665 218998
rect 145599 218933 145665 218934
rect 145407 51462 145473 51463
rect 145407 51398 145408 51462
rect 145472 51398 145473 51462
rect 145407 51397 145473 51398
rect 145602 51167 145662 218933
rect 181802 216660 193604 261204
rect 195968 248422 206088 269788
rect 208998 267922 209862 268102
rect 209016 267096 209598 267276
rect 209418 266750 209598 267096
rect 209682 266806 209862 267922
rect 210210 266410 210390 266516
rect 210474 266068 210654 270248
rect 290751 269170 290817 269171
rect 290751 269106 290752 269170
rect 290816 269106 290817 269170
rect 290751 269105 290817 269106
rect 316671 269170 316737 269171
rect 316671 269106 316672 269170
rect 316736 269106 316737 269170
rect 316671 269105 316737 269106
rect 347199 269170 347265 269171
rect 347199 269106 347200 269170
rect 347264 269106 347265 269170
rect 347199 269105 347265 269106
rect 347583 269170 347649 269171
rect 347583 269106 347584 269170
rect 347648 269106 347649 269170
rect 347583 269105 347649 269106
rect 290754 268431 290814 269105
rect 290751 268430 290817 268431
rect 290751 268366 290752 268430
rect 290816 268366 290817 268430
rect 290751 268365 290817 268366
rect 316674 268135 316734 269105
rect 292287 268134 292353 268135
rect 292287 268070 292288 268134
rect 292352 268070 292353 268134
rect 312447 268134 312513 268135
rect 292287 268069 292353 268070
rect 267903 267838 267969 267839
rect 267903 267774 267904 267838
rect 267968 267774 267969 267838
rect 267903 267773 267969 267774
rect 267906 267517 267966 267773
rect 292290 267517 292350 268069
rect 307842 268035 308478 268095
rect 312447 268070 312448 268134
rect 312512 268070 312513 268134
rect 312447 268069 312513 268070
rect 316671 268134 316737 268135
rect 316671 268070 316672 268134
rect 316736 268070 316737 268134
rect 316671 268069 316737 268070
rect 336447 268134 336513 268135
rect 336447 268070 336448 268134
rect 336512 268070 336513 268134
rect 336447 268069 336513 268070
rect 307842 267839 307902 268035
rect 308418 267839 308478 268035
rect 307839 267838 307905 267839
rect 307839 267774 307840 267838
rect 307904 267774 307905 267838
rect 307839 267773 307905 267774
rect 308415 267838 308481 267839
rect 308415 267774 308416 267838
rect 308480 267774 308481 267838
rect 308415 267773 308481 267774
rect 312450 267691 312510 268069
rect 336450 267691 336510 268069
rect 347202 267691 347262 269105
rect 347586 267691 347646 269105
rect 348546 268761 348606 270881
rect 369471 270650 369537 270651
rect 369471 270586 369472 270650
rect 369536 270586 369537 270650
rect 369471 270585 369537 270586
rect 369855 270586 369856 270611
rect 369920 270586 369921 270611
rect 369855 270585 369921 270586
rect 369474 270181 369534 270585
rect 384066 270181 384126 273249
rect 408255 273018 408321 273019
rect 408255 272954 408256 273018
rect 408320 272954 408321 273018
rect 408255 272953 408321 272954
rect 407871 271834 407937 271835
rect 407871 271770 407872 271834
rect 407936 271770 407937 271834
rect 407871 271769 407937 271770
rect 406143 271686 406209 271687
rect 406143 271622 406144 271686
rect 406208 271622 406209 271686
rect 406143 271621 406209 271622
rect 391743 270946 391809 270947
rect 391743 270882 391744 270946
rect 391808 270882 391809 270946
rect 391743 270881 391809 270882
rect 391746 270759 391806 270881
rect 391510 270699 391806 270759
rect 348354 268701 348606 268761
rect 348354 268431 348414 268701
rect 348351 268430 348417 268431
rect 348351 268366 348352 268430
rect 348416 268366 348417 268430
rect 348351 268365 348417 268366
rect 377535 268430 377601 268431
rect 377535 268366 377536 268430
rect 377600 268366 377601 268430
rect 377535 268365 377601 268366
rect 405951 268430 406017 268431
rect 405951 268366 405952 268430
rect 406016 268366 406017 268430
rect 405951 268365 406017 268366
rect 376578 268035 377022 268095
rect 376578 267839 376638 268035
rect 376575 267838 376641 267839
rect 376575 267774 376576 267838
rect 376640 267774 376641 267838
rect 376575 267773 376641 267774
rect 376962 267691 377022 268035
rect 312447 267690 312513 267691
rect 312447 267626 312448 267690
rect 312512 267626 312513 267690
rect 312447 267625 312513 267626
rect 336447 267690 336513 267691
rect 336447 267626 336448 267690
rect 336512 267626 336513 267690
rect 336447 267625 336513 267626
rect 347199 267690 347265 267691
rect 347199 267626 347200 267690
rect 347264 267626 347265 267690
rect 347199 267625 347265 267626
rect 347583 267690 347649 267691
rect 347583 267626 347584 267690
rect 347648 267626 347649 267690
rect 347583 267625 347649 267626
rect 376959 267690 377025 267691
rect 376959 267626 376960 267690
rect 377024 267626 377025 267690
rect 376959 267625 377025 267626
rect 377538 267517 377598 268365
rect 405375 267986 405441 267987
rect 405375 267922 405376 267986
rect 405440 267922 405441 267986
rect 405375 267921 405441 267922
rect 405759 267986 405825 267987
rect 405759 267922 405760 267986
rect 405824 267922 405825 267986
rect 405759 267921 405825 267922
rect 383679 267838 383745 267839
rect 383679 267774 383680 267838
rect 383744 267774 383745 267838
rect 383679 267773 383745 267774
rect 383682 267517 383742 267773
rect 210738 266372 211376 266552
rect 210738 265566 210918 266372
rect 405378 265431 405438 267921
rect 405378 265371 405630 265431
rect 211792 265166 212922 265206
rect 211792 261176 211832 265166
rect 212882 261176 212922 265166
rect 211792 261136 212922 261176
rect 206950 259514 209064 259554
rect 206950 256918 206990 259514
rect 209024 256918 209064 259514
rect 206950 256878 209064 256918
rect 206440 256334 209056 256374
rect 206440 256326 206480 256334
rect 206440 253276 206478 256326
rect 209016 253280 209056 256334
rect 208996 253276 209056 253280
rect 206440 253240 209056 253276
rect 194648 248416 206912 248422
rect 206854 240282 206912 248416
rect 207231 246970 207297 246971
rect 207231 246906 207232 246970
rect 207296 246906 207297 246970
rect 207231 246905 207297 246906
rect 207234 246231 207294 246905
rect 207231 246230 207297 246231
rect 207231 246166 207232 246230
rect 207296 246166 207297 246230
rect 207231 246165 207297 246166
rect 211530 245746 211710 246532
rect 211846 245954 215788 245994
rect 211846 245746 211886 245954
rect 211530 245566 211886 245746
rect 211846 244036 211886 245566
rect 215748 244036 215788 245954
rect 211846 243996 215788 244036
rect 210303 243714 210369 243715
rect 210303 243650 210304 243714
rect 210368 243650 210369 243714
rect 210303 243649 210369 243650
rect 211071 243714 211137 243715
rect 211071 243650 211072 243714
rect 211136 243650 211137 243714
rect 211071 243649 211137 243650
rect 194648 230162 206912 240282
rect 210306 233947 210366 243649
rect 210687 243122 210753 243123
rect 210687 243058 210688 243122
rect 210752 243058 210753 243122
rect 210687 243057 210753 243058
rect 210303 233946 210369 233947
rect 210303 233882 210304 233946
rect 210368 233882 210369 233946
rect 210303 233881 210369 233882
rect 210690 233651 210750 243057
rect 210687 233650 210753 233651
rect 210687 233586 210688 233650
rect 210752 233586 210753 233650
rect 210687 233585 210753 233586
rect 211074 233503 211134 243649
rect 405570 243567 405630 265371
rect 405762 247119 405822 267921
rect 405759 247118 405825 247119
rect 405759 247054 405760 247118
rect 405824 247054 405825 247118
rect 405759 247053 405825 247054
rect 405954 243567 406014 268365
rect 405567 243566 405633 243567
rect 405567 243502 405568 243566
rect 405632 243502 405633 243566
rect 405567 243501 405633 243502
rect 405951 243566 406017 243567
rect 405951 243502 405952 243566
rect 406016 243502 406017 243566
rect 405951 243501 406017 243502
rect 406146 242975 406206 271621
rect 407487 271538 407553 271539
rect 407487 271474 407488 271538
rect 407552 271474 407553 271538
rect 407487 271473 407553 271474
rect 406527 271242 406593 271243
rect 406527 271178 406528 271242
rect 406592 271178 406593 271242
rect 406527 271177 406593 271178
rect 406335 267986 406401 267987
rect 406335 267922 406336 267986
rect 406400 267922 406401 267986
rect 406335 267921 406401 267922
rect 406338 243419 406398 267921
rect 406530 246836 406590 271177
rect 406719 271094 406785 271095
rect 406719 271030 406720 271094
rect 406784 271030 406785 271094
rect 406719 271029 406785 271030
rect 406722 246971 406782 271029
rect 406911 270946 406977 270947
rect 406911 270882 406912 270946
rect 406976 270882 406977 270946
rect 406911 270881 406977 270882
rect 406719 246970 406785 246971
rect 406719 246906 406720 246970
rect 406784 246906 406785 246970
rect 406719 246905 406785 246906
rect 406518 246834 406600 246836
rect 406518 246758 406520 246834
rect 406598 246758 406600 246834
rect 406914 246823 406974 270881
rect 407091 264945 407175 264953
rect 407091 264875 407098 264945
rect 407168 264875 407175 264945
rect 407091 264867 407175 264875
rect 407295 264878 407361 264879
rect 407106 247267 407166 264867
rect 407295 264814 407296 264878
rect 407360 264814 407361 264878
rect 407295 264813 407361 264814
rect 407298 247563 407358 264813
rect 407490 247711 407550 271473
rect 407679 270798 407745 270799
rect 407679 270734 407680 270798
rect 407744 270734 407745 270798
rect 407679 270733 407745 270734
rect 407487 247710 407553 247711
rect 407487 247646 407488 247710
rect 407552 247646 407553 247710
rect 407487 247645 407553 247646
rect 407295 247562 407361 247563
rect 407295 247498 407296 247562
rect 407360 247498 407361 247562
rect 407295 247497 407361 247498
rect 407103 247266 407169 247267
rect 407103 247202 407104 247266
rect 407168 247202 407169 247266
rect 407103 247201 407169 247202
rect 407295 247266 407361 247267
rect 407295 247202 407296 247266
rect 407360 247202 407361 247266
rect 407295 247201 407361 247202
rect 407298 246971 407358 247201
rect 407682 247116 407742 270733
rect 407490 247056 407742 247116
rect 407295 246970 407361 246971
rect 407295 246906 407296 246970
rect 407360 246906 407361 246970
rect 407295 246905 407361 246906
rect 407490 246823 407550 247056
rect 407874 246968 407934 271769
rect 408108 264938 408180 264939
rect 408108 264935 408109 264938
rect 407682 246908 407934 246968
rect 408066 264868 408109 264935
rect 408179 264935 408180 264938
rect 408179 264875 408184 264935
rect 408179 264868 408180 264875
rect 408066 264867 408180 264868
rect 406518 246754 406600 246758
rect 406911 246822 406977 246823
rect 406911 246758 406912 246822
rect 406976 246758 406977 246822
rect 406911 246757 406977 246758
rect 407487 246822 407553 246823
rect 407487 246758 407488 246822
rect 407552 246758 407553 246822
rect 407487 246757 407553 246758
rect 406335 243418 406401 243419
rect 406335 243354 406336 243418
rect 406400 243354 406401 243418
rect 406335 243353 406401 243354
rect 407682 243271 407742 246908
rect 408066 246823 408126 264867
rect 408063 246822 408129 246823
rect 408063 246758 408064 246822
rect 408128 246758 408129 246822
rect 408063 246757 408129 246758
rect 408258 243567 408318 272953
rect 409215 271242 409281 271243
rect 409215 271178 409216 271242
rect 409280 271178 409281 271242
rect 409215 271177 409281 271178
rect 408447 247710 408513 247711
rect 408447 247646 408448 247710
rect 408512 247646 408513 247710
rect 408447 247645 408513 247646
rect 408639 247710 408705 247711
rect 408639 247646 408640 247710
rect 408704 247646 408705 247710
rect 408639 247645 408705 247646
rect 408450 246823 408510 247645
rect 408447 246822 408513 246823
rect 408447 246758 408448 246822
rect 408512 246758 408513 246822
rect 408642 246820 408702 247645
rect 409218 247449 409278 271177
rect 408834 247389 409278 247449
rect 408834 246971 408894 247389
rect 408831 246970 408897 246971
rect 408831 246906 408832 246970
rect 408896 246906 408897 246970
rect 408831 246905 408897 246906
rect 408831 246822 408897 246823
rect 408831 246820 408832 246822
rect 408642 246760 408832 246820
rect 408447 246757 408513 246758
rect 408831 246758 408832 246760
rect 408896 246758 408897 246822
rect 408831 246757 408897 246758
rect 409215 246822 409281 246823
rect 409215 246758 409216 246822
rect 409280 246820 409281 246822
rect 409410 246820 409470 273397
rect 409791 273314 409857 273315
rect 409791 273250 409792 273314
rect 409856 273250 409857 273314
rect 409791 273249 409857 273250
rect 409599 272722 409665 272723
rect 409599 272658 409600 272722
rect 409664 272658 409665 272722
rect 409599 272657 409665 272658
rect 409602 246823 409662 272657
rect 409794 247563 409854 273249
rect 410559 272870 410625 272871
rect 410559 272806 410560 272870
rect 410624 272806 410625 272870
rect 410559 272805 410625 272806
rect 410175 272278 410241 272279
rect 410175 272214 410176 272278
rect 410240 272214 410241 272278
rect 410175 272213 410241 272214
rect 409983 264730 410049 264731
rect 409983 264666 409984 264730
rect 410048 264666 410049 264730
rect 409983 264665 410049 264666
rect 409791 247562 409857 247563
rect 409791 247498 409792 247562
rect 409856 247498 409857 247562
rect 409791 247497 409857 247498
rect 409986 247267 410046 264665
rect 410178 247267 410238 272213
rect 410367 264878 410433 264879
rect 410367 264814 410368 264878
rect 410432 264814 410433 264878
rect 410367 264813 410433 264814
rect 410370 247415 410430 264813
rect 410562 264765 410622 272805
rect 410943 271982 411009 271983
rect 410943 271918 410944 271982
rect 411008 271918 411009 271982
rect 410943 271917 411009 271918
rect 410562 264731 410814 264765
rect 410562 264730 410817 264731
rect 410562 264705 410752 264730
rect 410751 264666 410752 264705
rect 410816 264666 410817 264730
rect 410751 264665 410817 264666
rect 410559 264582 410625 264583
rect 410559 264518 410560 264582
rect 410624 264518 410625 264582
rect 410559 264517 410625 264518
rect 410367 247414 410433 247415
rect 410367 247350 410368 247414
rect 410432 247350 410433 247414
rect 410367 247349 410433 247350
rect 409983 247266 410049 247267
rect 409983 247202 409984 247266
rect 410048 247202 410049 247266
rect 409983 247201 410049 247202
rect 410175 247266 410241 247267
rect 410175 247202 410176 247266
rect 410240 247202 410241 247266
rect 410175 247201 410241 247202
rect 410562 247119 410622 264517
rect 410751 247858 410817 247859
rect 410751 247794 410752 247858
rect 410816 247794 410817 247858
rect 410751 247793 410817 247794
rect 410754 247119 410814 247793
rect 410559 247118 410625 247119
rect 410559 247054 410560 247118
rect 410624 247054 410625 247118
rect 410559 247053 410625 247054
rect 410751 247118 410817 247119
rect 410751 247054 410752 247118
rect 410816 247054 410817 247118
rect 410751 247053 410817 247054
rect 410946 246971 411006 271917
rect 411135 271686 411201 271687
rect 411135 271622 411136 271686
rect 411200 271622 411201 271686
rect 411135 271621 411201 271622
rect 411138 247711 411198 271621
rect 411327 271538 411393 271539
rect 411327 271474 411328 271538
rect 411392 271474 411393 271538
rect 411327 271473 411393 271474
rect 411135 247710 411201 247711
rect 411135 247646 411136 247710
rect 411200 247646 411201 247710
rect 411135 247645 411201 247646
rect 411330 247415 411390 271473
rect 413886 269066 415028 269246
rect 411638 267970 412568 268010
rect 411638 265796 411678 267970
rect 412528 266564 412568 267970
rect 412528 266384 413010 266564
rect 412528 265796 412568 266384
rect 411638 265756 412568 265796
rect 412830 265302 413010 266384
rect 413094 265530 413274 267242
rect 413886 266360 414066 269066
rect 414150 268090 415068 268270
rect 414150 266570 414330 268090
rect 650628 266628 651228 279318
rect 654388 269618 654988 275470
rect 653130 269578 654988 269618
rect 653130 269026 653170 269578
rect 654946 269026 654988 269578
rect 653130 269006 654988 269026
rect 653130 268986 654986 269006
rect 655328 268554 655928 274538
rect 658682 273109 660572 317003
rect 658682 271927 659369 273109
rect 660551 271927 660572 273109
rect 654876 268526 656474 268554
rect 654876 267934 654916 268526
rect 656440 267934 656474 268526
rect 654876 267890 656474 267934
rect 649894 266624 652026 266628
rect 647060 266582 654386 266624
rect 647060 265124 647144 266582
rect 654338 265124 654386 266582
rect 647060 265036 654386 265124
rect 411519 264730 411585 264731
rect 411519 264666 411520 264730
rect 411584 264666 411585 264730
rect 411519 264665 411585 264666
rect 411522 247859 411582 264665
rect 424642 264332 424962 264684
rect 434642 264428 434962 264682
rect 432388 264388 436506 264428
rect 411832 264272 412460 264312
rect 411832 261174 411872 264272
rect 412420 261174 412460 264272
rect 422480 264292 426788 264332
rect 422480 261214 422520 264292
rect 426748 261214 426788 264292
rect 422480 261174 426788 261214
rect 411832 261134 412460 261174
rect 416314 259552 424246 259592
rect 416314 256926 416354 259552
rect 424206 256926 424246 259552
rect 416314 256886 424246 256926
rect 416408 256862 424200 256886
rect 416290 256398 424314 256438
rect 416290 253332 416330 256398
rect 424274 253332 424314 256398
rect 416290 253292 424314 253332
rect 411519 247858 411585 247859
rect 411519 247794 411520 247858
rect 411584 247794 411585 247858
rect 411519 247793 411585 247794
rect 411327 247414 411393 247415
rect 411327 247350 411328 247414
rect 411392 247350 411393 247414
rect 411327 247349 411393 247350
rect 410943 246970 411009 246971
rect 410943 246906 410944 246970
rect 411008 246906 411009 246970
rect 410943 246905 411009 246906
rect 409280 246760 409470 246820
rect 409599 246822 409665 246823
rect 409280 246758 409281 246760
rect 409215 246757 409281 246758
rect 409599 246758 409600 246822
rect 409664 246758 409665 246822
rect 409599 246757 409665 246758
rect 412566 244978 412746 248888
rect 409606 244938 412758 244978
rect 408255 243566 408321 243567
rect 408255 243502 408256 243566
rect 408320 243502 408321 243566
rect 408255 243501 408321 243502
rect 407679 243270 407745 243271
rect 407679 243206 407680 243270
rect 407744 243206 407745 243270
rect 407679 243205 407745 243206
rect 406143 242974 406209 242975
rect 406143 242910 406144 242974
rect 406208 242910 406209 242974
rect 406143 242909 406209 242910
rect 409606 242868 409646 244938
rect 412718 242868 412758 244938
rect 409606 242828 412758 242868
rect 328767 242826 328833 242827
rect 328767 242787 328768 242826
rect 328386 242762 328768 242787
rect 328832 242762 328833 242826
rect 328386 242761 328833 242762
rect 328386 242727 328830 242761
rect 328386 242383 328446 242727
rect 328383 242382 328449 242383
rect 328383 242318 328384 242382
rect 328448 242318 328449 242382
rect 328383 242317 328449 242318
rect 212031 242234 212097 242235
rect 212031 242170 212032 242234
rect 212096 242170 212097 242234
rect 212031 242169 212097 242170
rect 211455 237794 211521 237795
rect 211455 237730 211456 237794
rect 211520 237730 211521 237794
rect 211455 237729 211521 237730
rect 211071 233502 211137 233503
rect 211071 233438 211072 233502
rect 211136 233438 211137 233502
rect 211071 233437 211137 233438
rect 210687 233354 210753 233355
rect 210687 233290 210688 233354
rect 210752 233290 210753 233354
rect 210687 233289 210753 233290
rect 206846 224480 206912 230162
rect 145791 216482 145857 216483
rect 145791 216418 145792 216482
rect 145856 216418 145857 216482
rect 145791 216417 145857 216418
rect 145794 51315 145854 216417
rect 145983 214558 146049 214559
rect 145983 214494 145984 214558
rect 146048 214494 146049 214558
rect 145983 214493 146049 214494
rect 145791 51314 145857 51315
rect 145791 51250 145792 51314
rect 145856 51250 145857 51314
rect 145791 51249 145857 51250
rect 145599 51166 145665 51167
rect 145599 51102 145600 51166
rect 145664 51102 145665 51166
rect 145599 51101 145665 51102
rect 145986 51019 146046 214493
rect 193602 206248 193604 216660
rect 181802 185790 193604 206248
rect 194648 202814 206912 224480
rect 210690 223473 210750 233289
rect 210690 223413 211134 223473
rect 211074 207489 211134 223413
rect 210498 207429 211134 207489
rect 181802 174942 181814 185790
rect 193522 174942 193604 185790
rect 181802 155854 193604 174942
rect 193516 144926 193604 155854
rect 181802 127140 193604 144926
rect 194648 173320 206912 192744
rect 210111 190138 210177 190139
rect 210111 190074 210112 190138
rect 210176 190074 210177 190138
rect 210111 190073 210177 190074
rect 209919 175782 209985 175783
rect 209919 175718 209920 175782
rect 209984 175718 209985 175782
rect 209919 175717 209985 175718
rect 194648 163330 194714 173320
rect 209922 171343 209982 175717
rect 209919 171342 209985 171343
rect 209919 171278 209920 171342
rect 209984 171278 209985 171342
rect 209919 171277 209985 171278
rect 210114 170603 210174 190073
rect 210498 174855 210558 207429
rect 211458 206157 211518 237729
rect 211647 234686 211713 234687
rect 211647 234622 211648 234686
rect 211712 234622 211713 234686
rect 211647 234621 211713 234622
rect 210882 206097 211518 206157
rect 210882 195023 210942 206097
rect 211650 205491 211710 234621
rect 212034 233799 212094 242169
rect 241791 238534 241857 238535
rect 241791 238470 241792 238534
rect 241856 238470 241857 238534
rect 241791 238469 241857 238470
rect 241794 238239 241854 238469
rect 241791 238238 241857 238239
rect 241791 238174 241792 238238
rect 241856 238174 241857 238238
rect 241791 238173 241857 238174
rect 239103 236758 239169 236759
rect 239103 236694 239104 236758
rect 239168 236694 239169 236758
rect 239103 236693 239169 236694
rect 239106 236315 239166 236693
rect 239103 236314 239169 236315
rect 239103 236250 239104 236314
rect 239168 236250 239169 236314
rect 239103 236249 239169 236250
rect 212031 233798 212097 233799
rect 212031 233734 212032 233798
rect 212096 233734 212097 233798
rect 212031 233733 212097 233734
rect 212991 233798 213057 233799
rect 212991 233734 212992 233798
rect 213056 233734 213057 233798
rect 212991 233733 213057 233734
rect 212607 233650 212673 233651
rect 212607 233648 212608 233650
rect 212562 233586 212608 233648
rect 212672 233586 212673 233650
rect 212562 233585 212673 233586
rect 212223 233502 212289 233503
rect 212223 233438 212224 233502
rect 212288 233438 212289 233502
rect 212223 233437 212289 233438
rect 211266 205431 211710 205491
rect 211071 205086 211137 205087
rect 211071 205022 211072 205086
rect 211136 205084 211137 205086
rect 211266 205084 211326 205431
rect 211136 205024 211326 205084
rect 211136 205022 211137 205024
rect 211071 205021 211137 205022
rect 212226 195501 212286 233437
rect 212562 232131 212622 233585
rect 212799 233502 212865 233503
rect 212799 233438 212800 233502
rect 212864 233438 212865 233502
rect 212799 233437 212865 233438
rect 211074 195441 212286 195501
rect 212418 232071 212622 232131
rect 211074 195023 211134 195441
rect 210879 195022 210945 195023
rect 210879 194958 210880 195022
rect 210944 194958 210945 195022
rect 210879 194957 210945 194958
rect 211071 195022 211137 195023
rect 211071 194958 211072 195022
rect 211136 194958 211137 195022
rect 211071 194957 211137 194958
rect 212418 194835 212478 232071
rect 210306 174795 210558 174855
rect 210690 194775 212478 194835
rect 210306 174007 210366 174795
rect 210690 174451 210750 194775
rect 210879 194578 210945 194579
rect 210879 194514 210880 194578
rect 210944 194514 210945 194578
rect 210879 194513 210945 194514
rect 210687 174450 210753 174451
rect 210687 174386 210688 174450
rect 210752 174386 210753 174450
rect 210687 174385 210753 174386
rect 210882 174189 210942 194513
rect 211074 194135 212286 194169
rect 211071 194134 212286 194135
rect 211071 194070 211072 194134
rect 211136 194109 212286 194134
rect 211136 194070 211137 194109
rect 211071 194069 211137 194070
rect 212226 190173 212286 194109
rect 211074 190139 212286 190173
rect 211071 190138 212286 190139
rect 211071 190074 211072 190138
rect 211136 190113 212286 190138
rect 211136 190074 211137 190113
rect 211071 190073 211137 190074
rect 211071 175782 211137 175783
rect 211071 175718 211072 175782
rect 211136 175780 211137 175782
rect 212802 175780 212862 233437
rect 211136 175720 212862 175780
rect 211136 175718 211137 175720
rect 211071 175717 211137 175718
rect 211071 174450 211137 174451
rect 211071 174386 211072 174450
rect 211136 174448 211137 174450
rect 211136 174388 212862 174448
rect 211136 174386 211137 174388
rect 211071 174385 211137 174386
rect 210498 174129 210942 174189
rect 210303 174006 210369 174007
rect 210303 173942 210304 174006
rect 210368 173942 210369 174006
rect 210303 173941 210369 173942
rect 210111 170602 210177 170603
rect 210111 170538 210112 170602
rect 210176 170538 210177 170602
rect 210111 170537 210177 170538
rect 194648 141504 206912 163330
rect 210111 151954 210177 151955
rect 210111 151890 210112 151954
rect 210176 151890 210177 151954
rect 210111 151889 210177 151890
rect 206858 131594 206912 141504
rect 181802 115426 181900 127140
rect 193528 115426 193604 127140
rect 181802 98150 193604 115426
rect 194648 112852 206912 131594
rect 210114 121575 210174 151889
rect 210498 143553 210558 174129
rect 210879 174006 210945 174007
rect 210879 173942 210880 174006
rect 210944 173942 210945 174006
rect 210879 173941 210945 173942
rect 210882 151955 210942 173941
rect 211071 171342 211137 171343
rect 211071 171278 211072 171342
rect 211136 171278 211137 171342
rect 211071 171277 211137 171278
rect 211074 170859 211134 171277
rect 211074 170799 211518 170859
rect 211071 170602 211137 170603
rect 211071 170538 211072 170602
rect 211136 170600 211137 170602
rect 211136 170540 211326 170600
rect 211136 170538 211137 170540
rect 211071 170537 211137 170538
rect 211266 165531 211326 170540
rect 211458 167529 211518 170799
rect 211458 167469 212478 167529
rect 211266 165471 211902 165531
rect 211071 164238 211137 164239
rect 211071 164174 211072 164238
rect 211136 164199 211137 164238
rect 211136 164174 211326 164199
rect 211071 164173 211326 164174
rect 211074 164139 211326 164173
rect 210879 151954 210945 151955
rect 210879 151890 210880 151954
rect 210944 151890 210945 151954
rect 210879 151889 210945 151890
rect 210498 143493 211134 143553
rect 211074 138225 211134 143493
rect 210498 138165 211134 138225
rect 210303 137302 210369 137303
rect 210303 137238 210304 137302
rect 210368 137238 210369 137302
rect 210303 137237 210369 137238
rect 210306 124905 210366 137237
rect 210498 125167 210558 138165
rect 211266 137559 211326 164139
rect 211842 155541 211902 165471
rect 211074 137499 211326 137559
rect 211458 155481 211902 155541
rect 211074 137303 211134 137499
rect 211071 137302 211137 137303
rect 211071 137238 211072 137302
rect 211136 137238 211137 137302
rect 211071 137237 211137 137238
rect 211458 132897 211518 155481
rect 212418 154875 212478 167469
rect 212226 154815 212478 154875
rect 212226 151952 212286 154815
rect 211842 151892 212286 151952
rect 211842 150879 211902 151892
rect 212802 151545 212862 174388
rect 212418 151485 212862 151545
rect 211842 150819 212286 150879
rect 211074 132837 211518 132897
rect 210495 125166 210561 125167
rect 210495 125102 210496 125166
rect 210560 125102 210561 125166
rect 210495 125101 210561 125102
rect 210306 124845 210942 124905
rect 210303 123094 210369 123095
rect 210303 123030 210304 123094
rect 210368 123030 210369 123094
rect 210303 123029 210369 123030
rect 210306 121763 210366 123029
rect 210303 121762 210369 121763
rect 210303 121698 210304 121762
rect 210368 121698 210369 121762
rect 210303 121697 210369 121698
rect 210114 121515 210558 121575
rect 210111 121318 210177 121319
rect 210111 121254 210112 121318
rect 210176 121254 210177 121318
rect 210111 121253 210177 121254
rect 210303 121318 210369 121319
rect 210303 121254 210304 121318
rect 210368 121254 210369 121318
rect 210303 121253 210369 121254
rect 209727 106518 209793 106519
rect 209727 106454 209728 106518
rect 209792 106454 209793 106518
rect 209727 106453 209793 106454
rect 181802 86356 181900 98150
rect 181802 60778 193604 86356
rect 194648 83100 206912 100374
rect 206852 83060 206912 83100
rect 193566 54130 193604 60778
rect 145983 51018 146049 51019
rect 145983 50954 145984 51018
rect 146048 50954 146049 51018
rect 145983 50953 146049 50954
rect 144462 50648 144938 50716
rect 45558 49544 48232 49658
rect 45558 46014 45634 49544
rect 48118 46014 48232 49544
rect 144740 49132 144920 50648
rect 45558 45912 48232 46014
rect 45186 43052 45208 45628
rect 143440 42520 143620 48626
rect 143860 45500 144040 48622
rect 181802 45584 193604 54130
rect 194648 49686 206912 60770
rect 209730 53831 209790 106453
rect 210114 90979 210174 121253
rect 210306 118063 210366 121253
rect 210303 118062 210369 118063
rect 210303 117998 210304 118062
rect 210368 117998 210369 118062
rect 210303 117997 210369 117998
rect 210498 106519 210558 121515
rect 210495 106518 210561 106519
rect 210495 106454 210496 106518
rect 210560 106454 210561 106518
rect 210495 106453 210561 106454
rect 210111 90978 210177 90979
rect 210111 90914 210112 90978
rect 210176 90914 210177 90978
rect 210111 90913 210177 90914
rect 210495 90978 210561 90979
rect 210495 90914 210496 90978
rect 210560 90914 210561 90978
rect 210495 90913 210561 90914
rect 210111 90386 210177 90387
rect 210111 90322 210112 90386
rect 210176 90322 210177 90386
rect 210111 90321 210177 90322
rect 210114 82691 210174 90321
rect 210303 87722 210369 87723
rect 210303 87658 210304 87722
rect 210368 87658 210369 87722
rect 210303 87657 210369 87658
rect 210111 82690 210177 82691
rect 210111 82626 210112 82690
rect 210176 82626 210177 82690
rect 210111 82625 210177 82626
rect 210111 72922 210177 72923
rect 210111 72858 210112 72922
rect 210176 72858 210177 72922
rect 210111 72857 210177 72858
rect 210114 69627 210174 72857
rect 210306 70293 210366 87657
rect 210498 70959 210558 90913
rect 210687 89350 210753 89351
rect 210687 89286 210688 89350
rect 210752 89286 210753 89350
rect 210687 89285 210753 89286
rect 210690 87279 210750 89285
rect 210687 87278 210753 87279
rect 210687 87214 210688 87278
rect 210752 87214 210753 87278
rect 210687 87213 210753 87214
rect 210882 84945 210942 124845
rect 211074 123095 211134 132837
rect 211071 123094 211137 123095
rect 211071 123030 211072 123094
rect 211136 123030 211137 123094
rect 211071 123029 211137 123030
rect 212226 122241 212286 150819
rect 211842 122181 212286 122241
rect 211071 118062 211137 118063
rect 211071 117998 211072 118062
rect 211136 117998 211137 118062
rect 211071 117997 211137 117998
rect 211074 90387 211134 117997
rect 211842 117579 211902 122181
rect 212418 121316 212478 151485
rect 212418 121256 212670 121316
rect 211842 117519 212286 117579
rect 212226 102261 212286 117519
rect 211266 102201 212286 102261
rect 211071 90386 211137 90387
rect 211071 90322 211072 90386
rect 211136 90322 211137 90386
rect 211071 90321 211137 90322
rect 211266 89607 211326 102201
rect 212610 100263 212670 121256
rect 212994 100263 213054 233733
rect 424642 229466 424962 261174
rect 432388 261166 432428 264388
rect 436466 261166 436506 264388
rect 444642 264354 444962 264564
rect 454642 264358 454962 264664
rect 432388 261126 436506 261166
rect 442152 264314 446456 264354
rect 429642 248522 429962 249030
rect 428124 248482 431026 248522
rect 428124 242898 428164 248482
rect 430986 242898 431026 248482
rect 428124 242858 431026 242898
rect 429642 228810 429962 242858
rect 434642 230594 434962 261126
rect 442152 261084 442192 264314
rect 446416 261084 446456 264314
rect 452868 264318 457092 264358
rect 464642 264354 464962 264758
rect 474642 264354 474962 264800
rect 452868 261168 452908 264318
rect 457052 261168 457092 264318
rect 463502 264314 467226 264354
rect 463502 261250 463542 264314
rect 467186 261250 467226 264314
rect 463502 261210 467226 261250
rect 472646 264314 477196 264354
rect 452868 261128 457092 261168
rect 442152 261044 446456 261084
rect 439642 248350 439962 249308
rect 437704 248310 440526 248350
rect 437704 242806 437744 248310
rect 440486 242806 440526 248310
rect 437704 242766 440526 242806
rect 439642 230050 439962 242766
rect 444642 230164 444962 261044
rect 449642 248614 449962 249180
rect 448158 248574 451474 248614
rect 448158 242806 448198 248574
rect 451434 242806 451474 248574
rect 448158 242766 451474 242806
rect 449642 229358 449962 242766
rect 454642 228874 454962 261128
rect 459642 248626 459962 249180
rect 458290 248586 461526 248626
rect 458290 242898 458330 248586
rect 461486 242898 461526 248586
rect 458290 242858 461526 242898
rect 459642 229766 459962 242858
rect 464642 229506 464962 261210
rect 472646 261168 472686 264314
rect 477156 261168 477196 264314
rect 484642 264272 484962 264704
rect 494642 264396 494962 264900
rect 492504 264356 497138 264396
rect 482740 264232 488036 264272
rect 482740 261208 482780 264232
rect 487996 261208 488036 264232
rect 482740 261168 488036 261208
rect 492504 261168 492544 264356
rect 497098 261168 497138 264356
rect 504642 264314 504962 264710
rect 472646 261128 477196 261168
rect 469642 248592 469962 248636
rect 468330 248552 471486 248592
rect 468330 242944 468370 248552
rect 471446 242944 471486 248552
rect 468330 242904 471486 242944
rect 469642 230050 469962 242904
rect 474642 229506 474962 261128
rect 479642 248568 479962 248954
rect 478278 248528 481272 248568
rect 478278 242898 478318 248528
rect 481232 242898 481272 248528
rect 478278 242858 481272 242898
rect 479642 229630 479962 242858
rect 484642 229242 484962 261168
rect 492504 261128 497138 261168
rect 502518 264274 507730 264314
rect 489642 248706 489962 249162
rect 488272 248666 491126 248706
rect 488272 242852 488312 248666
rect 491086 242852 491126 248666
rect 488272 242812 491126 242852
rect 489642 229652 489962 242812
rect 494642 229890 494962 261128
rect 502518 261126 502558 264274
rect 507690 261126 507730 264274
rect 514642 264272 514962 264616
rect 524642 264354 524962 264810
rect 522748 264314 527382 264354
rect 534642 264314 534962 264716
rect 544642 264358 544962 264622
rect 542774 264318 547492 264358
rect 502518 261086 507730 261126
rect 511868 264232 517494 264272
rect 511868 261126 511908 264232
rect 517454 261126 517494 264232
rect 522748 261168 522788 264314
rect 527342 261168 527382 264314
rect 522748 261128 527382 261168
rect 532638 264274 537436 264314
rect 511868 261086 517494 261126
rect 499642 248626 499962 248982
rect 498772 248586 501546 248626
rect 498772 242852 498812 248586
rect 501506 242852 501546 248586
rect 498772 242812 501546 242852
rect 499642 230024 499962 242812
rect 504642 229962 504962 261086
rect 509642 248592 509962 248828
rect 508122 248552 510816 248592
rect 508122 242898 508162 248552
rect 510776 242898 510816 248552
rect 508122 242858 510816 242898
rect 509642 230434 509962 242858
rect 514642 229412 514962 261086
rect 519642 248568 519962 249346
rect 517884 248528 521754 248568
rect 517884 242852 517924 248528
rect 521714 242852 521754 248528
rect 517884 242812 521754 242852
rect 519642 230050 519962 242812
rect 524642 229450 524962 261128
rect 532638 261084 532678 264274
rect 537396 261084 537436 264274
rect 542774 261208 542814 264318
rect 547452 261208 547492 264318
rect 554642 264314 554962 264906
rect 542774 261168 547492 261208
rect 552496 264274 557876 264314
rect 552496 261208 552536 264274
rect 557836 261208 557876 264274
rect 564642 264190 564962 264716
rect 574642 264478 574962 264744
rect 573184 264438 577694 264478
rect 584642 264438 584962 264738
rect 594642 264438 594962 264644
rect 552496 261168 557876 261208
rect 562922 264150 567474 264190
rect 532638 261044 537436 261084
rect 529642 248442 529962 249066
rect 527878 248402 531668 248442
rect 527878 242806 527918 248402
rect 531628 242806 531668 248402
rect 527878 242766 531668 242806
rect 529642 229908 529962 242766
rect 534642 229890 534962 261044
rect 539642 248614 539962 249236
rect 538102 248574 541510 248614
rect 538102 242806 538142 248574
rect 541470 242806 541510 248574
rect 538102 242766 541510 242806
rect 539642 229918 539962 242766
rect 544642 229070 544962 261168
rect 549642 248580 549962 248814
rect 547774 248540 551102 248580
rect 547774 242852 547814 248540
rect 551062 242852 551102 248540
rect 547774 242812 551102 242852
rect 549642 230050 549962 242812
rect 554642 229356 554962 261168
rect 562922 261126 562962 264150
rect 567434 261126 567474 264150
rect 562922 261086 567474 261126
rect 573184 261126 573224 264438
rect 577654 261126 577694 264438
rect 573184 261086 577694 261126
rect 582782 264398 587748 264438
rect 559642 248568 559962 248886
rect 557170 248528 561268 248568
rect 557170 242898 557210 248528
rect 561228 242898 561268 248528
rect 557170 242858 561268 242898
rect 559642 230008 559962 242858
rect 564642 229890 564962 261086
rect 569642 248614 569962 249098
rect 567578 248574 571862 248614
rect 567578 242806 567618 248574
rect 571822 242806 571862 248574
rect 567578 242766 571862 242806
rect 569642 229346 569962 242766
rect 574642 230154 574962 261086
rect 582782 261084 582822 264398
rect 587708 261084 587748 264398
rect 592298 264398 596890 264438
rect 592298 261168 592338 264398
rect 596850 261168 596890 264398
rect 604642 264354 604962 264644
rect 592298 261128 596890 261168
rect 602600 264314 606820 264354
rect 582782 261044 587748 261084
rect 579642 248476 579962 249608
rect 577066 248436 581118 248476
rect 577066 242898 577106 248436
rect 581078 242898 581118 248436
rect 577066 242858 581118 242898
rect 579642 229450 579962 242858
rect 584642 229954 584962 261044
rect 589642 248614 589962 248722
rect 588210 248574 591756 248614
rect 588210 242898 588250 248574
rect 591716 242898 591756 248574
rect 588210 242858 591756 242898
rect 589642 229628 589962 242858
rect 594642 229890 594962 261128
rect 602600 261044 602640 264314
rect 606780 261044 606820 264314
rect 614642 264272 614962 264832
rect 624642 264314 624962 264832
rect 634642 264314 634962 264582
rect 622708 264274 626970 264314
rect 613192 264232 617412 264272
rect 613192 261250 613232 264232
rect 617372 261250 617412 264232
rect 613192 261210 617412 261250
rect 602600 261004 606820 261044
rect 599642 248568 599962 248988
rect 597606 248528 601474 248568
rect 597606 242898 597646 248528
rect 601434 242898 601474 248528
rect 597606 242858 601474 242898
rect 599642 229892 599962 242858
rect 604642 229890 604962 261004
rect 609642 248488 609962 249254
rect 607324 248448 611112 248488
rect 607324 242898 607364 248448
rect 611072 242898 611112 248448
rect 607324 242858 611112 242898
rect 609642 230434 609962 242858
rect 614642 229390 614962 261210
rect 622708 261168 622748 264274
rect 626930 261168 626970 264274
rect 622708 261128 626970 261168
rect 632430 264274 637562 264314
rect 632430 261168 632470 264274
rect 637522 261168 637562 264274
rect 632430 261128 637562 261168
rect 619642 248706 619962 248990
rect 618192 248666 621324 248706
rect 618192 242898 618232 248666
rect 621284 242898 621324 248666
rect 618192 242858 621324 242898
rect 619642 230434 619962 242858
rect 624642 229954 624962 261128
rect 629642 248568 629962 248970
rect 627864 248528 631594 248568
rect 627864 242852 627904 248528
rect 631554 242852 631594 248528
rect 627864 242812 631594 242852
rect 629642 230524 629962 242812
rect 634642 228802 634962 261128
rect 655328 252656 655928 267890
rect 658682 259624 660572 271927
rect 661102 990384 661196 992954
rect 664096 990384 664196 992954
rect 661102 947415 664196 990384
rect 661102 946233 662179 947415
rect 663361 946233 664196 947415
rect 661102 768629 664196 946233
rect 661102 767447 662179 768629
rect 663361 767447 664196 768629
rect 661102 723371 664196 767447
rect 661102 722189 662179 723371
rect 663361 722189 664196 723371
rect 661102 678967 664196 722189
rect 661102 677785 662179 678967
rect 663361 677785 664196 678967
rect 661102 633625 664196 677785
rect 661102 632443 662179 633625
rect 663361 632443 664196 633625
rect 661102 587355 664196 632443
rect 661102 586173 662179 587355
rect 663361 586173 664196 587355
rect 661102 543901 664196 586173
rect 661102 542719 662179 543901
rect 663361 542719 664196 543901
rect 661102 499413 664196 542719
rect 661102 498231 662179 499413
rect 663361 498231 664196 499413
rect 661102 411215 664196 498231
rect 665024 985912 668306 994456
rect 671662 994230 673462 994266
rect 671658 994178 673462 994230
rect 671658 991374 671690 994178
rect 673416 991374 673462 994178
rect 671658 991312 673462 991374
rect 665024 983950 665082 985912
rect 668280 983950 668306 985912
rect 665024 949401 668306 983950
rect 665024 948219 666067 949401
rect 667249 948219 668306 949401
rect 665024 770527 668306 948219
rect 669318 987294 670414 990652
rect 669318 986772 669334 987294
rect 670384 986772 670414 987294
rect 669318 832446 670414 986772
rect 671662 985060 673462 991312
rect 671662 981854 671718 985060
rect 672730 985058 673462 985060
rect 673374 981854 673462 985058
rect 671662 950872 673462 981854
rect 675711 967434 675777 967435
rect 675711 967370 675712 967434
rect 675776 967370 675777 967434
rect 675711 967369 675777 967370
rect 674367 965066 674433 965067
rect 674367 965002 674368 965066
rect 674432 965002 674433 965066
rect 674367 965001 674433 965002
rect 673983 956038 674049 956039
rect 673983 955974 673984 956038
rect 674048 955974 674049 956038
rect 673983 955973 674049 955974
rect 671662 949780 671683 950872
rect 672775 949780 673462 950872
rect 671662 917976 673462 949780
rect 673986 932655 674046 955973
rect 674370 937539 674430 965001
rect 675135 964918 675201 964919
rect 675135 964854 675136 964918
rect 675200 964854 675201 964918
rect 675135 964853 675201 964854
rect 674943 962846 675009 962847
rect 674943 962782 674944 962846
rect 675008 962782 675009 962846
rect 674943 962781 675009 962782
rect 674559 962550 674625 962551
rect 674559 962486 674560 962550
rect 674624 962486 674625 962550
rect 674559 962485 674625 962486
rect 674367 937538 674433 937539
rect 674367 937474 674368 937538
rect 674432 937474 674433 937538
rect 674367 937473 674433 937474
rect 674562 933987 674622 962485
rect 674751 961514 674817 961515
rect 674751 961450 674752 961514
rect 674816 961450 674817 961514
rect 674751 961449 674817 961450
rect 674559 933986 674625 933987
rect 674559 933922 674560 933986
rect 674624 933922 674625 933986
rect 674559 933921 674625 933922
rect 673983 932654 674049 932655
rect 673983 932590 673984 932654
rect 674048 932590 674049 932654
rect 673983 932589 674049 932590
rect 674754 931767 674814 961449
rect 674946 936059 675006 962781
rect 675138 936651 675198 964853
rect 675714 961071 675774 967369
rect 676095 965658 676161 965659
rect 676095 965594 676096 965658
rect 676160 965594 676161 965658
rect 676095 965593 676161 965594
rect 675711 961070 675777 961071
rect 675711 961006 675712 961070
rect 675776 961006 675777 961070
rect 675711 961005 675777 961006
rect 675327 959146 675393 959147
rect 675327 959082 675328 959146
rect 675392 959082 675393 959146
rect 675327 959081 675393 959082
rect 675135 936650 675201 936651
rect 675135 936586 675136 936650
rect 675200 936586 675201 936650
rect 675135 936585 675201 936586
rect 674943 936058 675009 936059
rect 674943 935994 674944 936058
rect 675008 935994 675009 936058
rect 674943 935993 675009 935994
rect 675330 935615 675390 959081
rect 675519 957666 675585 957667
rect 675519 957602 675520 957666
rect 675584 957602 675585 957666
rect 675519 957601 675585 957602
rect 675327 935614 675393 935615
rect 675327 935550 675328 935614
rect 675392 935550 675393 935614
rect 675327 935549 675393 935550
rect 675522 932359 675582 957601
rect 675519 932358 675585 932359
rect 675519 932294 675520 932358
rect 675584 932294 675585 932358
rect 675519 932293 675585 932294
rect 674751 931766 674817 931767
rect 674751 931702 674752 931766
rect 674816 931702 674817 931766
rect 674751 931701 674817 931702
rect 671662 917844 675044 917976
rect 671662 912320 671794 917844
rect 674916 912320 675044 917844
rect 671662 912226 675044 912320
rect 669318 832428 671202 832446
rect 668718 832382 671202 832428
rect 668718 819526 668858 832382
rect 670730 819526 671202 832382
rect 668718 819410 671202 819526
rect 665024 769345 666067 770527
rect 667249 769345 668306 770527
rect 665024 725405 668306 769345
rect 665024 724223 666067 725405
rect 667249 724223 668306 725405
rect 665024 680803 668306 724223
rect 665024 679621 666067 680803
rect 667249 679621 668306 680803
rect 665024 635485 668306 679621
rect 665024 634303 666067 635485
rect 667249 634303 668306 635485
rect 665024 589137 668306 634303
rect 665024 587955 666067 589137
rect 667249 587955 668306 589137
rect 665024 545495 668306 587955
rect 665024 544313 666067 545495
rect 667249 544313 668306 545495
rect 665024 501273 668306 544313
rect 665024 500091 666067 501273
rect 667249 500091 668306 501273
rect 665024 474086 668306 500091
rect 665000 473848 668306 474086
rect 665000 460522 665144 473848
rect 668046 460522 668306 473848
rect 665000 460284 668306 460522
rect 661102 410033 662179 411215
rect 663361 410033 664196 411215
rect 661102 366061 664196 410033
rect 661102 364879 662179 366061
rect 663361 364879 664196 366061
rect 661102 320471 664196 364879
rect 661102 319289 662179 320471
rect 663361 319289 664196 320471
rect 661102 275227 664196 319289
rect 661102 274045 662179 275227
rect 663361 274045 664196 275227
rect 661102 264314 664196 274045
rect 665024 412999 668306 460284
rect 665024 411817 666067 412999
rect 667249 411817 668306 412999
rect 665024 367915 668306 411817
rect 665024 366733 666067 367915
rect 667249 366733 668306 367915
rect 665024 322605 668306 366733
rect 665024 321423 666067 322605
rect 667249 321423 668306 322605
rect 665024 277999 668306 321423
rect 665024 276817 666067 277999
rect 667249 276817 668306 277999
rect 665024 275208 666084 276817
rect 667226 275208 668306 276817
rect 665024 267722 668306 275208
rect 669318 819382 671202 819410
rect 669318 518424 670414 819382
rect 671662 817994 673462 912226
rect 674751 877006 674817 877007
rect 674751 876942 674752 877006
rect 674816 876942 674817 877006
rect 674751 876941 674817 876942
rect 673983 876562 674049 876563
rect 673983 876498 673984 876562
rect 674048 876498 674049 876562
rect 673983 876497 674049 876498
rect 669318 518422 669372 518424
rect 669318 514106 669368 518422
rect 669318 504232 669372 514106
rect 670344 508462 670414 518424
rect 670350 504232 670414 508462
rect 669318 270706 670414 504232
rect 670882 771920 673462 817994
rect 670882 770828 671683 771920
rect 672775 770828 673462 771920
rect 670882 727724 673462 770828
rect 673986 755795 674046 876497
rect 674559 875822 674625 875823
rect 674559 875758 674560 875822
rect 674624 875758 674625 875822
rect 674559 875757 674625 875758
rect 674175 874194 674241 874195
rect 674175 874130 674176 874194
rect 674240 874130 674241 874194
rect 674175 874129 674241 874130
rect 674178 757423 674238 874129
rect 674367 872862 674433 872863
rect 674367 872798 674368 872862
rect 674432 872798 674433 872862
rect 674367 872797 674433 872798
rect 674175 757422 674241 757423
rect 674175 757358 674176 757422
rect 674240 757358 674241 757422
rect 674175 757357 674241 757358
rect 673983 755794 674049 755795
rect 673983 755730 673984 755794
rect 674048 755730 674049 755794
rect 673983 755729 674049 755730
rect 674370 754759 674430 872797
rect 674562 759347 674622 875757
rect 674559 759346 674625 759347
rect 674559 759282 674560 759346
rect 674624 759282 674625 759346
rect 674559 759281 674625 759282
rect 674754 758311 674814 876941
rect 675714 875971 675774 961005
rect 675903 960182 675969 960183
rect 675903 960118 675904 960182
rect 675968 960118 675969 960182
rect 675903 960117 675969 960118
rect 675711 875970 675777 875971
rect 675711 875906 675712 875970
rect 675776 875906 675777 875970
rect 675711 875905 675777 875906
rect 675906 875675 675966 960117
rect 676098 934579 676158 965593
rect 676287 962254 676353 962255
rect 676287 962190 676288 962254
rect 676352 962190 676353 962254
rect 676287 962189 676353 962190
rect 676095 934578 676161 934579
rect 676095 934514 676096 934578
rect 676160 934514 676161 934578
rect 676095 934513 676161 934514
rect 676290 933395 676350 962189
rect 677055 953522 677121 953523
rect 677055 953458 677056 953522
rect 677120 953458 677121 953522
rect 677055 953457 677121 953458
rect 676863 953374 676929 953375
rect 676863 953310 676864 953374
rect 676928 953310 676929 953374
rect 676863 953309 676929 953310
rect 676287 933394 676353 933395
rect 676287 933330 676288 933394
rect 676352 933330 676353 933394
rect 676287 933329 676353 933330
rect 676866 930731 676926 953309
rect 677058 931323 677118 953457
rect 699410 950873 700506 950874
rect 699410 949779 699411 950873
rect 700505 949779 700506 950873
rect 699410 949778 700506 949779
rect 699639 939824 699959 949778
rect 709355 949402 710541 949403
rect 709355 948218 709356 949402
rect 710540 948218 710541 949402
rect 709355 948217 710541 948218
rect 700959 947417 701279 947438
rect 700801 947416 701987 947417
rect 700801 946232 700802 947416
rect 701986 946232 701987 947416
rect 700801 946231 701987 946232
rect 700959 938506 701279 946231
rect 708037 945492 709223 945493
rect 708037 944308 708038 945492
rect 709222 944308 709223 945492
rect 708037 944307 709223 944308
rect 708583 938682 708903 944307
rect 709903 940030 710223 948217
rect 677055 931322 677121 931323
rect 677055 931258 677056 931322
rect 677120 931258 677121 931322
rect 677055 931257 677121 931258
rect 676863 930730 676929 930731
rect 676863 930666 676864 930730
rect 676928 930666 676929 930730
rect 676863 930665 676929 930666
rect 675903 875674 675969 875675
rect 675903 875610 675904 875674
rect 675968 875610 675969 875674
rect 675903 875609 675969 875610
rect 674943 873454 675009 873455
rect 674943 873390 674944 873454
rect 675008 873390 675009 873454
rect 674943 873389 675009 873390
rect 674751 758310 674817 758311
rect 674751 758246 674752 758310
rect 674816 758246 674817 758310
rect 674751 758245 674817 758246
rect 674946 755647 675006 873389
rect 675135 869902 675201 869903
rect 675135 869838 675136 869902
rect 675200 869838 675201 869902
rect 675135 869837 675201 869838
rect 675138 757275 675198 869837
rect 675327 864722 675393 864723
rect 675327 864658 675328 864722
rect 675392 864658 675393 864722
rect 675327 864657 675393 864658
rect 675330 758903 675390 864657
rect 675903 788058 675969 788059
rect 675903 787994 675904 788058
rect 675968 787994 675969 788058
rect 675903 787993 675969 787994
rect 675519 787170 675585 787171
rect 675519 787106 675520 787170
rect 675584 787106 675585 787170
rect 675519 787105 675585 787106
rect 675327 758902 675393 758903
rect 675327 758838 675328 758902
rect 675392 758838 675393 758902
rect 675327 758837 675393 758838
rect 675135 757274 675201 757275
rect 675135 757210 675136 757274
rect 675200 757210 675201 757274
rect 675135 757209 675201 757210
rect 674943 755646 675009 755647
rect 674943 755582 674944 755646
rect 675008 755582 675009 755646
rect 674943 755581 675009 755582
rect 674367 754758 674433 754759
rect 674367 754694 674368 754758
rect 674432 754694 674433 754758
rect 674367 754693 674433 754694
rect 674175 743214 674241 743215
rect 674175 743150 674176 743214
rect 674240 743150 674241 743214
rect 674175 743149 674241 743150
rect 673983 742474 674049 742475
rect 673983 742410 673984 742474
rect 674048 742410 674049 742474
rect 673983 742409 674049 742410
rect 670882 726632 671683 727724
rect 672775 726632 673462 727724
rect 670882 682316 673462 726632
rect 670882 681224 671683 682316
rect 672775 681224 673462 682316
rect 670882 636972 673462 681224
rect 673986 665663 674046 742409
rect 674178 667809 674238 743149
rect 674367 741734 674433 741735
rect 674367 741670 674368 741734
rect 674432 741670 674433 741734
rect 674367 741669 674433 741670
rect 674370 668919 674430 741669
rect 675135 740106 675201 740107
rect 675135 740042 675136 740106
rect 675200 740042 675201 740106
rect 675135 740041 675201 740042
rect 674943 739218 675009 739219
rect 674943 739154 674944 739218
rect 675008 739154 675009 739218
rect 674943 739153 675009 739154
rect 674751 738626 674817 738627
rect 674751 738562 674752 738626
rect 674816 738562 674817 738626
rect 674751 738561 674817 738562
rect 674559 694374 674625 694375
rect 674559 694310 674560 694374
rect 674624 694310 674625 694374
rect 674559 694309 674625 694310
rect 674367 668918 674433 668919
rect 674367 668854 674368 668918
rect 674432 668854 674433 668918
rect 674367 668853 674433 668854
rect 674175 667808 674241 667809
rect 674175 667744 674176 667808
rect 674240 667744 674241 667808
rect 674175 667743 674241 667744
rect 673983 665662 674049 665663
rect 673983 665598 673984 665662
rect 674048 665598 674049 665662
rect 673983 665597 674049 665598
rect 674175 652194 674241 652195
rect 674175 652130 674176 652194
rect 674240 652130 674241 652194
rect 674175 652129 674241 652130
rect 673983 649826 674049 649827
rect 673983 649762 673984 649826
rect 674048 649762 674049 649826
rect 673983 649761 674049 649762
rect 673986 641055 674046 649761
rect 670882 635880 671683 636972
rect 672775 635880 673462 636972
rect 670882 592642 673462 635880
rect 673794 640995 674046 641055
rect 673794 630883 673854 640995
rect 673983 640354 674049 640355
rect 673983 640290 673984 640354
rect 674048 640290 674049 640354
rect 673983 640289 674049 640290
rect 673791 630882 673857 630883
rect 673791 630818 673792 630882
rect 673856 630818 673857 630882
rect 673791 630817 673857 630818
rect 673986 613715 674046 640289
rect 673983 613714 674049 613715
rect 673983 613650 673984 613714
rect 674048 613650 674049 613714
rect 673983 613649 674049 613650
rect 673983 607794 674049 607795
rect 673983 607730 673984 607794
rect 674048 607730 674049 607794
rect 673983 607729 674049 607730
rect 670882 591550 671683 592642
rect 672775 591550 673462 592642
rect 670882 547150 673462 591550
rect 670882 546058 671683 547150
rect 672775 546058 673462 547150
rect 670882 503088 673462 546058
rect 673986 532611 674046 607729
rect 674178 575383 674238 652129
rect 674367 648938 674433 648939
rect 674367 648874 674368 648938
rect 674432 648874 674433 648938
rect 674367 648873 674433 648874
rect 674370 630735 674430 648873
rect 674367 630734 674433 630735
rect 674367 630670 674368 630734
rect 674432 630670 674433 630734
rect 674367 630669 674433 630670
rect 674562 620375 674622 694309
rect 674754 664923 674814 738561
rect 674946 665367 675006 739153
rect 675138 667587 675198 740041
rect 675327 734482 675393 734483
rect 675327 734418 675328 734482
rect 675392 734418 675393 734482
rect 675327 734417 675393 734418
rect 675330 697039 675390 734417
rect 675522 711099 675582 787105
rect 675711 784210 675777 784211
rect 675711 784146 675712 784210
rect 675776 784146 675777 784210
rect 675711 784145 675777 784146
rect 675519 711098 675585 711099
rect 675519 711034 675520 711098
rect 675584 711034 675585 711098
rect 675519 711033 675585 711034
rect 675714 710655 675774 784145
rect 675906 713319 675966 787993
rect 676095 786726 676161 786727
rect 676095 786662 676096 786726
rect 676160 786662 676161 786726
rect 676095 786661 676161 786662
rect 676098 714355 676158 786661
rect 676287 784950 676353 784951
rect 676287 784886 676288 784950
rect 676352 784886 676353 784950
rect 676287 784885 676353 784886
rect 676095 714354 676161 714355
rect 676095 714290 676096 714354
rect 676160 714290 676161 714354
rect 676095 714289 676161 714290
rect 675903 713318 675969 713319
rect 675903 713254 675904 713318
rect 675968 713254 675969 713318
rect 675903 713253 675969 713254
rect 676290 712727 676350 784885
rect 676671 781990 676737 781991
rect 676671 781926 676672 781990
rect 676736 781926 676737 781990
rect 676671 781925 676737 781926
rect 676479 780658 676545 780659
rect 676479 780594 676480 780658
rect 676544 780594 676545 780658
rect 676479 780593 676545 780594
rect 676287 712726 676353 712727
rect 676287 712662 676288 712726
rect 676352 712662 676353 712726
rect 676287 712661 676353 712662
rect 676482 712283 676542 780593
rect 676674 740403 676734 781925
rect 677058 777551 677502 777585
rect 677055 777550 677502 777551
rect 677055 777486 677056 777550
rect 677120 777525 677502 777550
rect 677120 777486 677121 777525
rect 677055 777485 677121 777486
rect 677055 776958 677121 776959
rect 677055 776894 677056 776958
rect 677120 776919 677121 776958
rect 677120 776894 677310 776919
rect 677055 776893 677310 776894
rect 677058 776859 677310 776893
rect 677055 776218 677121 776219
rect 677055 776154 677056 776218
rect 677120 776154 677121 776218
rect 677055 776153 677121 776154
rect 676863 774886 676929 774887
rect 676863 774822 676864 774886
rect 676928 774822 676929 774886
rect 676863 774821 676929 774822
rect 676866 756683 676926 774821
rect 677058 760383 677118 776153
rect 677055 760382 677121 760383
rect 677055 760318 677056 760382
rect 677120 760318 677121 760382
rect 677055 760317 677121 760318
rect 676863 756682 676929 756683
rect 676863 756618 676864 756682
rect 676928 756618 676929 756682
rect 676863 756617 676929 756618
rect 676863 756090 676929 756091
rect 676863 756026 676864 756090
rect 676928 756026 676929 756090
rect 676863 756025 676929 756026
rect 676866 744547 676926 756025
rect 677250 753427 677310 776859
rect 677442 754463 677502 777525
rect 677631 773110 677697 773111
rect 677631 773046 677632 773110
rect 677696 773046 677697 773110
rect 677631 773045 677697 773046
rect 677439 754462 677505 754463
rect 677439 754398 677440 754462
rect 677504 754398 677505 754462
rect 677439 754397 677505 754398
rect 677634 754019 677694 773045
rect 699639 771922 699959 771996
rect 699228 771921 700324 771922
rect 699228 770827 699229 771921
rect 700323 770827 700324 771921
rect 699228 770826 700324 770827
rect 699639 761526 699959 770826
rect 709903 770529 710223 770582
rect 709389 770528 710575 770529
rect 709389 769344 709390 770528
rect 710574 769344 710575 770528
rect 709389 769343 710575 769344
rect 700827 768630 702013 768631
rect 700827 767446 700828 768630
rect 702012 767446 702013 768630
rect 700827 767445 702013 767446
rect 700959 760316 701279 767445
rect 708583 766961 708903 767008
rect 707977 766960 709163 766961
rect 707977 765776 707978 766960
rect 709162 765776 709163 766960
rect 707977 765775 709163 765776
rect 708583 760372 708903 765775
rect 709903 761756 710223 769343
rect 677823 759938 677889 759939
rect 677823 759874 677824 759938
rect 677888 759874 677889 759938
rect 677823 759873 677889 759874
rect 677631 754018 677697 754019
rect 677631 753954 677632 754018
rect 677696 753954 677697 754018
rect 677631 753953 677697 753954
rect 677247 753426 677313 753427
rect 677247 753362 677248 753426
rect 677312 753362 677313 753426
rect 677247 753361 677313 753362
rect 677631 753426 677697 753427
rect 677631 753362 677632 753426
rect 677696 753362 677697 753426
rect 677631 753361 677697 753362
rect 676863 744546 676929 744547
rect 676863 744482 676864 744546
rect 676928 744482 676929 744546
rect 676863 744481 676929 744482
rect 677247 744546 677313 744547
rect 677247 744482 677248 744546
rect 677312 744482 677313 744546
rect 677247 744481 677313 744482
rect 676863 744398 676929 744399
rect 676863 744334 676864 744398
rect 676928 744334 676929 744398
rect 676863 744333 676929 744334
rect 676671 740402 676737 740403
rect 676671 740338 676672 740402
rect 676736 740338 676737 740402
rect 676671 740337 676737 740338
rect 676866 734295 676926 744333
rect 676674 734235 676926 734295
rect 676674 726047 676734 734235
rect 677250 733000 677310 744481
rect 677634 744399 677694 753361
rect 677826 752835 677886 759873
rect 677823 752834 677889 752835
rect 677823 752770 677824 752834
rect 677888 752770 677889 752834
rect 677823 752769 677889 752770
rect 677631 744398 677697 744399
rect 677631 744334 677632 744398
rect 677696 744334 677697 744398
rect 677631 744333 677697 744334
rect 676866 732940 677310 733000
rect 676671 726046 676737 726047
rect 676671 725982 676672 726046
rect 676736 725982 676737 726046
rect 676671 725981 676737 725982
rect 676866 715539 676926 732940
rect 677247 728118 677313 728119
rect 677247 728054 677248 728118
rect 677312 728054 677313 728118
rect 677247 728053 677313 728054
rect 676863 715538 676929 715539
rect 676863 715474 676864 715538
rect 676928 715474 676929 715538
rect 676863 715473 676929 715474
rect 677055 714354 677121 714355
rect 677055 714290 677056 714354
rect 677120 714290 677121 714354
rect 677055 714289 677121 714290
rect 676479 712282 676545 712283
rect 676479 712218 676480 712282
rect 676544 712218 676545 712282
rect 676479 712217 676545 712218
rect 675711 710654 675777 710655
rect 675711 710590 675712 710654
rect 675776 710590 675777 710654
rect 675711 710589 675777 710590
rect 675519 697926 675585 697927
rect 675519 697862 675520 697926
rect 675584 697862 675585 697926
rect 675519 697861 675585 697862
rect 675327 697038 675393 697039
rect 675327 696974 675328 697038
rect 675392 696974 675393 697038
rect 675327 696973 675393 696974
rect 675327 696890 675393 696891
rect 675327 696826 675328 696890
rect 675392 696826 675393 696890
rect 675327 696825 675393 696826
rect 675135 667586 675201 667587
rect 675135 667522 675136 667586
rect 675200 667522 675201 667586
rect 675135 667521 675201 667522
rect 674943 665366 675009 665367
rect 674943 665302 674944 665366
rect 675008 665302 675009 665366
rect 674943 665301 675009 665302
rect 674751 664922 674817 664923
rect 674751 664858 674752 664922
rect 674816 664858 674817 664922
rect 674751 664857 674817 664858
rect 674751 652638 674817 652639
rect 674751 652574 674752 652638
rect 674816 652574 674817 652638
rect 674751 652573 674817 652574
rect 674754 649827 674814 652573
rect 675135 651454 675201 651455
rect 675135 651390 675136 651454
rect 675200 651390 675201 651454
rect 675135 651389 675201 651390
rect 674751 649826 674817 649827
rect 674751 649762 674752 649826
rect 674816 649762 674817 649826
rect 674751 649761 674817 649762
rect 674751 649678 674817 649679
rect 674751 649614 674752 649678
rect 674816 649614 674817 649678
rect 674751 649613 674817 649614
rect 674559 620374 674625 620375
rect 674559 620310 674560 620374
rect 674624 620310 674625 620374
rect 674559 620309 674625 620310
rect 674559 619930 674625 619931
rect 674559 619866 674560 619930
rect 674624 619866 674625 619930
rect 674559 619865 674625 619866
rect 674367 604834 674433 604835
rect 674367 604770 674368 604834
rect 674432 604770 674433 604834
rect 674367 604769 674433 604770
rect 674175 575382 674241 575383
rect 674175 575318 674176 575382
rect 674240 575318 674241 575382
rect 674175 575317 674241 575318
rect 674175 562062 674241 562063
rect 674175 561998 674176 562062
rect 674240 561998 674241 562062
rect 674175 561997 674241 561998
rect 673983 532610 674049 532611
rect 673983 532546 673984 532610
rect 674048 532546 674049 532610
rect 673983 532545 674049 532546
rect 670882 501996 671683 503088
rect 672775 501996 673462 503088
rect 670882 414948 673462 501996
rect 674178 486435 674238 561997
rect 674370 532019 674430 604769
rect 674562 590627 674622 619865
rect 674754 613863 674814 649613
rect 674943 630882 675009 630883
rect 674943 630818 674944 630882
rect 675008 630818 675009 630882
rect 674943 630817 675009 630818
rect 674946 621075 675006 630817
rect 675138 630735 675198 651389
rect 675135 630734 675201 630735
rect 675135 630670 675136 630734
rect 675200 630670 675201 630734
rect 675135 630669 675201 630670
rect 675330 624223 675390 696825
rect 675327 624222 675393 624223
rect 675327 624158 675328 624222
rect 675392 624158 675393 624222
rect 675327 624157 675393 624158
rect 675522 623187 675582 697861
rect 676671 697334 676737 697335
rect 676671 697270 676672 697334
rect 676736 697270 676737 697334
rect 676671 697269 676737 697270
rect 676287 697038 676353 697039
rect 676287 696974 676288 697038
rect 676352 696974 676353 697038
rect 676287 696973 676353 696974
rect 675711 694818 675777 694819
rect 675711 694754 675712 694818
rect 675776 694754 675777 694818
rect 675711 694753 675777 694754
rect 675519 623186 675585 623187
rect 675519 623122 675520 623186
rect 675584 623122 675585 623186
rect 675519 623121 675585 623122
rect 675714 622595 675774 694753
rect 675903 689194 675969 689195
rect 675903 689130 675904 689194
rect 675968 689130 675969 689194
rect 675903 689129 675969 689130
rect 675711 622594 675777 622595
rect 675711 622530 675712 622594
rect 675776 622530 675777 622594
rect 675711 622529 675777 622530
rect 674946 621015 675390 621075
rect 674943 620818 675009 620819
rect 674943 620754 674944 620818
rect 675008 620754 675009 620818
rect 674943 620753 675009 620754
rect 674751 613862 674817 613863
rect 674751 613798 674752 613862
rect 674816 613798 674817 613862
rect 674751 613797 674817 613798
rect 674751 594770 674817 594771
rect 674751 594706 674752 594770
rect 674816 594706 674817 594770
rect 674751 594705 674817 594706
rect 674559 590626 674625 590627
rect 674559 590562 674560 590626
rect 674624 590562 674625 590626
rect 674559 590561 674625 590562
rect 674559 590330 674625 590331
rect 674559 590266 674560 590330
rect 674624 590266 674625 590330
rect 674754 590328 674814 594705
rect 674946 590923 675006 620753
rect 675135 607202 675201 607203
rect 675135 607138 675136 607202
rect 675200 607138 675201 607202
rect 675135 607137 675201 607138
rect 674943 590922 675009 590923
rect 674943 590858 674944 590922
rect 675008 590858 675009 590922
rect 674943 590857 675009 590858
rect 675138 590331 675198 607137
rect 675330 606611 675390 621015
rect 675906 618747 675966 689129
rect 676095 688306 676161 688307
rect 676095 688242 676096 688306
rect 676160 688242 676161 688306
rect 676095 688241 676161 688242
rect 676098 619931 676158 688241
rect 676290 663739 676350 696973
rect 676479 692006 676545 692007
rect 676479 691942 676480 692006
rect 676544 691942 676545 692006
rect 676479 691941 676545 691942
rect 676287 663738 676353 663739
rect 676287 663674 676288 663738
rect 676352 663674 676353 663738
rect 676287 663673 676353 663674
rect 676482 653675 676542 691941
rect 676479 653674 676545 653675
rect 676479 653610 676480 653674
rect 676544 653610 676545 653674
rect 676479 653609 676545 653610
rect 676287 645386 676353 645387
rect 676287 645322 676288 645386
rect 676352 645322 676353 645386
rect 676287 645321 676353 645322
rect 676095 619930 676161 619931
rect 676095 619866 676096 619930
rect 676160 619866 676161 619930
rect 676095 619865 676161 619866
rect 675903 618746 675969 618747
rect 675903 618682 675904 618746
rect 675968 618682 675969 618746
rect 675903 618681 675969 618682
rect 676095 613862 676161 613863
rect 676095 613798 676096 613862
rect 676160 613798 676161 613862
rect 676095 613797 676161 613798
rect 675519 613714 675585 613715
rect 675519 613650 675520 613714
rect 675584 613650 675585 613714
rect 675519 613649 675585 613650
rect 675327 606610 675393 606611
rect 675327 606546 675328 606610
rect 675392 606546 675393 606610
rect 675327 606545 675393 606546
rect 675327 606462 675393 606463
rect 675327 606398 675328 606462
rect 675392 606398 675393 606462
rect 675327 606397 675393 606398
rect 675135 590330 675201 590331
rect 674754 590268 675006 590328
rect 674559 590265 674625 590266
rect 674367 532018 674433 532019
rect 674367 531954 674368 532018
rect 674432 531954 674433 532018
rect 674367 531953 674433 531954
rect 674562 530687 674622 590265
rect 674751 590182 674817 590183
rect 674751 590118 674752 590182
rect 674816 590118 674817 590182
rect 674751 590117 674817 590118
rect 674754 575235 674814 590117
rect 674946 577899 675006 590268
rect 675135 590266 675136 590330
rect 675200 590266 675201 590330
rect 675135 590265 675201 590266
rect 675135 590034 675201 590035
rect 675135 589970 675136 590034
rect 675200 589970 675201 590034
rect 675135 589969 675201 589970
rect 674943 577898 675009 577899
rect 674943 577834 674944 577898
rect 675008 577834 675009 577898
rect 674943 577833 675009 577834
rect 675138 576271 675198 589969
rect 675135 576270 675201 576271
rect 675135 576206 675136 576270
rect 675200 576206 675201 576270
rect 675135 576205 675201 576206
rect 674751 575234 674817 575235
rect 674751 575170 674752 575234
rect 674816 575170 674817 575234
rect 674751 575169 674817 575170
rect 674943 562506 675009 562507
rect 674943 562442 674944 562506
rect 675008 562442 675009 562506
rect 674943 562441 675009 562442
rect 674751 558954 674817 558955
rect 674751 558890 674752 558954
rect 674816 558890 674817 558954
rect 674751 558889 674817 558890
rect 674559 530686 674625 530687
rect 674559 530622 674560 530686
rect 674624 530622 674625 530686
rect 674559 530621 674625 530622
rect 674175 486434 674241 486435
rect 674175 486370 674176 486434
rect 674240 486370 674241 486434
rect 674175 486369 674241 486370
rect 674754 486139 674814 558889
rect 674946 488951 675006 562441
rect 675135 561470 675201 561471
rect 675135 561406 675136 561470
rect 675200 561406 675201 561470
rect 675135 561405 675201 561406
rect 675138 489987 675198 561405
rect 675330 533943 675390 606397
rect 675522 600543 675582 613649
rect 675903 606610 675969 606611
rect 675903 606546 675904 606610
rect 675968 606546 675969 606610
rect 675903 606545 675969 606546
rect 675519 600542 675585 600543
rect 675519 600478 675520 600542
rect 675584 600478 675585 600542
rect 675519 600477 675585 600478
rect 675906 594771 675966 606545
rect 676098 595511 676158 613797
rect 676095 595510 676161 595511
rect 676095 595446 676096 595510
rect 676160 595446 676161 595510
rect 676095 595445 676161 595446
rect 676095 595362 676161 595363
rect 676095 595298 676096 595362
rect 676160 595298 676161 595362
rect 676095 595297 676161 595298
rect 675903 594770 675969 594771
rect 675903 594706 675904 594770
rect 675968 594706 675969 594770
rect 675903 594705 675969 594706
rect 675903 593438 675969 593439
rect 675903 593374 675904 593438
rect 675968 593374 675969 593438
rect 675903 593373 675969 593374
rect 675711 590478 675777 590479
rect 675711 590414 675712 590478
rect 675776 590414 675777 590478
rect 675711 590413 675777 590414
rect 675519 590330 675585 590331
rect 675519 590266 675520 590330
rect 675584 590266 675585 590330
rect 675519 590265 675585 590266
rect 675522 577307 675582 590265
rect 675519 577306 675585 577307
rect 675519 577242 675520 577306
rect 675584 577242 675585 577306
rect 675519 577241 675585 577242
rect 675327 533942 675393 533943
rect 675327 533878 675328 533942
rect 675392 533878 675393 533942
rect 675327 533877 675393 533878
rect 675714 531871 675774 590413
rect 675711 531870 675777 531871
rect 675711 531806 675712 531870
rect 675776 531806 675777 531870
rect 675711 531805 675777 531806
rect 675906 531279 675966 593373
rect 676098 533499 676158 595297
rect 676290 576863 676350 645321
rect 676479 638578 676545 638579
rect 676479 638514 676480 638578
rect 676544 638514 676545 638578
rect 676479 638513 676545 638514
rect 676482 590035 676542 638513
rect 676674 620967 676734 697269
rect 677058 669659 677118 714289
rect 677250 711691 677310 728053
rect 699639 727726 699959 727798
rect 699314 727725 700410 727726
rect 699314 726631 699315 727725
rect 700409 726631 700410 727725
rect 699314 726630 700410 726631
rect 677439 725898 677505 725899
rect 677439 725834 677440 725898
rect 677504 725834 677505 725898
rect 677439 725833 677505 725834
rect 677442 718977 677502 725833
rect 677442 718917 677694 718977
rect 677634 714947 677694 718917
rect 699639 716578 699959 726630
rect 709903 725407 710223 725448
rect 709349 725406 710535 725407
rect 709349 724222 709350 725406
rect 710534 724222 710535 725406
rect 709349 724221 710535 724222
rect 700685 723372 701871 723373
rect 700685 722188 700686 723372
rect 701870 722188 701871 723372
rect 700685 722187 701871 722188
rect 700959 715078 701279 722187
rect 708583 721283 708903 721286
rect 708075 721282 709261 721283
rect 708075 720098 708076 721282
rect 709260 720098 709261 721282
rect 708075 720097 709261 720098
rect 708583 715418 708903 720097
rect 709903 716266 710223 724221
rect 677439 714946 677505 714947
rect 677439 714882 677440 714946
rect 677504 714882 677505 714946
rect 677439 714881 677505 714882
rect 677631 714946 677697 714947
rect 677631 714882 677632 714946
rect 677696 714882 677697 714946
rect 677631 714881 677697 714882
rect 677247 711690 677313 711691
rect 677247 711626 677248 711690
rect 677312 711626 677313 711690
rect 677247 711625 677313 711626
rect 677442 670251 677502 714881
rect 699120 682317 700216 682318
rect 699120 681223 699121 682317
rect 700215 681223 700216 682317
rect 699120 681222 700216 681223
rect 699639 671100 699959 681222
rect 709903 680805 710223 680814
rect 709417 680804 710603 680805
rect 709417 679620 709418 680804
rect 710602 679620 710603 680804
rect 709417 679619 710603 679620
rect 700497 678968 701683 678969
rect 700497 677784 700498 678968
rect 701682 677784 701683 678968
rect 700497 677783 701683 677784
rect 677247 670250 677313 670251
rect 677247 670186 677248 670250
rect 677312 670186 677313 670250
rect 677247 670185 677313 670186
rect 677439 670250 677505 670251
rect 677439 670186 677440 670250
rect 677504 670186 677505 670250
rect 677439 670185 677505 670186
rect 677055 669658 677121 669659
rect 677055 669594 677056 669658
rect 677120 669594 677121 669658
rect 677055 669593 677121 669594
rect 677058 624667 677118 669593
rect 677250 626443 677310 670185
rect 677247 626442 677313 626443
rect 677247 626378 677248 626442
rect 677312 626378 677313 626442
rect 677247 626377 677313 626378
rect 677442 625222 677502 670185
rect 700959 669678 701279 677783
rect 708583 677245 708903 677384
rect 708329 677244 709515 677245
rect 708329 676060 708330 677244
rect 709514 676060 709515 677244
rect 708329 676059 709515 676060
rect 708583 670626 708903 676059
rect 709903 671238 710223 679619
rect 699639 636974 699959 637076
rect 699308 636973 700404 636974
rect 699308 635879 699309 636973
rect 700403 635879 700404 636973
rect 699308 635878 700404 635879
rect 699639 626174 699959 635878
rect 709903 635487 710223 635496
rect 709373 635486 710559 635487
rect 709373 634302 709374 635486
rect 710558 634302 710559 635486
rect 709373 634301 710559 634302
rect 700959 633627 701279 633724
rect 700649 633626 701835 633627
rect 700649 632442 700650 633626
rect 701834 632442 701835 633626
rect 700649 632441 701835 632442
rect 677439 625221 677505 625222
rect 677439 625157 677440 625221
rect 677504 625157 677505 625221
rect 677439 625156 677505 625157
rect 700959 624844 701279 632441
rect 708583 630017 708903 630096
rect 708127 630016 709313 630017
rect 708127 628832 708128 630016
rect 709312 628832 709313 630016
rect 708127 628831 709313 628832
rect 708583 625592 708903 628831
rect 709903 626146 710223 634301
rect 677055 624666 677121 624667
rect 677055 624602 677056 624666
rect 677120 624602 677121 624666
rect 677055 624601 677121 624602
rect 676671 620966 676737 620967
rect 676671 620902 676672 620966
rect 676736 620902 676737 620966
rect 676671 620901 676737 620902
rect 676671 600542 676737 600543
rect 676671 600478 676672 600542
rect 676736 600478 676737 600542
rect 676671 600477 676737 600478
rect 676674 591105 676734 600477
rect 699394 592643 700490 592644
rect 699394 591549 699395 592643
rect 700489 591549 700490 592643
rect 699394 591548 700490 591549
rect 676674 591045 676926 591105
rect 676671 590922 676737 590923
rect 676671 590858 676672 590922
rect 676736 590858 676737 590922
rect 676671 590857 676737 590858
rect 676479 590034 676545 590035
rect 676479 589970 676480 590034
rect 676544 589970 676545 590034
rect 676479 589969 676545 589970
rect 676479 589886 676545 589887
rect 676479 589822 676480 589886
rect 676544 589822 676545 589886
rect 676479 589821 676545 589822
rect 676482 578491 676542 589821
rect 676674 578935 676734 590857
rect 676866 589887 676926 591045
rect 676863 589886 676929 589887
rect 676863 589822 676864 589886
rect 676928 589822 676929 589886
rect 676863 589821 676929 589822
rect 699639 581092 699959 591548
rect 709903 589139 710223 589352
rect 709313 589138 710499 589139
rect 709313 587954 709314 589138
rect 710498 587954 710499 589138
rect 709313 587953 710499 587954
rect 700959 587357 701279 587402
rect 700809 587356 701995 587357
rect 700809 586172 700810 587356
rect 701994 586172 701995 587356
rect 700809 586171 701995 586172
rect 700959 580014 701279 586171
rect 708583 585087 708903 585234
rect 708067 585086 709253 585087
rect 708067 583902 708068 585086
rect 709252 583902 709253 585086
rect 708067 583901 709253 583902
rect 708583 580312 708903 583901
rect 709903 580906 710223 587953
rect 677247 579526 677313 579527
rect 677247 579462 677248 579526
rect 677312 579462 677313 579526
rect 677247 579461 677313 579462
rect 677055 579082 677121 579083
rect 677055 579018 677056 579082
rect 677120 579018 677121 579082
rect 677055 579017 677121 579018
rect 676671 578934 676737 578935
rect 676671 578870 676672 578934
rect 676736 578870 676737 578934
rect 676671 578869 676737 578870
rect 676479 578490 676545 578491
rect 676479 578426 676480 578490
rect 676544 578426 676545 578490
rect 676479 578425 676545 578426
rect 676287 576862 676353 576863
rect 676287 576798 676288 576862
rect 676352 576798 676353 576862
rect 676287 576797 676353 576798
rect 676863 554514 676929 554515
rect 676863 554450 676864 554514
rect 676928 554450 676929 554514
rect 676863 554449 676929 554450
rect 676095 533498 676161 533499
rect 676095 533434 676096 533498
rect 676160 533434 676161 533498
rect 676095 533433 676161 533434
rect 675903 531278 675969 531279
rect 675903 531214 675904 531278
rect 675968 531214 675969 531278
rect 675903 531213 675969 531214
rect 675135 489986 675201 489987
rect 675135 489922 675136 489986
rect 675200 489922 675201 489986
rect 675135 489921 675201 489922
rect 674943 488950 675009 488951
rect 674943 488886 674944 488950
rect 675008 488886 675009 488950
rect 674943 488885 675009 488886
rect 674751 486138 674817 486139
rect 674751 486074 674752 486138
rect 674816 486074 674817 486138
rect 674751 486073 674817 486074
rect 676866 483475 676926 554449
rect 677058 534535 677118 579017
rect 677250 535127 677310 579461
rect 699204 547151 700300 547152
rect 699204 546057 699205 547151
rect 700299 546057 700300 547151
rect 699204 546056 700300 546057
rect 699639 536080 699959 546056
rect 709903 545497 710223 545596
rect 709417 545496 710603 545497
rect 709417 544312 709418 545496
rect 710602 544312 710603 545496
rect 709417 544311 710603 544312
rect 700959 543903 701279 543948
rect 700595 543902 701781 543903
rect 700595 542718 700596 543902
rect 701780 542718 701781 543902
rect 700595 542717 701781 542718
rect 677247 535126 677313 535127
rect 677247 535062 677248 535126
rect 677312 535062 677313 535126
rect 677247 535061 677313 535062
rect 700959 534752 701279 542717
rect 708583 541883 708903 541980
rect 707929 541882 709115 541883
rect 707929 540698 707930 541882
rect 709114 540698 709115 541882
rect 707929 540697 709115 540698
rect 708583 535230 708903 540697
rect 709903 535814 710223 544311
rect 677055 534534 677121 534535
rect 677055 534470 677056 534534
rect 677120 534470 677121 534534
rect 677055 534469 677121 534470
rect 699152 503089 700248 503090
rect 699152 501995 699153 503089
rect 700247 501995 700248 503089
rect 699152 501994 700248 501995
rect 699639 491912 699959 501994
rect 709903 501275 710223 501532
rect 709151 501274 710337 501275
rect 709151 500090 709152 501274
rect 710336 500090 710337 501274
rect 709151 500089 710337 500090
rect 700595 499414 701781 499415
rect 700595 498230 700596 499414
rect 701780 498230 701781 499414
rect 700595 498229 701781 498230
rect 677823 491022 677889 491023
rect 677823 490958 677824 491022
rect 677888 490958 677889 491022
rect 677823 490957 677889 490958
rect 677631 490578 677697 490579
rect 677631 490514 677632 490578
rect 677696 490514 677697 490578
rect 677631 490513 677697 490514
rect 677439 489986 677505 489987
rect 677439 489922 677440 489986
rect 677504 489922 677505 489986
rect 677439 489921 677505 489922
rect 676863 483474 676929 483475
rect 676863 483410 676864 483474
rect 676928 483410 676929 483474
rect 676863 483409 676929 483410
rect 670882 413856 671683 414948
rect 672775 413856 673462 414948
rect 670882 369980 673462 413856
rect 677442 402223 677502 489921
rect 677634 402815 677694 490513
rect 677826 403999 677886 490957
rect 700959 490688 701279 498229
rect 708035 497500 709221 497501
rect 708035 496316 708036 497500
rect 709220 496316 709221 497500
rect 708035 496315 709221 496316
rect 708583 491432 708903 496315
rect 709903 492230 710223 500089
rect 699208 414949 700304 414950
rect 699208 413855 699209 414949
rect 700303 413855 700304 414949
rect 699208 413854 700304 413855
rect 677823 403998 677889 403999
rect 677823 403934 677824 403998
rect 677888 403934 677889 403998
rect 677823 403933 677889 403934
rect 699639 403380 699959 413854
rect 709903 413001 710223 413106
rect 709365 413000 710551 413001
rect 709365 411816 709366 413000
rect 710550 411816 710551 413000
rect 709365 411815 710551 411816
rect 700719 411216 701905 411217
rect 700719 410032 700720 411216
rect 701904 410032 701905 411216
rect 700719 410031 701905 410032
rect 677631 402814 677697 402815
rect 677631 402750 677632 402814
rect 677696 402750 677697 402814
rect 677631 402749 677697 402750
rect 700959 402716 701279 410031
rect 708099 409432 709285 409433
rect 708099 408248 708100 409432
rect 709284 408248 709285 409432
rect 708099 408247 709285 408248
rect 708583 403032 708903 408247
rect 709903 403770 710223 411815
rect 677439 402222 677505 402223
rect 677439 402158 677440 402222
rect 677504 402158 677505 402222
rect 677439 402157 677505 402158
rect 674559 400594 674625 400595
rect 674559 400530 674560 400594
rect 674624 400530 674625 400594
rect 674559 400529 674625 400530
rect 674367 399262 674433 399263
rect 674367 399198 674368 399262
rect 674432 399198 674433 399262
rect 674367 399197 674433 399198
rect 674175 398818 674241 398819
rect 674175 398754 674176 398818
rect 674240 398754 674241 398818
rect 674175 398753 674241 398754
rect 674178 372031 674238 398753
rect 674370 378839 674430 399197
rect 674367 378838 674433 378839
rect 674367 378774 674368 378838
rect 674432 378774 674433 378838
rect 674367 378773 674433 378774
rect 674562 373955 674622 400529
rect 675327 374546 675393 374547
rect 675327 374482 675328 374546
rect 675392 374482 675393 374546
rect 675327 374481 675393 374482
rect 674559 373954 674625 373955
rect 674559 373890 674560 373954
rect 674624 373890 674625 373954
rect 674559 373889 674625 373890
rect 674175 372030 674241 372031
rect 674175 371966 674176 372030
rect 674240 371966 674241 372030
rect 674175 371965 674241 371966
rect 670882 368888 671683 369980
rect 672775 368888 673462 369980
rect 670882 324236 673462 368888
rect 673983 355750 674049 355751
rect 673983 355686 673984 355750
rect 674048 355686 674049 355750
rect 673983 355685 674049 355686
rect 673986 328371 674046 355685
rect 675330 335031 675390 374481
rect 677055 374398 677121 374399
rect 677055 374334 677056 374398
rect 677120 374334 677121 374398
rect 677055 374333 677121 374334
rect 675519 374102 675585 374103
rect 675519 374038 675520 374102
rect 675584 374038 675585 374102
rect 675519 374037 675585 374038
rect 675327 335030 675393 335031
rect 675327 334966 675328 335030
rect 675392 334966 675393 335030
rect 675327 334965 675393 334966
rect 675522 333847 675582 374037
rect 677058 373989 677118 374333
rect 677058 373929 677310 373989
rect 677055 373066 677121 373067
rect 677055 373002 677056 373066
rect 677120 373002 677121 373066
rect 677055 373001 677121 373002
rect 677058 357675 677118 373001
rect 676863 357674 676929 357675
rect 676863 357610 676864 357674
rect 676928 357610 676929 357674
rect 676863 357609 676929 357610
rect 677055 357674 677121 357675
rect 677055 357610 677056 357674
rect 677120 357610 677121 357674
rect 677055 357609 677121 357610
rect 676479 345538 676545 345539
rect 676479 345474 676480 345538
rect 676544 345474 676545 345538
rect 676479 345473 676545 345474
rect 675519 333846 675585 333847
rect 675519 333782 675520 333846
rect 675584 333782 675585 333846
rect 675519 333781 675585 333782
rect 675327 329554 675393 329555
rect 675327 329490 675328 329554
rect 675392 329490 675393 329554
rect 675327 329489 675393 329490
rect 673983 328370 674049 328371
rect 673983 328306 673984 328370
rect 674048 328306 674049 328370
rect 673983 328305 674049 328306
rect 670882 323144 671683 324236
rect 672775 323144 673462 324236
rect 670882 280948 673462 323144
rect 673983 310758 674049 310759
rect 673983 310694 673984 310758
rect 674048 310694 674049 310758
rect 673983 310693 674049 310694
rect 673986 283675 674046 310693
rect 675330 290039 675390 329489
rect 675327 290038 675393 290039
rect 675327 289974 675328 290038
rect 675392 289974 675393 290038
rect 675327 289973 675393 289974
rect 675522 289595 675582 333781
rect 676482 330591 676542 345473
rect 676671 345390 676737 345391
rect 676671 345326 676672 345390
rect 676736 345326 676737 345390
rect 676671 345325 676737 345326
rect 676479 330590 676545 330591
rect 676479 330526 676480 330590
rect 676544 330526 676545 330590
rect 676479 330525 676545 330526
rect 676674 326891 676734 345325
rect 676671 326890 676737 326891
rect 676671 326826 676672 326890
rect 676736 326826 676737 326890
rect 676671 326825 676737 326826
rect 676866 313719 676926 357609
rect 676863 313718 676929 313719
rect 676863 313654 676864 313718
rect 676928 313654 676929 313718
rect 676863 313653 676929 313654
rect 677058 312091 677118 357609
rect 677250 356673 677310 373929
rect 699639 369982 699959 370026
rect 699306 369981 700402 369982
rect 699306 368887 699307 369981
rect 700401 368887 700402 369981
rect 699306 368886 700402 368887
rect 699639 358922 699959 368886
rect 709903 367917 710223 367928
rect 709267 367916 710453 367917
rect 709267 366732 709268 367916
rect 710452 366732 710453 367916
rect 709267 366731 710453 366732
rect 700567 366062 701753 366063
rect 700567 364878 700568 366062
rect 701752 364878 701753 366062
rect 700567 364877 701753 364878
rect 700959 357368 701279 364877
rect 707887 364312 709073 364313
rect 707887 363128 707888 364312
rect 709072 363128 709073 364312
rect 707887 363127 709073 363128
rect 708583 358068 708903 363127
rect 709903 359208 710223 366731
rect 677250 356613 677502 356673
rect 677442 356491 677502 356613
rect 677439 356490 677505 356491
rect 677439 356426 677440 356490
rect 677504 356426 677505 356490
rect 677439 356425 677505 356426
rect 677247 312534 677313 312535
rect 677247 312470 677248 312534
rect 677312 312470 677313 312534
rect 677247 312469 677313 312470
rect 677055 312090 677121 312091
rect 677055 312026 677056 312090
rect 677120 312026 677121 312090
rect 677055 312025 677121 312026
rect 676863 311498 676929 311499
rect 676863 311434 676864 311498
rect 676928 311434 676929 311498
rect 676863 311433 676929 311434
rect 675903 299510 675969 299511
rect 675903 299446 675904 299510
rect 675968 299446 675969 299510
rect 675903 299445 675969 299446
rect 675519 289594 675585 289595
rect 675519 289530 675520 289594
rect 675584 289530 675585 289594
rect 675519 289529 675585 289530
rect 674559 285006 674625 285007
rect 674559 284942 674560 285006
rect 674624 284942 674625 285006
rect 674559 284941 674625 284942
rect 674367 284858 674433 284859
rect 674367 284794 674368 284858
rect 674432 284794 674433 284858
rect 674367 284793 674433 284794
rect 673983 283674 674049 283675
rect 673983 283610 673984 283674
rect 674048 283610 674049 283674
rect 673983 283609 674049 283610
rect 670882 279568 671708 280948
rect 670882 278476 671683 279568
rect 670882 275858 671708 278476
rect 673376 275858 673462 280948
rect 669304 270666 670416 270706
rect 669304 268850 669344 270666
rect 670376 268850 670416 270666
rect 669304 268810 670416 268850
rect 669318 268540 670414 268810
rect 665024 267072 665026 267722
rect 668262 267072 668306 267722
rect 661092 264274 664206 264314
rect 661092 261240 661132 264274
rect 664166 261240 664206 264274
rect 661092 261200 664206 261240
rect 656786 259369 660572 259624
rect 641148 252616 656268 252656
rect 641148 249422 641188 252616
rect 656228 252608 656268 252616
rect 656228 249422 656316 252608
rect 641148 249382 656316 249422
rect 641196 249286 656316 249382
rect 656786 248522 660558 259369
rect 656722 248516 660622 248522
rect 656700 248482 660622 248516
rect 656700 248476 656762 248482
rect 656700 244612 656740 248476
rect 656700 244572 656762 244612
rect 656722 242888 656762 244572
rect 660582 242888 660622 248482
rect 656722 242848 660622 242888
rect 656780 241434 660558 242848
rect 638822 234498 644382 234540
rect 638822 234446 652594 234498
rect 656780 234446 660552 241434
rect 638822 234294 660552 234446
rect 636927 233946 636993 233947
rect 636927 233882 636928 233946
rect 636992 233882 636993 233946
rect 636927 233881 636993 233882
rect 212418 100203 212670 100263
rect 212802 100203 213054 100263
rect 212418 99597 212478 100203
rect 211074 89547 211326 89607
rect 211458 99537 212478 99597
rect 211074 89351 211134 89547
rect 211071 89350 211137 89351
rect 211071 89286 211072 89350
rect 211136 89286 211137 89350
rect 211071 89285 211137 89286
rect 211071 87722 211137 87723
rect 211071 87658 211072 87722
rect 211136 87720 211137 87722
rect 211458 87720 211518 99537
rect 211136 87660 211518 87720
rect 211136 87658 211137 87660
rect 211071 87657 211137 87658
rect 212802 87609 212862 100203
rect 212802 87549 213054 87609
rect 211071 87278 211137 87279
rect 211071 87214 211072 87278
rect 211136 87214 211137 87278
rect 211071 87213 211137 87214
rect 211074 86943 211134 87213
rect 211074 86883 212478 86943
rect 210882 84885 211326 84945
rect 210879 82690 210945 82691
rect 210879 82626 210880 82690
rect 210944 82626 210945 82690
rect 210879 82625 210945 82626
rect 210882 71625 210942 82625
rect 211266 74955 211326 84885
rect 212418 76953 212478 86883
rect 212034 76893 212478 76953
rect 212034 74955 212094 76893
rect 212994 74955 213054 87549
rect 211266 74895 211902 74955
rect 212034 74895 212286 74955
rect 211842 72957 211902 74895
rect 211074 72923 211902 72957
rect 211071 72922 211902 72923
rect 211071 72858 211072 72922
rect 211136 72897 211902 72922
rect 211136 72858 211137 72897
rect 211071 72857 211137 72858
rect 210882 71565 211902 71625
rect 210498 70899 211710 70959
rect 210306 70233 211518 70293
rect 210114 69567 210750 69627
rect 209919 62858 209985 62859
rect 209919 62794 209920 62858
rect 209984 62794 209985 62858
rect 209919 62793 209985 62794
rect 209922 54127 209982 62793
rect 210303 62562 210369 62563
rect 210303 62498 210304 62562
rect 210368 62498 210369 62562
rect 210303 62497 210369 62498
rect 210306 54275 210366 62497
rect 210690 55063 210750 69567
rect 211071 58270 211137 58271
rect 211071 58206 211072 58270
rect 211136 58206 211137 58270
rect 211071 58205 211137 58206
rect 210303 54274 210369 54275
rect 210303 54210 210304 54274
rect 210368 54210 210369 54274
rect 210303 54209 210369 54210
rect 209919 54126 209985 54127
rect 209919 54062 209920 54126
rect 209984 54062 209985 54126
rect 209919 54061 209985 54062
rect 211074 53979 211134 58205
rect 211071 53978 211137 53979
rect 211071 53914 211072 53978
rect 211136 53914 211137 53978
rect 211071 53913 211137 53914
rect 209727 53830 209793 53831
rect 209727 53766 209728 53830
rect 209792 53766 209793 53830
rect 209727 53765 209793 53766
rect 211458 53239 211518 70233
rect 211650 54275 211710 70899
rect 211842 54975 211902 71565
rect 212226 64965 212286 74895
rect 212610 74895 213054 74955
rect 212610 74289 212670 74895
rect 212610 74229 212862 74289
rect 212226 64905 212478 64965
rect 211842 54915 212286 54975
rect 211647 54274 211713 54275
rect 211647 54210 211648 54274
rect 211712 54210 211713 54274
rect 211647 54209 211713 54210
rect 212226 53683 212286 54915
rect 212223 53682 212289 53683
rect 212223 53618 212224 53682
rect 212288 53618 212289 53682
rect 212223 53617 212289 53618
rect 212418 53387 212478 64905
rect 212802 54127 212862 74229
rect 212994 55581 213438 55641
rect 212799 54126 212865 54127
rect 212799 54062 212800 54126
rect 212864 54062 212865 54126
rect 212799 54061 212865 54062
rect 212994 53535 213054 55581
rect 213378 55063 213438 55581
rect 212991 53534 213057 53535
rect 212991 53470 212992 53534
rect 213056 53470 213057 53534
rect 212991 53469 213057 53470
rect 212415 53386 212481 53387
rect 212415 53322 212416 53386
rect 212480 53322 212481 53386
rect 212415 53321 212481 53322
rect 211455 53238 211521 53239
rect 211455 53174 211456 53238
rect 211520 53174 211521 53238
rect 211455 53173 211521 53174
rect 205416 46158 205456 46166
rect 143770 45200 143858 45310
rect 143770 43084 143852 45200
rect 181802 43114 181926 45584
rect 143770 43054 143858 43084
rect 214642 45548 214962 56300
rect 219642 49564 219962 56616
rect 218490 49524 220886 49564
rect 218490 46206 218530 49524
rect 220846 46206 220886 49524
rect 218490 46166 220886 46206
rect 213090 45508 216424 45548
rect 143770 43028 144386 43054
rect 213090 43030 213130 45508
rect 216384 43030 216424 45508
rect 224642 45112 224962 56118
rect 229642 49524 229962 56530
rect 229642 46174 229962 46228
rect 234642 45192 234962 56162
rect 239642 49544 239962 56616
rect 244642 45272 244962 56206
rect 249642 49544 249962 56186
rect 245726 46184 245756 47758
rect 251524 47018 251542 47758
rect 251524 46272 251570 47018
rect 251512 46184 251570 46272
rect 213090 42990 216424 43030
rect 214642 42850 214962 42990
rect 224642 42734 224962 43120
rect 234642 42876 234962 43120
rect 244642 42688 244962 43120
rect 143180 42494 143926 42520
rect 245726 42388 251570 46184
rect 254642 45352 254962 56050
rect 259642 49566 259962 56444
rect 264642 45336 264962 56206
rect 269642 49530 269962 56444
rect 274642 45464 274962 56118
rect 279642 49588 279962 56570
rect 254642 42828 254962 43120
rect 284642 45402 284962 56050
rect 289642 49552 289962 56096
rect 294642 45434 294962 56118
rect 299642 49544 299962 56484
rect 299642 46058 299962 46292
rect 264642 42822 264962 43024
rect 274642 42728 274962 43072
rect 284642 42446 284962 42930
rect 304642 45162 304962 56162
rect 309642 49524 309962 56096
rect 309642 46100 309962 46228
rect 314642 45338 314962 56050
rect 319642 49524 319962 56354
rect 319642 46100 319962 46228
rect 324642 45480 324962 56050
rect 329642 49566 329962 56312
rect 329642 46014 329962 46228
rect 294642 42822 294962 42882
rect 304642 42540 304962 43024
rect 314642 42540 314962 43120
rect 334642 45290 334962 56050
rect 339642 49524 339962 56054
rect 339642 46058 339962 46206
rect 344642 45386 344962 56162
rect 349642 49544 349962 56050
rect 349642 46058 349962 46248
rect 324642 42916 324962 42976
rect 354642 45320 354962 56162
rect 359642 49524 359962 56182
rect 364642 45258 364962 56294
rect 369642 49544 369962 56140
rect 369642 46058 369962 46248
rect 374642 45386 374962 56206
rect 379642 49588 379962 56096
rect 379642 46144 379962 46248
rect 384642 45290 384962 56206
rect 389642 49524 389962 56050
rect 389642 46014 389962 46248
rect 394642 45290 394962 56050
rect 399642 49588 399962 56182
rect 399642 46058 399962 46184
rect 404642 45290 404962 56050
rect 409642 49524 409962 56050
rect 409642 46014 409962 46270
rect 414642 45242 414962 56074
rect 419642 49544 419962 56140
rect 419642 45886 419962 46248
rect 424642 45226 424962 56050
rect 429642 49544 429962 56440
rect 429642 45972 429962 46228
rect 434642 45258 434962 56074
rect 439642 49566 439962 56096
rect 439642 46100 439962 46228
rect 444642 45338 444962 56118
rect 449642 49588 449962 56182
rect 449642 45886 449962 46248
rect 454642 45210 454962 56074
rect 459642 49544 459962 56268
rect 459642 45756 459962 46228
rect 464642 45314 464962 56118
rect 469642 49544 469962 56226
rect 471039 49094 471105 49095
rect 471039 49030 471040 49094
rect 471104 49030 471105 49094
rect 471039 49029 471105 49030
rect 469642 45972 469962 46270
rect 189951 41842 190017 41843
rect 189951 41778 189952 41842
rect 190016 41778 190017 41842
rect 189951 41777 190017 41778
rect 189954 40659 190014 41777
rect 245754 41678 251570 42388
rect 471042 42139 471102 49029
rect 474642 45242 474962 56294
rect 479642 49544 479962 56226
rect 479642 46100 479962 46248
rect 484642 45290 484962 56162
rect 489642 49524 489962 56140
rect 494642 45290 494962 56050
rect 499642 49566 499962 56140
rect 499642 45756 499962 46270
rect 504642 45332 504962 56250
rect 509642 49502 509962 56140
rect 509642 45370 509962 46248
rect 514642 45332 514962 56074
rect 519642 49676 519962 56312
rect 519642 45456 519962 46184
rect 474642 42540 474962 43104
rect 524642 45266 524962 56206
rect 529642 49480 529962 56312
rect 521343 45098 521409 45099
rect 521343 45034 521344 45098
rect 521408 45034 521409 45098
rect 521343 45033 521409 45034
rect 521346 43323 521406 45033
rect 521343 43322 521409 43323
rect 521343 43258 521344 43322
rect 521408 43258 521409 43322
rect 521343 43257 521409 43258
rect 529642 45240 529962 46184
rect 534642 45204 534962 56162
rect 539642 49544 539962 56096
rect 539642 45240 539962 46228
rect 544642 45332 544962 56050
rect 594642 45410 594962 56068
rect 599642 49634 599962 56068
rect 604642 45490 604962 56050
rect 609642 49500 609962 56122
rect 614642 45624 614962 56284
rect 619642 49420 619962 56050
rect 619642 45990 619962 46298
rect 527103 44950 527169 44951
rect 527103 44886 527104 44950
rect 527168 44886 527169 44950
rect 527103 44885 527169 44886
rect 527106 43323 527166 44885
rect 527103 43322 527169 43323
rect 527103 43258 527104 43322
rect 527168 43258 527169 43322
rect 527103 43257 527169 43258
rect 504642 42874 504962 42996
rect 514642 42494 514962 43090
rect 524642 42778 524962 43184
rect 624642 45596 624962 56050
rect 629642 49580 629962 56230
rect 629642 45882 629962 46244
rect 634642 45622 634962 56050
rect 636930 51611 636990 233881
rect 637695 233798 637761 233799
rect 637695 233734 637696 233798
rect 637760 233734 637761 233798
rect 637695 233733 637761 233734
rect 637119 233650 637185 233651
rect 637119 233586 637120 233650
rect 637184 233586 637185 233650
rect 637119 233585 637185 233586
rect 637503 233650 637569 233651
rect 637503 233586 637504 233650
rect 637568 233586 637569 233650
rect 637503 233585 637569 233586
rect 637122 51759 637182 233585
rect 637311 233502 637377 233503
rect 637311 233438 637312 233502
rect 637376 233438 637377 233502
rect 637311 233437 637377 233438
rect 637314 52351 637374 233437
rect 637311 52350 637377 52351
rect 637311 52286 637312 52350
rect 637376 52286 637377 52350
rect 637311 52285 637377 52286
rect 637506 52055 637566 233585
rect 637503 52054 637569 52055
rect 637503 51990 637504 52054
rect 637568 51990 637569 52054
rect 637503 51989 637569 51990
rect 637698 51907 637758 233733
rect 637887 233502 637953 233503
rect 637887 233438 637888 233502
rect 637952 233438 637953 233502
rect 637887 233437 637953 233438
rect 637890 52203 637950 233437
rect 644294 233636 660552 234294
rect 644294 228076 660654 233636
rect 661102 230916 664196 261200
rect 665024 256444 668306 267072
rect 670882 266716 673462 275858
rect 670882 262940 671666 266716
rect 673392 262940 673462 266716
rect 674175 264138 674241 264139
rect 674175 264074 674176 264138
rect 674240 264074 674241 264138
rect 674175 264073 674241 264074
rect 670882 259546 673462 262940
rect 673983 260882 674049 260883
rect 673983 260818 673984 260882
rect 674048 260818 674049 260882
rect 673983 260817 674049 260818
rect 670582 259506 673462 259546
rect 670582 256906 670622 259506
rect 673366 256906 673462 259506
rect 670582 256866 673462 256906
rect 664958 256404 668374 256444
rect 664958 253308 664998 256404
rect 668334 253308 668374 256404
rect 664958 253268 668374 253308
rect 661100 229652 664196 230916
rect 661084 229055 664196 229652
rect 644294 226138 644382 228076
rect 638822 225131 641093 226138
rect 643327 225131 644382 226138
rect 661084 227873 662179 229055
rect 663361 227873 664196 229055
rect 661084 225562 664196 227873
rect 638822 198466 644382 225131
rect 645382 219024 664196 225562
rect 645388 215738 664196 219024
rect 645392 215654 651070 215738
rect 660442 215696 664196 215738
rect 665024 231435 668306 253268
rect 670882 249204 673462 256866
rect 670882 249174 673414 249204
rect 665024 230253 666067 231435
rect 667249 230253 668306 231435
rect 644292 194640 644382 198466
rect 638822 183191 644382 194640
rect 645392 185881 651070 210840
rect 645392 184342 645421 185881
rect 647655 184342 651070 185881
rect 665024 187433 668306 230253
rect 670842 248872 673414 249174
rect 670842 233636 673412 248872
rect 673986 242087 674046 260817
rect 674178 243567 674238 264073
rect 674370 244751 674430 284793
rect 674562 276423 674622 284941
rect 675906 284859 675966 299445
rect 676671 299362 676737 299363
rect 676671 299298 676672 299362
rect 676736 299298 676737 299362
rect 676671 299297 676737 299298
rect 675903 284858 675969 284859
rect 675903 284794 675904 284858
rect 675968 284794 675969 284858
rect 675903 284793 675969 284794
rect 676674 281899 676734 299297
rect 676671 281898 676737 281899
rect 676671 281834 676672 281898
rect 676736 281834 676737 281898
rect 676671 281833 676737 281834
rect 674559 276422 674625 276423
rect 674559 276358 674560 276422
rect 674624 276358 674625 276422
rect 674559 276357 674625 276358
rect 674562 246823 674622 276357
rect 676866 267099 676926 311433
rect 677058 267099 677118 312025
rect 677250 268727 677310 312469
rect 677442 312091 677502 356425
rect 699639 324238 699959 324276
rect 699294 324237 700390 324238
rect 699294 323143 699295 324237
rect 700389 323143 700390 324237
rect 699294 323142 700390 323143
rect 699639 313680 699959 323142
rect 709501 322606 710687 322607
rect 709501 321422 709502 322606
rect 710686 321422 710687 322606
rect 709501 321421 710687 321422
rect 700627 320472 701813 320473
rect 700627 319288 700628 320472
rect 701812 319288 701813 320472
rect 700627 319287 701813 319288
rect 700959 312276 701279 319287
rect 708583 318187 708903 318258
rect 707919 318186 709105 318187
rect 707919 317002 707920 318186
rect 709104 317002 709105 318186
rect 707919 317001 709105 317002
rect 708583 312966 708903 317001
rect 709903 314394 710223 321421
rect 677439 312090 677505 312091
rect 677439 312026 677440 312090
rect 677504 312026 677505 312090
rect 677439 312025 677505 312026
rect 699639 279570 699959 279582
rect 699328 279569 700424 279570
rect 699328 278475 699329 279569
rect 700423 278475 700424 279569
rect 699328 278474 700424 278475
rect 699639 268802 699959 278474
rect 709903 278001 710223 278142
rect 709389 278000 710575 278001
rect 709389 276816 709390 278000
rect 710574 276816 710575 278000
rect 709389 276815 710575 276816
rect 700623 275228 701809 275229
rect 700623 274044 700624 275228
rect 701808 274044 701809 275228
rect 700623 274043 701809 274044
rect 677247 268726 677313 268727
rect 677247 268662 677248 268726
rect 677312 268662 677313 268726
rect 677247 268661 677313 268662
rect 677439 267690 677505 267691
rect 677439 267626 677440 267690
rect 677504 267626 677505 267690
rect 677439 267625 677505 267626
rect 676863 267098 676929 267099
rect 676863 267034 676864 267098
rect 676928 267034 676929 267098
rect 676863 267033 676929 267034
rect 677055 267098 677121 267099
rect 677055 267034 677056 267098
rect 677120 267034 677121 267098
rect 677055 267033 677121 267034
rect 676866 256773 676926 267033
rect 676482 256713 676926 256773
rect 675903 251706 675969 251707
rect 675903 251642 675904 251706
rect 675968 251642 675969 251706
rect 675903 251641 675969 251642
rect 675711 251558 675777 251559
rect 675711 251494 675712 251558
rect 675776 251494 675777 251558
rect 675711 251493 675777 251494
rect 674559 246822 674625 246823
rect 674559 246758 674560 246822
rect 674624 246758 674625 246822
rect 674559 246757 674625 246758
rect 674562 245935 674622 246757
rect 674559 245934 674625 245935
rect 674559 245870 674560 245934
rect 674624 245870 674625 245934
rect 674559 245869 674625 245870
rect 674367 244750 674433 244751
rect 674367 244686 674368 244750
rect 674432 244686 674433 244750
rect 674367 244685 674433 244686
rect 675327 244750 675393 244751
rect 675327 244686 675328 244750
rect 675392 244686 675393 244750
rect 675327 244685 675393 244686
rect 674370 243863 674430 244685
rect 674367 243862 674433 243863
rect 674367 243798 674368 243862
rect 674432 243798 674433 243862
rect 674367 243797 674433 243798
rect 674175 243566 674241 243567
rect 674175 243502 674176 243566
rect 674240 243502 674241 243566
rect 674175 243501 674241 243502
rect 673983 242086 674049 242087
rect 673983 242022 673984 242086
rect 674048 242022 674049 242086
rect 673983 242021 674049 242022
rect 670842 232544 671683 233636
rect 672775 232544 673412 233636
rect 670842 207568 673412 232544
rect 674175 220552 674241 220553
rect 674175 220488 674176 220552
rect 674240 220488 674241 220552
rect 674175 220487 674241 220488
rect 665024 186251 666067 187433
rect 667249 186251 668306 187433
rect 638822 180957 641093 183191
rect 643327 180957 644382 183191
rect 638822 168156 644382 180957
rect 644302 164250 644382 168156
rect 638822 137703 644382 164250
rect 645392 154070 651070 179608
rect 650942 149416 651070 154070
rect 638822 137000 641093 137703
rect 643327 137000 644382 137703
rect 638822 133408 638896 137000
rect 644302 133408 644382 137000
rect 638822 107164 644382 133408
rect 645392 139451 651070 149416
rect 645392 137217 645421 139451
rect 647655 137217 651070 139451
rect 665024 141405 668306 186251
rect 665024 140223 666067 141405
rect 667249 140223 668306 141405
rect 670784 189502 673412 207568
rect 674178 193543 674238 220487
rect 675330 200055 675390 244685
rect 675519 238978 675585 238979
rect 675519 238914 675520 238978
rect 675584 238914 675585 238978
rect 675519 238913 675585 238914
rect 675327 200054 675393 200055
rect 675327 199990 675328 200054
rect 675392 199990 675393 200054
rect 675327 199989 675393 199990
rect 675522 199611 675582 238913
rect 675714 238683 675774 251493
rect 675711 238682 675777 238683
rect 675711 238618 675712 238682
rect 675776 238618 675777 238682
rect 675711 238617 675777 238618
rect 675906 236907 675966 251641
rect 676482 237795 676542 256713
rect 676479 237794 676545 237795
rect 676479 237730 676480 237794
rect 676544 237730 676545 237794
rect 676479 237729 676545 237730
rect 675903 236906 675969 236907
rect 675903 236842 675904 236906
rect 675968 236842 675969 236906
rect 675903 236841 675969 236842
rect 676482 236315 676542 237729
rect 677058 237647 677118 267033
rect 677055 237646 677121 237647
rect 677055 237582 677056 237646
rect 677120 237582 677121 237646
rect 677055 237581 677121 237582
rect 676479 236314 676545 236315
rect 676479 236250 676480 236314
rect 676544 236250 676545 236314
rect 676479 236249 676545 236250
rect 676863 236314 676929 236315
rect 676863 236250 676864 236314
rect 676928 236250 676929 236314
rect 676863 236249 676929 236250
rect 676866 221367 676926 236249
rect 677058 222551 677118 237581
rect 677442 223587 677502 267625
rect 700959 267262 701279 274043
rect 707923 273110 709109 273111
rect 707923 271926 707924 273110
rect 709108 271926 709109 273110
rect 707923 271925 709109 271926
rect 708583 267968 708903 271925
rect 709903 269130 710223 276815
rect 684954 254778 685638 254934
rect 684954 251802 685012 254778
rect 685600 251802 685638 254778
rect 684954 251718 685638 251802
rect 709243 233638 709563 233760
rect 708936 233637 710032 233638
rect 708936 232543 708937 233637
rect 710031 232543 710032 233637
rect 708936 232542 710032 232543
rect 698979 231437 699299 231440
rect 698421 231436 699607 231437
rect 698421 230252 698422 231436
rect 699606 230252 699607 231436
rect 698421 230251 699607 230252
rect 698979 223860 699299 230251
rect 707213 229000 708399 229001
rect 707213 227816 707214 229000
rect 708398 227816 708399 229000
rect 707213 227815 708399 227816
rect 699853 227314 701039 227315
rect 699853 226130 699854 227314
rect 701038 226130 701039 227314
rect 699853 226129 701039 226130
rect 677439 223586 677505 223587
rect 677439 223522 677440 223586
rect 677504 223522 677505 223586
rect 677439 223521 677505 223522
rect 700299 222674 700619 226129
rect 677055 222550 677121 222551
rect 677055 222486 677056 222550
rect 677120 222486 677121 222550
rect 677055 222485 677121 222486
rect 676863 221366 676929 221367
rect 676863 221302 676864 221366
rect 676928 221302 676929 221366
rect 676863 221301 676929 221302
rect 675711 207750 675777 207751
rect 675711 207686 675712 207750
rect 675776 207686 675777 207750
rect 675711 207685 675777 207686
rect 675519 199610 675585 199611
rect 675519 199546 675520 199610
rect 675584 199546 675585 199610
rect 675519 199545 675585 199546
rect 674175 193542 674241 193543
rect 674175 193478 674176 193542
rect 674240 193478 674241 193542
rect 674175 193477 674241 193478
rect 675327 193098 675393 193099
rect 675327 193034 675328 193098
rect 675392 193034 675393 193098
rect 675327 193033 675393 193034
rect 670784 188410 671683 189502
rect 672775 188410 673412 189502
rect 670784 143722 673412 188410
rect 673983 171194 674049 171195
rect 673983 171130 673984 171194
rect 674048 171130 674049 171194
rect 673983 171129 674049 171130
rect 673986 150327 674046 171129
rect 675330 155211 675390 193033
rect 675327 155210 675393 155211
rect 675327 155146 675328 155210
rect 675392 155146 675393 155210
rect 675327 155145 675393 155146
rect 673983 150326 674049 150327
rect 673983 150262 673984 150326
rect 674048 150262 674049 150326
rect 673983 150261 674049 150262
rect 670784 142630 671683 143722
rect 672775 142630 673412 143722
rect 670784 140766 673412 142630
rect 665024 139140 668306 140223
rect 670720 139250 673424 140766
rect 645392 123540 651070 137217
rect 673983 128718 674049 128719
rect 673983 128654 673984 128718
rect 674048 128654 674049 128718
rect 673983 128653 674049 128654
rect 650914 118966 651070 123540
rect 644346 103406 644382 107164
rect 645392 105666 651070 118966
rect 673986 108147 674046 128653
rect 674175 126054 674241 126055
rect 674175 125990 674176 126054
rect 674240 125990 674241 126054
rect 674175 125989 674241 125990
rect 673983 108146 674049 108147
rect 673983 108082 673984 108146
rect 674048 108082 674049 108146
rect 673983 108081 674049 108082
rect 638822 85142 644382 103406
rect 650836 101988 651070 105666
rect 638822 81544 638908 85142
rect 644344 81544 644382 85142
rect 638822 76240 644382 81544
rect 644378 72698 644382 76240
rect 637887 52202 637953 52203
rect 637887 52138 637888 52202
rect 637952 52138 637953 52202
rect 637887 52137 637953 52138
rect 637695 51906 637761 51907
rect 637695 51842 637696 51906
rect 637760 51842 637761 51906
rect 637695 51841 637761 51842
rect 637119 51758 637185 51759
rect 637119 51694 637120 51758
rect 637184 51694 637185 51758
rect 637119 51693 637185 51694
rect 636927 51610 636993 51611
rect 636927 51546 636928 51610
rect 636992 51546 636993 51610
rect 636927 51545 636993 51546
rect 638822 49474 644382 72698
rect 645392 92904 651070 101988
rect 645392 88410 645508 92904
rect 651042 88410 651070 92904
rect 645392 83008 651070 88410
rect 645392 79336 645426 83008
rect 650912 79336 651070 83008
rect 645392 60958 651070 79336
rect 650986 57944 651070 60958
rect 638822 46262 639000 49474
rect 644086 46262 644382 49474
rect 645392 46688 651070 57944
rect 651746 105627 653180 105634
rect 651746 105227 654584 105627
rect 638822 46218 644382 46262
rect 640686 46198 644054 46218
rect 641092 46186 643328 46198
rect 534642 42968 534962 43042
rect 594642 42846 594962 43046
rect 604642 42630 604962 43046
rect 614642 42954 614962 43100
rect 624642 42792 624962 42992
rect 645256 43036 645270 45460
rect 645256 43026 645372 43036
rect 650996 43026 651104 43036
rect 645256 42962 651104 43026
rect 573608 42492 579178 42522
rect 573608 42478 573714 42492
rect 471039 42138 471105 42139
rect 471039 42074 471040 42138
rect 471104 42074 471105 42138
rect 471039 42073 471105 42074
rect 245694 41648 251570 41678
rect 189951 40658 190017 40659
rect 189951 40594 189952 40658
rect 190016 40594 190017 40658
rect 189951 40593 190017 40594
rect 245694 40136 245742 41648
rect 251484 40136 251570 41648
rect 469314 40929 469566 40989
rect 469314 40659 469374 40929
rect 469506 40807 469566 40929
rect 469503 40806 469569 40807
rect 469503 40742 469504 40806
rect 469568 40742 469569 40806
rect 469503 40741 469569 40742
rect 469311 40658 469377 40659
rect 469311 40594 469312 40658
rect 469376 40594 469377 40658
rect 469311 40593 469377 40594
rect 573608 40312 573642 42478
rect 579078 40344 579178 42492
rect 651746 42488 653188 105227
rect 674178 105187 674238 125989
rect 675330 110071 675390 155145
rect 675522 154471 675582 199545
rect 675714 198427 675774 207685
rect 676671 207602 676737 207603
rect 676671 207538 676672 207602
rect 676736 207538 676737 207602
rect 676671 207537 676737 207538
rect 676479 207454 676545 207455
rect 676479 207390 676480 207454
rect 676544 207390 676545 207454
rect 676479 207389 676545 207390
rect 675711 198426 675777 198427
rect 675711 198362 675712 198426
rect 675776 198362 675777 198426
rect 675711 198361 675777 198362
rect 676482 195319 676542 207389
rect 676479 195318 676545 195319
rect 676479 195254 676480 195318
rect 676544 195254 676545 195318
rect 676479 195253 676545 195254
rect 676674 191619 676734 207537
rect 676671 191618 676737 191619
rect 676671 191554 676672 191618
rect 676736 191554 676737 191618
rect 676671 191553 676737 191554
rect 677058 177411 677118 222485
rect 677439 222402 677505 222403
rect 677439 222338 677440 222402
rect 677504 222338 677505 222402
rect 677439 222337 677505 222338
rect 677247 221366 677313 221367
rect 677247 221302 677248 221366
rect 677312 221302 677313 221366
rect 677247 221301 677313 221302
rect 677055 177410 677121 177411
rect 677055 177346 677056 177410
rect 677120 177346 677121 177410
rect 677055 177345 677121 177346
rect 675711 161574 675777 161575
rect 675711 161510 675712 161574
rect 675776 161510 675777 161574
rect 675711 161509 675777 161510
rect 675519 154470 675585 154471
rect 675519 154406 675520 154470
rect 675584 154406 675585 154470
rect 675519 154405 675585 154406
rect 675327 110070 675393 110071
rect 675327 110006 675328 110070
rect 675392 110006 675393 110070
rect 675327 110005 675393 110006
rect 675522 109331 675582 154405
rect 675714 148551 675774 161509
rect 676671 161426 676737 161427
rect 676671 161362 676672 161426
rect 676736 161362 676737 161426
rect 676671 161361 676737 161362
rect 675711 148550 675777 148551
rect 675711 148486 675712 148550
rect 675776 148486 675777 148550
rect 675711 148485 675777 148486
rect 676674 146627 676734 161361
rect 676671 146626 676737 146627
rect 676671 146562 676672 146626
rect 676736 146562 676737 146626
rect 676671 146561 676737 146562
rect 677058 132271 677118 177345
rect 677250 176375 677310 221301
rect 677442 178447 677502 222337
rect 707923 222180 708243 227815
rect 709243 223316 709563 232542
rect 709243 189504 709563 189652
rect 708776 189503 709872 189504
rect 708776 188409 708777 189503
rect 709871 188409 709872 189503
rect 708776 188408 709872 188409
rect 698979 187435 699299 187462
rect 698513 187434 699699 187435
rect 698513 186250 698514 187434
rect 699698 186250 699699 187434
rect 698513 186249 699699 186250
rect 698979 179066 699299 186249
rect 700959 185085 701279 185128
rect 700655 185084 701841 185085
rect 700655 183900 700656 185084
rect 701840 183900 701841 185084
rect 700655 183899 701841 183900
rect 677439 178446 677505 178447
rect 677439 178382 677440 178446
rect 677504 178382 677505 178446
rect 677439 178381 677505 178382
rect 677439 177410 677505 177411
rect 677439 177346 677440 177410
rect 677504 177346 677505 177410
rect 677439 177345 677505 177346
rect 677247 176374 677313 176375
rect 677247 176310 677248 176374
rect 677312 176310 677313 176374
rect 677247 176309 677313 176310
rect 677055 132270 677121 132271
rect 677055 132206 677056 132270
rect 677120 132206 677121 132270
rect 677055 132205 677121 132206
rect 677250 131827 677310 176309
rect 677442 133455 677502 177345
rect 700959 177072 701279 183899
rect 706103 182394 707289 182395
rect 706103 181210 706104 182394
rect 707288 181868 707289 182394
rect 707288 181548 708903 181868
rect 707288 181210 707289 181548
rect 706103 181209 707289 181210
rect 708583 177168 708903 181548
rect 709243 178142 709563 188408
rect 709243 143724 709563 143788
rect 708742 143723 709838 143724
rect 708742 142629 708743 143723
rect 709837 142629 709838 143723
rect 708742 142628 709838 142629
rect 698401 141406 699587 141407
rect 698401 140222 698402 141406
rect 699586 140222 699587 141406
rect 698401 140221 699587 140222
rect 698979 134034 699299 140221
rect 700959 138677 701279 138732
rect 700549 138676 701735 138677
rect 700549 137492 700550 138676
rect 701734 137492 701735 138676
rect 700549 137491 701735 137492
rect 677439 133454 677505 133455
rect 677439 133390 677440 133454
rect 677504 133390 677505 133454
rect 677439 133389 677505 133390
rect 700959 131956 701279 137491
rect 706921 136690 708107 136691
rect 706921 135506 706922 136690
rect 708106 136342 708107 136690
rect 708106 136022 708903 136342
rect 708106 135506 708107 136022
rect 706921 135505 708107 135506
rect 708583 132618 708903 136022
rect 709243 133476 709563 142628
rect 677247 131826 677313 131827
rect 677247 131762 677248 131826
rect 677312 131762 677313 131826
rect 677247 131761 677313 131762
rect 676479 118062 676545 118063
rect 676479 117998 676480 118062
rect 676544 117998 676545 118062
rect 676479 117997 676545 117998
rect 675903 117914 675969 117915
rect 675903 117850 675904 117914
rect 675968 117850 675969 117914
rect 675903 117849 675969 117850
rect 675519 109330 675585 109331
rect 675519 109266 675520 109330
rect 675584 109266 675585 109330
rect 675519 109265 675585 109266
rect 674175 105186 674241 105187
rect 674175 105122 674176 105186
rect 674240 105122 674241 105186
rect 674175 105121 674241 105122
rect 653454 104900 653914 104906
rect 653454 104596 654236 104900
rect 653454 103828 654118 104596
rect 653454 103724 655012 103828
rect 653458 53866 655012 103724
rect 664997 103712 665326 104920
rect 675906 103263 675966 117849
rect 675903 103262 675969 103263
rect 675903 103198 675904 103262
rect 675968 103198 675969 103262
rect 675903 103197 675969 103198
rect 676482 101487 676542 117997
rect 676479 101486 676545 101487
rect 676479 101422 676480 101486
rect 676544 101422 676545 101486
rect 676479 101421 676545 101422
rect 654866 50706 655012 53866
rect 653550 50680 654476 50706
rect 653814 50610 654118 50680
rect 651746 42484 653462 42488
rect 579070 40312 579178 40344
rect 573608 40270 579178 40312
rect 245694 40088 251570 40136
rect 245754 40046 251570 40088
<< via4 >>
rect 54718 996198 56068 997038
rect 53140 994938 54504 995752
rect 51620 993544 52878 994554
rect 49664 992148 51396 993104
rect 44866 989600 45466 990200
rect 41134 988042 42390 988148
rect 41134 984584 41196 988042
rect 41196 984584 42102 988042
rect 42102 984584 42390 988042
rect 41134 984514 42390 984584
rect 43290 983126 44470 985550
rect 46142 988556 46742 989156
rect 43906 275482 44432 277114
rect 47268 985814 49228 986974
rect 47242 269828 49208 275552
rect 46142 267794 46742 268394
rect 44912 266996 45430 267378
rect 43870 266248 44470 266848
rect 49020 262254 51400 265720
rect 48262 256860 54378 259448
rect 125358 996172 125910 996724
rect 124030 994918 124582 995470
rect 122840 993746 123392 994298
rect 121382 992366 121934 992918
rect 177484 996172 178036 996724
rect 176228 994918 176780 995470
rect 174544 993746 175096 994298
rect 173292 992366 173844 992918
rect 228798 996172 229350 996724
rect 227348 994918 227900 995470
rect 225508 993746 226060 994298
rect 223930 992366 224482 992918
rect 278946 996172 279498 996724
rect 277804 994918 278356 995470
rect 276398 993746 276950 994298
rect 274904 992366 275456 992918
rect 332460 996172 333012 996724
rect 330912 994918 331464 995470
rect 329356 993746 329908 994298
rect 327798 992366 328350 992918
rect 381572 996172 382124 996724
rect 380104 994918 380656 995470
rect 378554 993746 379106 994298
rect 377220 992366 377772 992918
rect 415946 996172 416498 996724
rect 414382 994918 414934 995470
rect 412172 993746 412724 994298
rect 410170 992366 410722 992918
rect 496120 996172 496672 996724
rect 494606 994918 495158 995470
rect 493094 993746 493646 994298
rect 491674 992366 492226 992918
rect 573470 996172 574022 996724
rect 580186 997072 585676 997096
rect 580186 996004 580256 997072
rect 580256 996004 585666 997072
rect 585666 996004 585676 997072
rect 580186 995988 585676 996004
rect 651576 996024 656490 996686
rect 655360 996022 655902 996024
rect 571858 994918 572410 995470
rect 650578 994470 653584 995000
rect 570352 993746 570904 994298
rect 648716 993536 651292 994070
rect 568202 992366 568754 992918
rect 665102 994456 668240 996748
rect 659386 992298 660564 993070
rect 59102 270210 61054 270606
rect 57688 267890 59474 268836
rect 56474 267052 58874 267312
rect 208550 270178 208870 270498
rect 60476 266096 62762 266660
rect 181826 261204 193584 265614
rect 45536 247120 47756 248490
rect 45520 244696 47756 247120
rect 45536 244520 47756 244696
rect 43732 239408 44458 239410
rect 43722 239398 44458 239408
rect 43714 239366 44458 239398
rect 42530 237972 45096 239366
rect 45600 232804 47800 233890
rect 43698 229082 44424 229084
rect 43688 229072 44424 229082
rect 43680 229040 44424 229072
rect 42496 227646 45062 229040
rect 45588 222882 47788 223968
rect 43720 218756 44446 218758
rect 43710 218746 44446 218756
rect 43702 218714 44446 218746
rect 42518 217320 45084 218714
rect 50568 253286 56050 256282
rect 45614 212904 47814 213990
rect 43744 209076 44470 209078
rect 43734 209066 44470 209076
rect 43726 209034 44470 209066
rect 42542 207640 45108 209034
rect 43722 199136 44448 199138
rect 43712 199126 44448 199136
rect 43704 199094 44448 199126
rect 42520 197700 45086 199094
rect 43726 189048 44452 189050
rect 43716 189038 44452 189048
rect 43708 189006 44452 189038
rect 42524 187612 45090 189006
rect 45614 202576 47814 203662
rect 45614 192792 47814 193878
rect 45614 183006 47814 184092
rect 43738 179100 44464 179102
rect 43728 179090 44464 179100
rect 43720 179058 44464 179090
rect 42536 177664 45102 179058
rect 43726 169174 44452 169176
rect 43716 169132 44452 169174
rect 42524 167738 45090 169132
rect 43714 159044 44440 159088
rect 42512 157650 45078 159044
rect 42502 147666 45068 149060
rect 42512 137844 45078 139238
rect 42502 127976 45068 129370
rect 42528 117936 45094 119330
rect 45614 172678 47814 173764
rect 45614 162894 47814 163980
rect 45614 153110 47814 154196
rect 45614 142782 47814 143868
rect 45614 132996 47814 134082
rect 45614 122668 47814 123754
rect 45682 113088 47882 114174
rect 43666 109050 44392 109052
rect 43656 109040 44392 109050
rect 43648 109008 44392 109040
rect 42464 107614 45030 109008
rect 45682 102760 47882 103846
rect 43690 98964 44416 98966
rect 43680 98954 44416 98964
rect 43672 98922 44416 98954
rect 42488 97528 45054 98922
rect 45670 92782 47870 93868
rect 43720 89140 44446 89142
rect 43714 89138 44446 89140
rect 43704 89128 44446 89138
rect 43696 89096 44446 89128
rect 42512 87702 45078 89096
rect 40888 77556 40974 79288
rect 40974 77556 45006 79288
rect 45006 77556 45134 79288
rect 45698 82830 47898 83916
rect 45668 72892 47790 73834
rect 40900 69066 40974 69384
rect 40974 69066 45006 69384
rect 45006 69066 45180 69384
rect 40900 67906 45180 69066
rect 40844 57596 45106 59078
rect 45694 63064 47816 64006
rect 48426 52944 50830 55910
rect 48426 50656 50852 52944
rect 144490 50716 144898 51598
rect 208678 267852 208998 268172
rect 208696 267026 209016 267346
rect 369770 270650 370006 270847
rect 369770 270611 369856 270650
rect 369856 270611 369920 270650
rect 369920 270611 370006 270650
rect 391274 270611 391510 270847
rect 369386 269945 369622 270181
rect 383978 269945 384214 270181
rect 267818 267281 268054 267517
rect 292202 267281 292438 267517
rect 377450 267281 377686 267517
rect 383594 267281 383830 267517
rect 211376 266302 211696 266622
rect 211832 261176 212882 265166
rect 206990 259496 209024 259514
rect 206990 256926 206998 259496
rect 206998 256926 209004 259496
rect 209004 256926 209024 259496
rect 206990 256918 209024 256926
rect 206480 256326 209016 256334
rect 206480 253280 208996 256326
rect 208996 253280 209016 256326
rect 194614 240282 206854 248416
rect 211886 244036 215748 245954
rect 411678 265796 412528 267970
rect 413024 267242 413344 267562
rect 415028 268996 415348 269316
rect 415068 268020 415388 268340
rect 653170 269026 654946 269578
rect 654916 267934 656440 268526
rect 647144 265124 654338 266582
rect 411872 261174 412420 264272
rect 422520 261214 426748 264292
rect 416354 259382 424206 259552
rect 416354 256980 416548 259382
rect 416548 256980 423896 259382
rect 423896 256980 424206 259382
rect 416354 256926 424206 256980
rect 416330 256270 424274 256398
rect 416330 253412 416506 256270
rect 416506 253412 424074 256270
rect 424074 253412 424274 256270
rect 416330 253332 424274 253412
rect 409646 242868 412718 244938
rect 194542 224480 206846 230162
rect 181728 206248 193602 216660
rect 194542 192744 206932 202814
rect 181814 174942 193522 185790
rect 181728 144926 193516 155854
rect 194714 163330 207024 173320
rect 194628 131594 206858 141504
rect 181900 115426 193528 127140
rect 194456 100374 206932 112852
rect 181900 86356 193608 98150
rect 194456 83060 206852 83100
rect 194456 70702 207022 83060
rect 181674 54130 193566 60778
rect 194520 60770 207022 70702
rect 48426 50098 50830 50656
rect 45634 46014 48118 49544
rect 40802 40944 45186 45628
rect 432428 261166 436466 264388
rect 428164 242898 430986 248482
rect 442192 261084 446416 264314
rect 452908 261168 457052 264318
rect 463542 261250 467186 264314
rect 437744 242806 440486 248310
rect 448198 242806 451434 248574
rect 458330 242898 461486 248586
rect 472686 261168 477156 264314
rect 482780 261208 487996 264232
rect 492544 261168 497098 264356
rect 468370 242944 471446 248552
rect 478318 242898 481232 248528
rect 488312 242852 491086 248666
rect 502558 261126 507690 264274
rect 511908 261126 517454 264232
rect 522788 261168 527342 264314
rect 498812 242852 501506 248586
rect 508162 242898 510776 248552
rect 517924 242852 521714 248528
rect 532678 261084 537396 264274
rect 542814 261208 547452 264318
rect 552536 261208 557836 264274
rect 527918 242806 531628 248402
rect 538142 242806 541470 248574
rect 547814 242852 551062 248540
rect 562962 261126 567434 264150
rect 573224 261126 577654 264438
rect 557210 242898 561228 248528
rect 567618 242806 571822 248574
rect 582822 261084 587708 264398
rect 592338 261168 596850 264398
rect 577106 242898 581078 248436
rect 588250 242898 591716 248574
rect 602640 261044 606780 264314
rect 613232 261250 617372 264232
rect 597646 242898 601434 248528
rect 607364 242898 611072 248448
rect 622748 261168 626930 264274
rect 632470 261168 637522 264274
rect 618232 242898 621284 248666
rect 627904 242852 631554 248528
rect 661196 990384 664096 992954
rect 671690 991374 673416 994178
rect 665082 983950 668280 985912
rect 669334 986772 670384 987294
rect 671718 985058 672730 985060
rect 671718 981854 673374 985058
rect 666084 276817 667226 277424
rect 666084 275208 667226 276817
rect 671708 279568 673376 280948
rect 671708 278476 672775 279568
rect 672775 278476 673376 279568
rect 671708 275858 673376 278476
rect 669344 268850 670376 270666
rect 665026 267072 668262 267722
rect 661132 261240 664166 264274
rect 641188 252222 656228 252616
rect 641188 249864 641918 252222
rect 641918 249864 655400 252222
rect 655400 249864 656228 252222
rect 641188 249422 656228 249864
rect 656762 248476 660582 248482
rect 656740 244612 660582 248476
rect 656762 242888 660582 244612
rect 210602 54827 210838 55063
rect 213290 54827 213526 55063
rect 194648 46166 207040 49686
rect 198642 46158 205416 46166
rect 143858 45200 145810 45500
rect 143852 43084 145810 45200
rect 143858 43054 145810 43084
rect 181926 43070 195992 45584
rect 218530 46206 220846 49524
rect 213130 43030 216384 45508
rect 228244 46228 231018 49524
rect 238350 46228 240972 49544
rect 245756 48302 251512 49544
rect 245756 46272 251524 48302
rect 245756 46184 251512 46272
rect 223370 43120 226464 45112
rect 232944 43120 236118 45192
rect 241992 43120 245246 45272
rect 142006 40624 143984 42494
rect 258084 46184 260922 49566
rect 253530 43120 256864 45352
rect 268168 46228 270926 49530
rect 278448 46184 280676 49588
rect 262720 43024 266134 45336
rect 273300 43072 276794 45464
rect 288444 46228 290592 49552
rect 298376 46292 300998 49544
rect 282922 42930 286496 45402
rect 293024 42882 296678 45434
rect 308178 46228 311320 49524
rect 317934 46228 321622 49524
rect 327976 46228 331228 49566
rect 303508 43024 306174 45162
rect 313416 43120 316162 45338
rect 323470 42976 326550 45480
rect 337972 46206 341202 49524
rect 348100 46248 351788 49544
rect 332518 43072 335980 45290
rect 343002 42930 346272 45386
rect 357988 46228 361524 49524
rect 353150 43024 355926 45320
rect 368138 46248 371608 49544
rect 378112 46248 381518 49588
rect 363012 42882 365868 45258
rect 373208 42930 376144 45386
rect 388110 46248 391296 49524
rect 397954 46184 401250 49588
rect 407602 46270 411270 49524
rect 382878 43072 386244 45290
rect 393218 42976 396250 45290
rect 402410 42976 405824 45290
rect 417382 46248 421222 49544
rect 413372 42930 416212 45242
rect 427924 46228 431634 49544
rect 437420 46228 441260 49566
rect 447896 46248 451540 49588
rect 423090 43072 425914 45226
rect 433192 43024 436096 45258
rect 443100 43024 446084 45338
rect 458372 46228 461516 49544
rect 468020 46270 470336 49544
rect 453344 43120 456344 45210
rect 463500 43010 465734 45314
rect 478650 46248 481074 49544
rect 488580 46184 490810 49524
rect 498360 46270 501308 49566
rect 508314 46248 511566 49502
rect 517832 46184 521324 49676
rect 473898 43104 475988 45242
rect 483074 43120 486056 45290
rect 492934 43120 496014 45290
rect 503498 42996 506214 45332
rect 513212 43138 516308 45332
rect 527784 46184 531408 49480
rect 523684 43184 525578 45266
rect 537586 46228 541362 49544
rect 598014 46352 601404 49634
rect 607988 46298 611298 49500
rect 618342 46298 621572 49420
rect 513734 43090 515548 43138
rect 533968 43042 535942 45204
rect 543776 43090 545830 45332
rect 592974 43046 596096 45410
rect 603056 43046 606258 45490
rect 613356 43100 616638 45624
rect 628262 46244 631652 49580
rect 638808 227365 644294 234294
rect 671666 262940 673392 266716
rect 670622 256906 673366 259506
rect 664998 253308 668334 256404
rect 638808 226138 641093 227365
rect 641093 226138 643327 227365
rect 643327 226138 644294 227365
rect 645352 210840 651206 215654
rect 638712 194640 644292 198466
rect 645352 183647 645421 184342
rect 645421 183647 647655 184342
rect 647655 183647 651126 184342
rect 645352 179608 651126 183647
rect 638642 164250 644302 168156
rect 645248 149416 650942 154070
rect 638896 135469 641093 137000
rect 641093 135469 643327 137000
rect 643327 135469 644302 137000
rect 638896 133408 644302 135469
rect 645300 118966 650914 123540
rect 638750 103406 644346 107164
rect 645320 101988 650836 105666
rect 638908 81544 644344 85142
rect 638806 72698 644378 76240
rect 645508 88410 651042 92904
rect 645426 79336 650912 83008
rect 645390 57944 650986 60958
rect 639000 46262 644086 49474
rect 623220 42992 626582 45596
rect 633196 42938 636638 45622
rect 645270 43036 651352 46688
rect 645372 43026 650996 43036
rect 573714 42478 579078 42492
rect 573714 40344 579070 42478
rect 579070 40344 579078 42478
rect 663816 101994 665508 103712
rect 653458 50706 654866 53866
rect 651706 39978 653730 42484
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 54684 997038 56092 997236
rect 54684 996198 54718 997038
rect 56068 996748 56092 997038
rect 580160 997096 585714 997134
rect 56068 996724 578714 996748
rect 56068 996198 125358 996724
rect 54684 996172 125358 996198
rect 125910 996172 177484 996724
rect 178036 996172 228798 996724
rect 229350 996172 278946 996724
rect 279498 996172 332460 996724
rect 333012 996172 381572 996724
rect 382124 996172 415946 996724
rect 416498 996172 496120 996724
rect 496672 996172 573470 996724
rect 574022 996172 578714 996724
rect 54684 996148 578714 996172
rect 54684 996138 56092 996148
rect 53092 995752 54538 995806
rect 53092 994938 53140 995752
rect 54504 995494 54538 995752
rect 54504 995488 576298 995494
rect 54504 995470 576456 995488
rect 54504 994938 124030 995470
rect 53092 994918 124030 994938
rect 124582 994918 176228 995470
rect 176780 994918 227348 995470
rect 227900 994918 277804 995470
rect 278356 994918 330912 995470
rect 331464 994918 380104 995470
rect 380656 994918 414382 995470
rect 414934 994918 494606 995470
rect 495158 994918 571858 995470
rect 572410 994918 576456 995470
rect 53092 994894 576456 994918
rect 53092 994884 54538 994894
rect 51584 994554 52910 994596
rect 51584 994542 51620 994554
rect 51558 993544 51620 994542
rect 52878 994542 52910 994554
rect 52878 994298 575178 994542
rect 52878 993746 122840 994298
rect 123392 993746 174544 994298
rect 175096 993746 225508 994298
rect 226060 993746 276398 994298
rect 276950 993746 329356 994298
rect 329908 993746 378554 994298
rect 379106 993746 412172 994298
rect 412724 993746 493094 994298
rect 493646 993746 570352 994298
rect 570904 993746 575178 994298
rect 52878 993544 575178 993746
rect 51558 993506 575178 993544
rect 49570 993104 51456 993180
rect 574142 993134 575178 993506
rect 575856 994094 576456 994894
rect 578114 995034 578714 996148
rect 580160 995988 580186 997096
rect 585676 996588 585714 997096
rect 665028 996748 668306 996830
rect 651552 996686 656548 996746
rect 651552 996588 651576 996686
rect 585676 996024 651576 996588
rect 656490 996024 656548 996686
rect 585676 996022 655360 996024
rect 655902 996022 656548 996024
rect 585676 995988 656548 996022
rect 580160 995962 585714 995988
rect 651552 995984 656548 995988
rect 665028 995034 665102 996748
rect 578114 995000 665102 995034
rect 578114 994470 650578 995000
rect 653584 994470 665102 995000
rect 578114 994456 665102 994470
rect 668240 994456 668306 996748
rect 578114 994434 668306 994456
rect 665028 994430 668306 994434
rect 671652 994178 673472 994302
rect 671652 994094 671690 994178
rect 575856 994070 671690 994094
rect 575856 993536 648716 994070
rect 651292 993536 671690 994070
rect 575856 993494 671690 993536
rect 49570 992148 49664 993104
rect 51396 992942 51456 993104
rect 574120 993070 660601 993134
rect 51396 992918 573712 992942
rect 51396 992366 121382 992918
rect 121934 992366 173292 992918
rect 173844 992366 223930 992918
rect 224482 992366 274904 992918
rect 275456 992366 327798 992918
rect 328350 992366 377220 992918
rect 377772 992366 410170 992918
rect 410722 992366 491674 992918
rect 492226 992366 568202 992918
rect 568754 992366 573712 992918
rect 51396 992342 573712 992366
rect 51396 992148 51456 992342
rect 49570 992096 51456 992148
rect 573112 991882 573712 992342
rect 574120 992298 659386 993070
rect 660564 992298 660601 993070
rect 574120 992272 660601 992298
rect 661102 992954 664178 993016
rect 661102 991882 661196 992954
rect 573112 991282 661196 991882
rect 661102 990384 661196 991282
rect 664096 990384 664178 992954
rect 671652 991374 671690 993494
rect 673416 991374 673472 994178
rect 671652 991298 673472 991374
rect 661102 990303 664178 990384
rect 44842 990200 45490 990224
rect 44842 990158 44866 990200
rect 44612 989600 44866 990158
rect 45466 990158 45490 990200
rect 45466 989600 58892 990158
rect 44612 989558 58892 989600
rect 45956 989156 59494 989218
rect 45956 988618 46142 989156
rect 46118 988556 46142 988618
rect 46742 988618 59494 989156
rect 46742 988556 46766 988618
rect 46118 988532 46766 988556
rect 41094 988148 42430 988188
rect 41094 984514 41134 988148
rect 42390 986667 42430 988148
rect 651596 987294 670986 987338
rect 47232 986974 49272 987022
rect 47232 986667 47268 986974
rect 42390 986137 47268 986667
rect 42390 984514 42430 986137
rect 46936 985814 47268 986137
rect 49228 986398 49272 986974
rect 651596 986772 669334 987294
rect 670384 986772 670986 987294
rect 651596 986738 670986 986772
rect 49228 985814 61862 986398
rect 46936 985798 61862 985814
rect 665026 985912 668316 985948
rect 47232 985786 49272 985798
rect 41094 984474 42430 984514
rect 43264 985550 44498 985646
rect 43264 983126 43290 985550
rect 44470 985458 44498 985550
rect 44470 984858 63004 985458
rect 44470 983126 44498 984858
rect 665026 984518 665082 985912
rect 650488 983950 665082 984518
rect 668280 983950 668316 985912
rect 671666 985106 673444 985126
rect 650488 983922 668316 983950
rect 671662 985060 673444 985106
rect 650488 983918 667846 983922
rect 671662 983578 671718 985060
rect 672730 985058 673444 985060
rect 43264 983082 44498 983126
rect 648614 982978 671718 983578
rect 671662 981854 671718 982978
rect 673374 981854 673444 985058
rect 671662 981798 673444 981854
rect 671666 981766 673444 981798
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 671642 280948 673476 281048
rect 671642 278394 671708 280948
rect 649042 277794 671708 278394
rect 666044 277454 667266 277464
rect 649560 277424 667370 277454
rect 43866 277114 44472 277154
rect 43866 276514 43906 277114
rect 43852 275914 43906 276514
rect 43866 275482 43906 275914
rect 44432 276514 44472 277114
rect 649560 276854 666084 277424
rect 44432 275914 62828 276514
rect 44432 275482 44472 275914
rect 43866 275442 44472 275482
rect 47196 275584 48322 275590
rect 47196 275574 49260 275584
rect 47196 275552 63184 275574
rect 47196 269828 47242 275552
rect 49208 274974 63184 275552
rect 666044 275208 666084 276854
rect 667226 276854 667370 277424
rect 667226 275208 667266 276854
rect 671642 275858 671708 277794
rect 673376 275858 673476 280948
rect 671642 275776 673476 275858
rect 666044 275168 667266 275208
rect 49208 270498 49260 274974
rect 369728 270847 391552 270889
rect 59062 270606 61094 270646
rect 59062 270498 59102 270606
rect 49208 270210 59102 270498
rect 61054 270498 61094 270606
rect 369728 270611 369770 270847
rect 370006 270611 391274 270847
rect 391510 270611 391552 270847
rect 369728 270569 391552 270611
rect 669304 270666 670416 270706
rect 208526 270498 208894 270522
rect 61054 270210 208550 270498
rect 49208 270178 208550 270210
rect 208870 270178 208894 270498
rect 49208 269828 49260 270178
rect 59062 270170 61094 270178
rect 208526 270154 208894 270178
rect 369344 270181 384256 270223
rect 369344 269945 369386 270181
rect 369622 269945 383978 270181
rect 384214 269945 384256 270181
rect 369344 269903 384256 269945
rect 47196 269792 49260 269828
rect 47222 269752 49260 269792
rect 653130 269578 654986 269618
rect 415004 269316 415372 269340
rect 653130 269316 653170 269578
rect 415004 268996 415028 269316
rect 415348 269026 653170 269316
rect 654946 269316 654986 269578
rect 669304 269316 669344 270666
rect 654946 269026 669344 269316
rect 415348 268996 669344 269026
rect 415004 268972 415372 268996
rect 653130 268986 654986 268996
rect 57648 268836 59514 268876
rect 46118 268394 46766 268418
rect 46118 268172 46142 268394
rect 46050 267852 46142 268172
rect 46118 267794 46142 267852
rect 46742 268172 46766 268394
rect 57648 268172 57688 268836
rect 46742 267890 57688 268172
rect 59474 268172 59514 268836
rect 669304 268850 669344 268996
rect 670376 268850 670416 270666
rect 669304 268810 670416 268850
rect 654876 268526 656474 268554
rect 415044 268340 415412 268364
rect 654876 268340 654916 268526
rect 208654 268172 209022 268196
rect 59474 267890 208678 268172
rect 46742 267852 208678 267890
rect 208998 267852 209022 268172
rect 415044 268020 415068 268340
rect 415388 268020 654916 268340
rect 46742 267794 46766 267852
rect 57648 267850 59514 267852
rect 208654 267828 209022 267852
rect 411638 267970 412568 268010
rect 415044 267996 415412 268020
rect 46118 267770 46766 267794
rect 267776 267517 292480 267559
rect 44864 267378 45462 267410
rect 44864 267346 44912 267378
rect 44838 267026 44912 267346
rect 44864 266996 44912 267026
rect 45430 267346 45462 267378
rect 208672 267346 209040 267370
rect 45430 267312 208696 267346
rect 45430 267052 56474 267312
rect 58874 267052 208696 267312
rect 45430 267026 208696 267052
rect 209016 267026 209040 267346
rect 267776 267281 267818 267517
rect 268054 267281 292202 267517
rect 292438 267281 292480 267517
rect 267776 267239 292480 267281
rect 377408 267517 383872 267559
rect 377408 267281 377450 267517
rect 377686 267281 383594 267517
rect 383830 267281 383872 267517
rect 377408 267239 383872 267281
rect 45430 266996 45462 267026
rect 208672 267002 209040 267026
rect 44864 266966 45462 266996
rect 43846 266848 44494 266872
rect 43846 266622 43870 266848
rect 43842 266302 43870 266622
rect 43846 266248 43870 266302
rect 44470 266622 44494 266848
rect 60436 266660 62802 266700
rect 60436 266622 60476 266660
rect 44470 266302 60476 266622
rect 44470 266248 44494 266302
rect 43846 266224 44494 266248
rect 60436 266096 60476 266302
rect 62762 266622 62802 266660
rect 211352 266622 211720 266646
rect 62762 266302 211376 266622
rect 211696 266302 211720 266622
rect 62762 266096 62802 266302
rect 211352 266278 211720 266302
rect 60436 266056 62802 266096
rect 411638 265796 411678 267970
rect 412528 266634 412568 267970
rect 654876 267934 654916 268020
rect 656440 268340 656474 268526
rect 656440 268020 656688 268340
rect 656440 267934 656474 268020
rect 654876 267890 656474 267934
rect 664994 267722 668300 267752
rect 413000 267562 413368 267586
rect 664994 267562 665026 267722
rect 413000 267242 413024 267562
rect 413344 267242 665026 267562
rect 413000 267218 413368 267242
rect 664994 267072 665026 267242
rect 668262 267562 668300 267722
rect 668262 267242 668488 267562
rect 668262 267072 668300 267242
rect 664994 267024 668300 267072
rect 666054 267016 667246 267024
rect 671660 266798 673470 266830
rect 671658 266786 673470 266798
rect 671578 266716 673470 266786
rect 671578 266634 671666 266716
rect 412528 266582 671666 266634
rect 412528 265796 647144 266582
rect 48980 265720 51440 265760
rect 48980 262254 49020 265720
rect 51400 265626 51440 265720
rect 181786 265644 193624 265654
rect 181786 265626 197682 265644
rect 51400 265614 406762 265626
rect 51400 262254 181826 265614
rect 48980 262214 181826 262254
rect 49574 262188 181826 262214
rect 181420 261204 181826 262188
rect 193584 265166 406762 265614
rect 193584 261204 211832 265166
rect 181420 261176 211832 261204
rect 212882 264300 406762 265166
rect 411638 265124 647144 265796
rect 654338 265124 671666 266582
rect 411638 265070 671666 265124
rect 411638 265064 412568 265070
rect 573184 264438 577694 264478
rect 432388 264388 436506 264428
rect 411832 264300 412460 264312
rect 422480 264300 426788 264332
rect 432388 264300 432428 264388
rect 212882 264292 432428 264300
rect 212882 264272 422520 264292
rect 212882 261176 411872 264272
rect 181420 261174 411872 261176
rect 412420 261214 422520 264272
rect 426748 261214 432428 264292
rect 412420 261174 432428 261214
rect 181420 261166 432428 261174
rect 436466 264300 436506 264388
rect 442152 264314 446456 264354
rect 442152 264300 442192 264314
rect 436466 261166 442192 264300
rect 181420 261130 442192 261166
rect 432388 261126 436506 261130
rect 442152 261084 442192 261130
rect 446416 264300 446456 264314
rect 452868 264318 457092 264358
rect 492504 264356 497138 264396
rect 452868 264300 452908 264318
rect 446416 261168 452908 264300
rect 457052 264300 457092 264318
rect 463502 264314 467226 264354
rect 463502 264300 463542 264314
rect 457052 261250 463542 264300
rect 467186 264300 467226 264314
rect 472646 264314 477196 264354
rect 472646 264300 472686 264314
rect 467186 261250 472686 264300
rect 457052 261168 472686 261250
rect 477156 264300 477196 264314
rect 492504 264300 492544 264356
rect 477156 264232 492544 264300
rect 477156 261208 482780 264232
rect 487996 261208 492544 264232
rect 477156 261168 492544 261208
rect 497098 264300 497138 264356
rect 522748 264314 527382 264354
rect 542774 264318 547492 264358
rect 502518 264300 507730 264314
rect 522748 264300 522788 264314
rect 497098 264274 522788 264300
rect 497098 261168 502558 264274
rect 446416 261130 502558 261168
rect 446416 261084 446456 261130
rect 452868 261128 457092 261130
rect 472646 261128 477196 261130
rect 492504 261128 497138 261130
rect 502518 261126 502558 261130
rect 507690 264232 522788 264274
rect 507690 261130 511908 264232
rect 507690 261126 507730 261130
rect 502518 261086 507730 261126
rect 511868 261126 511908 261130
rect 517454 261168 522788 264232
rect 527342 264300 527382 264314
rect 532638 264300 537436 264314
rect 542774 264300 542814 264318
rect 527342 264274 542814 264300
rect 527342 261168 532678 264274
rect 517454 261130 532678 261168
rect 517454 261126 517494 261130
rect 522748 261128 527382 261130
rect 511868 261086 517494 261126
rect 442152 261044 446456 261084
rect 532638 261084 532678 261130
rect 537396 261208 542814 264274
rect 547452 264300 547492 264318
rect 552496 264300 557876 264314
rect 573184 264300 573224 264438
rect 547452 264274 573224 264300
rect 547452 261208 552536 264274
rect 557836 264150 573224 264274
rect 557836 261208 562962 264150
rect 537396 261130 562962 261208
rect 537396 261084 537436 261130
rect 562922 261126 562962 261130
rect 567434 261130 573224 264150
rect 567434 261126 567474 261130
rect 562922 261086 567474 261126
rect 573184 261126 573224 261130
rect 577654 264300 577694 264438
rect 582782 264398 587748 264438
rect 582782 264300 582822 264398
rect 577654 261130 582822 264300
rect 577654 261126 577694 261130
rect 573184 261086 577694 261126
rect 532638 261044 537436 261084
rect 582782 261084 582822 261130
rect 587708 264300 587748 264398
rect 592298 264398 596890 264438
rect 592298 264300 592338 264398
rect 587708 261168 592338 264300
rect 596850 264300 596890 264398
rect 602600 264314 606820 264354
rect 602600 264300 602640 264314
rect 596850 261168 602640 264300
rect 587708 261130 602640 261168
rect 587708 261084 587748 261130
rect 592298 261128 596890 261130
rect 582782 261044 587748 261084
rect 602600 261044 602640 261130
rect 606780 264300 606820 264314
rect 622708 264300 626970 264314
rect 632430 264300 637562 264314
rect 661092 264300 664206 264314
rect 606780 264274 664513 264300
rect 606780 264232 622748 264274
rect 606780 261250 613232 264232
rect 617372 261250 622748 264232
rect 606780 261168 622748 261250
rect 626930 261168 632470 264274
rect 637522 261240 661132 264274
rect 664166 261240 664513 264274
rect 671578 262940 671666 265070
rect 673392 262940 673470 266716
rect 671578 262850 673470 262940
rect 671660 262816 673470 262850
rect 637522 261168 664513 261240
rect 606780 261130 664513 261168
rect 606780 261044 606820 261130
rect 622708 261128 626970 261130
rect 632430 261128 637562 261130
rect 602600 261004 606820 261044
rect 206950 259534 209064 259554
rect 416314 259552 424246 259592
rect 416314 259534 416354 259552
rect 48262 259514 416354 259534
rect 48262 259488 206990 259514
rect 48222 259448 206990 259488
rect 48222 256860 48262 259448
rect 54378 256918 206990 259448
rect 209024 256926 416354 259514
rect 424206 259534 424246 259552
rect 670582 259534 673406 259546
rect 424206 259506 673547 259534
rect 424206 256926 670622 259506
rect 209024 256918 670622 256926
rect 54378 256906 670622 256918
rect 673366 256906 673547 259506
rect 54378 256860 673547 256906
rect 48222 256820 54418 256860
rect 416290 256398 424314 256438
rect 206440 256368 209056 256374
rect 416290 256368 416330 256398
rect 50528 256334 416330 256368
rect 50528 256282 206480 256334
rect 50528 253286 50568 256282
rect 56050 253286 206480 256282
rect 50528 253280 206480 253286
rect 209016 253332 416330 256334
rect 424274 256368 424314 256398
rect 664958 256404 668374 256444
rect 664958 256368 664998 256404
rect 424274 253332 664998 256368
rect 209016 253308 664998 253332
rect 668334 256368 668374 256404
rect 668334 253308 668733 256368
rect 209016 253280 668733 253308
rect 50528 253246 668733 253280
rect 206440 253240 209056 253246
rect 641148 252616 656268 252656
rect 641148 249422 641188 252616
rect 656228 249422 656268 252616
rect 641148 249382 656268 249422
rect 488272 248666 491126 248706
rect 448158 248574 451474 248614
rect 45496 248490 47796 248530
rect 428124 248514 431026 248522
rect 448158 248514 448198 248574
rect 45496 248484 45536 248490
rect 45376 247120 45536 248484
rect 47756 248484 47796 248490
rect 194548 248484 448198 248514
rect 47756 248482 448198 248484
rect 47756 248416 428164 248482
rect 45376 244696 45520 247120
rect 45376 244520 45536 244696
rect 47756 244520 194614 248416
rect 45376 244450 194614 244520
rect 194574 240282 194614 244450
rect 206854 245954 428164 248416
rect 206854 244560 211886 245954
rect 206854 240282 206894 244560
rect 211846 244036 211886 244560
rect 215748 244938 428164 245954
rect 215748 244560 409646 244938
rect 215748 244036 215788 244560
rect 211846 243996 215788 244036
rect 409606 242868 409646 244560
rect 412718 242898 428164 244938
rect 430986 248310 448198 248482
rect 430986 242898 437744 248310
rect 412718 242868 437744 242898
rect 409606 242854 437744 242868
rect 409606 242844 413448 242854
rect 409606 242828 412758 242844
rect 437704 242806 437744 242854
rect 440486 242854 448198 248310
rect 440486 242806 440526 242854
rect 437704 242766 440526 242806
rect 448158 242806 448198 242854
rect 451434 248514 451474 248574
rect 458290 248586 461526 248626
rect 458290 248514 458330 248586
rect 451434 242898 458330 248514
rect 461486 248514 461526 248586
rect 468330 248552 471486 248592
rect 468330 248514 468370 248552
rect 461486 242944 468370 248514
rect 471446 248514 471486 248552
rect 478278 248528 481272 248568
rect 478278 248514 478318 248528
rect 471446 242944 478318 248514
rect 461486 242898 478318 242944
rect 481232 248514 481272 248528
rect 488272 248514 488312 248666
rect 481232 242898 488312 248514
rect 451434 242854 488312 242898
rect 451434 242806 451474 242854
rect 488272 242852 488312 242854
rect 491086 248514 491126 248666
rect 618192 248666 621324 248706
rect 498772 248586 501546 248626
rect 498772 248514 498812 248586
rect 491086 242854 498812 248514
rect 491086 242852 491126 242854
rect 488272 242812 491126 242852
rect 498772 242852 498812 242854
rect 501506 248514 501546 248586
rect 508122 248552 510816 248592
rect 538102 248574 541510 248614
rect 508122 248514 508162 248552
rect 501506 242898 508162 248514
rect 510776 248514 510816 248552
rect 517884 248528 521754 248568
rect 517884 248514 517924 248528
rect 510776 242898 517924 248514
rect 501506 242854 517924 242898
rect 501506 242852 501546 242854
rect 498772 242812 501546 242852
rect 517884 242852 517924 242854
rect 521714 248514 521754 248528
rect 538102 248514 538142 248574
rect 521714 248402 538142 248514
rect 521714 242854 527918 248402
rect 521714 242852 521754 242854
rect 517884 242812 521754 242852
rect 448158 242766 451474 242806
rect 527878 242806 527918 242854
rect 531628 242854 538142 248402
rect 531628 242806 531668 242854
rect 527878 242766 531668 242806
rect 538102 242806 538142 242854
rect 541470 248514 541510 248574
rect 547774 248540 551102 248580
rect 567578 248574 571862 248614
rect 547774 248514 547814 248540
rect 541470 242854 547814 248514
rect 541470 242806 541510 242854
rect 547774 242852 547814 242854
rect 551062 248514 551102 248540
rect 557170 248528 561268 248568
rect 557170 248514 557210 248528
rect 551062 242898 557210 248514
rect 561228 248514 561268 248528
rect 567578 248514 567618 248574
rect 561228 242898 567618 248514
rect 551062 242854 567618 242898
rect 551062 242852 551102 242854
rect 547774 242812 551102 242852
rect 538102 242766 541510 242806
rect 567578 242806 567618 242854
rect 571822 248514 571862 248574
rect 588210 248574 591756 248614
rect 588210 248514 588250 248574
rect 571822 248436 588250 248514
rect 571822 242898 577106 248436
rect 581078 242898 588250 248436
rect 591716 248514 591756 248574
rect 597606 248528 601474 248568
rect 597606 248514 597646 248528
rect 591716 242898 597646 248514
rect 601434 248514 601474 248528
rect 618192 248514 618232 248666
rect 601434 248448 618232 248514
rect 601434 242898 607364 248448
rect 611072 242898 618232 248448
rect 621284 248514 621324 248666
rect 627864 248528 631594 248568
rect 627864 248514 627904 248528
rect 621284 242898 627904 248514
rect 571822 242854 627904 242898
rect 571822 242806 571862 242854
rect 627864 242852 627904 242854
rect 631554 248514 631594 248528
rect 656722 248516 660622 248522
rect 656700 248514 660622 248516
rect 631554 248482 660631 248514
rect 631554 248476 656762 248482
rect 631554 244612 656740 248476
rect 631554 242888 656762 244612
rect 660582 244560 660631 248482
rect 660582 242888 660622 244560
rect 631554 242854 660622 242888
rect 631554 242852 631594 242854
rect 627864 242812 631594 242852
rect 656722 242848 660622 242854
rect 567578 242766 571862 242806
rect 194574 240242 206894 240282
rect 6598 227040 19088 239560
rect 42488 239410 45170 239658
rect 42488 239408 43732 239410
rect 42488 239398 43722 239408
rect 42488 239366 43714 239398
rect 44458 239366 45170 239410
rect 42488 237972 42530 239366
rect 45096 238568 45170 239366
rect 45096 238248 52450 238568
rect 45096 237972 45170 238248
rect 42488 237850 45170 237972
rect 698512 236640 711002 249160
rect 638768 234294 644334 234334
rect 45544 233890 47826 233928
rect 45544 232804 45600 233890
rect 47800 233568 47826 233890
rect 47800 233248 53596 233568
rect 47800 232804 47826 233248
rect 45544 232746 47826 232804
rect 194502 230162 206886 230202
rect 42454 229084 45136 229332
rect 42454 229082 43698 229084
rect 42454 229072 43688 229082
rect 42454 229040 43680 229072
rect 44424 229040 45136 229084
rect 42454 227646 42496 229040
rect 45062 228568 45136 229040
rect 45062 228248 52574 228568
rect 45062 227646 45136 228248
rect 194502 227718 194542 230162
rect 42454 227524 45136 227646
rect 194072 227398 194542 227718
rect 194502 224480 194542 227398
rect 206846 227718 206886 230162
rect 638768 227718 638808 234294
rect 206846 227398 215992 227718
rect 638640 227398 638808 227718
rect 206846 224480 206886 227398
rect 638768 226138 638808 227398
rect 644294 226138 644334 234294
rect 638768 226098 644334 226138
rect 194502 224440 206886 224480
rect 45532 223968 47814 224006
rect 45532 222882 45588 223968
rect 47788 223568 47814 223968
rect 47788 223248 53852 223568
rect 47788 222882 47814 223248
rect 45532 222824 47814 222882
rect 42476 218758 45158 219006
rect 42476 218756 43720 218758
rect 42476 218746 43710 218756
rect 42476 218714 43702 218746
rect 44446 218714 45158 218758
rect 42476 217320 42518 218714
rect 45084 218568 45158 218714
rect 45084 218248 52574 218568
rect 45084 217320 45158 218248
rect 42476 217198 45158 217320
rect 181688 216660 193642 216700
rect 45558 213990 47854 214028
rect 45558 212904 45614 213990
rect 47814 213642 47854 213990
rect 47814 213568 47860 213642
rect 47814 213248 52526 213568
rect 47814 212904 47854 213248
rect 45558 212846 47854 212904
rect 181688 212400 181728 216660
rect 180840 212080 181728 212400
rect 42500 209078 45182 209326
rect 42500 209076 43744 209078
rect 42500 209066 43734 209076
rect 42500 209034 43726 209066
rect 44470 209034 45182 209078
rect 42500 207640 42542 209034
rect 45108 208568 45182 209034
rect 45108 208248 52658 208568
rect 45108 207640 45182 208248
rect 42500 207518 45182 207640
rect 181688 206248 181728 212080
rect 193602 212400 193642 216660
rect 645312 215654 651246 215694
rect 645312 212400 645352 215654
rect 193602 212080 216852 212400
rect 638806 212080 645352 212400
rect 193602 206248 193642 212080
rect 645312 210840 645352 212080
rect 651206 210840 651246 215654
rect 645312 210800 651246 210840
rect 181688 206208 193642 206248
rect 45558 203662 47854 203700
rect 45558 202576 45614 203662
rect 47814 203568 47854 203662
rect 47814 203248 52568 203568
rect 47814 202994 47860 203248
rect 47814 202576 47854 202994
rect 45558 202518 47854 202576
rect 194502 202814 206972 202854
rect 42478 199138 45160 199386
rect 42478 199136 43722 199138
rect 42478 199126 43712 199136
rect 42478 199094 43704 199126
rect 44448 199094 45160 199138
rect 42478 197700 42520 199094
rect 45086 198568 45160 199094
rect 45086 198248 52658 198568
rect 45086 197700 45160 198248
rect 42478 197578 45160 197700
rect 194502 197082 194542 202814
rect 194170 196762 194542 197082
rect 6598 183840 19088 196360
rect 45558 193878 47854 193916
rect 45558 192792 45614 193878
rect 47814 193568 47854 193878
rect 47814 193248 52740 193568
rect 47814 193210 47860 193248
rect 47814 192792 47854 193210
rect 45558 192734 47854 192792
rect 194502 192744 194542 196762
rect 206932 197082 206972 202814
rect 638672 198466 644332 198506
rect 638672 197082 638712 198466
rect 206932 196762 216680 197082
rect 638340 196762 638712 197082
rect 206932 192744 206972 196762
rect 638672 194640 638712 196762
rect 644292 194640 644332 198466
rect 638672 194600 644332 194640
rect 194502 192704 206972 192744
rect 698512 191440 711002 203960
rect 42442 189050 45924 189298
rect 42442 189048 43726 189050
rect 42442 189038 43716 189048
rect 42442 189006 43708 189038
rect 44452 189006 45924 189050
rect 42442 187612 42524 189006
rect 45090 188568 45924 189006
rect 45090 188248 52782 188568
rect 45090 187612 45924 188248
rect 42442 187490 45924 187612
rect 181774 185790 193562 185830
rect 45558 184092 47854 184130
rect 45558 183006 45614 184092
rect 47814 183744 47854 184092
rect 47814 183568 47860 183744
rect 47814 183248 52482 183568
rect 47814 183006 47854 183248
rect 45558 182948 47854 183006
rect 181774 181764 181814 185790
rect 181098 181444 181814 181764
rect 43690 179104 44490 179134
rect 42498 179102 45172 179104
rect 42498 179100 43738 179102
rect 42498 179090 43728 179100
rect 42498 179058 43720 179090
rect 44464 179058 45172 179102
rect 42498 177664 42536 179058
rect 45102 178568 45172 179058
rect 45102 178248 52450 178568
rect 45102 177976 45174 178248
rect 45102 177664 45172 177976
rect 42498 177584 45172 177664
rect 181774 174942 181814 181444
rect 193522 181764 193562 185790
rect 645312 184342 651166 184382
rect 645312 181764 645352 184342
rect 193522 181444 215992 181764
rect 635556 181444 645352 181764
rect 193522 174942 193562 181444
rect 645312 179608 645352 181444
rect 651126 179608 651166 184342
rect 645312 179568 651166 179608
rect 181774 174902 193562 174942
rect 45558 173764 47854 173802
rect 45558 172678 45614 173764
rect 47814 173568 47854 173764
rect 47814 173248 52610 173568
rect 194674 173320 207064 173360
rect 47814 173096 47860 173248
rect 47814 172678 47854 173096
rect 45558 172620 47854 172678
rect 43686 169178 44486 169218
rect 42486 169176 45160 169178
rect 42486 169174 43726 169176
rect 42486 169132 43716 169174
rect 44452 169132 45160 169176
rect 42486 167738 42524 169132
rect 45090 168568 45160 169132
rect 45090 168248 52574 168568
rect 45090 168050 45162 168248
rect 45090 167738 45160 168050
rect 42486 167658 45160 167738
rect 194674 166446 194714 173320
rect 194170 166126 194714 166446
rect 45558 163980 47854 164018
rect 45558 162894 45614 163980
rect 47814 163632 47854 163980
rect 47814 163568 47860 163632
rect 47814 163248 52610 163568
rect 194674 163330 194714 166126
rect 207024 166446 207064 173320
rect 638602 168156 644342 168196
rect 638602 166446 638642 168156
rect 207024 166126 216508 166446
rect 638550 166126 638642 166446
rect 207024 163330 207064 166126
rect 638602 164250 638642 166126
rect 644302 166446 644342 168156
rect 644302 166126 644442 166446
rect 644302 164250 644342 166126
rect 638602 164210 644342 164250
rect 194674 163290 207064 163330
rect 47814 162894 47854 163248
rect 45558 162836 47854 162894
rect 43684 159090 44484 159132
rect 42474 159088 45148 159090
rect 42474 159044 43714 159088
rect 44440 159044 45148 159088
rect 42474 157650 42512 159044
rect 45078 158568 45148 159044
rect 45078 158248 52450 158568
rect 45078 157962 45150 158248
rect 45078 157650 45148 157962
rect 42474 157570 45148 157650
rect 181688 155854 193556 155894
rect 45558 154196 47854 154234
rect 45558 153110 45614 154196
rect 47814 153848 47854 154196
rect 47814 153568 47860 153848
rect 47814 153248 52526 153568
rect 47814 153110 47854 153248
rect 45558 153052 47854 153110
rect 181688 151128 181728 155854
rect 181184 150808 181728 151128
rect 42464 149060 45138 149106
rect 42464 147666 42502 149060
rect 45068 148568 45138 149060
rect 45068 148248 52490 148568
rect 45068 147978 45140 148248
rect 45068 147666 45138 147978
rect 42464 147586 45138 147666
rect 181688 144926 181728 150808
rect 193516 151128 193556 155854
rect 645208 154070 650982 154110
rect 645208 151128 645248 154070
rect 193516 150808 216422 151128
rect 635824 150808 645248 151128
rect 193516 144926 193556 150808
rect 645208 149416 645248 150808
rect 650942 151128 650982 154070
rect 650942 150808 651098 151128
rect 650942 149416 650982 150808
rect 645208 149376 650982 149416
rect 698512 146440 711002 158960
rect 181688 144886 193556 144926
rect 45558 143868 47854 143906
rect 45558 142782 45614 143868
rect 47814 143568 47854 143868
rect 47814 143248 52526 143568
rect 47814 143200 47860 143248
rect 47814 142782 47854 143200
rect 45558 142724 47854 142782
rect 194588 141504 206898 141544
rect 42474 139238 45148 139284
rect 42474 137844 42512 139238
rect 45078 138568 45148 139238
rect 45078 138248 52490 138568
rect 45078 138156 45150 138248
rect 45078 137844 45148 138156
rect 42474 137764 45148 137844
rect 194588 135810 194628 141504
rect 194170 135490 194628 135810
rect 45558 134082 47854 134120
rect 45558 132996 45614 134082
rect 47814 133734 47854 134082
rect 47814 133568 47860 133734
rect 47814 133248 52526 133568
rect 47814 132996 47854 133248
rect 45558 132938 47854 132996
rect 194588 131594 194628 135490
rect 206858 135810 206898 141504
rect 638856 137000 644342 137040
rect 638856 135810 638896 137000
rect 206858 135490 215390 135810
rect 638604 135490 638896 135810
rect 206858 131594 206898 135490
rect 638856 133408 638896 135490
rect 644302 135810 644342 137000
rect 644302 135490 644390 135810
rect 644302 133408 644342 135490
rect 638856 133368 644342 133408
rect 194588 131554 206898 131594
rect 42464 129370 45138 129416
rect 42464 127976 42502 129370
rect 45068 128608 45138 129370
rect 45068 128568 45140 128608
rect 45068 128248 52658 128568
rect 45068 127976 45138 128248
rect 42464 127896 45138 127976
rect 181860 127140 193568 127180
rect 45558 123754 47854 123792
rect 45558 122668 45614 123754
rect 47814 123568 47854 123754
rect 47814 123248 52610 123568
rect 47814 123086 47860 123248
rect 47814 122668 47854 123086
rect 45558 122610 47854 122668
rect 181860 120492 181900 127140
rect 181270 120172 181900 120492
rect 42470 119330 45164 119376
rect 42470 117936 42528 119330
rect 45094 118568 45164 119330
rect 45094 118248 52574 118568
rect 45094 117936 45164 118248
rect 42470 117856 45164 117936
rect 181860 115426 181900 120172
rect 193528 120492 193568 127140
rect 645260 123540 650954 123580
rect 645260 120492 645300 123540
rect 193528 120172 216766 120492
rect 635772 120172 645300 120492
rect 193528 115426 193568 120172
rect 645260 118966 645300 120172
rect 650914 120492 650954 123540
rect 650914 120172 651148 120492
rect 650914 118966 650954 120172
rect 645260 118926 650954 118966
rect 181860 115386 193568 115426
rect 45626 114174 47922 114212
rect 45626 113568 45682 114174
rect 45524 113248 45682 113568
rect 45626 113088 45682 113248
rect 47882 113826 47922 114174
rect 47882 113568 47928 113826
rect 47882 113248 52610 113568
rect 47882 113088 47922 113248
rect 45626 113030 47922 113088
rect 194416 112852 206972 112892
rect 42422 109052 45104 109300
rect 42422 109050 43666 109052
rect 42422 109040 43656 109050
rect 42422 109008 43648 109040
rect 44392 109008 45104 109052
rect 42422 107614 42464 109008
rect 45030 108568 45104 109008
rect 45030 108248 52490 108568
rect 45030 107614 45104 108248
rect 42422 107492 45104 107614
rect 194416 105174 194456 112852
rect 194084 104854 194456 105174
rect 45626 103846 47922 103884
rect 45626 102760 45682 103846
rect 47882 103568 47922 103846
rect 47882 103248 52568 103568
rect 47882 103178 47928 103248
rect 47882 102760 47922 103178
rect 45626 102702 47922 102760
rect 194416 100374 194456 104854
rect 206932 105174 206972 112852
rect 638710 107164 644386 107204
rect 638710 105174 638750 107164
rect 206932 104854 217282 105174
rect 638288 104854 638750 105174
rect 206932 100374 206972 104854
rect 638710 103406 638750 104854
rect 644346 105174 644386 107164
rect 645280 105666 650876 105706
rect 644346 104854 644390 105174
rect 644346 103406 644386 104854
rect 638710 103366 644386 103406
rect 645280 101988 645320 105666
rect 650836 103700 650876 105666
rect 663776 103712 665548 103752
rect 663776 103700 663816 103712
rect 650836 101994 663816 103700
rect 665508 101994 665548 103712
rect 650836 101988 665548 101994
rect 645280 101954 665548 101988
rect 645280 101948 650876 101954
rect 698512 101240 711002 113760
rect 194416 100334 206972 100374
rect 42446 98966 45128 99214
rect 42446 98964 43690 98966
rect 42446 98954 43680 98964
rect 42446 98922 43672 98954
rect 44416 98922 45128 98966
rect 42446 97528 42488 98922
rect 45054 98568 45128 98922
rect 45054 98248 52782 98568
rect 45054 97528 45128 98248
rect 42446 97406 45128 97528
rect 181860 98150 193648 98190
rect 45614 93868 47910 93906
rect 45614 92782 45670 93868
rect 47870 93568 47910 93868
rect 47870 93248 52610 93568
rect 47870 93200 47916 93248
rect 47870 92782 47910 93200
rect 45614 92724 47910 92782
rect 181860 89856 181900 98150
rect 180926 89536 181900 89856
rect 42470 89142 45152 89388
rect 42470 89140 43720 89142
rect 42470 89138 43714 89140
rect 42470 89128 43704 89138
rect 42470 89096 43696 89128
rect 44446 89096 45152 89142
rect 42470 87702 42512 89096
rect 45078 88568 45152 89096
rect 45078 88248 52782 88568
rect 45078 87702 45152 88248
rect 42470 87580 45152 87702
rect 181860 86356 181900 89536
rect 193608 89856 193648 98150
rect 645468 92904 651082 92944
rect 645468 89856 645508 92904
rect 193608 89536 216078 89856
rect 638096 89536 645508 89856
rect 193608 86356 193648 89536
rect 645468 88410 645508 89536
rect 651042 88410 651082 92904
rect 645468 88370 651082 88410
rect 181860 86316 193648 86356
rect 638868 85142 644384 85182
rect 45642 83916 47938 83960
rect 45642 83568 45698 83916
rect 45566 83248 45698 83568
rect 45642 82830 45698 83248
rect 47898 83568 47938 83916
rect 47898 83248 52568 83568
rect 47898 82830 47938 83248
rect 45642 82772 47938 82830
rect 194416 83100 206892 83140
rect 6167 70054 19620 80934
rect 42382 79346 45064 79358
rect 40820 79288 45192 79346
rect 40820 77556 40888 79288
rect 45134 78568 45192 79288
rect 45134 78248 52866 78568
rect 45134 77556 45192 78248
rect 40820 77498 45192 77556
rect 194416 74538 194456 83100
rect 206852 83060 207062 83100
rect 194170 74218 194456 74538
rect 45628 73834 47894 73936
rect 45628 73568 45668 73834
rect 45566 73248 45668 73568
rect 45628 72892 45668 73248
rect 47790 73568 47894 73834
rect 47790 73248 52954 73568
rect 47790 73076 47914 73248
rect 47790 72892 47894 73076
rect 45628 72808 47894 72892
rect 194416 70702 194456 74218
rect 207022 74538 207062 83060
rect 638868 81544 638908 85142
rect 644344 83758 644384 85142
rect 644344 83438 658056 83758
rect 644344 81544 644384 83438
rect 645386 83008 650952 83048
rect 645386 82942 645426 83008
rect 645282 82622 645426 82942
rect 638868 81504 644384 81544
rect 645386 79336 645426 82622
rect 650912 82942 650952 83008
rect 650912 82622 658048 82942
rect 650912 79336 650952 82622
rect 645386 79296 650952 79336
rect 638766 76240 644418 76280
rect 207022 74218 217368 74538
rect 194416 70662 194520 70702
rect 40818 69384 45226 69476
rect 40818 67906 40900 69384
rect 45180 68568 45226 69384
rect 45180 68248 57696 68568
rect 45180 67906 45226 68248
rect 40818 67826 45226 67906
rect 45592 64006 47920 64108
rect 45592 63568 45694 64006
rect 45586 63248 45694 63568
rect 45592 63064 45694 63248
rect 47816 63568 47920 64006
rect 194480 63568 194520 70662
rect 47816 63248 52496 63568
rect 138920 63248 194520 63568
rect 47816 63064 47920 63248
rect 45592 62980 47920 63064
rect 181634 60778 193606 60818
rect 40728 59078 45176 59148
rect 40728 57596 40844 59078
rect 45106 58568 45176 59078
rect 181634 58568 181674 60778
rect 45106 58248 52462 58568
rect 137208 58248 181674 58568
rect 45106 57596 45176 58248
rect 40728 57480 45176 57596
rect 48386 55910 50870 55950
rect 48386 50098 48426 55910
rect 50830 55816 50870 55910
rect 50830 53272 180738 55816
rect 181634 54130 181674 58248
rect 193566 59220 193606 60778
rect 194480 60770 194520 63248
rect 207022 63568 207062 74218
rect 638766 72698 638806 76240
rect 644378 72698 644418 76240
rect 638766 72658 644418 72698
rect 207022 63248 207310 63568
rect 207022 60770 207062 63248
rect 194480 60730 207062 60770
rect 645350 60958 651026 60998
rect 645350 59220 645390 60958
rect 193566 58900 216336 59220
rect 638828 58900 645390 59220
rect 193566 54130 193606 58900
rect 645350 57944 645390 58900
rect 650986 57944 651026 60958
rect 645350 57904 651026 57944
rect 210560 55063 213568 55105
rect 210560 54827 210602 55063
rect 210838 54827 213290 55063
rect 213526 54827 213568 55063
rect 210560 54785 213568 54827
rect 181634 54090 193606 54130
rect 653418 53868 654906 53906
rect 194576 53866 654912 53868
rect 194576 53318 653458 53866
rect 192636 53272 653458 53318
rect 50830 52944 653458 53272
rect 50852 51598 653458 52944
rect 50852 50716 144490 51598
rect 144898 50716 653458 51598
rect 50852 50706 653458 50716
rect 654866 50706 654912 53866
rect 50852 50698 654912 50706
rect 50852 50666 654906 50698
rect 50852 50656 654836 50666
rect 50830 50098 194166 50656
rect 223428 50594 226328 50656
rect 48386 50058 194166 50098
rect 48422 50014 194166 50058
rect 180076 49978 194166 50014
rect 194608 49686 207080 49726
rect 45558 49566 48232 49658
rect 194608 49566 194648 49686
rect 45558 49544 194648 49566
rect 45558 46014 45634 49544
rect 48118 46198 194648 49544
rect 48118 46014 48232 46198
rect 194608 46166 194648 46198
rect 207040 49566 207080 49686
rect 517792 49676 521364 49716
rect 238310 49566 241012 49584
rect 245716 49566 251552 49584
rect 258044 49566 260962 49606
rect 278408 49588 280716 49628
rect 268128 49566 270966 49570
rect 278408 49566 278448 49588
rect 207040 49544 258084 49566
rect 207040 49524 238350 49544
rect 207040 46206 218530 49524
rect 220846 46228 228244 49524
rect 231018 46228 238350 49524
rect 240972 46228 245756 49544
rect 251512 48302 258084 49544
rect 251524 46272 258084 48302
rect 220846 46206 245756 46228
rect 207040 46198 245756 46206
rect 207040 46166 207080 46198
rect 218490 46166 220886 46198
rect 228204 46188 231058 46198
rect 238310 46188 241012 46198
rect 245716 46184 245756 46198
rect 251512 46198 258084 46272
rect 251512 46184 251552 46198
rect 194608 46158 198642 46166
rect 205416 46158 207080 46166
rect 194608 46126 207080 46158
rect 245716 46144 251552 46184
rect 258044 46184 258084 46198
rect 260922 49530 278448 49566
rect 260922 46228 268168 49530
rect 270926 46228 278448 49530
rect 260922 46198 278448 46228
rect 260922 46184 260962 46198
rect 268128 46188 270966 46198
rect 258044 46144 260962 46184
rect 278408 46184 278448 46198
rect 280676 49566 280716 49588
rect 288404 49566 290632 49592
rect 298336 49566 301038 49584
rect 327936 49566 331268 49606
rect 378072 49588 381558 49628
rect 348060 49566 351828 49584
rect 368098 49566 371648 49584
rect 378072 49566 378112 49588
rect 280676 49552 327976 49566
rect 280676 46228 288444 49552
rect 290592 49544 327976 49552
rect 290592 46292 298376 49544
rect 300998 49524 327976 49544
rect 300998 46292 308178 49524
rect 290592 46228 308178 46292
rect 311320 46228 317934 49524
rect 321622 46228 327976 49524
rect 331228 49544 378112 49566
rect 331228 49524 348100 49544
rect 331228 46228 337972 49524
rect 280676 46206 337972 46228
rect 341202 46248 348100 49524
rect 351788 49524 368138 49544
rect 351788 46248 357988 49524
rect 341202 46228 357988 46248
rect 361524 46248 368138 49524
rect 371608 46248 378112 49544
rect 381518 49566 381558 49588
rect 397914 49588 401290 49628
rect 397914 49566 397954 49588
rect 381518 49524 397954 49566
rect 381518 46248 388110 49524
rect 391296 46248 397954 49524
rect 361524 46228 397954 46248
rect 341202 46206 397954 46228
rect 280676 46198 397954 46206
rect 280676 46184 280716 46198
rect 288404 46188 290632 46198
rect 308138 46188 311360 46198
rect 317894 46188 321662 46198
rect 327936 46188 331268 46198
rect 278408 46144 280716 46184
rect 337932 46166 341242 46198
rect 357948 46188 361564 46198
rect 397914 46184 397954 46198
rect 401250 49566 401290 49588
rect 417342 49566 421262 49584
rect 427884 49566 431674 49584
rect 437380 49566 441300 49606
rect 447856 49588 451580 49628
rect 447856 49566 447896 49588
rect 401250 49544 437420 49566
rect 401250 49524 417382 49544
rect 401250 46270 407602 49524
rect 411270 46270 417382 49524
rect 401250 46248 417382 46270
rect 421222 46248 427924 49544
rect 401250 46228 427924 46248
rect 431634 46228 437420 49544
rect 441260 46248 447896 49566
rect 451540 49566 451580 49588
rect 458332 49566 461556 49584
rect 467980 49566 470376 49584
rect 478610 49566 481114 49584
rect 498320 49566 501348 49606
rect 517792 49566 517832 49676
rect 451540 49544 498360 49566
rect 451540 46248 458372 49544
rect 441260 46228 458372 46248
rect 461516 46270 468020 49544
rect 470336 46270 478650 49544
rect 461516 46248 478650 46270
rect 481074 49524 498360 49544
rect 481074 46248 488580 49524
rect 461516 46228 488580 46248
rect 401250 46198 488580 46228
rect 401250 46184 401290 46198
rect 427884 46188 431674 46198
rect 437380 46188 441300 46198
rect 458332 46188 461556 46198
rect 397914 46144 401290 46184
rect 488540 46184 488580 46198
rect 490810 46270 498360 49524
rect 501308 49502 517832 49566
rect 501308 46270 508314 49502
rect 490810 46248 508314 46270
rect 511566 46248 517832 49502
rect 490810 46198 517832 46248
rect 490810 46184 490850 46198
rect 488540 46144 490850 46184
rect 517792 46184 517832 46198
rect 521324 49566 521364 49676
rect 597974 49634 601444 49674
rect 537546 49566 541402 49584
rect 597974 49566 598014 49634
rect 521324 49544 598014 49566
rect 521324 49480 537586 49544
rect 521324 46198 527784 49480
rect 521324 46184 521364 46198
rect 517792 46144 521364 46184
rect 527744 46184 527784 46198
rect 531408 46228 537586 49480
rect 541362 46352 598014 49544
rect 601404 49566 601444 49634
rect 628222 49580 631692 49620
rect 628222 49566 628262 49580
rect 601404 49500 628262 49566
rect 601404 46352 607988 49500
rect 541362 46298 607988 46352
rect 611298 49420 628262 49500
rect 611298 46298 618342 49420
rect 621572 46298 628262 49420
rect 541362 46244 628262 46298
rect 631652 49566 631692 49580
rect 638922 49566 644408 49578
rect 631652 49474 644408 49566
rect 631652 46262 639000 49474
rect 644086 46262 644408 49474
rect 631652 46244 644408 46262
rect 541362 46228 644408 46244
rect 531408 46210 644408 46228
rect 645230 46688 651392 46728
rect 531408 46198 644054 46210
rect 531408 46184 531448 46198
rect 537546 46188 541402 46198
rect 527744 46144 531448 46184
rect 198602 46118 205456 46126
rect 45558 45912 48232 46014
rect 40806 45668 45186 45740
rect 40762 45628 45226 45668
rect 40762 40944 40802 45628
rect 45186 45526 45226 45628
rect 613316 45624 616678 45664
rect 181886 45584 196032 45624
rect 143818 45526 145850 45540
rect 181886 45526 181926 45584
rect 45186 45500 181926 45526
rect 45186 45200 143858 45500
rect 45186 43084 143852 45200
rect 45186 43054 143858 43084
rect 145810 43070 181926 45500
rect 195992 45526 196032 45584
rect 213090 45526 216424 45548
rect 603016 45526 606298 45530
rect 613316 45526 613356 45624
rect 195992 45508 613356 45526
rect 195992 43070 213130 45508
rect 145810 43054 213130 43070
rect 45186 43030 213130 43054
rect 216384 45490 613356 45508
rect 216384 45480 603056 45490
rect 216384 45464 323470 45480
rect 216384 45352 273300 45464
rect 216384 45272 253530 45352
rect 216384 45192 241992 45272
rect 216384 45112 232944 45192
rect 216384 43120 223370 45112
rect 226464 43120 232944 45112
rect 236118 43120 241992 45192
rect 245246 43120 253530 45272
rect 256864 45336 273300 45352
rect 256864 43120 262720 45336
rect 216384 43030 262720 43120
rect 45186 43024 262720 43030
rect 266134 43072 273300 45336
rect 276794 45434 323470 45464
rect 276794 45402 293024 45434
rect 276794 43072 282922 45402
rect 266134 43024 282922 43072
rect 45186 43020 282922 43024
rect 45186 40944 140470 43020
rect 143818 43014 145850 43020
rect 213090 42990 216424 43020
rect 262680 42984 266174 43020
rect 282882 42930 282922 43020
rect 286496 43020 293024 45402
rect 286496 42930 286536 43020
rect 282882 42890 286536 42930
rect 292984 42882 293024 43020
rect 296678 45338 323470 45434
rect 296678 45162 313416 45338
rect 296678 43024 303508 45162
rect 306174 43120 313416 45162
rect 316162 43120 323470 45338
rect 306174 43024 323470 43120
rect 296678 43020 323470 43024
rect 296678 42882 296718 43020
rect 303468 42984 306214 43020
rect 323430 42976 323470 43020
rect 326550 45410 603056 45480
rect 326550 45386 592974 45410
rect 326550 45290 343002 45386
rect 326550 43072 332518 45290
rect 335980 43072 343002 45290
rect 326550 43020 343002 43072
rect 326550 42976 326590 43020
rect 323430 42936 326590 42976
rect 342962 42930 343002 43020
rect 346272 45320 373208 45386
rect 346272 43024 353150 45320
rect 355926 45258 373208 45320
rect 355926 43024 363012 45258
rect 346272 43020 363012 43024
rect 346272 42930 346312 43020
rect 353110 42984 355966 43020
rect 342962 42890 346312 42930
rect 292984 42842 296718 42882
rect 362972 42882 363012 43020
rect 365868 43020 373208 45258
rect 365868 42882 365908 43020
rect 373168 42930 373208 43020
rect 376144 45338 592974 45386
rect 376144 45290 443100 45338
rect 376144 43072 382878 45290
rect 386244 43072 393218 45290
rect 376144 43020 393218 43072
rect 376144 42930 376184 43020
rect 393178 42976 393218 43020
rect 396250 43020 402410 45290
rect 396250 42976 396290 43020
rect 393178 42936 396290 42976
rect 402370 42976 402410 43020
rect 405824 45258 443100 45290
rect 405824 45242 433192 45258
rect 405824 43020 413372 45242
rect 405824 42976 405864 43020
rect 402370 42936 405864 42976
rect 373168 42890 376184 42930
rect 413332 42930 413372 43020
rect 416212 45226 433192 45242
rect 416212 43072 423090 45226
rect 425914 43072 433192 45226
rect 416212 43024 433192 43072
rect 436096 43024 443100 45258
rect 446084 45332 592974 45338
rect 446084 45314 503498 45332
rect 446084 45210 463500 45314
rect 446084 43120 453344 45210
rect 456344 43120 463500 45210
rect 446084 43024 463500 43120
rect 416212 43020 463500 43024
rect 416212 42930 416252 43020
rect 433152 42984 436136 43020
rect 443060 42984 446124 43020
rect 463460 43010 463500 43020
rect 465734 45290 503498 45314
rect 465734 45242 483074 45290
rect 465734 43104 473898 45242
rect 475988 43120 483074 45242
rect 486056 43120 492934 45290
rect 496014 43120 503498 45290
rect 475988 43104 503498 43120
rect 465734 43020 503498 43104
rect 465734 43010 465774 43020
rect 463460 42970 465774 43010
rect 503458 42996 503498 43020
rect 506214 43138 513212 45332
rect 516308 45266 543776 45332
rect 516308 43184 523684 45266
rect 525578 45204 543776 45266
rect 525578 43184 533968 45204
rect 516308 43138 533968 43184
rect 506214 43090 513734 43138
rect 515548 43090 533968 43138
rect 506214 43042 533968 43090
rect 535942 43090 543776 45204
rect 545830 43090 592974 45332
rect 535942 43046 592974 43090
rect 596096 43046 603056 45410
rect 606258 43100 613356 45490
rect 616638 45526 616678 45624
rect 623180 45596 626622 45636
rect 623180 45526 623220 45596
rect 616638 43100 623220 45526
rect 606258 43046 623220 43100
rect 535942 43042 623220 43046
rect 506214 43020 623220 43042
rect 506214 42996 506254 43020
rect 533928 43002 535982 43020
rect 592934 43006 596136 43020
rect 603016 43006 606298 43020
rect 503458 42956 506254 42996
rect 623180 42992 623220 43020
rect 626582 45526 626622 45596
rect 633156 45622 636678 45662
rect 633156 45526 633196 45622
rect 626582 43020 633196 45526
rect 626582 42992 626622 43020
rect 623180 42952 626622 42992
rect 413332 42890 416252 42930
rect 633156 42938 633196 43020
rect 636638 45526 636678 45622
rect 645230 45526 645270 46688
rect 636638 43036 645270 45526
rect 651352 43036 651392 46688
rect 636638 43026 645372 43036
rect 650996 43026 651392 43036
rect 636638 43020 651392 43026
rect 636638 42938 636678 43020
rect 645230 42972 651392 43020
rect 645256 42962 651104 42972
rect 633156 42898 636678 42938
rect 362972 42842 365908 42882
rect 40762 40942 140470 40944
rect 141966 42510 144024 42534
rect 573604 42510 579176 42556
rect 651666 42510 653770 42524
rect 141966 42494 653770 42510
rect 40762 40904 45226 40942
rect 141966 40624 142006 42494
rect 143984 42492 653770 42494
rect 143984 40714 573714 42492
rect 143984 40624 239404 40714
rect 141966 40584 239404 40624
rect 141972 39934 239404 40584
rect 241412 40344 573714 40714
rect 579078 42484 653770 42492
rect 579078 40344 651706 42484
rect 241412 39978 651706 40344
rect 653730 39978 653770 42484
rect 241412 39938 653770 39978
rect 241412 39934 653756 39938
rect 154784 39924 173378 39934
rect 80222 6811 92390 18976
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 624222 6811 636390 18976
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use copyright_block  copyright_block_0
timestamp 1608325192
transform 1 0 149582 0 1 16298
box -262 -9464 35048 2764
use storage  storage
timestamp 1613304178
transform 1 0 52032 0 1 53156
box 0 0 88934 189234
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1608587411
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use open_source  open_source_0
timestamp 1613162426
transform 1 0 205230 0 1 2174
box 752 5164 29030 16242
use user_id_programming  user_id_value
timestamp 1606755340
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use simple_por  por
timestamp 1606688983
transform 1 0 654146 0 -1 112882
box 0 0 11344 8338
use gpio_control_block  gpio_control_bidir\[0\]
timestamp 1611581575
transform -1 0 708603 0 1 121000
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_bidir\[1\]
timestamp 1611581575
transform -1 0 708603 0 1 166200
box -1664 -364 34000 13964
use mgmt_core  soc
timestamp 1608935209
transform 1 0 210434 0 1 53602
box 0 0 430000 180000
use gpio_control_block  gpio_control_in\[37\]
timestamp 1611581575
transform 1 0 8567 0 1 202600
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[36\]
timestamp 1611581575
transform 1 0 8567 0 1 245800
box -1664 -364 34000 13964
use mgmt_protect  mgmt_buffers
timestamp 1608143532
transform 1 0 212180 0 1 246836
box -2762 -2778 202678 20730
use gpio_control_block  gpio_control_in\[3\]
timestamp 1611581575
transform -1 0 708603 0 1 256400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[2\]
timestamp 1611581575
transform -1 0 708603 0 1 211200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[35\]
timestamp 1611581575
transform 1 0 8567 0 1 289000
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[34\]
timestamp 1611581575
transform 1 0 8567 0 1 332200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[33\]
timestamp 1611581575
transform 1 0 8567 0 1 375400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[5\]
timestamp 1611581575
transform -1 0 708603 0 1 346400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[4\]
timestamp 1611581575
transform -1 0 708603 0 1 301400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[7\]
timestamp 1611581575
transform -1 0 708603 0 1 479800
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[6\]
timestamp 1611581575
transform -1 0 708603 0 1 391600
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[32\]
timestamp 1611581575
transform 1 0 8567 0 1 418600
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[31\]
timestamp 1611581575
transform 1 0 8567 0 1 546200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[30\]
timestamp 1611581575
transform 1 0 8567 0 1 589400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[29\]
timestamp 1611581575
transform 1 0 8567 0 1 632600
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[9\]
timestamp 1611581575
transform -1 0 708603 0 1 568800
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[8\]
timestamp 1611581575
transform -1 0 708603 0 1 523800
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[10\]
timestamp 1611581575
transform -1 0 708603 0 1 614000
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[28\]
timestamp 1611581575
transform 1 0 8567 0 1 675800
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[27\]
timestamp 1611581575
transform 1 0 8567 0 1 719000
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[26\]
timestamp 1611581575
transform 1 0 8567 0 1 762200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[13\]
timestamp 1611581575
transform -1 0 708603 0 1 749200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[12\]
timestamp 1611581575
transform -1 0 708603 0 1 704200
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[11\]
timestamp 1611581575
transform -1 0 708603 0 1 659000
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[25\]
timestamp 1611581575
transform 1 0 8567 0 1 805400
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[24\]
timestamp 1611581575
transform 1 0 8567 0 1 931224
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[23\]
timestamp 1611581575
transform 0 1 97200 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[22\]
timestamp 1611581575
transform 0 1 148600 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[21\]
timestamp 1611581575
transform 0 1 200000 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[20\]
timestamp 1611581575
transform 0 1 251400 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[19\]
timestamp 1611581575
transform 0 1 303000 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[18\]
timestamp 1611581575
transform 0 1 353400 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[17\]
timestamp 1611581575
transform 0 1 420800 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[16\]
timestamp 1611581575
transform 0 1 497800 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[15\]
timestamp 1611581575
transform 0 1 549200 -1 0 1029813
box -1664 -364 34000 13964
use gpio_control_block  gpio_control_in\[14\]
timestamp 1611581575
transform -1 0 708603 0 1 927600
box -1664 -364 34000 13964
use chip_io  padframe
timestamp 1613148814
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_project_wrapper  mprj
timestamp 1610388215
transform 1 0 65308 0 1 278718
box -8576 -7506 592500 711442
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 44 nsew signal input
rlabel metal3 s 39593 120278 39999 125058 6 vddio
port 54 nsew signal bidirectional
rlabel metal2 s 225172 53602 225228 54402 6 pwr_ctrl_out[0]
port 59 nsew signal tristate
rlabel metal2 s 225540 53602 225596 54402 6 pwr_ctrl_out[1]
port 60 nsew signal tristate
rlabel metal2 s 225908 53602 225964 54402 6 pwr_ctrl_out[2]
port 61 nsew signal tristate
rlabel metal2 s 226276 53602 226332 54402 6 pwr_ctrl_out[3]
port 62 nsew signal tristate
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 80222 6811 92390 18976 1 vssa
port 63 n
rlabel metal5 243266 6167 254146 19620 1 vssd
port 64 n
rlabel metal5 624222 6811 636390 18976 1 vdda
port 65 n
rlabel metal5 697980 461866 711433 472746 1 vssd1
port 66 n
rlabel metal5 698624 819822 710789 831990 1 vdda1
port 67 n
rlabel metal5 697980 909666 711433 920546 1 vccd1
port 68 n
rlabel metal5 577010 1018624 589178 1030789 1 vssa1
port 69 n
rlabel metal5 334810 1018624 346978 1030789 1 vssio
port 70 n
rlabel metal5 6167 914054 19620 924934 1 vccd2
port 71 n
rlabel metal5 6811 829010 18976 841178 1 vssa2
port 72 n
rlabel metal5 6811 484410 18976 496578 1 vdda2
port 73 n
rlabel metal5 6167 442854 19620 453734 1 vssd2
port 74 n
rlabel metal5 6167 70054 19620 80934 1 vccd
port 75 n
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
