magic
tech micross
magscale 1 2
timestamp 1611856895
<< checkpaint >>
rect -26897 -26897 38184 26897
<< rdl >>
tri -6988 26080 -2353 26897 se
rect -2353 26080 2353 26897
tri 2353 26080 6988 26897 sw
tri -11411 24470 -6988 26080 se
rect -6988 24470 6988 26080
tri 6988 24470 11411 26080 sw
tri -15487 22117 -11411 24470 se
rect -11411 22117 11411 24470
tri 11411 22117 15487 24470 sw
tri -15626 22000 -15487 22117 se
rect -15487 22000 15487 22117
tri 15487 22000 15626 22117 sw
tri -16024 21666 -15626 22000 se
rect -15626 21666 -3820 22000
tri -3820 21666 0 22000 nw
tri 0 21666 3820 22000 ne
rect 3820 21666 15626 22000
tri 15626 21666 16024 22000 sw
tri -17208 20673 -16024 21666 se
rect -16024 20673 -7524 21666
tri -7524 20673 -3820 21666 nw
tri 3820 20673 7524 21666 ne
rect 7524 20673 16024 21666
tri 16024 20673 17207 21666 sw
tri -19092 19092 -17208 20673 se
rect -17208 19092 -10916 20673
tri -10916 19092 -7524 20673 nw
tri 7524 19092 10916 20673 ne
rect 10916 19092 17207 20673
tri 17207 19092 19092 20673 sw
tri -19125 19053 -19092 19092 se
rect -19092 19053 -11000 19092
tri -11000 19053 -10916 19092 nw
tri 10916 19053 11000 19092 ne
rect 11000 19053 19092 19092
tri 19092 19053 19131 19092 sw
tri -20971 16853 -19125 19053 se
rect -19125 16853 -14141 19053
tri -14141 16853 -11000 19053 nw
tri 11000 16853 14141 19053 ne
rect 14141 16853 19131 19053
tri 19131 16853 21331 19053 sw
tri -22117 15487 -20971 16853 se
rect -20971 15487 -15507 16853
tri -15507 15487 -14141 16853 nw
tri 14141 15487 15507 16853 ne
rect 15507 15487 21331 16853
tri -22894 14141 -22117 15487 se
rect -22117 14141 -16853 15487
tri -16853 14141 -15507 15487 nw
tri 15507 14141 16853 15487 ne
rect 16853 14141 21331 15487
tri 21331 14141 24043 16853 sw
tri -24470 11411 -22894 14141 se
rect -22894 11411 -18765 14141
tri -18765 11411 -16853 14141 nw
tri 16853 11411 18765 14141 ne
rect 18765 11411 24043 14141
tri -24620 11000 -24470 11411 se
rect -24470 11000 -19053 11411
tri -19053 11000 -18765 11411 nw
tri 18765 11000 19053 11411 ne
rect 19053 11000 24043 11411
tri 24043 11000 27184 14141 sw
tri -25885 7524 -24620 10999 se
rect -24620 7524 -20673 11000
tri -20673 7524 -19053 11000 nw
tri 19053 10916 19092 11000 ne
rect 19092 10916 27184 11000
tri 27184 10916 27268 11000 sw
tri 19092 7524 20673 10916 ne
rect 20673 7524 27268 10916
tri 27268 7524 30660 10916 sw
tri -26080 6988 -25885 7524 se
rect -25885 6988 -20817 7524
tri -20817 6988 -20673 7524 nw
tri -26638 3822 -26080 6988 se
rect -26080 3822 -21666 6988
rect -26638 3820 -21666 3822
tri -21666 3820 -20817 6988 nw
tri 20673 3820 21666 7524 ne
rect 21666 3820 30660 7524
tri 30660 3820 34364 7524 sw
tri -26897 2353 -26638 3820 se
rect -26638 2353 -21794 3820
tri -21794 2353 -21666 3820 nw
rect -26897 -2353 -22000 2353
tri -22000 0 -21794 2353 nw
tri -22000 -2353 -21794 0 sw
tri 21666 0 22000 3820 ne
tri -26897 -3817 -26639 -2353 ne
rect -26639 -3820 -21794 -2353
tri -21794 -3820 -21666 -2353 sw
tri 21666 -3820 22000 0 se
rect 22000 -3820 34364 3820
tri 34364 0 38184 3820 sw
tri 34364 -3820 38184 0 nw
tri -26639 -6988 -26080 -3820 ne
rect -26080 -6988 -21666 -3820
tri -21666 -6988 -20817 -3820 sw
tri -26080 -7524 -25885 -6988 ne
rect -25885 -7524 -20817 -6988
tri -20817 -7524 -20673 -6988 sw
tri 20673 -7524 21666 -3820 se
rect 21666 -7524 30660 -3820
tri 30660 -7524 34364 -3820 nw
tri -25885 -10999 -24620 -7524 ne
rect -24620 -11000 -20673 -7524
tri -20673 -11000 -19053 -7524 sw
tri 19092 -10916 20673 -7524 se
rect 20673 -10916 27268 -7524
tri 27268 -10916 30660 -7524 nw
tri 19053 -11000 19092 -10916 se
rect 19092 -11000 27184 -10916
tri 27184 -11000 27268 -10916 nw
tri -24620 -11411 -24470 -11000 ne
rect -24470 -11411 -19053 -11000
tri -19053 -11411 -18765 -11000 sw
tri 18765 -11411 19053 -11000 se
rect 19053 -11411 24043 -11000
tri -24470 -14140 -22895 -11411 ne
rect -22895 -14141 -18765 -11411
tri -18765 -14141 -16853 -11411 sw
tri 16853 -14141 18765 -11411 se
rect 18765 -14141 24043 -11411
tri 24043 -14141 27184 -11000 nw
tri -22895 -15487 -22117 -14141 ne
rect -22117 -15487 -16853 -14141
tri -16853 -15487 -15507 -14141 sw
tri 15507 -15487 16853 -14141 se
rect 16853 -15487 21331 -14141
tri -22117 -16853 -20971 -15487 ne
rect -20971 -16853 -15507 -15487
tri -15507 -16853 -14141 -15487 sw
tri 14141 -16853 15507 -15487 se
rect 15507 -16853 21331 -15487
tri 21331 -16853 24043 -14141 nw
tri -20971 -19053 -19125 -16853 ne
rect -19125 -19053 -14141 -16853
tri -14141 -19053 -11000 -16853 sw
tri 11000 -19053 14141 -16853 se
rect 14141 -19053 19131 -16853
tri 19131 -19053 21331 -16853 nw
tri -19125 -19092 -19092 -19053 ne
rect -19092 -19092 -11000 -19053
tri -11000 -19092 -10916 -19053 sw
tri 10916 -19092 11000 -19053 se
rect 11000 -19092 19092 -19053
tri 19092 -19092 19131 -19053 nw
tri -19092 -20673 -17208 -19092 ne
rect -17208 -20673 -10916 -19092
tri -10916 -20673 -7524 -19092 sw
tri 7524 -20673 10916 -19092 se
rect 10916 -20673 17208 -19092
tri 17208 -20673 19092 -19092 nw
tri -17208 -21666 -16025 -20673 ne
rect -16025 -21666 -7524 -20673
tri -7524 -21666 -3820 -20673 sw
tri 3820 -21666 7524 -20673 se
rect 7524 -21666 16024 -20673
tri 16024 -21666 17208 -20673 nw
tri -16025 -22000 -15627 -21666 ne
rect -15627 -22000 -3820 -21666
tri -3820 -22000 0 -21666 sw
tri 0 -22000 3820 -21666 se
rect 3820 -22000 15626 -21666
tri 15626 -22000 16024 -21666 nw
tri -15627 -22117 -15487 -22000 ne
rect -15487 -22117 15487 -22000
tri 15487 -22117 15626 -22000 nw
tri -15487 -24470 -11411 -22117 ne
rect -11411 -24470 11411 -22117
tri 11411 -24470 15487 -22117 nw
tri -11411 -26080 -6988 -24470 ne
rect -6988 -26080 6988 -24470
tri 6988 -26080 11411 -24470 nw
tri -6988 -26897 -2353 -26080 ne
rect -2353 -26897 2353 -26080
tri 2353 -26897 6988 -26080 nw
<< pi2 >>
tri -3820 21666 0 22000 se
tri 0 21666 3820 22000 sw
tri -7524 20673 -3820 21666 se
rect -3820 20673 3820 21666
tri 3820 20673 7524 21666 sw
tri -10916 19092 -7524 20673 se
rect -7524 19092 7524 20673
tri 7524 19092 10916 20673 sw
tri -11000 19053 -10916 19092 se
rect -10916 19053 10916 19092
tri 10916 19053 11000 19092 sw
tri -14141 16853 -11000 19053 se
rect -11000 16853 11000 19053
tri 11000 16853 14141 19053 sw
tri -15507 15487 -14141 16853 se
rect -14141 15487 14141 16853
tri 14141 15487 15507 16853 sw
tri -16853 14141 -15507 15487 se
rect -15507 14141 15507 15487
tri 15507 14141 16853 15487 sw
tri -18765 11411 -16853 14141 se
rect -16853 11411 16853 14141
tri 16853 11411 18765 14141 sw
tri -19053 11000 -18765 11411 se
rect -18765 11000 18765 11411
tri 18765 11000 19053 11411 sw
tri -20673 7524 -19053 11000 se
rect -19053 10916 19053 11000
tri 19053 10916 19092 11000 sw
rect -19053 7524 19092 10916
tri 19092 7524 20673 10916 sw
tri -20817 6988 -20673 7524 se
rect -20673 6988 20673 7524
tri -21666 3820 -20817 6988 se
rect -20817 3820 20673 6988
tri 20673 3820 21666 7524 sw
tri -21794 2353 -21666 3820 se
rect -21666 2353 21666 3820
tri -22000 0 -21794 2353 se
tri -22000 -2353 -21794 0 ne
rect -21794 -2353 21666 2353
tri 21666 0 22000 3820 sw
tri -21794 -3820 -21666 -2353 ne
rect -21666 -3820 21666 -2353
tri 21666 -3820 22000 0 nw
tri -21666 -6988 -20817 -3820 ne
rect -20817 -6988 20673 -3820
tri -20817 -7524 -20673 -6988 ne
rect -20673 -7524 20673 -6988
tri 20673 -7524 21666 -3820 nw
tri -20673 -11000 -19053 -7524 ne
rect -19053 -10916 19092 -7524
tri 19092 -10916 20673 -7524 nw
rect -19053 -11000 19053 -10916
tri 19053 -11000 19092 -10916 nw
tri -19053 -11411 -18765 -11000 ne
rect -18765 -11411 18765 -11000
tri 18765 -11411 19053 -11000 nw
tri -18765 -14141 -16853 -11411 ne
rect -16853 -14141 16853 -11411
tri 16853 -14141 18765 -11411 nw
tri -16853 -15487 -15507 -14141 ne
rect -15507 -15487 15507 -14141
tri 15507 -15487 16853 -14141 nw
tri -15507 -16853 -14141 -15487 ne
rect -14141 -16853 14141 -15487
tri 14141 -16853 15507 -15487 nw
tri -14141 -19053 -11000 -16853 ne
rect -11000 -19053 11000 -16853
tri 11000 -19053 14141 -16853 nw
tri -11000 -19092 -10916 -19053 ne
rect -10916 -19092 10916 -19053
tri 10916 -19092 11000 -19053 nw
tri -10916 -20673 -7524 -19092 ne
rect -7524 -20673 7524 -19092
tri 7524 -20673 10916 -19092 nw
tri -7524 -21666 -3820 -20673 ne
rect -3820 -21666 3820 -20673
tri 3820 -21666 7524 -20673 nw
tri -3820 -22000 0 -21666 ne
tri 0 -22000 3820 -21666 nw
<< ubm >>
tri -4341 24620 0 25000 se
tri 0 24620 4341 25000 sw
tri -8551 23492 -4341 24620 se
rect -4341 23492 4341 24620
tri 4341 23492 8551 24620 sw
tri -12500 21651 -8551 23492 se
rect -8551 22000 8551 23492
rect -8551 21666 -3820 22000
tri -3820 21666 0 22000 nw
tri 0 21666 3820 22000 ne
rect 3820 21666 8551 22000
rect -8551 21651 -3876 21666
tri -3876 21651 -3820 21666 nw
tri 3820 21651 3875 21666 ne
rect 3875 21651 8551 21666
tri 8551 21651 12500 23492 sw
tri -16070 19151 -12500 21651 se
rect -12500 20673 -7524 21651
tri -7524 20673 -3876 21651 nw
tri 3875 20673 7524 21651 ne
rect 7524 20673 12500 21651
rect -12500 19151 -10790 20673
tri -10790 19151 -7524 20673 nw
tri 7524 19151 10789 20673 ne
rect 10789 19151 12500 20673
tri 12500 19151 16070 21651 sw
tri -18368 16853 -16070 19151 se
rect -16070 19053 -11000 19151
tri -11000 19053 -10790 19151 nw
tri 10789 19053 11000 19151 ne
rect 11000 19053 16070 19151
rect -16070 16853 -14141 19053
tri -14141 16853 -11000 19053 nw
tri 11000 16853 14141 19053 ne
rect 14141 16853 16070 19053
tri 16070 16853 18368 19151 sw
tri -19151 16070 -18368 16853 se
rect -18368 16070 -14924 16853
tri -14924 16070 -14141 16853 nw
tri 14141 16070 14924 16853 ne
rect 14924 16070 18368 16853
tri 18368 16070 19151 16853 sw
tri -21651 12500 -19151 16070 se
rect -19151 14141 -16853 16070
tri -16853 14141 -14924 16070 nw
tri 14924 14141 16853 16070 ne
rect 16853 14141 19151 16070
rect -19151 12500 -18002 14141
tri -18002 12501 -16853 14141 nw
tri 16853 12500 18002 14141 ne
rect 18002 12500 19151 14141
tri 19151 12500 21651 16070 sw
tri -23492 8551 -21651 12500 se
rect -21651 11000 -19053 12500
tri -19053 11000 -18002 12500 nw
tri 18002 11000 19053 12500 ne
rect 19053 11000 21651 12500
rect -21651 8551 -20194 11000
tri -20194 8552 -19053 11000 nw
tri 19053 8551 20194 11000 ne
rect 20194 8551 21651 11000
tri 21651 8551 23492 12500 sw
tri -24620 4341 -23492 8551 se
rect -23492 7524 -20673 8551
tri -20673 7524 -20194 8551 nw
tri 20194 7524 20673 8551 ne
rect 20673 7524 23492 8551
rect -23492 4341 -21526 7524
tri -21526 4342 -20673 7524 nw
tri 20673 4342 21526 7524 ne
tri -25000 0 -24620 4341 se
rect -24620 3820 -21666 4341
tri -21666 3820 -21526 4341 nw
rect 21526 4341 23492 7524
tri 23492 4341 24620 8551 sw
tri 21526 3820 21666 4341 ne
rect 21666 3820 24620 4341
tri -25000 -4341 -24620 0 ne
rect -24620 -3820 -22000 3820
tri -22000 0 -21666 3820 nw
tri -22000 -3820 -21666 0 sw
tri 21666 0 22000 3820 ne
tri 21666 -3820 22000 0 se
rect 22000 -3820 24620 3820
tri 24620 0 25000 4341 sw
rect -24620 -4339 -21666 -3820
tri -21666 -4339 -21527 -3820 sw
rect -24620 -4341 -21527 -4339
tri 21526 -4341 21666 -3820 se
rect 21666 -4341 24620 -3820
tri 24620 -4341 25000 0 nw
tri -24620 -8551 -23492 -4341 ne
rect -23492 -7524 -21527 -4341
tri -21527 -7524 -20673 -4341 sw
tri 20673 -7524 21526 -4342 se
rect 21526 -7524 23492 -4341
rect -23492 -8550 -20673 -7524
tri -20673 -8550 -20195 -7524 sw
rect -23492 -8551 -20195 -8550
tri 20194 -8551 20673 -7524 se
rect 20673 -8551 23492 -7524
tri 23492 -8551 24620 -4341 nw
tri -23492 -12500 -21651 -8551 ne
rect -21651 -11000 -20195 -8551
tri -20195 -11000 -19053 -8551 sw
tri 19053 -11000 20194 -8552 se
rect 20194 -11000 21651 -8551
rect -21651 -12500 -19053 -11000
tri -19053 -12500 -18003 -11000 sw
tri 18002 -12500 19053 -11000 se
rect 19053 -12500 21651 -11000
tri 21651 -12500 23492 -8551 nw
tri -21651 -16070 -19151 -12500 ne
rect -19151 -14141 -18003 -12500
tri -18003 -14141 -16853 -12500 sw
tri 16853 -14141 18002 -12501 se
rect 18002 -14141 19151 -12500
rect -19151 -16070 -16853 -14141
tri -16853 -16070 -14924 -14141 sw
tri 14924 -16070 16853 -14141 se
rect 16853 -16070 19151 -14141
tri 19151 -16070 21651 -12500 nw
tri -19151 -16853 -18368 -16070 ne
rect -18368 -16853 -14924 -16070
tri -14924 -16853 -14141 -16070 sw
tri 14141 -16853 14924 -16070 se
rect 14924 -16853 18368 -16070
tri 18368 -16853 19151 -16070 nw
tri -18368 -19151 -16070 -16853 ne
rect -16070 -19053 -14141 -16853
tri -14141 -19053 -11000 -16853 sw
tri 11000 -19053 14141 -16853 se
rect 14141 -19053 16070 -16853
rect -16070 -19151 -11000 -19053
tri -11000 -19151 -10790 -19053 sw
tri 10790 -19151 11000 -19053 se
rect 11000 -19151 16070 -19053
tri 16070 -19151 18368 -16853 nw
tri -16070 -21651 -12500 -19151 ne
rect -12500 -20673 -10790 -19151
tri -10790 -20673 -7524 -19151 sw
tri 7524 -20673 10790 -19151 se
rect 10790 -20673 12500 -19151
rect -12500 -21651 -7524 -20673
tri -7524 -21651 -3876 -20673 sw
tri 3876 -21651 7524 -20673 se
rect 7524 -21651 12500 -20673
tri 12500 -21651 16070 -19151 nw
tri -12500 -23492 -8551 -21651 ne
rect -8551 -21666 -3876 -21651
tri -3876 -21666 -3820 -21651 sw
tri 3820 -21666 3876 -21651 se
rect 3876 -21666 8551 -21651
rect -8551 -22000 -3820 -21666
tri -3820 -22000 0 -21666 sw
tri 0 -22000 3820 -21666 se
rect 3820 -22000 8551 -21666
rect -8551 -23492 8551 -22000
tri 8551 -23492 12500 -21651 nw
tri -8551 -24620 -4341 -23492 ne
rect -4341 -24620 4341 -23492
tri 4341 -24620 8551 -23492 nw
tri -4341 -25000 0 -24620 ne
tri 0 -25000 4341 -24620 nw
<< properties >>
string FIXED_BBOX -27000 -27000 27000 27000
<< end >>
