* NGSPICE file created from mprj2_logic_high.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_1_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_213 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_1
XFILLER_1_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_0 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_4 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_5 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_6 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_7 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_8 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_10 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_11 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_212 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__fill_2
Xinst vssd2 vssd2 vccd2 vccd2 HI inst/LO sky130_fd_sc_hd__conb_1
XFILLER_0_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_14 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_15 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_16 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XPHY_17 vssd2 vccd2 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
.ends

