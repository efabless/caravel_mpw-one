magic
tech sky130A
magscale 1 2
timestamp 1622561372
<< viali >>
rect 4353 4437 4387 4471
rect 2145 4233 2179 4267
rect 3801 4233 3835 4267
rect 5549 4233 5583 4267
rect 2053 4165 2087 4199
rect 4169 4165 4203 4199
rect 4629 4029 4663 4063
rect 4905 4029 4939 4063
rect 1685 3553 1719 3587
rect 2145 3553 2179 3587
rect 2697 3553 2731 3587
rect 5365 3553 5399 3587
rect 1593 3485 1627 3519
rect 4077 3485 4111 3519
rect 2421 3417 2455 3451
rect 4537 3349 4571 3383
rect 4813 3349 4847 3383
rect 3341 3145 3375 3179
rect 4721 3009 4755 3043
rect 3985 2941 4019 2975
rect 1685 2465 1719 2499
rect 5549 2465 5583 2499
rect 1593 2397 1627 2431
rect 1685 2057 1719 2091
rect 2973 2057 3007 2091
rect 1961 1853 1995 1887
rect 2145 1309 2179 1343
rect 2789 1309 2823 1343
rect 4905 1309 4939 1343
rect 2237 1241 2271 1275
rect 2881 1173 2915 1207
rect 5365 1173 5399 1207
<< metal1 >>
rect 1104 5466 5888 5488
rect 1104 5414 1780 5466
rect 1832 5414 1844 5466
rect 1896 5414 1908 5466
rect 1960 5414 1972 5466
rect 2024 5414 3378 5466
rect 3430 5414 3442 5466
rect 3494 5414 3506 5466
rect 3558 5414 3570 5466
rect 3622 5414 4975 5466
rect 5027 5414 5039 5466
rect 5091 5414 5103 5466
rect 5155 5414 5167 5466
rect 5219 5414 5888 5466
rect 1104 5392 5888 5414
rect 1104 4922 5888 4944
rect 1104 4870 2579 4922
rect 2631 4870 2643 4922
rect 2695 4870 2707 4922
rect 2759 4870 2771 4922
rect 2823 4870 4176 4922
rect 4228 4870 4240 4922
rect 4292 4870 4304 4922
rect 4356 4870 4368 4922
rect 4420 4870 5888 4922
rect 1104 4848 5888 4870
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 5350 4536 5356 4548
rect 4120 4508 5356 4536
rect 4120 4496 4126 4508
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4614 4468 4620 4480
rect 4387 4440 4620 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 1104 4378 5888 4400
rect 1104 4326 1780 4378
rect 1832 4326 1844 4378
rect 1896 4326 1908 4378
rect 1960 4326 1972 4378
rect 2024 4326 3378 4378
rect 3430 4326 3442 4378
rect 3494 4326 3506 4378
rect 3558 4326 3570 4378
rect 3622 4326 4975 4378
rect 5027 4326 5039 4378
rect 5091 4326 5103 4378
rect 5155 4326 5167 4378
rect 5219 4326 5888 4378
rect 1104 4304 5888 4326
rect 934 4224 940 4276
rect 992 4264 998 4276
rect 2133 4267 2191 4273
rect 2133 4264 2145 4267
rect 992 4236 2145 4264
rect 992 4224 998 4236
rect 2133 4233 2145 4236
rect 2179 4233 2191 4267
rect 2133 4227 2191 4233
rect 3789 4267 3847 4273
rect 3789 4233 3801 4267
rect 3835 4264 3847 4267
rect 5534 4264 5540 4276
rect 3835 4236 4936 4264
rect 5495 4236 5540 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 2041 4199 2099 4205
rect 2041 4165 2053 4199
rect 2087 4196 2099 4199
rect 2406 4196 2412 4208
rect 2087 4168 2412 4196
rect 2087 4165 2099 4168
rect 2041 4159 2099 4165
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 4157 4199 4215 4205
rect 4157 4196 4169 4199
rect 2832 4168 4169 4196
rect 2832 4156 2838 4168
rect 4157 4165 4169 4168
rect 4203 4165 4215 4199
rect 4908 4196 4936 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5994 4196 6000 4208
rect 4908 4168 6000 4196
rect 4157 4159 4215 4165
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 4617 4063 4675 4069
rect 4617 4060 4629 4063
rect 992 4032 4629 4060
rect 992 4020 998 4032
rect 4617 4029 4629 4032
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5258 4060 5264 4072
rect 4939 4032 5264 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 6454 3924 6460 3936
rect 2280 3896 6460 3924
rect 2280 3884 2286 3896
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 1104 3834 5888 3856
rect 1104 3782 2579 3834
rect 2631 3782 2643 3834
rect 2695 3782 2707 3834
rect 2759 3782 2771 3834
rect 2823 3782 4176 3834
rect 4228 3782 4240 3834
rect 4292 3782 4304 3834
rect 4356 3782 4368 3834
rect 4420 3782 5888 3834
rect 1104 3760 5888 3782
rect 5994 3720 6000 3732
rect 2700 3692 6000 3720
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1452 3556 1685 3584
rect 1452 3544 1458 3556
rect 1673 3553 1685 3556
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 2222 3584 2228 3596
rect 2179 3556 2228 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2700 3593 2728 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 4706 3652 4712 3664
rect 2884 3624 4712 3652
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3553 2743 3587
rect 2685 3547 2743 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2884 3516 2912 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 3016 3556 5365 3584
rect 3016 3544 3022 3556
rect 5353 3553 5365 3556
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 1627 3488 2912 3516
rect 4065 3519 4123 3525
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4798 3516 4804 3528
rect 4111 3488 4804 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 2409 3451 2467 3457
rect 2409 3417 2421 3451
rect 2455 3448 2467 3451
rect 4154 3448 4160 3460
rect 2455 3420 4160 3448
rect 2455 3417 2467 3420
rect 2409 3411 2467 3417
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4890 3448 4896 3460
rect 4816 3420 4896 3448
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4706 3380 4712 3392
rect 4571 3352 4712 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 4816 3389 4844 3420
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 1104 3290 5888 3312
rect 1104 3238 1780 3290
rect 1832 3238 1844 3290
rect 1896 3238 1908 3290
rect 1960 3238 1972 3290
rect 2024 3238 3378 3290
rect 3430 3238 3442 3290
rect 3494 3238 3506 3290
rect 3558 3238 3570 3290
rect 3622 3238 4975 3290
rect 5027 3238 5039 3290
rect 5091 3238 5103 3290
rect 5155 3238 5167 3290
rect 5219 3238 5888 3290
rect 1104 3216 5888 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 3329 3179 3387 3185
rect 3329 3176 3341 3179
rect 2188 3148 3341 3176
rect 2188 3136 2194 3148
rect 3329 3145 3341 3148
rect 3375 3145 3387 3179
rect 3329 3139 3387 3145
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 4709 3043 4767 3049
rect 4709 3040 4721 3043
rect 3752 3012 4721 3040
rect 3752 3000 3758 3012
rect 4709 3009 4721 3012
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 1394 2932 1400 2984
rect 1452 2972 1458 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 1452 2944 3985 2972
rect 1452 2932 1458 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 1104 2746 5888 2768
rect 1104 2694 2579 2746
rect 2631 2694 2643 2746
rect 2695 2694 2707 2746
rect 2759 2694 2771 2746
rect 2823 2694 4176 2746
rect 4228 2694 4240 2746
rect 4292 2694 4304 2746
rect 4356 2694 4368 2746
rect 4420 2694 5888 2746
rect 1104 2672 5888 2694
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 5626 2428 5632 2440
rect 1627 2400 5632 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 1104 2202 5888 2224
rect 1104 2150 1780 2202
rect 1832 2150 1844 2202
rect 1896 2150 1908 2202
rect 1960 2150 1972 2202
rect 2024 2150 3378 2202
rect 3430 2150 3442 2202
rect 3494 2150 3506 2202
rect 3558 2150 3570 2202
rect 3622 2150 4975 2202
rect 5027 2150 5039 2202
rect 5091 2150 5103 2202
rect 5155 2150 5167 2202
rect 5219 2150 5888 2202
rect 1104 2128 5888 2150
rect 1673 2091 1731 2097
rect 1673 2057 1685 2091
rect 1719 2088 1731 2091
rect 2314 2088 2320 2100
rect 1719 2060 2320 2088
rect 1719 2057 1731 2060
rect 1673 2051 1731 2057
rect 2314 2048 2320 2060
rect 2372 2048 2378 2100
rect 2961 2091 3019 2097
rect 2961 2057 2973 2091
rect 3007 2088 3019 2091
rect 4522 2088 4528 2100
rect 3007 2060 4528 2088
rect 3007 2057 3019 2060
rect 2961 2051 3019 2057
rect 4522 2048 4528 2060
rect 4580 2048 4586 2100
rect 2774 1980 2780 2032
rect 2832 2020 2838 2032
rect 5258 2020 5264 2032
rect 2832 1992 5264 2020
rect 2832 1980 2838 1992
rect 5258 1980 5264 1992
rect 5316 1980 5322 2032
rect 1946 1884 1952 1896
rect 1907 1856 1952 1884
rect 1946 1844 1952 1856
rect 2004 1844 2010 1896
rect 1104 1658 5888 1680
rect 1104 1606 2579 1658
rect 2631 1606 2643 1658
rect 2695 1606 2707 1658
rect 2759 1606 2771 1658
rect 2823 1606 4176 1658
rect 4228 1606 4240 1658
rect 4292 1606 4304 1658
rect 4356 1606 4368 1658
rect 4420 1606 5888 1658
rect 1104 1584 5888 1606
rect 2133 1343 2191 1349
rect 2133 1309 2145 1343
rect 2179 1340 2191 1343
rect 2777 1343 2835 1349
rect 2179 1312 2728 1340
rect 2179 1309 2191 1312
rect 2133 1303 2191 1309
rect 474 1232 480 1284
rect 532 1272 538 1284
rect 2225 1275 2283 1281
rect 2225 1272 2237 1275
rect 532 1244 2237 1272
rect 532 1232 538 1244
rect 2225 1241 2237 1244
rect 2271 1241 2283 1275
rect 2700 1272 2728 1312
rect 2777 1309 2789 1343
rect 2823 1340 2835 1343
rect 2866 1340 2872 1352
rect 2823 1312 2872 1340
rect 2823 1309 2835 1312
rect 2777 1303 2835 1309
rect 2866 1300 2872 1312
rect 2924 1300 2930 1352
rect 4893 1343 4951 1349
rect 4893 1309 4905 1343
rect 4939 1340 4951 1343
rect 5350 1340 5356 1352
rect 4939 1312 5356 1340
rect 4939 1309 4951 1312
rect 4893 1303 4951 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 3234 1272 3240 1284
rect 2700 1244 3240 1272
rect 2225 1235 2283 1241
rect 3234 1232 3240 1244
rect 3292 1232 3298 1284
rect 2314 1164 2320 1216
rect 2372 1204 2378 1216
rect 2869 1207 2927 1213
rect 2869 1204 2881 1207
rect 2372 1176 2881 1204
rect 2372 1164 2378 1176
rect 2869 1173 2881 1176
rect 2915 1173 2927 1207
rect 2869 1167 2927 1173
rect 5353 1207 5411 1213
rect 5353 1173 5365 1207
rect 5399 1204 5411 1207
rect 5534 1204 5540 1216
rect 5399 1176 5540 1204
rect 5399 1173 5411 1176
rect 5353 1167 5411 1173
rect 5534 1164 5540 1176
rect 5592 1164 5598 1216
rect 1104 1114 5888 1136
rect 1104 1062 1780 1114
rect 1832 1062 1844 1114
rect 1896 1062 1908 1114
rect 1960 1062 1972 1114
rect 2024 1062 3378 1114
rect 3430 1062 3442 1114
rect 3494 1062 3506 1114
rect 3558 1062 3570 1114
rect 3622 1062 4975 1114
rect 5027 1062 5039 1114
rect 5091 1062 5103 1114
rect 5155 1062 5167 1114
rect 5219 1062 5888 1114
rect 1104 1040 5888 1062
<< via1 >>
rect 1780 5414 1832 5466
rect 1844 5414 1896 5466
rect 1908 5414 1960 5466
rect 1972 5414 2024 5466
rect 3378 5414 3430 5466
rect 3442 5414 3494 5466
rect 3506 5414 3558 5466
rect 3570 5414 3622 5466
rect 4975 5414 5027 5466
rect 5039 5414 5091 5466
rect 5103 5414 5155 5466
rect 5167 5414 5219 5466
rect 2579 4870 2631 4922
rect 2643 4870 2695 4922
rect 2707 4870 2759 4922
rect 2771 4870 2823 4922
rect 4176 4870 4228 4922
rect 4240 4870 4292 4922
rect 4304 4870 4356 4922
rect 4368 4870 4420 4922
rect 4068 4496 4120 4548
rect 5356 4496 5408 4548
rect 4620 4428 4672 4480
rect 1780 4326 1832 4378
rect 1844 4326 1896 4378
rect 1908 4326 1960 4378
rect 1972 4326 2024 4378
rect 3378 4326 3430 4378
rect 3442 4326 3494 4378
rect 3506 4326 3558 4378
rect 3570 4326 3622 4378
rect 4975 4326 5027 4378
rect 5039 4326 5091 4378
rect 5103 4326 5155 4378
rect 5167 4326 5219 4378
rect 940 4224 992 4276
rect 5540 4267 5592 4276
rect 2412 4156 2464 4208
rect 2780 4156 2832 4208
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 6000 4156 6052 4208
rect 940 4020 992 4072
rect 5264 4020 5316 4072
rect 2228 3884 2280 3936
rect 6460 3884 6512 3936
rect 2579 3782 2631 3834
rect 2643 3782 2695 3834
rect 2707 3782 2759 3834
rect 2771 3782 2823 3834
rect 4176 3782 4228 3834
rect 4240 3782 4292 3834
rect 4304 3782 4356 3834
rect 4368 3782 4420 3834
rect 1400 3544 1452 3596
rect 2228 3544 2280 3596
rect 6000 3680 6052 3732
rect 4712 3612 4764 3664
rect 2964 3544 3016 3596
rect 4804 3476 4856 3528
rect 4160 3408 4212 3460
rect 4712 3340 4764 3392
rect 4896 3408 4948 3460
rect 1780 3238 1832 3290
rect 1844 3238 1896 3290
rect 1908 3238 1960 3290
rect 1972 3238 2024 3290
rect 3378 3238 3430 3290
rect 3442 3238 3494 3290
rect 3506 3238 3558 3290
rect 3570 3238 3622 3290
rect 4975 3238 5027 3290
rect 5039 3238 5091 3290
rect 5103 3238 5155 3290
rect 5167 3238 5219 3290
rect 2136 3136 2188 3188
rect 3700 3000 3752 3052
rect 1400 2932 1452 2984
rect 2579 2694 2631 2746
rect 2643 2694 2695 2746
rect 2707 2694 2759 2746
rect 2771 2694 2823 2746
rect 4176 2694 4228 2746
rect 4240 2694 4292 2746
rect 4304 2694 4356 2746
rect 4368 2694 4420 2746
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 5632 2388 5684 2440
rect 1780 2150 1832 2202
rect 1844 2150 1896 2202
rect 1908 2150 1960 2202
rect 1972 2150 2024 2202
rect 3378 2150 3430 2202
rect 3442 2150 3494 2202
rect 3506 2150 3558 2202
rect 3570 2150 3622 2202
rect 4975 2150 5027 2202
rect 5039 2150 5091 2202
rect 5103 2150 5155 2202
rect 5167 2150 5219 2202
rect 2320 2048 2372 2100
rect 4528 2048 4580 2100
rect 2780 1980 2832 2032
rect 5264 1980 5316 2032
rect 1952 1887 2004 1896
rect 1952 1853 1961 1887
rect 1961 1853 1995 1887
rect 1995 1853 2004 1887
rect 1952 1844 2004 1853
rect 2579 1606 2631 1658
rect 2643 1606 2695 1658
rect 2707 1606 2759 1658
rect 2771 1606 2823 1658
rect 4176 1606 4228 1658
rect 4240 1606 4292 1658
rect 4304 1606 4356 1658
rect 4368 1606 4420 1658
rect 480 1232 532 1284
rect 2872 1300 2924 1352
rect 5356 1300 5408 1352
rect 3240 1232 3292 1284
rect 2320 1164 2372 1216
rect 5540 1164 5592 1216
rect 1780 1062 1832 1114
rect 1844 1062 1896 1114
rect 1908 1062 1960 1114
rect 1972 1062 2024 1114
rect 3378 1062 3430 1114
rect 3442 1062 3494 1114
rect 3506 1062 3558 1114
rect 3570 1062 3622 1114
rect 4975 1062 5027 1114
rect 5039 1062 5091 1114
rect 5103 1062 5155 1114
rect 5167 1062 5219 1114
<< metal2 >>
rect 938 6200 994 7000
rect 1398 6200 1454 7000
rect 1858 6200 1914 7000
rect 2778 6200 2834 7000
rect 3238 6200 3294 7000
rect 4158 6200 4214 7000
rect 4618 6200 4674 7000
rect 4802 6216 4858 6225
rect 952 4282 980 6200
rect 940 4276 992 4282
rect 940 4218 992 4224
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 480 1284 532 1290
rect 480 1226 532 1232
rect 492 800 520 1226
rect 952 800 980 4014
rect 1412 3602 1440 6200
rect 1872 5658 1900 6200
rect 1872 5630 2176 5658
rect 1754 5468 2050 5488
rect 1810 5466 1834 5468
rect 1890 5466 1914 5468
rect 1970 5466 1994 5468
rect 1832 5414 1834 5466
rect 1896 5414 1908 5466
rect 1970 5414 1972 5466
rect 1810 5412 1834 5414
rect 1890 5412 1914 5414
rect 1970 5412 1994 5414
rect 1754 5392 2050 5412
rect 1754 4380 2050 4400
rect 1810 4378 1834 4380
rect 1890 4378 1914 4380
rect 1970 4378 1994 4380
rect 1832 4326 1834 4378
rect 1896 4326 1908 4378
rect 1970 4326 1972 4378
rect 1810 4324 1834 4326
rect 1890 4324 1914 4326
rect 1970 4324 1994 4326
rect 1754 4304 2050 4324
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 800 1440 2926
rect 1688 2514 1716 3431
rect 1754 3292 2050 3312
rect 1810 3290 1834 3292
rect 1890 3290 1914 3292
rect 1970 3290 1994 3292
rect 1832 3238 1834 3290
rect 1896 3238 1908 3290
rect 1970 3238 1972 3290
rect 1810 3236 1834 3238
rect 1890 3236 1914 3238
rect 1970 3236 1994 3238
rect 1754 3216 2050 3236
rect 2148 3194 2176 5630
rect 2318 5264 2374 5273
rect 2318 5199 2374 5208
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3602 2268 3878
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1754 2204 2050 2224
rect 1810 2202 1834 2204
rect 1890 2202 1914 2204
rect 1970 2202 1994 2204
rect 1832 2150 1834 2202
rect 1896 2150 1908 2202
rect 1970 2150 1972 2202
rect 1810 2148 1834 2150
rect 1890 2148 1914 2150
rect 1970 2148 1994 2150
rect 1754 2128 2050 2148
rect 2332 2106 2360 5199
rect 2792 5114 2820 6200
rect 2792 5086 2912 5114
rect 2553 4924 2849 4944
rect 2609 4922 2633 4924
rect 2689 4922 2713 4924
rect 2769 4922 2793 4924
rect 2631 4870 2633 4922
rect 2695 4870 2707 4922
rect 2769 4870 2771 4922
rect 2609 4868 2633 4870
rect 2689 4868 2713 4870
rect 2769 4868 2793 4870
rect 2553 4848 2849 4868
rect 2412 4208 2464 4214
rect 2780 4208 2832 4214
rect 2412 4150 2464 4156
rect 2778 4176 2780 4185
rect 2832 4176 2834 4185
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 1964 1465 1992 1838
rect 2424 1465 2452 4150
rect 2778 4111 2834 4120
rect 2553 3836 2849 3856
rect 2609 3834 2633 3836
rect 2689 3834 2713 3836
rect 2769 3834 2793 3836
rect 2631 3782 2633 3834
rect 2695 3782 2707 3834
rect 2769 3782 2771 3834
rect 2609 3780 2633 3782
rect 2689 3780 2713 3782
rect 2769 3780 2793 3782
rect 2553 3760 2849 3780
rect 2553 2748 2849 2768
rect 2609 2746 2633 2748
rect 2689 2746 2713 2748
rect 2769 2746 2793 2748
rect 2631 2694 2633 2746
rect 2695 2694 2707 2746
rect 2769 2694 2771 2746
rect 2609 2692 2633 2694
rect 2689 2692 2713 2694
rect 2769 2692 2793 2694
rect 2553 2672 2849 2692
rect 2780 2032 2832 2038
rect 2778 2000 2780 2009
rect 2832 2000 2834 2009
rect 2778 1935 2834 1944
rect 2553 1660 2849 1680
rect 2609 1658 2633 1660
rect 2689 1658 2713 1660
rect 2769 1658 2793 1660
rect 2631 1606 2633 1658
rect 2695 1606 2707 1658
rect 2769 1606 2771 1658
rect 2609 1604 2633 1606
rect 2689 1604 2713 1606
rect 2769 1604 2793 1606
rect 2553 1584 2849 1604
rect 1950 1456 2006 1465
rect 1950 1391 2006 1400
rect 2410 1456 2466 1465
rect 2410 1391 2466 1400
rect 2884 1358 2912 5086
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 2320 1216 2372 1222
rect 2976 1170 3004 3538
rect 3252 1290 3280 6200
rect 3352 5468 3648 5488
rect 3408 5466 3432 5468
rect 3488 5466 3512 5468
rect 3568 5466 3592 5468
rect 3430 5414 3432 5466
rect 3494 5414 3506 5466
rect 3568 5414 3570 5466
rect 3408 5412 3432 5414
rect 3488 5412 3512 5414
rect 3568 5412 3592 5414
rect 3352 5392 3648 5412
rect 4066 5128 4122 5137
rect 4172 5114 4200 6200
rect 4172 5086 4568 5114
rect 4066 5063 4122 5072
rect 4080 4554 4108 5063
rect 4150 4924 4446 4944
rect 4206 4922 4230 4924
rect 4286 4922 4310 4924
rect 4366 4922 4390 4924
rect 4228 4870 4230 4922
rect 4292 4870 4304 4922
rect 4366 4870 4368 4922
rect 4206 4868 4230 4870
rect 4286 4868 4310 4870
rect 4366 4868 4390 4870
rect 4150 4848 4446 4868
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3352 4380 3648 4400
rect 3408 4378 3432 4380
rect 3488 4378 3512 4380
rect 3568 4378 3592 4380
rect 3430 4326 3432 4378
rect 3494 4326 3506 4378
rect 3568 4326 3570 4378
rect 3408 4324 3432 4326
rect 3488 4324 3512 4326
rect 3568 4324 3592 4326
rect 3352 4304 3648 4324
rect 4150 3836 4446 3856
rect 4206 3834 4230 3836
rect 4286 3834 4310 3836
rect 4366 3834 4390 3836
rect 4228 3782 4230 3834
rect 4292 3782 4304 3834
rect 4366 3782 4368 3834
rect 4206 3780 4230 3782
rect 4286 3780 4310 3782
rect 4366 3780 4390 3782
rect 4150 3760 4446 3780
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3352 3292 3648 3312
rect 3408 3290 3432 3292
rect 3488 3290 3512 3292
rect 3568 3290 3592 3292
rect 3430 3238 3432 3290
rect 3494 3238 3506 3290
rect 3568 3238 3570 3290
rect 3408 3236 3432 3238
rect 3488 3236 3512 3238
rect 3568 3236 3592 3238
rect 3352 3216 3648 3236
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3352 2204 3648 2224
rect 3408 2202 3432 2204
rect 3488 2202 3512 2204
rect 3568 2202 3592 2204
rect 3430 2150 3432 2202
rect 3494 2150 3506 2202
rect 3568 2150 3570 2202
rect 3408 2148 3432 2150
rect 3488 2148 3512 2150
rect 3568 2148 3592 2150
rect 3352 2128 3648 2148
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 2320 1158 2372 1164
rect 1754 1116 2050 1136
rect 1810 1114 1834 1116
rect 1890 1114 1914 1116
rect 1970 1114 1994 1116
rect 1832 1062 1834 1114
rect 1896 1062 1908 1114
rect 1970 1062 1972 1114
rect 1810 1060 1834 1062
rect 1890 1060 1914 1062
rect 1970 1060 1994 1062
rect 1754 1040 2050 1060
rect 2332 800 2360 1158
rect 2792 1142 3004 1170
rect 2792 800 2820 1142
rect 3352 1116 3648 1136
rect 3408 1114 3432 1116
rect 3488 1114 3512 1116
rect 3568 1114 3592 1116
rect 3430 1062 3432 1114
rect 3494 1062 3506 1114
rect 3568 1062 3570 1114
rect 3408 1060 3432 1062
rect 3488 1060 3512 1062
rect 3568 1060 3592 1062
rect 3352 1040 3648 1060
rect 3712 800 3740 2994
rect 4172 2938 4200 3402
rect 4080 2910 4200 2938
rect 4080 2530 4108 2910
rect 4150 2748 4446 2768
rect 4206 2746 4230 2748
rect 4286 2746 4310 2748
rect 4366 2746 4390 2748
rect 4228 2694 4230 2746
rect 4292 2694 4304 2746
rect 4366 2694 4368 2746
rect 4206 2692 4230 2694
rect 4286 2692 4310 2694
rect 4366 2692 4390 2694
rect 4150 2672 4446 2692
rect 4080 2502 4200 2530
rect 4172 1850 4200 2502
rect 4540 2106 4568 5086
rect 4632 4570 4660 6200
rect 5538 6200 5594 7000
rect 5998 6200 6054 7000
rect 6458 6200 6514 7000
rect 4802 6151 4858 6160
rect 4632 4542 4752 4570
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 2825 4660 4422
rect 4724 3670 4752 4542
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4816 3618 4844 6151
rect 4949 5468 5245 5488
rect 5005 5466 5029 5468
rect 5085 5466 5109 5468
rect 5165 5466 5189 5468
rect 5027 5414 5029 5466
rect 5091 5414 5103 5466
rect 5165 5414 5167 5466
rect 5005 5412 5029 5414
rect 5085 5412 5109 5414
rect 5165 5412 5189 5414
rect 4949 5392 5245 5412
rect 5552 4978 5580 6200
rect 5552 4950 5672 4978
rect 5538 4856 5594 4865
rect 5538 4791 5594 4800
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 4949 4380 5245 4400
rect 5005 4378 5029 4380
rect 5085 4378 5109 4380
rect 5165 4378 5189 4380
rect 5027 4326 5029 4378
rect 5091 4326 5103 4378
rect 5165 4326 5167 4378
rect 5005 4324 5029 4326
rect 5085 4324 5109 4326
rect 5165 4324 5189 4326
rect 4949 4304 5245 4324
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 4816 3590 4936 3618
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4080 1822 4200 1850
rect 4080 1442 4108 1822
rect 4150 1660 4446 1680
rect 4206 1658 4230 1660
rect 4286 1658 4310 1660
rect 4366 1658 4390 1660
rect 4228 1606 4230 1658
rect 4292 1606 4304 1658
rect 4366 1606 4368 1658
rect 4206 1604 4230 1606
rect 4286 1604 4310 1606
rect 4366 1604 4390 1606
rect 4150 1584 4446 1604
rect 4080 1414 4200 1442
rect 4172 800 4200 1414
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4724 785 4752 3334
rect 4816 898 4844 3470
rect 4908 3466 4936 3590
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4949 3292 5245 3312
rect 5005 3290 5029 3292
rect 5085 3290 5109 3292
rect 5165 3290 5189 3292
rect 5027 3238 5029 3290
rect 5091 3238 5103 3290
rect 5165 3238 5167 3290
rect 5005 3236 5029 3238
rect 5085 3236 5109 3238
rect 5165 3236 5189 3238
rect 4949 3216 5245 3236
rect 4949 2204 5245 2224
rect 5005 2202 5029 2204
rect 5085 2202 5109 2204
rect 5165 2202 5189 2204
rect 5027 2150 5029 2202
rect 5091 2150 5103 2202
rect 5165 2150 5167 2202
rect 5005 2148 5029 2150
rect 5085 2148 5109 2150
rect 5165 2148 5189 2150
rect 4949 2128 5245 2148
rect 5276 2038 5304 4014
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5368 1358 5396 4490
rect 5552 4282 5580 4791
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5552 2514 5580 3431
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5644 2446 5672 4950
rect 6012 4214 6040 6200
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6472 3942 6500 6200
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5540 1216 5592 1222
rect 5540 1158 5592 1164
rect 4949 1116 5245 1136
rect 5005 1114 5029 1116
rect 5085 1114 5109 1116
rect 5165 1114 5189 1116
rect 5027 1062 5029 1114
rect 5091 1062 5103 1114
rect 5165 1062 5167 1114
rect 5005 1060 5029 1062
rect 5085 1060 5109 1062
rect 5165 1060 5189 1062
rect 4949 1040 5245 1060
rect 4816 870 5120 898
rect 5092 800 5120 870
rect 5552 800 5580 1158
rect 6012 800 6040 3674
rect 4710 776 4766 785
rect 4710 711 4766 720
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
<< via2 >>
rect 1754 5466 1810 5468
rect 1834 5466 1890 5468
rect 1914 5466 1970 5468
rect 1994 5466 2050 5468
rect 1754 5414 1780 5466
rect 1780 5414 1810 5466
rect 1834 5414 1844 5466
rect 1844 5414 1890 5466
rect 1914 5414 1960 5466
rect 1960 5414 1970 5466
rect 1994 5414 2024 5466
rect 2024 5414 2050 5466
rect 1754 5412 1810 5414
rect 1834 5412 1890 5414
rect 1914 5412 1970 5414
rect 1994 5412 2050 5414
rect 1754 4378 1810 4380
rect 1834 4378 1890 4380
rect 1914 4378 1970 4380
rect 1994 4378 2050 4380
rect 1754 4326 1780 4378
rect 1780 4326 1810 4378
rect 1834 4326 1844 4378
rect 1844 4326 1890 4378
rect 1914 4326 1960 4378
rect 1960 4326 1970 4378
rect 1994 4326 2024 4378
rect 2024 4326 2050 4378
rect 1754 4324 1810 4326
rect 1834 4324 1890 4326
rect 1914 4324 1970 4326
rect 1994 4324 2050 4326
rect 1674 3440 1730 3496
rect 1754 3290 1810 3292
rect 1834 3290 1890 3292
rect 1914 3290 1970 3292
rect 1994 3290 2050 3292
rect 1754 3238 1780 3290
rect 1780 3238 1810 3290
rect 1834 3238 1844 3290
rect 1844 3238 1890 3290
rect 1914 3238 1960 3290
rect 1960 3238 1970 3290
rect 1994 3238 2024 3290
rect 2024 3238 2050 3290
rect 1754 3236 1810 3238
rect 1834 3236 1890 3238
rect 1914 3236 1970 3238
rect 1994 3236 2050 3238
rect 2318 5208 2374 5264
rect 1754 2202 1810 2204
rect 1834 2202 1890 2204
rect 1914 2202 1970 2204
rect 1994 2202 2050 2204
rect 1754 2150 1780 2202
rect 1780 2150 1810 2202
rect 1834 2150 1844 2202
rect 1844 2150 1890 2202
rect 1914 2150 1960 2202
rect 1960 2150 1970 2202
rect 1994 2150 2024 2202
rect 2024 2150 2050 2202
rect 1754 2148 1810 2150
rect 1834 2148 1890 2150
rect 1914 2148 1970 2150
rect 1994 2148 2050 2150
rect 2553 4922 2609 4924
rect 2633 4922 2689 4924
rect 2713 4922 2769 4924
rect 2793 4922 2849 4924
rect 2553 4870 2579 4922
rect 2579 4870 2609 4922
rect 2633 4870 2643 4922
rect 2643 4870 2689 4922
rect 2713 4870 2759 4922
rect 2759 4870 2769 4922
rect 2793 4870 2823 4922
rect 2823 4870 2849 4922
rect 2553 4868 2609 4870
rect 2633 4868 2689 4870
rect 2713 4868 2769 4870
rect 2793 4868 2849 4870
rect 2778 4156 2780 4176
rect 2780 4156 2832 4176
rect 2832 4156 2834 4176
rect 2778 4120 2834 4156
rect 2553 3834 2609 3836
rect 2633 3834 2689 3836
rect 2713 3834 2769 3836
rect 2793 3834 2849 3836
rect 2553 3782 2579 3834
rect 2579 3782 2609 3834
rect 2633 3782 2643 3834
rect 2643 3782 2689 3834
rect 2713 3782 2759 3834
rect 2759 3782 2769 3834
rect 2793 3782 2823 3834
rect 2823 3782 2849 3834
rect 2553 3780 2609 3782
rect 2633 3780 2689 3782
rect 2713 3780 2769 3782
rect 2793 3780 2849 3782
rect 2553 2746 2609 2748
rect 2633 2746 2689 2748
rect 2713 2746 2769 2748
rect 2793 2746 2849 2748
rect 2553 2694 2579 2746
rect 2579 2694 2609 2746
rect 2633 2694 2643 2746
rect 2643 2694 2689 2746
rect 2713 2694 2759 2746
rect 2759 2694 2769 2746
rect 2793 2694 2823 2746
rect 2823 2694 2849 2746
rect 2553 2692 2609 2694
rect 2633 2692 2689 2694
rect 2713 2692 2769 2694
rect 2793 2692 2849 2694
rect 2778 1980 2780 2000
rect 2780 1980 2832 2000
rect 2832 1980 2834 2000
rect 2778 1944 2834 1980
rect 2553 1658 2609 1660
rect 2633 1658 2689 1660
rect 2713 1658 2769 1660
rect 2793 1658 2849 1660
rect 2553 1606 2579 1658
rect 2579 1606 2609 1658
rect 2633 1606 2643 1658
rect 2643 1606 2689 1658
rect 2713 1606 2759 1658
rect 2759 1606 2769 1658
rect 2793 1606 2823 1658
rect 2823 1606 2849 1658
rect 2553 1604 2609 1606
rect 2633 1604 2689 1606
rect 2713 1604 2769 1606
rect 2793 1604 2849 1606
rect 1950 1400 2006 1456
rect 2410 1400 2466 1456
rect 3352 5466 3408 5468
rect 3432 5466 3488 5468
rect 3512 5466 3568 5468
rect 3592 5466 3648 5468
rect 3352 5414 3378 5466
rect 3378 5414 3408 5466
rect 3432 5414 3442 5466
rect 3442 5414 3488 5466
rect 3512 5414 3558 5466
rect 3558 5414 3568 5466
rect 3592 5414 3622 5466
rect 3622 5414 3648 5466
rect 3352 5412 3408 5414
rect 3432 5412 3488 5414
rect 3512 5412 3568 5414
rect 3592 5412 3648 5414
rect 4066 5072 4122 5128
rect 4150 4922 4206 4924
rect 4230 4922 4286 4924
rect 4310 4922 4366 4924
rect 4390 4922 4446 4924
rect 4150 4870 4176 4922
rect 4176 4870 4206 4922
rect 4230 4870 4240 4922
rect 4240 4870 4286 4922
rect 4310 4870 4356 4922
rect 4356 4870 4366 4922
rect 4390 4870 4420 4922
rect 4420 4870 4446 4922
rect 4150 4868 4206 4870
rect 4230 4868 4286 4870
rect 4310 4868 4366 4870
rect 4390 4868 4446 4870
rect 3352 4378 3408 4380
rect 3432 4378 3488 4380
rect 3512 4378 3568 4380
rect 3592 4378 3648 4380
rect 3352 4326 3378 4378
rect 3378 4326 3408 4378
rect 3432 4326 3442 4378
rect 3442 4326 3488 4378
rect 3512 4326 3558 4378
rect 3558 4326 3568 4378
rect 3592 4326 3622 4378
rect 3622 4326 3648 4378
rect 3352 4324 3408 4326
rect 3432 4324 3488 4326
rect 3512 4324 3568 4326
rect 3592 4324 3648 4326
rect 4150 3834 4206 3836
rect 4230 3834 4286 3836
rect 4310 3834 4366 3836
rect 4390 3834 4446 3836
rect 4150 3782 4176 3834
rect 4176 3782 4206 3834
rect 4230 3782 4240 3834
rect 4240 3782 4286 3834
rect 4310 3782 4356 3834
rect 4356 3782 4366 3834
rect 4390 3782 4420 3834
rect 4420 3782 4446 3834
rect 4150 3780 4206 3782
rect 4230 3780 4286 3782
rect 4310 3780 4366 3782
rect 4390 3780 4446 3782
rect 3352 3290 3408 3292
rect 3432 3290 3488 3292
rect 3512 3290 3568 3292
rect 3592 3290 3648 3292
rect 3352 3238 3378 3290
rect 3378 3238 3408 3290
rect 3432 3238 3442 3290
rect 3442 3238 3488 3290
rect 3512 3238 3558 3290
rect 3558 3238 3568 3290
rect 3592 3238 3622 3290
rect 3622 3238 3648 3290
rect 3352 3236 3408 3238
rect 3432 3236 3488 3238
rect 3512 3236 3568 3238
rect 3592 3236 3648 3238
rect 3352 2202 3408 2204
rect 3432 2202 3488 2204
rect 3512 2202 3568 2204
rect 3592 2202 3648 2204
rect 3352 2150 3378 2202
rect 3378 2150 3408 2202
rect 3432 2150 3442 2202
rect 3442 2150 3488 2202
rect 3512 2150 3558 2202
rect 3558 2150 3568 2202
rect 3592 2150 3622 2202
rect 3622 2150 3648 2202
rect 3352 2148 3408 2150
rect 3432 2148 3488 2150
rect 3512 2148 3568 2150
rect 3592 2148 3648 2150
rect 1754 1114 1810 1116
rect 1834 1114 1890 1116
rect 1914 1114 1970 1116
rect 1994 1114 2050 1116
rect 1754 1062 1780 1114
rect 1780 1062 1810 1114
rect 1834 1062 1844 1114
rect 1844 1062 1890 1114
rect 1914 1062 1960 1114
rect 1960 1062 1970 1114
rect 1994 1062 2024 1114
rect 2024 1062 2050 1114
rect 1754 1060 1810 1062
rect 1834 1060 1890 1062
rect 1914 1060 1970 1062
rect 1994 1060 2050 1062
rect 3352 1114 3408 1116
rect 3432 1114 3488 1116
rect 3512 1114 3568 1116
rect 3592 1114 3648 1116
rect 3352 1062 3378 1114
rect 3378 1062 3408 1114
rect 3432 1062 3442 1114
rect 3442 1062 3488 1114
rect 3512 1062 3558 1114
rect 3558 1062 3568 1114
rect 3592 1062 3622 1114
rect 3622 1062 3648 1114
rect 3352 1060 3408 1062
rect 3432 1060 3488 1062
rect 3512 1060 3568 1062
rect 3592 1060 3648 1062
rect 4150 2746 4206 2748
rect 4230 2746 4286 2748
rect 4310 2746 4366 2748
rect 4390 2746 4446 2748
rect 4150 2694 4176 2746
rect 4176 2694 4206 2746
rect 4230 2694 4240 2746
rect 4240 2694 4286 2746
rect 4310 2694 4356 2746
rect 4356 2694 4366 2746
rect 4390 2694 4420 2746
rect 4420 2694 4446 2746
rect 4150 2692 4206 2694
rect 4230 2692 4286 2694
rect 4310 2692 4366 2694
rect 4390 2692 4446 2694
rect 4802 6160 4858 6216
rect 4949 5466 5005 5468
rect 5029 5466 5085 5468
rect 5109 5466 5165 5468
rect 5189 5466 5245 5468
rect 4949 5414 4975 5466
rect 4975 5414 5005 5466
rect 5029 5414 5039 5466
rect 5039 5414 5085 5466
rect 5109 5414 5155 5466
rect 5155 5414 5165 5466
rect 5189 5414 5219 5466
rect 5219 5414 5245 5466
rect 4949 5412 5005 5414
rect 5029 5412 5085 5414
rect 5109 5412 5165 5414
rect 5189 5412 5245 5414
rect 5538 4800 5594 4856
rect 4949 4378 5005 4380
rect 5029 4378 5085 4380
rect 5109 4378 5165 4380
rect 5189 4378 5245 4380
rect 4949 4326 4975 4378
rect 4975 4326 5005 4378
rect 5029 4326 5039 4378
rect 5039 4326 5085 4378
rect 5109 4326 5155 4378
rect 5155 4326 5165 4378
rect 5189 4326 5219 4378
rect 5219 4326 5245 4378
rect 4949 4324 5005 4326
rect 5029 4324 5085 4326
rect 5109 4324 5165 4326
rect 5189 4324 5245 4326
rect 4618 2760 4674 2816
rect 4150 1658 4206 1660
rect 4230 1658 4286 1660
rect 4310 1658 4366 1660
rect 4390 1658 4446 1660
rect 4150 1606 4176 1658
rect 4176 1606 4206 1658
rect 4230 1606 4240 1658
rect 4240 1606 4286 1658
rect 4310 1606 4356 1658
rect 4356 1606 4366 1658
rect 4390 1606 4420 1658
rect 4420 1606 4446 1658
rect 4150 1604 4206 1606
rect 4230 1604 4286 1606
rect 4310 1604 4366 1606
rect 4390 1604 4446 1606
rect 4949 3290 5005 3292
rect 5029 3290 5085 3292
rect 5109 3290 5165 3292
rect 5189 3290 5245 3292
rect 4949 3238 4975 3290
rect 4975 3238 5005 3290
rect 5029 3238 5039 3290
rect 5039 3238 5085 3290
rect 5109 3238 5155 3290
rect 5155 3238 5165 3290
rect 5189 3238 5219 3290
rect 5219 3238 5245 3290
rect 4949 3236 5005 3238
rect 5029 3236 5085 3238
rect 5109 3236 5165 3238
rect 5189 3236 5245 3238
rect 4949 2202 5005 2204
rect 5029 2202 5085 2204
rect 5109 2202 5165 2204
rect 5189 2202 5245 2204
rect 4949 2150 4975 2202
rect 4975 2150 5005 2202
rect 5029 2150 5039 2202
rect 5039 2150 5085 2202
rect 5109 2150 5155 2202
rect 5155 2150 5165 2202
rect 5189 2150 5219 2202
rect 5219 2150 5245 2202
rect 4949 2148 5005 2150
rect 5029 2148 5085 2150
rect 5109 2148 5165 2150
rect 5189 2148 5245 2150
rect 5538 3440 5594 3496
rect 4949 1114 5005 1116
rect 5029 1114 5085 1116
rect 5109 1114 5165 1116
rect 5189 1114 5245 1116
rect 4949 1062 4975 1114
rect 4975 1062 5005 1114
rect 5029 1062 5039 1114
rect 5039 1062 5085 1114
rect 5109 1062 5155 1114
rect 5155 1062 5165 1114
rect 5189 1062 5219 1114
rect 5219 1062 5245 1114
rect 4949 1060 5005 1062
rect 5029 1060 5085 1062
rect 5109 1060 5165 1062
rect 5189 1060 5245 1062
rect 4710 720 4766 776
<< metal3 >>
rect 0 6218 800 6248
rect 4797 6218 4863 6221
rect 0 6216 4863 6218
rect 0 6160 4802 6216
rect 4858 6160 4863 6216
rect 0 6158 4863 6160
rect 0 6128 800 6158
rect 4797 6155 4863 6158
rect 0 5538 800 5568
rect 6200 5538 7000 5568
rect 0 5478 1594 5538
rect 0 5448 800 5478
rect 1534 5130 1594 5478
rect 5398 5478 7000 5538
rect 1742 5472 2062 5473
rect 1742 5408 1750 5472
rect 1814 5408 1830 5472
rect 1894 5408 1910 5472
rect 1974 5408 1990 5472
rect 2054 5408 2062 5472
rect 1742 5407 2062 5408
rect 3340 5472 3660 5473
rect 3340 5408 3348 5472
rect 3412 5408 3428 5472
rect 3492 5408 3508 5472
rect 3572 5408 3588 5472
rect 3652 5408 3660 5472
rect 3340 5407 3660 5408
rect 4937 5472 5257 5473
rect 4937 5408 4945 5472
rect 5009 5408 5025 5472
rect 5089 5408 5105 5472
rect 5169 5408 5185 5472
rect 5249 5408 5257 5472
rect 4937 5407 5257 5408
rect 2313 5266 2379 5269
rect 5398 5266 5458 5478
rect 6200 5448 7000 5478
rect 2313 5264 5458 5266
rect 2313 5208 2318 5264
rect 2374 5208 5458 5264
rect 2313 5206 5458 5208
rect 2313 5203 2379 5206
rect 4061 5130 4127 5133
rect 1534 5128 4127 5130
rect 1534 5072 4066 5128
rect 4122 5072 4127 5128
rect 1534 5070 4127 5072
rect 4061 5067 4127 5070
rect 2541 4928 2861 4929
rect 2541 4864 2549 4928
rect 2613 4864 2629 4928
rect 2693 4864 2709 4928
rect 2773 4864 2789 4928
rect 2853 4864 2861 4928
rect 2541 4863 2861 4864
rect 4138 4928 4458 4929
rect 4138 4864 4146 4928
rect 4210 4864 4226 4928
rect 4290 4864 4306 4928
rect 4370 4864 4386 4928
rect 4450 4864 4458 4928
rect 4138 4863 4458 4864
rect 5533 4858 5599 4861
rect 6200 4858 7000 4888
rect 5533 4856 7000 4858
rect 5533 4800 5538 4856
rect 5594 4800 7000 4856
rect 5533 4798 7000 4800
rect 5533 4795 5599 4798
rect 6200 4768 7000 4798
rect 1742 4384 2062 4385
rect 1742 4320 1750 4384
rect 1814 4320 1830 4384
rect 1894 4320 1910 4384
rect 1974 4320 1990 4384
rect 2054 4320 2062 4384
rect 1742 4319 2062 4320
rect 3340 4384 3660 4385
rect 3340 4320 3348 4384
rect 3412 4320 3428 4384
rect 3492 4320 3508 4384
rect 3572 4320 3588 4384
rect 3652 4320 3660 4384
rect 3340 4319 3660 4320
rect 4937 4384 5257 4385
rect 4937 4320 4945 4384
rect 5009 4320 5025 4384
rect 5089 4320 5105 4384
rect 5169 4320 5185 4384
rect 5249 4320 5257 4384
rect 4937 4319 5257 4320
rect 0 4178 800 4208
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4088 800 4118
rect 2773 4115 2839 4118
rect 2541 3840 2861 3841
rect 2541 3776 2549 3840
rect 2613 3776 2629 3840
rect 2693 3776 2709 3840
rect 2773 3776 2789 3840
rect 2853 3776 2861 3840
rect 2541 3775 2861 3776
rect 4138 3840 4458 3841
rect 4138 3776 4146 3840
rect 4210 3776 4226 3840
rect 4290 3776 4306 3840
rect 4370 3776 4386 3840
rect 4450 3776 4458 3840
rect 4138 3775 4458 3776
rect 0 3498 800 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 800 3438
rect 1669 3435 1735 3438
rect 5533 3498 5599 3501
rect 6200 3498 7000 3528
rect 5533 3496 7000 3498
rect 5533 3440 5538 3496
rect 5594 3440 7000 3496
rect 5533 3438 7000 3440
rect 5533 3435 5599 3438
rect 6200 3408 7000 3438
rect 1742 3296 2062 3297
rect 1742 3232 1750 3296
rect 1814 3232 1830 3296
rect 1894 3232 1910 3296
rect 1974 3232 1990 3296
rect 2054 3232 2062 3296
rect 1742 3231 2062 3232
rect 3340 3296 3660 3297
rect 3340 3232 3348 3296
rect 3412 3232 3428 3296
rect 3492 3232 3508 3296
rect 3572 3232 3588 3296
rect 3652 3232 3660 3296
rect 3340 3231 3660 3232
rect 4937 3296 5257 3297
rect 4937 3232 4945 3296
rect 5009 3232 5025 3296
rect 5089 3232 5105 3296
rect 5169 3232 5185 3296
rect 5249 3232 5257 3296
rect 4937 3231 5257 3232
rect 4613 2818 4679 2821
rect 6200 2818 7000 2848
rect 4613 2816 7000 2818
rect 4613 2760 4618 2816
rect 4674 2760 7000 2816
rect 4613 2758 7000 2760
rect 4613 2755 4679 2758
rect 2541 2752 2861 2753
rect 2541 2688 2549 2752
rect 2613 2688 2629 2752
rect 2693 2688 2709 2752
rect 2773 2688 2789 2752
rect 2853 2688 2861 2752
rect 2541 2687 2861 2688
rect 4138 2752 4458 2753
rect 4138 2688 4146 2752
rect 4210 2688 4226 2752
rect 4290 2688 4306 2752
rect 4370 2688 4386 2752
rect 4450 2688 4458 2752
rect 6200 2728 7000 2758
rect 4138 2687 4458 2688
rect 1742 2208 2062 2209
rect 0 2138 800 2168
rect 1742 2144 1750 2208
rect 1814 2144 1830 2208
rect 1894 2144 1910 2208
rect 1974 2144 1990 2208
rect 2054 2144 2062 2208
rect 1742 2143 2062 2144
rect 3340 2208 3660 2209
rect 3340 2144 3348 2208
rect 3412 2144 3428 2208
rect 3492 2144 3508 2208
rect 3572 2144 3588 2208
rect 3652 2144 3660 2208
rect 3340 2143 3660 2144
rect 4937 2208 5257 2209
rect 4937 2144 4945 2208
rect 5009 2144 5025 2208
rect 5089 2144 5105 2208
rect 5169 2144 5185 2208
rect 5249 2144 5257 2208
rect 4937 2143 5257 2144
rect 0 2078 1594 2138
rect 0 2048 800 2078
rect 1534 2002 1594 2078
rect 2773 2002 2839 2005
rect 1534 2000 2839 2002
rect 1534 1944 2778 2000
rect 2834 1944 2839 2000
rect 1534 1942 2839 1944
rect 2773 1939 2839 1942
rect 2541 1664 2861 1665
rect 2541 1600 2549 1664
rect 2613 1600 2629 1664
rect 2693 1600 2709 1664
rect 2773 1600 2789 1664
rect 2853 1600 2861 1664
rect 2541 1599 2861 1600
rect 4138 1664 4458 1665
rect 4138 1600 4146 1664
rect 4210 1600 4226 1664
rect 4290 1600 4306 1664
rect 4370 1600 4386 1664
rect 4450 1600 4458 1664
rect 4138 1599 4458 1600
rect 0 1458 800 1488
rect 1945 1458 2011 1461
rect 0 1456 2011 1458
rect 0 1400 1950 1456
rect 2006 1400 2011 1456
rect 0 1398 2011 1400
rect 0 1368 800 1398
rect 1945 1395 2011 1398
rect 2405 1458 2471 1461
rect 6200 1458 7000 1488
rect 2405 1456 7000 1458
rect 2405 1400 2410 1456
rect 2466 1400 7000 1456
rect 2405 1398 7000 1400
rect 2405 1395 2471 1398
rect 6200 1368 7000 1398
rect 1742 1120 2062 1121
rect 1742 1056 1750 1120
rect 1814 1056 1830 1120
rect 1894 1056 1910 1120
rect 1974 1056 1990 1120
rect 2054 1056 2062 1120
rect 1742 1055 2062 1056
rect 3340 1120 3660 1121
rect 3340 1056 3348 1120
rect 3412 1056 3428 1120
rect 3492 1056 3508 1120
rect 3572 1056 3588 1120
rect 3652 1056 3660 1120
rect 3340 1055 3660 1056
rect 4937 1120 5257 1121
rect 4937 1056 4945 1120
rect 5009 1056 5025 1120
rect 5089 1056 5105 1120
rect 5169 1056 5185 1120
rect 5249 1056 5257 1120
rect 4937 1055 5257 1056
rect 4705 778 4771 781
rect 6200 778 7000 808
rect 4705 776 7000 778
rect 4705 720 4710 776
rect 4766 720 7000 776
rect 4705 718 7000 720
rect 4705 715 4771 718
rect 6200 688 7000 718
<< via3 >>
rect 1750 5468 1814 5472
rect 1750 5412 1754 5468
rect 1754 5412 1810 5468
rect 1810 5412 1814 5468
rect 1750 5408 1814 5412
rect 1830 5468 1894 5472
rect 1830 5412 1834 5468
rect 1834 5412 1890 5468
rect 1890 5412 1894 5468
rect 1830 5408 1894 5412
rect 1910 5468 1974 5472
rect 1910 5412 1914 5468
rect 1914 5412 1970 5468
rect 1970 5412 1974 5468
rect 1910 5408 1974 5412
rect 1990 5468 2054 5472
rect 1990 5412 1994 5468
rect 1994 5412 2050 5468
rect 2050 5412 2054 5468
rect 1990 5408 2054 5412
rect 3348 5468 3412 5472
rect 3348 5412 3352 5468
rect 3352 5412 3408 5468
rect 3408 5412 3412 5468
rect 3348 5408 3412 5412
rect 3428 5468 3492 5472
rect 3428 5412 3432 5468
rect 3432 5412 3488 5468
rect 3488 5412 3492 5468
rect 3428 5408 3492 5412
rect 3508 5468 3572 5472
rect 3508 5412 3512 5468
rect 3512 5412 3568 5468
rect 3568 5412 3572 5468
rect 3508 5408 3572 5412
rect 3588 5468 3652 5472
rect 3588 5412 3592 5468
rect 3592 5412 3648 5468
rect 3648 5412 3652 5468
rect 3588 5408 3652 5412
rect 4945 5468 5009 5472
rect 4945 5412 4949 5468
rect 4949 5412 5005 5468
rect 5005 5412 5009 5468
rect 4945 5408 5009 5412
rect 5025 5468 5089 5472
rect 5025 5412 5029 5468
rect 5029 5412 5085 5468
rect 5085 5412 5089 5468
rect 5025 5408 5089 5412
rect 5105 5468 5169 5472
rect 5105 5412 5109 5468
rect 5109 5412 5165 5468
rect 5165 5412 5169 5468
rect 5105 5408 5169 5412
rect 5185 5468 5249 5472
rect 5185 5412 5189 5468
rect 5189 5412 5245 5468
rect 5245 5412 5249 5468
rect 5185 5408 5249 5412
rect 2549 4924 2613 4928
rect 2549 4868 2553 4924
rect 2553 4868 2609 4924
rect 2609 4868 2613 4924
rect 2549 4864 2613 4868
rect 2629 4924 2693 4928
rect 2629 4868 2633 4924
rect 2633 4868 2689 4924
rect 2689 4868 2693 4924
rect 2629 4864 2693 4868
rect 2709 4924 2773 4928
rect 2709 4868 2713 4924
rect 2713 4868 2769 4924
rect 2769 4868 2773 4924
rect 2709 4864 2773 4868
rect 2789 4924 2853 4928
rect 2789 4868 2793 4924
rect 2793 4868 2849 4924
rect 2849 4868 2853 4924
rect 2789 4864 2853 4868
rect 4146 4924 4210 4928
rect 4146 4868 4150 4924
rect 4150 4868 4206 4924
rect 4206 4868 4210 4924
rect 4146 4864 4210 4868
rect 4226 4924 4290 4928
rect 4226 4868 4230 4924
rect 4230 4868 4286 4924
rect 4286 4868 4290 4924
rect 4226 4864 4290 4868
rect 4306 4924 4370 4928
rect 4306 4868 4310 4924
rect 4310 4868 4366 4924
rect 4366 4868 4370 4924
rect 4306 4864 4370 4868
rect 4386 4924 4450 4928
rect 4386 4868 4390 4924
rect 4390 4868 4446 4924
rect 4446 4868 4450 4924
rect 4386 4864 4450 4868
rect 1750 4380 1814 4384
rect 1750 4324 1754 4380
rect 1754 4324 1810 4380
rect 1810 4324 1814 4380
rect 1750 4320 1814 4324
rect 1830 4380 1894 4384
rect 1830 4324 1834 4380
rect 1834 4324 1890 4380
rect 1890 4324 1894 4380
rect 1830 4320 1894 4324
rect 1910 4380 1974 4384
rect 1910 4324 1914 4380
rect 1914 4324 1970 4380
rect 1970 4324 1974 4380
rect 1910 4320 1974 4324
rect 1990 4380 2054 4384
rect 1990 4324 1994 4380
rect 1994 4324 2050 4380
rect 2050 4324 2054 4380
rect 1990 4320 2054 4324
rect 3348 4380 3412 4384
rect 3348 4324 3352 4380
rect 3352 4324 3408 4380
rect 3408 4324 3412 4380
rect 3348 4320 3412 4324
rect 3428 4380 3492 4384
rect 3428 4324 3432 4380
rect 3432 4324 3488 4380
rect 3488 4324 3492 4380
rect 3428 4320 3492 4324
rect 3508 4380 3572 4384
rect 3508 4324 3512 4380
rect 3512 4324 3568 4380
rect 3568 4324 3572 4380
rect 3508 4320 3572 4324
rect 3588 4380 3652 4384
rect 3588 4324 3592 4380
rect 3592 4324 3648 4380
rect 3648 4324 3652 4380
rect 3588 4320 3652 4324
rect 4945 4380 5009 4384
rect 4945 4324 4949 4380
rect 4949 4324 5005 4380
rect 5005 4324 5009 4380
rect 4945 4320 5009 4324
rect 5025 4380 5089 4384
rect 5025 4324 5029 4380
rect 5029 4324 5085 4380
rect 5085 4324 5089 4380
rect 5025 4320 5089 4324
rect 5105 4380 5169 4384
rect 5105 4324 5109 4380
rect 5109 4324 5165 4380
rect 5165 4324 5169 4380
rect 5105 4320 5169 4324
rect 5185 4380 5249 4384
rect 5185 4324 5189 4380
rect 5189 4324 5245 4380
rect 5245 4324 5249 4380
rect 5185 4320 5249 4324
rect 2549 3836 2613 3840
rect 2549 3780 2553 3836
rect 2553 3780 2609 3836
rect 2609 3780 2613 3836
rect 2549 3776 2613 3780
rect 2629 3836 2693 3840
rect 2629 3780 2633 3836
rect 2633 3780 2689 3836
rect 2689 3780 2693 3836
rect 2629 3776 2693 3780
rect 2709 3836 2773 3840
rect 2709 3780 2713 3836
rect 2713 3780 2769 3836
rect 2769 3780 2773 3836
rect 2709 3776 2773 3780
rect 2789 3836 2853 3840
rect 2789 3780 2793 3836
rect 2793 3780 2849 3836
rect 2849 3780 2853 3836
rect 2789 3776 2853 3780
rect 4146 3836 4210 3840
rect 4146 3780 4150 3836
rect 4150 3780 4206 3836
rect 4206 3780 4210 3836
rect 4146 3776 4210 3780
rect 4226 3836 4290 3840
rect 4226 3780 4230 3836
rect 4230 3780 4286 3836
rect 4286 3780 4290 3836
rect 4226 3776 4290 3780
rect 4306 3836 4370 3840
rect 4306 3780 4310 3836
rect 4310 3780 4366 3836
rect 4366 3780 4370 3836
rect 4306 3776 4370 3780
rect 4386 3836 4450 3840
rect 4386 3780 4390 3836
rect 4390 3780 4446 3836
rect 4446 3780 4450 3836
rect 4386 3776 4450 3780
rect 1750 3292 1814 3296
rect 1750 3236 1754 3292
rect 1754 3236 1810 3292
rect 1810 3236 1814 3292
rect 1750 3232 1814 3236
rect 1830 3292 1894 3296
rect 1830 3236 1834 3292
rect 1834 3236 1890 3292
rect 1890 3236 1894 3292
rect 1830 3232 1894 3236
rect 1910 3292 1974 3296
rect 1910 3236 1914 3292
rect 1914 3236 1970 3292
rect 1970 3236 1974 3292
rect 1910 3232 1974 3236
rect 1990 3292 2054 3296
rect 1990 3236 1994 3292
rect 1994 3236 2050 3292
rect 2050 3236 2054 3292
rect 1990 3232 2054 3236
rect 3348 3292 3412 3296
rect 3348 3236 3352 3292
rect 3352 3236 3408 3292
rect 3408 3236 3412 3292
rect 3348 3232 3412 3236
rect 3428 3292 3492 3296
rect 3428 3236 3432 3292
rect 3432 3236 3488 3292
rect 3488 3236 3492 3292
rect 3428 3232 3492 3236
rect 3508 3292 3572 3296
rect 3508 3236 3512 3292
rect 3512 3236 3568 3292
rect 3568 3236 3572 3292
rect 3508 3232 3572 3236
rect 3588 3292 3652 3296
rect 3588 3236 3592 3292
rect 3592 3236 3648 3292
rect 3648 3236 3652 3292
rect 3588 3232 3652 3236
rect 4945 3292 5009 3296
rect 4945 3236 4949 3292
rect 4949 3236 5005 3292
rect 5005 3236 5009 3292
rect 4945 3232 5009 3236
rect 5025 3292 5089 3296
rect 5025 3236 5029 3292
rect 5029 3236 5085 3292
rect 5085 3236 5089 3292
rect 5025 3232 5089 3236
rect 5105 3292 5169 3296
rect 5105 3236 5109 3292
rect 5109 3236 5165 3292
rect 5165 3236 5169 3292
rect 5105 3232 5169 3236
rect 5185 3292 5249 3296
rect 5185 3236 5189 3292
rect 5189 3236 5245 3292
rect 5245 3236 5249 3292
rect 5185 3232 5249 3236
rect 2549 2748 2613 2752
rect 2549 2692 2553 2748
rect 2553 2692 2609 2748
rect 2609 2692 2613 2748
rect 2549 2688 2613 2692
rect 2629 2748 2693 2752
rect 2629 2692 2633 2748
rect 2633 2692 2689 2748
rect 2689 2692 2693 2748
rect 2629 2688 2693 2692
rect 2709 2748 2773 2752
rect 2709 2692 2713 2748
rect 2713 2692 2769 2748
rect 2769 2692 2773 2748
rect 2709 2688 2773 2692
rect 2789 2748 2853 2752
rect 2789 2692 2793 2748
rect 2793 2692 2849 2748
rect 2849 2692 2853 2748
rect 2789 2688 2853 2692
rect 4146 2748 4210 2752
rect 4146 2692 4150 2748
rect 4150 2692 4206 2748
rect 4206 2692 4210 2748
rect 4146 2688 4210 2692
rect 4226 2748 4290 2752
rect 4226 2692 4230 2748
rect 4230 2692 4286 2748
rect 4286 2692 4290 2748
rect 4226 2688 4290 2692
rect 4306 2748 4370 2752
rect 4306 2692 4310 2748
rect 4310 2692 4366 2748
rect 4366 2692 4370 2748
rect 4306 2688 4370 2692
rect 4386 2748 4450 2752
rect 4386 2692 4390 2748
rect 4390 2692 4446 2748
rect 4446 2692 4450 2748
rect 4386 2688 4450 2692
rect 1750 2204 1814 2208
rect 1750 2148 1754 2204
rect 1754 2148 1810 2204
rect 1810 2148 1814 2204
rect 1750 2144 1814 2148
rect 1830 2204 1894 2208
rect 1830 2148 1834 2204
rect 1834 2148 1890 2204
rect 1890 2148 1894 2204
rect 1830 2144 1894 2148
rect 1910 2204 1974 2208
rect 1910 2148 1914 2204
rect 1914 2148 1970 2204
rect 1970 2148 1974 2204
rect 1910 2144 1974 2148
rect 1990 2204 2054 2208
rect 1990 2148 1994 2204
rect 1994 2148 2050 2204
rect 2050 2148 2054 2204
rect 1990 2144 2054 2148
rect 3348 2204 3412 2208
rect 3348 2148 3352 2204
rect 3352 2148 3408 2204
rect 3408 2148 3412 2204
rect 3348 2144 3412 2148
rect 3428 2204 3492 2208
rect 3428 2148 3432 2204
rect 3432 2148 3488 2204
rect 3488 2148 3492 2204
rect 3428 2144 3492 2148
rect 3508 2204 3572 2208
rect 3508 2148 3512 2204
rect 3512 2148 3568 2204
rect 3568 2148 3572 2204
rect 3508 2144 3572 2148
rect 3588 2204 3652 2208
rect 3588 2148 3592 2204
rect 3592 2148 3648 2204
rect 3648 2148 3652 2204
rect 3588 2144 3652 2148
rect 4945 2204 5009 2208
rect 4945 2148 4949 2204
rect 4949 2148 5005 2204
rect 5005 2148 5009 2204
rect 4945 2144 5009 2148
rect 5025 2204 5089 2208
rect 5025 2148 5029 2204
rect 5029 2148 5085 2204
rect 5085 2148 5089 2204
rect 5025 2144 5089 2148
rect 5105 2204 5169 2208
rect 5105 2148 5109 2204
rect 5109 2148 5165 2204
rect 5165 2148 5169 2204
rect 5105 2144 5169 2148
rect 5185 2204 5249 2208
rect 5185 2148 5189 2204
rect 5189 2148 5245 2204
rect 5245 2148 5249 2204
rect 5185 2144 5249 2148
rect 2549 1660 2613 1664
rect 2549 1604 2553 1660
rect 2553 1604 2609 1660
rect 2609 1604 2613 1660
rect 2549 1600 2613 1604
rect 2629 1660 2693 1664
rect 2629 1604 2633 1660
rect 2633 1604 2689 1660
rect 2689 1604 2693 1660
rect 2629 1600 2693 1604
rect 2709 1660 2773 1664
rect 2709 1604 2713 1660
rect 2713 1604 2769 1660
rect 2769 1604 2773 1660
rect 2709 1600 2773 1604
rect 2789 1660 2853 1664
rect 2789 1604 2793 1660
rect 2793 1604 2849 1660
rect 2849 1604 2853 1660
rect 2789 1600 2853 1604
rect 4146 1660 4210 1664
rect 4146 1604 4150 1660
rect 4150 1604 4206 1660
rect 4206 1604 4210 1660
rect 4146 1600 4210 1604
rect 4226 1660 4290 1664
rect 4226 1604 4230 1660
rect 4230 1604 4286 1660
rect 4286 1604 4290 1660
rect 4226 1600 4290 1604
rect 4306 1660 4370 1664
rect 4306 1604 4310 1660
rect 4310 1604 4366 1660
rect 4366 1604 4370 1660
rect 4306 1600 4370 1604
rect 4386 1660 4450 1664
rect 4386 1604 4390 1660
rect 4390 1604 4446 1660
rect 4446 1604 4450 1660
rect 4386 1600 4450 1604
rect 1750 1116 1814 1120
rect 1750 1060 1754 1116
rect 1754 1060 1810 1116
rect 1810 1060 1814 1116
rect 1750 1056 1814 1060
rect 1830 1116 1894 1120
rect 1830 1060 1834 1116
rect 1834 1060 1890 1116
rect 1890 1060 1894 1116
rect 1830 1056 1894 1060
rect 1910 1116 1974 1120
rect 1910 1060 1914 1116
rect 1914 1060 1970 1116
rect 1970 1060 1974 1116
rect 1910 1056 1974 1060
rect 1990 1116 2054 1120
rect 1990 1060 1994 1116
rect 1994 1060 2050 1116
rect 2050 1060 2054 1116
rect 1990 1056 2054 1060
rect 3348 1116 3412 1120
rect 3348 1060 3352 1116
rect 3352 1060 3408 1116
rect 3408 1060 3412 1116
rect 3348 1056 3412 1060
rect 3428 1116 3492 1120
rect 3428 1060 3432 1116
rect 3432 1060 3488 1116
rect 3488 1060 3492 1116
rect 3428 1056 3492 1060
rect 3508 1116 3572 1120
rect 3508 1060 3512 1116
rect 3512 1060 3568 1116
rect 3568 1060 3572 1116
rect 3508 1056 3572 1060
rect 3588 1116 3652 1120
rect 3588 1060 3592 1116
rect 3592 1060 3648 1116
rect 3648 1060 3652 1116
rect 3588 1056 3652 1060
rect 4945 1116 5009 1120
rect 4945 1060 4949 1116
rect 4949 1060 5005 1116
rect 5005 1060 5009 1116
rect 4945 1056 5009 1060
rect 5025 1116 5089 1120
rect 5025 1060 5029 1116
rect 5029 1060 5085 1116
rect 5085 1060 5089 1116
rect 5025 1056 5089 1060
rect 5105 1116 5169 1120
rect 5105 1060 5109 1116
rect 5109 1060 5165 1116
rect 5165 1060 5169 1116
rect 5105 1056 5169 1060
rect 5185 1116 5249 1120
rect 5185 1060 5189 1116
rect 5189 1060 5245 1116
rect 5245 1060 5249 1116
rect 5185 1056 5249 1060
<< metal4 >>
rect 1742 5472 2063 5488
rect 1742 5408 1750 5472
rect 1814 5408 1830 5472
rect 1894 5408 1910 5472
rect 1974 5408 1990 5472
rect 2054 5408 2063 5472
rect 1742 5178 2063 5408
rect 1742 4942 1784 5178
rect 2020 4942 2063 5178
rect 1742 4384 2063 4942
rect 1742 4320 1750 4384
rect 1814 4320 1830 4384
rect 1894 4320 1910 4384
rect 1974 4320 1990 4384
rect 2054 4320 2063 4384
rect 1742 3570 2063 4320
rect 1742 3334 1784 3570
rect 2020 3334 2063 3570
rect 1742 3296 2063 3334
rect 1742 3232 1750 3296
rect 1814 3232 1830 3296
rect 1894 3232 1910 3296
rect 1974 3232 1990 3296
rect 2054 3232 2063 3296
rect 1742 2208 2063 3232
rect 1742 2144 1750 2208
rect 1814 2144 1830 2208
rect 1894 2144 1910 2208
rect 1974 2144 1990 2208
rect 2054 2144 2063 2208
rect 1742 1962 2063 2144
rect 1742 1726 1784 1962
rect 2020 1726 2063 1962
rect 1742 1120 2063 1726
rect 1742 1056 1750 1120
rect 1814 1056 1830 1120
rect 1894 1056 1910 1120
rect 1974 1056 1990 1120
rect 2054 1056 2063 1120
rect 1742 1040 2063 1056
rect 2541 4928 2861 5488
rect 2541 4864 2549 4928
rect 2613 4864 2629 4928
rect 2693 4864 2709 4928
rect 2773 4864 2789 4928
rect 2853 4864 2861 4928
rect 2541 4374 2861 4864
rect 2541 4138 2583 4374
rect 2819 4138 2861 4374
rect 2541 3840 2861 4138
rect 2541 3776 2549 3840
rect 2613 3776 2629 3840
rect 2693 3776 2709 3840
rect 2773 3776 2789 3840
rect 2853 3776 2861 3840
rect 2541 2766 2861 3776
rect 2541 2752 2583 2766
rect 2819 2752 2861 2766
rect 2541 2688 2549 2752
rect 2853 2688 2861 2752
rect 2541 2530 2583 2688
rect 2819 2530 2861 2688
rect 2541 1664 2861 2530
rect 2541 1600 2549 1664
rect 2613 1600 2629 1664
rect 2693 1600 2709 1664
rect 2773 1600 2789 1664
rect 2853 1600 2861 1664
rect 2541 1040 2861 1600
rect 3340 5472 3660 5488
rect 3340 5408 3348 5472
rect 3412 5408 3428 5472
rect 3492 5408 3508 5472
rect 3572 5408 3588 5472
rect 3652 5408 3660 5472
rect 3340 5178 3660 5408
rect 3340 4942 3382 5178
rect 3618 4942 3660 5178
rect 3340 4384 3660 4942
rect 3340 4320 3348 4384
rect 3412 4320 3428 4384
rect 3492 4320 3508 4384
rect 3572 4320 3588 4384
rect 3652 4320 3660 4384
rect 3340 3570 3660 4320
rect 3340 3334 3382 3570
rect 3618 3334 3660 3570
rect 3340 3296 3660 3334
rect 3340 3232 3348 3296
rect 3412 3232 3428 3296
rect 3492 3232 3508 3296
rect 3572 3232 3588 3296
rect 3652 3232 3660 3296
rect 3340 2208 3660 3232
rect 3340 2144 3348 2208
rect 3412 2144 3428 2208
rect 3492 2144 3508 2208
rect 3572 2144 3588 2208
rect 3652 2144 3660 2208
rect 3340 1962 3660 2144
rect 3340 1726 3382 1962
rect 3618 1726 3660 1962
rect 3340 1120 3660 1726
rect 3340 1056 3348 1120
rect 3412 1056 3428 1120
rect 3492 1056 3508 1120
rect 3572 1056 3588 1120
rect 3652 1056 3660 1120
rect 3340 1040 3660 1056
rect 4138 4928 4459 5488
rect 4138 4864 4146 4928
rect 4210 4864 4226 4928
rect 4290 4864 4306 4928
rect 4370 4864 4386 4928
rect 4450 4864 4459 4928
rect 4138 4374 4459 4864
rect 4138 4138 4180 4374
rect 4416 4138 4459 4374
rect 4138 3840 4459 4138
rect 4138 3776 4146 3840
rect 4210 3776 4226 3840
rect 4290 3776 4306 3840
rect 4370 3776 4386 3840
rect 4450 3776 4459 3840
rect 4138 2766 4459 3776
rect 4138 2752 4180 2766
rect 4416 2752 4459 2766
rect 4138 2688 4146 2752
rect 4450 2688 4459 2752
rect 4138 2530 4180 2688
rect 4416 2530 4459 2688
rect 4138 1664 4459 2530
rect 4138 1600 4146 1664
rect 4210 1600 4226 1664
rect 4290 1600 4306 1664
rect 4370 1600 4386 1664
rect 4450 1600 4459 1664
rect 4138 1040 4459 1600
rect 4937 5472 5257 5488
rect 4937 5408 4945 5472
rect 5009 5408 5025 5472
rect 5089 5408 5105 5472
rect 5169 5408 5185 5472
rect 5249 5408 5257 5472
rect 4937 5178 5257 5408
rect 4937 4942 4979 5178
rect 5215 4942 5257 5178
rect 4937 4384 5257 4942
rect 4937 4320 4945 4384
rect 5009 4320 5025 4384
rect 5089 4320 5105 4384
rect 5169 4320 5185 4384
rect 5249 4320 5257 4384
rect 4937 3570 5257 4320
rect 4937 3334 4979 3570
rect 5215 3334 5257 3570
rect 4937 3296 5257 3334
rect 4937 3232 4945 3296
rect 5009 3232 5025 3296
rect 5089 3232 5105 3296
rect 5169 3232 5185 3296
rect 5249 3232 5257 3296
rect 4937 2208 5257 3232
rect 4937 2144 4945 2208
rect 5009 2144 5025 2208
rect 5089 2144 5105 2208
rect 5169 2144 5185 2208
rect 5249 2144 5257 2208
rect 4937 1962 5257 2144
rect 4937 1726 4979 1962
rect 5215 1726 5257 1962
rect 4937 1120 5257 1726
rect 4937 1056 4945 1120
rect 5009 1056 5025 1120
rect 5089 1056 5105 1120
rect 5169 1056 5185 1120
rect 5249 1056 5257 1120
rect 4937 1040 5257 1056
<< via4 >>
rect 1784 4942 2020 5178
rect 1784 3334 2020 3570
rect 1784 1726 2020 1962
rect 2583 4138 2819 4374
rect 2583 2752 2819 2766
rect 2583 2688 2613 2752
rect 2613 2688 2629 2752
rect 2629 2688 2693 2752
rect 2693 2688 2709 2752
rect 2709 2688 2773 2752
rect 2773 2688 2789 2752
rect 2789 2688 2819 2752
rect 2583 2530 2819 2688
rect 3382 4942 3618 5178
rect 3382 3334 3618 3570
rect 3382 1726 3618 1962
rect 4180 4138 4416 4374
rect 4180 2752 4416 2766
rect 4180 2688 4210 2752
rect 4210 2688 4226 2752
rect 4226 2688 4290 2752
rect 4290 2688 4306 2752
rect 4306 2688 4370 2752
rect 4370 2688 4386 2752
rect 4386 2688 4416 2752
rect 4180 2530 4416 2688
rect 4979 4942 5215 5178
rect 4979 3334 5215 3570
rect 4979 1726 5215 1962
<< metal5 >>
rect 1104 5178 5888 5220
rect 1104 4942 1784 5178
rect 2020 4942 3382 5178
rect 3618 4942 4979 5178
rect 5215 4942 5888 5178
rect 1104 4900 5888 4942
rect 1104 4374 5888 4416
rect 1104 4138 2583 4374
rect 2819 4138 4180 4374
rect 4416 4138 5888 4374
rect 1104 4096 5888 4138
rect 1104 3570 5888 3612
rect 1104 3334 1784 3570
rect 2020 3334 3382 3570
rect 3618 3334 4979 3570
rect 5215 3334 5888 3570
rect 1104 3292 5888 3334
rect 1104 2766 5888 2808
rect 1104 2530 2583 2766
rect 2819 2530 4180 2766
rect 4416 2530 5888 2766
rect 1104 2488 5888 2530
rect 1104 1962 5888 2004
rect 1104 1726 1784 1962
rect 2020 1726 3382 1962
rect 3618 1726 4979 1962
rect 5215 1726 5888 1962
rect 1104 1684 5888 1726
use sky130_fd_sc_hd__fill_1  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 1380 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1622467964
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[23\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 1472 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 1748 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[28\]
timestamp 1622467964
transform -1 0 2484 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[1\]
timestamp 1622467964
transform -1 0 2208 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[15\]
timestamp 1622467964
transform 1 0 1932 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 2208 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 1622467964
transform 1 0 1380 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[11\]
timestamp 1622467964
transform 1 0 2576 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[21\]
timestamp 1622467964
transform -1 0 3128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[7\]
timestamp 1622467964
transform 1 0 2760 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15
timestamp 1622467964
transform 1 0 2484 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1622467964
transform 1 0 3128 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 3036 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 3772 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1622467964
transform 1 0 3680 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 3864 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp 1622467964
transform 1 0 4600 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_33
timestamp 1622467964
transform 1 0 4140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[25\]
timestamp 1622467964
transform 1 0 5152 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[9\]
timestamp 1622467964
transform -1 0 5152 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1622467964
transform -1 0 5888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1622467964
transform -1 0 5888 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47
timestamp 1622467964
transform 1 0 5428 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1622467964
transform 1 0 5244 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[12\]
timestamp 1622467964
transform -1 0 1932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[17\]
timestamp 1622467964
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1622467964
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_9
timestamp 1622467964
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1622467964
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1622467964
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1622467964
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[8\]
timestamp 1622467964
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1622467964
transform -1 0 5888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1622467964
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1622467964
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1622467964
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[16\]
timestamp 1622467964
transform -1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1622467964
transform 1 0 2484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 1622467964
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[4\]
timestamp 1622467964
transform -1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1622467964
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1622467964
transform 1 0 4232 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1622467964
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[13\]
timestamp 1622467964
transform -1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1622467964
transform -1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_42
timestamp 1622467964
transform 1 0 4968 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1622467964
transform 1 0 5520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[10\]
timestamp 1622467964
transform -1 0 1932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[18\]
timestamp 1622467964
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[2\]
timestamp 1622467964
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[31\]
timestamp 1622467964
transform 1 0 2208 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1622467964
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[14\]
timestamp 1622467964
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1622467964
transform 1 0 2760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[22\]
timestamp 1622467964
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[24\]
timestamp 1622467964
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1622467964
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_26
timestamp 1622467964
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_33
timestamp 1622467964
transform 1 0 4140 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_38
timestamp 1622467964
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[20\]
timestamp 1622467964
transform -1 0 5060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[27\]
timestamp 1622467964
transform -1 0 5612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1622467964
transform -1 0 5888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_43
timestamp 1622467964
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[29\]
timestamp 1622467964
transform 1 0 1840 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[5\]
timestamp 1622467964
transform -1 0 2392 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1622467964
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1622467964
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1622467964
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_14
timestamp 1622467964
transform 1 0 2392 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[0\]
timestamp 1622467964
transform -1 0 4876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[3\]
timestamp 1622467964
transform -1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[6\]
timestamp 1622467964
transform 1 0 3588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1622467964
transform 1 0 3496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp 1622467964
transform 1 0 3864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1622467964
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[19\]
timestamp 1622467964
transform -1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[26\]
timestamp 1622467964
transform 1 0 5336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1622467964
transform -1 0 5888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1622467964
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1622467964
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1622467964
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1622467964
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1622467964
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1622467964
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1622467964
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[30\]
timestamp 1622467964
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1622467964
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1622467964
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1622467964
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_30
timestamp 1622467964
transform 1 0 3864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_36
timestamp 1622467964
transform 1 0 4416 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1622467964
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1622467964
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1622467964
transform -1 0 5888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1622467964
transform -1 0 5888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1622467964
transform 1 0 5520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_42
timestamp 1622467964
transform 1 0 4968 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_48
timestamp 1622467964
transform 1 0 5520 0 1 4896
box -38 -48 130 592
<< labels >>
rlabel metal2 s 938 0 994 800 6 mask_rev[0]
port 0 nsew signal tristate
rlabel metal2 s 1398 6200 1454 7000 6 mask_rev[10]
port 1 nsew signal tristate
rlabel metal2 s 2778 6200 2834 7000 6 mask_rev[11]
port 2 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 mask_rev[12]
port 3 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 mask_rev[13]
port 4 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 mask_rev[14]
port 5 nsew signal tristate
rlabel metal2 s 3238 6200 3294 7000 6 mask_rev[15]
port 6 nsew signal tristate
rlabel metal2 s 1858 6200 1914 7000 6 mask_rev[16]
port 7 nsew signal tristate
rlabel metal2 s 5538 6200 5594 7000 6 mask_rev[17]
port 8 nsew signal tristate
rlabel metal2 s 4618 6200 4674 7000 6 mask_rev[18]
port 9 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 mask_rev[19]
port 10 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 mask_rev[1]
port 11 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 mask_rev[20]
port 12 nsew signal tristate
rlabel metal2 s 2318 0 2374 800 6 mask_rev[21]
port 13 nsew signal tristate
rlabel metal3 s 6200 688 7000 808 6 mask_rev[22]
port 14 nsew signal tristate
rlabel metal3 s 6200 5448 7000 5568 6 mask_rev[23]
port 15 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 mask_rev[24]
port 16 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 mask_rev[25]
port 17 nsew signal tristate
rlabel metal3 s 6200 4768 7000 4888 6 mask_rev[26]
port 18 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 mask_rev[27]
port 19 nsew signal tristate
rlabel metal2 s 478 0 534 800 6 mask_rev[28]
port 20 nsew signal tristate
rlabel metal3 s 6200 1368 7000 1488 6 mask_rev[29]
port 21 nsew signal tristate
rlabel metal2 s 6458 6200 6514 7000 6 mask_rev[2]
port 22 nsew signal tristate
rlabel metal3 s 6200 2728 7000 2848 6 mask_rev[30]
port 23 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 mask_rev[31]
port 24 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 mask_rev[3]
port 25 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 mask_rev[4]
port 26 nsew signal tristate
rlabel metal2 s 938 6200 994 7000 6 mask_rev[5]
port 27 nsew signal tristate
rlabel metal2 s 5998 6200 6054 7000 6 mask_rev[6]
port 28 nsew signal tristate
rlabel metal2 s 4158 6200 4214 7000 6 mask_rev[7]
port 29 nsew signal tristate
rlabel metal3 s 6200 3408 7000 3528 6 mask_rev[8]
port 30 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 mask_rev[9]
port 31 nsew signal tristate
rlabel metal4 s 4937 1040 5257 5488 6 VPWR
port 32 nsew power bidirectional
rlabel metal4 s 3340 1040 3660 5488 6 VPWR
port 33 nsew power bidirectional
rlabel metal4 s 1743 1040 2063 5488 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1104 4900 5888 5220 6 VPWR
port 35 nsew power bidirectional
rlabel metal5 s 1104 3292 5888 3612 6 VPWR
port 36 nsew power bidirectional
rlabel metal5 s 1104 1684 5888 2004 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 4139 1040 4459 5488 6 VGND
port 38 nsew ground bidirectional
rlabel metal4 s 2541 1040 2861 5488 6 VGND
port 39 nsew ground bidirectional
rlabel metal5 s 1104 4096 5888 4416 6 VGND
port 40 nsew ground bidirectional
rlabel metal5 s 1104 2488 5888 2808 6 VGND
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7000 7000
<< end >>
