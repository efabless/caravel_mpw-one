* SKY130 Spice File.
* Number of bins: 1
.param
+ sky130_fd_pr__special_nfet_pass_flash__tox_mult = 0.9635
+ sky130_fd_pr__special_nfet_pass_flash__ajunction_mult = 8.4039e-1
+ sky130_fd_pr__special_nfet_pass_flash__pjunction_mult = 8.6147e-1
+ sky130_fd_pr__special_nfet_pass_flash__overlap_mult = 0.80232
+ sky130_fd_pr__special_nfet_pass_flash__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_pass_flash__wint_diff = -2.252e-8
+ sky130_fd_pr__special_nfet_pass_flash__dwg_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nlx_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt1l_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dlc_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_pass_flash__dwc_diff = -2.252e-8
*
* sky130_fd_pr__special_nfet_pass_flash, Bin 000, W = 0.45, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0 = -2.5324e-1
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_0 = 9.901e-2
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_0 = -0.00069863
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0 = -17497.0
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0 = -0.37718
*
* sky130_fd_pr__special_nfet_pass_flash, Bin 001, W = 0.35, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1 = -1.7722e-1
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1 = 2.9082e-2
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_1 = -8.7697e-3
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1 = -1.0357e+4
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1 = -2.4437e-1
* Number of bins: 1
.param
+ sky130_fd_pr__special_nfet_pass__tox_mult = 0.9635
+ sky130_fd_pr__special_nfet_pass__ajunction_mult = 8.4039e-1
+ sky130_fd_pr__special_nfet_pass__pjunction_mult = 8.6147e-1
+ sky130_fd_pr__special_nfet_pass__overlap_mult = 0.95013
+ sky130_fd_pr__special_nfet_pass__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_pass__wint_diff = -2.252e-8
+ sky130_fd_pr__special_nfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__kt1l_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__dlc_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_pass__dwc_diff = -2.252e-8
*
* sky130_fd_pr__special_nfet_pass, Bin 000, W = 0.14, L = 0.15
* ----------------------------------
+ sky130_fd_pr__special_nfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__u0_diff_0 = -0.0094635
+ sky130_fd_pr__special_nfet_pass__vth0_diff_0 = -0.14783
+ sky130_fd_pr__special_nfet_pass__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__voff_diff_0 = 0.0
* Number of bins: 1
.param
+ sky130_fd_pr__special_nfet_latch__tox_mult = 0.9635
+ sky130_fd_pr__special_nfet_latch__ajunction_mult = 8.4039e-1
+ sky130_fd_pr__special_nfet_latch__pjunction_mult = 8.6147e-1
+ sky130_fd_pr__special_nfet_latch__overlap_mult = 0.95013
+ sky130_fd_pr__special_nfet_latch__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_latch__wint_diff = -2.252e-8
+ sky130_fd_pr__special_nfet_latch__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__dvt1_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__dlc_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_latch__dwc_diff = -2.252e-8
*
* sky130_fd_pr__special_nfet_latch, Bin 000, W = 0.21, L = 0.15
* --------------------------------
+ sky130_fd_pr__special_nfet_latch__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__u0_diff_0 = -0.0088858
+ sky130_fd_pr__special_nfet_latch__vth0_diff_0 = -0.10936
+ sky130_fd_pr__special_nfet_latch__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__nfactor_diff_0 = 0.0
* Number of bins: 1
.param
+ sky130_fd_pr__special_pfet_pass__tox_mult = 0.9635
+ sky130_fd_pr__special_pfet_pass__ajunction_mult = 9.3001e-1
+ sky130_fd_pr__special_pfet_pass__pjunction_mult = 9.3439e-1
+ sky130_fd_pr__special_pfet_pass__overlap_mult = 8.8516e-1
+ sky130_fd_pr__special_pfet_pass__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_pfet_pass__wint_diff = -2.252e-8
+ sky130_fd_pr__special_pfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__dvt0_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cit_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cdsc_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cdscb_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cdscd_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__kt2_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__kt1l_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__dlc_diff = 1.21275e-8
+ sky130_fd_pr__special_pfet_pass__dwc_diff = -2.252e-8
*
* sky130_fd_pr__special_pfet_pass, Bin 000, W = 0.14, L = 0.15
* --------------------------------
+ sky130_fd_pr__special_pfet_pass__voff_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__vth0_diff_0 = 0.19102
+ sky130_fd_pr__special_pfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__u0_diff_0 = -0.001847
+ sky130_fd_pr__special_pfet_pass__rdsw_diff_0 = 0.0
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_latch__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_flash__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_pfet_pass__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_lvt__ff.corner.spice"
